magic
tech sky130A
magscale 1 2
timestamp 1682557711
<< viali >>
rect 25789 24361 25823 24395
rect 49433 24361 49467 24395
rect 27169 24293 27203 24327
rect 36645 24293 36679 24327
rect 37013 24293 37047 24327
rect 3249 24225 3283 24259
rect 5825 24225 5859 24259
rect 8217 24225 8251 24259
rect 13553 24225 13587 24259
rect 16129 24225 16163 24259
rect 20913 24225 20947 24259
rect 22477 24225 22511 24259
rect 25237 24225 25271 24259
rect 26341 24225 26375 24259
rect 27721 24225 27755 24259
rect 29009 24225 29043 24259
rect 29745 24225 29779 24259
rect 42625 24225 42659 24259
rect 45845 24225 45879 24259
rect 2237 24157 2271 24191
rect 4169 24157 4203 24191
rect 4813 24157 4847 24191
rect 6561 24157 6595 24191
rect 7297 24157 7331 24191
rect 9045 24157 9079 24191
rect 9321 24157 9355 24191
rect 9781 24157 9815 24191
rect 11621 24157 11655 24191
rect 11897 24157 11931 24191
rect 12541 24157 12575 24191
rect 14473 24157 14507 24191
rect 14933 24157 14967 24191
rect 16865 24157 16899 24191
rect 19625 24157 19659 24191
rect 20085 24157 20119 24191
rect 22201 24157 22235 24191
rect 25053 24157 25087 24191
rect 27629 24157 27663 24191
rect 28365 24157 28399 24191
rect 30021 24157 30055 24191
rect 31033 24157 31067 24191
rect 32321 24157 32355 24191
rect 32965 24157 32999 24191
rect 33425 24157 33459 24191
rect 34345 24157 34379 24191
rect 34897 24157 34931 24191
rect 36001 24157 36035 24191
rect 37473 24157 37507 24191
rect 38577 24157 38611 24191
rect 40049 24157 40083 24191
rect 41245 24157 41279 24191
rect 41521 24157 41555 24191
rect 42901 24157 42935 24191
rect 43913 24157 43947 24191
rect 45201 24157 45235 24191
rect 46581 24157 46615 24191
rect 47777 24157 47811 24191
rect 48881 24157 48915 24191
rect 1593 24089 1627 24123
rect 10977 24089 11011 24123
rect 17141 24089 17175 24123
rect 23857 24089 23891 24123
rect 24961 24089 24995 24123
rect 34069 24089 34103 24123
rect 35541 24089 35575 24123
rect 38117 24089 38151 24123
rect 46121 24089 46155 24123
rect 1777 24021 1811 24055
rect 3985 24021 4019 24055
rect 9137 24021 9171 24055
rect 11713 24021 11747 24055
rect 14289 24021 14323 24055
rect 18613 24021 18647 24055
rect 19073 24021 19107 24055
rect 19441 24021 19475 24055
rect 24593 24021 24627 24055
rect 26157 24021 26191 24055
rect 26249 24021 26283 24055
rect 27537 24021 27571 24055
rect 29285 24021 29319 24055
rect 31677 24021 31711 24055
rect 39221 24021 39255 24055
rect 39497 24021 39531 24055
rect 40693 24021 40727 24055
rect 44557 24021 44591 24055
rect 47225 24021 47259 24055
rect 48421 24021 48455 24055
rect 49065 24021 49099 24055
rect 21557 23817 21591 23851
rect 23765 23817 23799 23851
rect 32965 23817 32999 23851
rect 34437 23817 34471 23851
rect 40325 23817 40359 23851
rect 47041 23817 47075 23851
rect 48421 23817 48455 23851
rect 10977 23749 11011 23783
rect 12265 23749 12299 23783
rect 12357 23749 12391 23783
rect 14289 23749 14323 23783
rect 18153 23749 18187 23783
rect 21373 23749 21407 23783
rect 24225 23749 24259 23783
rect 25145 23749 25179 23783
rect 34069 23749 34103 23783
rect 42717 23749 42751 23783
rect 42901 23749 42935 23783
rect 47225 23749 47259 23783
rect 49433 23749 49467 23783
rect 1961 23681 1995 23715
rect 2973 23681 3007 23715
rect 3985 23681 4019 23715
rect 4629 23681 4663 23715
rect 6561 23681 6595 23715
rect 6837 23681 6871 23715
rect 8033 23681 8067 23715
rect 9873 23681 9907 23715
rect 11713 23681 11747 23715
rect 13277 23681 13311 23715
rect 14933 23681 14967 23715
rect 17141 23681 17175 23715
rect 21005 23681 21039 23715
rect 29377 23681 29411 23715
rect 30849 23681 30883 23715
rect 32321 23681 32355 23715
rect 33425 23681 33459 23715
rect 34897 23681 34931 23715
rect 36001 23681 36035 23715
rect 37473 23681 37507 23715
rect 38577 23681 38611 23715
rect 39681 23681 39715 23715
rect 40785 23681 40819 23715
rect 42073 23681 42107 23715
rect 43177 23681 43211 23715
rect 43545 23681 43579 23715
rect 44833 23681 44867 23715
rect 46213 23681 46247 23715
rect 47777 23681 47811 23715
rect 48881 23681 48915 23715
rect 2053 23613 2087 23647
rect 2237 23613 2271 23647
rect 5457 23613 5491 23647
rect 9137 23613 9171 23647
rect 12541 23613 12575 23647
rect 16129 23613 16163 23647
rect 18797 23613 18831 23647
rect 19073 23613 19107 23647
rect 22017 23613 22051 23647
rect 22293 23613 22327 23647
rect 24869 23613 24903 23647
rect 27169 23613 27203 23647
rect 27445 23613 27479 23647
rect 29653 23613 29687 23647
rect 31585 23613 31619 23647
rect 35541 23613 35575 23647
rect 43821 23613 43855 23647
rect 45937 23613 45971 23647
rect 11621 23545 11655 23579
rect 21189 23545 21223 23579
rect 26617 23545 26651 23579
rect 28917 23545 28951 23579
rect 34529 23545 34563 23579
rect 38117 23545 38151 23579
rect 41429 23545 41463 23579
rect 41889 23545 41923 23579
rect 1593 23477 1627 23511
rect 11897 23477 11931 23511
rect 20545 23477 20579 23511
rect 30481 23477 30515 23511
rect 36645 23477 36679 23511
rect 37105 23477 37139 23511
rect 39221 23477 39255 23511
rect 45477 23477 45511 23511
rect 49065 23477 49099 23511
rect 18889 23273 18923 23307
rect 32965 23273 32999 23307
rect 36645 23273 36679 23307
rect 40693 23273 40727 23307
rect 41797 23273 41831 23307
rect 44005 23273 44039 23307
rect 44465 23273 44499 23307
rect 49341 23273 49375 23307
rect 3617 23205 3651 23239
rect 13921 23205 13955 23239
rect 29101 23205 29135 23239
rect 31953 23205 31987 23239
rect 34069 23205 34103 23239
rect 42901 23205 42935 23239
rect 46121 23205 46155 23239
rect 3433 23137 3467 23171
rect 4261 23137 4295 23171
rect 6101 23137 6135 23171
rect 7849 23137 7883 23171
rect 10517 23137 10551 23171
rect 17141 23137 17175 23171
rect 17417 23137 17451 23171
rect 20085 23137 20119 23171
rect 22293 23137 22327 23171
rect 22569 23137 22603 23171
rect 25237 23137 25271 23171
rect 26341 23137 26375 23171
rect 27353 23137 27387 23171
rect 27629 23137 27663 23171
rect 30021 23137 30055 23171
rect 37749 23137 37783 23171
rect 48237 23137 48271 23171
rect 1777 23069 1811 23103
rect 3985 23069 4019 23103
rect 5457 23069 5491 23103
rect 7389 23069 7423 23103
rect 9505 23069 9539 23103
rect 11161 23069 11195 23103
rect 14657 23069 14691 23103
rect 15485 23069 15519 23103
rect 16405 23069 16439 23103
rect 26249 23069 26283 23103
rect 29745 23069 29779 23103
rect 32321 23069 32355 23103
rect 33425 23069 33459 23103
rect 34897 23069 34931 23103
rect 36001 23069 36035 23103
rect 37289 23069 37323 23103
rect 40049 23069 40083 23103
rect 41153 23069 41187 23103
rect 42257 23069 42291 23103
rect 43361 23069 43395 23103
rect 44649 23069 44683 23103
rect 45201 23069 45235 23103
rect 46489 23069 46523 23103
rect 47593 23069 47627 23103
rect 48697 23069 48731 23103
rect 2789 23001 2823 23035
rect 11437 23001 11471 23035
rect 13185 23001 13219 23035
rect 13553 23001 13587 23035
rect 20361 23001 20395 23035
rect 24961 23001 24995 23035
rect 35541 23001 35575 23035
rect 38025 23001 38059 23035
rect 9045 22933 9079 22967
rect 13737 22933 13771 22967
rect 14289 22933 14323 22967
rect 14749 22933 14783 22967
rect 19441 22933 19475 22967
rect 21833 22933 21867 22967
rect 24041 22933 24075 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 25789 22933 25823 22967
rect 26157 22933 26191 22967
rect 26893 22933 26927 22967
rect 26985 22933 27019 22967
rect 31493 22933 31527 22967
rect 31861 22933 31895 22967
rect 34345 22933 34379 22967
rect 37105 22933 37139 22967
rect 39497 22933 39531 22967
rect 45845 22933 45879 22967
rect 47133 22933 47167 22967
rect 3893 22729 3927 22763
rect 4353 22729 4387 22763
rect 25329 22729 25363 22763
rect 31953 22729 31987 22763
rect 34345 22729 34379 22763
rect 35541 22729 35575 22763
rect 36645 22729 36679 22763
rect 36921 22729 36955 22763
rect 38117 22729 38151 22763
rect 41429 22729 41463 22763
rect 47225 22729 47259 22763
rect 6653 22661 6687 22695
rect 8585 22661 8619 22695
rect 9505 22661 9539 22695
rect 11989 22661 12023 22695
rect 12541 22661 12575 22695
rect 14473 22661 14507 22695
rect 16129 22661 16163 22695
rect 17141 22661 17175 22695
rect 19993 22661 20027 22695
rect 28733 22661 28767 22695
rect 31125 22661 31159 22695
rect 47041 22661 47075 22695
rect 47869 22661 47903 22695
rect 1777 22593 1811 22627
rect 3341 22593 3375 22627
rect 3801 22593 3835 22627
rect 4629 22593 4663 22627
rect 7573 22593 7607 22627
rect 12265 22593 12299 22627
rect 14933 22593 14967 22627
rect 22017 22593 22051 22627
rect 23121 22593 23155 22627
rect 25697 22593 25731 22627
rect 27629 22593 27663 22627
rect 28457 22593 28491 22627
rect 31033 22593 31067 22627
rect 32321 22593 32355 22627
rect 33425 22593 33459 22627
rect 34069 22593 34103 22627
rect 34897 22593 34931 22627
rect 36001 22593 36035 22627
rect 37473 22593 37507 22627
rect 38577 22593 38611 22627
rect 39221 22593 39255 22627
rect 39681 22593 39715 22627
rect 40785 22593 40819 22627
rect 42901 22593 42935 22627
rect 43913 22593 43947 22627
rect 45017 22593 45051 22627
rect 45753 22593 45787 22627
rect 46489 22593 46523 22627
rect 48697 22593 48731 22627
rect 2237 22525 2271 22559
rect 4077 22525 4111 22559
rect 5089 22525 5123 22559
rect 6837 22525 6871 22559
rect 9229 22525 9263 22559
rect 16865 22525 16899 22559
rect 19073 22525 19107 22559
rect 19717 22525 19751 22559
rect 21465 22525 21499 22559
rect 23397 22525 23431 22559
rect 25789 22525 25823 22559
rect 25973 22525 26007 22559
rect 26341 22525 26375 22559
rect 27721 22525 27755 22559
rect 27905 22525 27939 22559
rect 31309 22525 31343 22559
rect 41889 22525 41923 22559
rect 42625 22525 42659 22559
rect 48421 22525 48455 22559
rect 11621 22457 11655 22491
rect 24869 22457 24903 22491
rect 27261 22457 27295 22491
rect 32965 22457 32999 22491
rect 34621 22457 34655 22491
rect 45937 22457 45971 22491
rect 3433 22389 3467 22423
rect 10977 22389 11011 22423
rect 11345 22389 11379 22423
rect 11713 22389 11747 22423
rect 14013 22389 14047 22423
rect 14657 22389 14691 22423
rect 18613 22389 18647 22423
rect 22661 22389 22695 22423
rect 26617 22389 26651 22423
rect 26801 22389 26835 22423
rect 30205 22389 30239 22423
rect 30665 22389 30699 22423
rect 31769 22389 31803 22423
rect 40325 22389 40359 22423
rect 44557 22389 44591 22423
rect 45201 22389 45235 22423
rect 46673 22389 46707 22423
rect 47961 22389 47995 22423
rect 49341 22389 49375 22423
rect 17404 22185 17438 22219
rect 26046 22185 26080 22219
rect 29101 22185 29135 22219
rect 29285 22185 29319 22219
rect 29745 22185 29779 22219
rect 46673 22185 46707 22219
rect 23305 22117 23339 22151
rect 46857 22117 46891 22151
rect 2053 22049 2087 22083
rect 4445 22049 4479 22083
rect 7297 22049 7331 22083
rect 9781 22049 9815 22083
rect 9965 22049 9999 22083
rect 11253 22049 11287 22083
rect 13461 22049 13495 22083
rect 15669 22049 15703 22083
rect 17141 22049 17175 22083
rect 20821 22049 20855 22083
rect 22845 22049 22879 22083
rect 23949 22049 23983 22083
rect 25145 22049 25179 22083
rect 27537 22049 27571 22083
rect 30389 22049 30423 22083
rect 31861 22049 31895 22083
rect 34069 22049 34103 22083
rect 37013 22049 37047 22083
rect 39221 22049 39255 22083
rect 40325 22049 40359 22083
rect 41613 22049 41647 22083
rect 49341 22049 49375 22083
rect 1593 21981 1627 22015
rect 3985 21981 4019 22015
rect 6101 21981 6135 22015
rect 6929 21981 6963 22015
rect 8585 21981 8619 22015
rect 10701 21981 10735 22015
rect 12541 21981 12575 22015
rect 14565 21981 14599 22015
rect 14749 21981 14783 22015
rect 15209 21981 15243 22015
rect 19472 21981 19506 22015
rect 20361 21981 20395 22015
rect 22201 21981 22235 22015
rect 23765 21981 23799 22015
rect 25789 21981 25823 22015
rect 27997 21981 28031 22015
rect 30113 21981 30147 22015
rect 30941 21981 30975 22015
rect 31585 21981 31619 22015
rect 32321 21981 32355 22015
rect 33425 21981 33459 22015
rect 34897 21981 34931 22015
rect 36001 21981 36035 22015
rect 37473 21981 37507 22015
rect 38577 21981 38611 22015
rect 40049 21981 40083 22015
rect 41337 21981 41371 22015
rect 42625 21981 42659 22015
rect 43729 21981 43763 22015
rect 44373 21981 44407 22015
rect 45201 21981 45235 22015
rect 45937 21981 45971 22015
rect 46489 21981 46523 22015
rect 47225 21981 47259 22015
rect 47961 21981 47995 22015
rect 48697 21981 48731 22015
rect 3433 21913 3467 21947
rect 9045 21913 9079 21947
rect 19717 21913 19751 21947
rect 24961 21913 24995 21947
rect 32965 21913 32999 21947
rect 37105 21913 37139 21947
rect 3525 21845 3559 21879
rect 5825 21845 5859 21879
rect 6285 21845 6319 21879
rect 8769 21845 8803 21879
rect 9321 21845 9355 21879
rect 9689 21845 9723 21879
rect 14197 21845 14231 21879
rect 18889 21845 18923 21879
rect 23673 21845 23707 21879
rect 24593 21845 24627 21879
rect 25053 21845 25087 21879
rect 28641 21845 28675 21879
rect 28917 21845 28951 21879
rect 30205 21845 30239 21879
rect 34345 21845 34379 21879
rect 35541 21845 35575 21879
rect 36645 21845 36679 21879
rect 38117 21845 38151 21879
rect 39497 21845 39531 21879
rect 43269 21845 43303 21879
rect 44649 21845 44683 21879
rect 45385 21845 45419 21879
rect 46121 21845 46155 21879
rect 47409 21845 47443 21879
rect 48145 21845 48179 21879
rect 5181 21641 5215 21675
rect 5733 21641 5767 21675
rect 6469 21641 6503 21675
rect 6929 21641 6963 21675
rect 11713 21641 11747 21675
rect 12173 21641 12207 21675
rect 15301 21641 15335 21675
rect 26617 21641 26651 21675
rect 27629 21641 27663 21675
rect 27721 21641 27755 21675
rect 32965 21641 32999 21675
rect 34345 21641 34379 21675
rect 36645 21641 36679 21675
rect 44097 21641 44131 21675
rect 45201 21641 45235 21675
rect 45569 21641 45603 21675
rect 45753 21641 45787 21675
rect 47041 21641 47075 21675
rect 47685 21641 47719 21675
rect 7021 21573 7055 21607
rect 9965 21573 9999 21607
rect 15117 21573 15151 21607
rect 18981 21573 19015 21607
rect 21097 21573 21131 21607
rect 23673 21573 23707 21607
rect 25973 21573 26007 21607
rect 26157 21573 26191 21607
rect 26249 21573 26283 21607
rect 28733 21573 28767 21607
rect 31769 21573 31803 21607
rect 1685 21505 1719 21539
rect 3617 21505 3651 21539
rect 5641 21505 5675 21539
rect 10241 21505 10275 21539
rect 12081 21505 12115 21539
rect 15945 21505 15979 21539
rect 17049 21505 17083 21539
rect 22017 21505 22051 21539
rect 28457 21505 28491 21539
rect 31033 21505 31067 21539
rect 31125 21505 31159 21539
rect 32321 21505 32355 21539
rect 33425 21505 33459 21539
rect 34897 21505 34931 21539
rect 36001 21505 36035 21539
rect 37749 21505 37783 21539
rect 38761 21505 38795 21539
rect 39865 21505 39899 21539
rect 40969 21505 41003 21539
rect 42717 21505 42751 21539
rect 43453 21505 43487 21539
rect 44281 21505 44315 21539
rect 44925 21505 44959 21539
rect 45385 21505 45419 21539
rect 47225 21505 47259 21539
rect 47961 21505 47995 21539
rect 2789 21437 2823 21471
rect 4169 21437 4203 21471
rect 5917 21437 5951 21471
rect 7205 21437 7239 21471
rect 7757 21437 7791 21471
rect 8033 21437 8067 21471
rect 10977 21437 11011 21471
rect 12265 21437 12299 21471
rect 12909 21437 12943 21471
rect 13185 21437 13219 21471
rect 16037 21437 16071 21471
rect 16221 21437 16255 21471
rect 17325 21437 17359 21471
rect 18705 21437 18739 21471
rect 22753 21437 22787 21471
rect 23397 21437 23431 21471
rect 27813 21437 27847 21471
rect 30205 21437 30239 21471
rect 31217 21437 31251 21471
rect 37473 21437 37507 21471
rect 41613 21437 41647 21471
rect 49157 21437 49191 21471
rect 9505 21369 9539 21403
rect 20453 21369 20487 21403
rect 25145 21369 25179 21403
rect 42073 21369 42107 21403
rect 5273 21301 5307 21335
rect 6561 21301 6595 21335
rect 14657 21301 14691 21335
rect 15577 21301 15611 21335
rect 21373 21301 21407 21335
rect 25697 21301 25731 21335
rect 27261 21301 27295 21335
rect 30665 21301 30699 21335
rect 31861 21301 31895 21335
rect 34069 21301 34103 21335
rect 34621 21301 34655 21335
rect 35541 21301 35575 21335
rect 37013 21301 37047 21335
rect 39405 21301 39439 21335
rect 40509 21301 40543 21335
rect 41889 21301 41923 21335
rect 42809 21301 42843 21335
rect 43545 21301 43579 21335
rect 44741 21301 44775 21335
rect 10977 21097 11011 21131
rect 14565 21097 14599 21131
rect 15761 21097 15795 21131
rect 27721 21097 27755 21131
rect 29101 21097 29135 21131
rect 35081 21097 35115 21131
rect 38853 21097 38887 21131
rect 40693 21097 40727 21131
rect 41337 21097 41371 21131
rect 44649 21097 44683 21131
rect 48421 21097 48455 21131
rect 49341 21097 49375 21131
rect 3525 21029 3559 21063
rect 14289 21029 14323 21063
rect 21465 21029 21499 21063
rect 28825 21029 28859 21063
rect 31217 21029 31251 21063
rect 44005 21029 44039 21063
rect 2053 20961 2087 20995
rect 4445 20961 4479 20995
rect 8401 20961 8435 20995
rect 10057 20961 10091 20995
rect 11529 20961 11563 20995
rect 12817 20961 12851 20995
rect 15117 20961 15151 20995
rect 16221 20961 16255 20995
rect 16313 20961 16347 20995
rect 17509 20961 17543 20995
rect 18613 20961 18647 20995
rect 18797 20961 18831 20995
rect 22293 20961 22327 20995
rect 22477 20961 22511 20995
rect 23673 20961 23707 20995
rect 25237 20961 25271 20995
rect 31861 20961 31895 20995
rect 35817 20961 35851 20995
rect 36093 20961 36127 20995
rect 1777 20893 1811 20927
rect 4077 20893 4111 20927
rect 6193 20893 6227 20927
rect 9321 20893 9355 20927
rect 11989 20893 12023 20927
rect 13829 20893 13863 20927
rect 17325 20893 17359 20927
rect 18521 20893 18555 20927
rect 19441 20893 19475 20927
rect 22201 20893 22235 20927
rect 23489 20893 23523 20927
rect 24225 20893 24259 20927
rect 25973 20893 26007 20927
rect 28181 20893 28215 20927
rect 31585 20893 31619 20927
rect 31677 20893 31711 20927
rect 32413 20893 32447 20927
rect 33517 20893 33551 20927
rect 34529 20893 34563 20927
rect 37105 20893 37139 20927
rect 38209 20893 38243 20927
rect 39497 20893 39531 20927
rect 40049 20893 40083 20927
rect 41981 20893 42015 20927
rect 43545 20893 43579 20927
rect 44189 20893 44223 20927
rect 44465 20893 44499 20927
rect 48697 20893 48731 20927
rect 6469 20825 6503 20859
rect 11161 20825 11195 20859
rect 13737 20825 13771 20859
rect 15025 20825 15059 20859
rect 19717 20825 19751 20859
rect 25053 20825 25087 20859
rect 26249 20825 26283 20859
rect 29837 20825 29871 20859
rect 30665 20825 30699 20859
rect 33057 20825 33091 20859
rect 34989 20825 35023 20859
rect 35541 20825 35575 20859
rect 41245 20825 41279 20859
rect 42717 20825 42751 20859
rect 42901 20825 42935 20859
rect 3433 20757 3467 20791
rect 5733 20757 5767 20791
rect 5917 20757 5951 20791
rect 7941 20757 7975 20791
rect 11345 20757 11379 20791
rect 11713 20757 11747 20791
rect 14933 20757 14967 20791
rect 16129 20757 16163 20791
rect 16957 20757 16991 20791
rect 17417 20757 17451 20791
rect 18153 20757 18187 20791
rect 21189 20757 21223 20791
rect 21741 20757 21775 20791
rect 21833 20757 21867 20791
rect 23029 20757 23063 20791
rect 23397 20757 23431 20791
rect 24685 20757 24719 20791
rect 25145 20757 25179 20791
rect 29285 20757 29319 20791
rect 34161 20757 34195 20791
rect 37749 20757 37783 20791
rect 39313 20757 39347 20791
rect 42073 20757 42107 20791
rect 43361 20757 43395 20791
rect 47777 20757 47811 20791
rect 11713 20553 11747 20587
rect 12357 20553 12391 20587
rect 16865 20553 16899 20587
rect 17601 20553 17635 20587
rect 18245 20553 18279 20587
rect 23581 20553 23615 20587
rect 24133 20553 24167 20587
rect 26157 20553 26191 20587
rect 26801 20553 26835 20587
rect 34621 20553 34655 20587
rect 35541 20553 35575 20587
rect 43453 20553 43487 20587
rect 49433 20553 49467 20587
rect 3709 20485 3743 20519
rect 8493 20485 8527 20519
rect 8953 20485 8987 20519
rect 12725 20485 12759 20519
rect 13829 20485 13863 20519
rect 16037 20485 16071 20519
rect 18889 20485 18923 20519
rect 31769 20485 31803 20519
rect 36645 20485 36679 20519
rect 49249 20485 49283 20519
rect 1593 20417 1627 20451
rect 3525 20417 3559 20451
rect 6745 20417 6779 20451
rect 10977 20417 11011 20451
rect 11897 20417 11931 20451
rect 16221 20417 16255 20451
rect 17509 20417 17543 20451
rect 18981 20417 19015 20451
rect 19717 20417 19751 20451
rect 22017 20417 22051 20451
rect 23489 20417 23523 20451
rect 26525 20417 26559 20451
rect 27537 20417 27571 20451
rect 28457 20417 28491 20451
rect 31033 20417 31067 20451
rect 32321 20417 32355 20451
rect 33425 20417 33459 20451
rect 34897 20417 34931 20451
rect 36001 20417 36035 20451
rect 37749 20417 37783 20451
rect 38761 20417 38795 20451
rect 39037 20417 39071 20451
rect 40049 20417 40083 20451
rect 40325 20417 40359 20451
rect 41245 20417 41279 20451
rect 42809 20417 42843 20451
rect 43085 20417 43119 20451
rect 2053 20349 2087 20383
rect 4261 20349 4295 20383
rect 4537 20349 4571 20383
rect 6009 20349 6043 20383
rect 7021 20349 7055 20383
rect 8677 20349 8711 20383
rect 12817 20349 12851 20383
rect 13001 20349 13035 20383
rect 13553 20349 13587 20383
rect 15301 20349 15335 20383
rect 17693 20349 17727 20383
rect 19073 20349 19107 20383
rect 19993 20349 20027 20383
rect 21465 20349 21499 20383
rect 22845 20349 22879 20383
rect 24409 20349 24443 20383
rect 24685 20349 24719 20383
rect 27629 20349 27663 20383
rect 27813 20349 27847 20383
rect 28733 20349 28767 20383
rect 31125 20349 31159 20383
rect 31309 20349 31343 20383
rect 34069 20349 34103 20383
rect 34345 20349 34379 20383
rect 37473 20349 37507 20383
rect 41521 20349 41555 20383
rect 11161 20281 11195 20315
rect 30665 20281 30699 20315
rect 43269 20281 43303 20315
rect 8401 20213 8435 20247
rect 10425 20213 10459 20247
rect 15669 20213 15703 20247
rect 17141 20213 17175 20247
rect 18521 20213 18555 20247
rect 27169 20213 27203 20247
rect 30205 20213 30239 20247
rect 31953 20213 31987 20247
rect 32965 20213 32999 20247
rect 37013 20213 37047 20247
rect 40785 20213 40819 20247
rect 42625 20213 42659 20247
rect 43637 20213 43671 20247
rect 3617 20009 3651 20043
rect 3893 20009 3927 20043
rect 9045 20009 9079 20043
rect 12449 20009 12483 20043
rect 19717 20009 19751 20043
rect 23949 20009 23983 20043
rect 27629 20009 27663 20043
rect 29009 20009 29043 20043
rect 35541 20009 35575 20043
rect 38853 20009 38887 20043
rect 41981 20009 42015 20043
rect 42349 20009 42383 20043
rect 12725 19941 12759 19975
rect 22293 19941 22327 19975
rect 22569 19941 22603 19975
rect 31585 19941 31619 19975
rect 40325 19941 40359 19975
rect 2053 19873 2087 19907
rect 3985 19873 4019 19907
rect 6837 19873 6871 19907
rect 13185 19873 13219 19907
rect 13277 19873 13311 19907
rect 17509 19873 17543 19907
rect 18797 19873 18831 19907
rect 23305 19873 23339 19907
rect 23489 19873 23523 19907
rect 25237 19873 25271 19907
rect 26157 19873 26191 19907
rect 29377 19873 29411 19907
rect 30297 19873 30331 19907
rect 31861 19873 31895 19907
rect 1593 19805 1627 19839
rect 4629 19805 4663 19839
rect 9413 19805 9447 19839
rect 10057 19805 10091 19839
rect 13829 19805 13863 19839
rect 14381 19805 14415 19839
rect 16681 19805 16715 19839
rect 17325 19805 17359 19839
rect 17417 19805 17451 19839
rect 19625 19805 19659 19839
rect 20269 19805 20303 19839
rect 23213 19805 23247 19839
rect 25145 19805 25179 19839
rect 25881 19805 25915 19839
rect 28089 19805 28123 19839
rect 30941 19805 30975 19839
rect 32321 19805 32355 19839
rect 32965 19805 32999 19839
rect 33425 19805 33459 19839
rect 34897 19805 34931 19839
rect 36001 19805 36035 19839
rect 37105 19805 37139 19839
rect 38209 19805 38243 19839
rect 39497 19805 39531 19839
rect 40877 19805 40911 19839
rect 41705 19805 41739 19839
rect 42165 19805 42199 19839
rect 4905 19737 4939 19771
rect 7113 19737 7147 19771
rect 10333 19737 10367 19771
rect 13093 19737 13127 19771
rect 14657 19737 14691 19771
rect 20545 19737 20579 19771
rect 28733 19737 28767 19771
rect 40141 19737 40175 19771
rect 3433 19669 3467 19703
rect 6377 19669 6411 19703
rect 8585 19669 8619 19703
rect 9505 19669 9539 19703
rect 11805 19669 11839 19703
rect 12265 19669 12299 19703
rect 16129 19669 16163 19703
rect 16957 19669 16991 19703
rect 18153 19669 18187 19703
rect 18521 19669 18555 19703
rect 18613 19669 18647 19703
rect 22017 19669 22051 19703
rect 22845 19669 22879 19703
rect 24225 19669 24259 19703
rect 24685 19669 24719 19703
rect 25053 19669 25087 19703
rect 29745 19669 29779 19703
rect 30113 19669 30147 19703
rect 30205 19669 30239 19703
rect 34069 19669 34103 19703
rect 34529 19669 34563 19703
rect 36645 19669 36679 19703
rect 37749 19669 37783 19703
rect 39313 19669 39347 19703
rect 40969 19669 41003 19703
rect 41521 19669 41555 19703
rect 42533 19669 42567 19703
rect 5273 19465 5307 19499
rect 5733 19465 5767 19499
rect 9229 19465 9263 19499
rect 9597 19465 9631 19499
rect 10425 19465 10459 19499
rect 10793 19465 10827 19499
rect 17601 19465 17635 19499
rect 19257 19465 19291 19499
rect 21465 19465 21499 19499
rect 22017 19465 22051 19499
rect 22477 19465 22511 19499
rect 23765 19465 23799 19499
rect 27169 19465 27203 19499
rect 27537 19465 27571 19499
rect 30113 19465 30147 19499
rect 31217 19465 31251 19499
rect 36645 19465 36679 19499
rect 41337 19465 41371 19499
rect 4353 19397 4387 19431
rect 6837 19397 6871 19431
rect 13553 19397 13587 19431
rect 14749 19397 14783 19431
rect 24961 19397 24995 19431
rect 26433 19397 26467 19431
rect 28641 19397 28675 19431
rect 38853 19397 38887 19431
rect 40141 19397 40175 19431
rect 40693 19397 40727 19431
rect 41153 19397 41187 19431
rect 1777 19329 1811 19363
rect 3617 19329 3651 19363
rect 5641 19329 5675 19363
rect 6561 19329 6595 19363
rect 8769 19329 8803 19363
rect 10885 19329 10919 19363
rect 11713 19329 11747 19363
rect 12357 19329 12391 19363
rect 12817 19329 12851 19363
rect 14657 19329 14691 19363
rect 15853 19329 15887 19363
rect 16957 19329 16991 19363
rect 18429 19329 18463 19363
rect 19717 19329 19751 19363
rect 22385 19329 22419 19363
rect 24133 19329 24167 19363
rect 24225 19329 24259 19363
rect 30573 19329 30607 19363
rect 31585 19329 31619 19363
rect 32321 19329 32355 19363
rect 33425 19329 33459 19363
rect 34069 19329 34103 19363
rect 34897 19329 34931 19363
rect 35541 19329 35575 19363
rect 36001 19329 36035 19363
rect 37749 19329 37783 19363
rect 39681 19329 39715 19363
rect 2053 19261 2087 19295
rect 5825 19261 5859 19295
rect 9689 19261 9723 19295
rect 9873 19261 9907 19295
rect 10977 19261 11011 19295
rect 14841 19261 14875 19295
rect 15945 19261 15979 19295
rect 16037 19261 16071 19295
rect 18521 19261 18555 19295
rect 18613 19261 18647 19295
rect 19993 19261 20027 19295
rect 22661 19261 22695 19295
rect 23305 19261 23339 19295
rect 24409 19261 24443 19295
rect 25789 19261 25823 19295
rect 27629 19261 27663 19295
rect 27721 19261 27755 19295
rect 28365 19261 28399 19295
rect 37473 19261 37507 19295
rect 39037 19261 39071 19295
rect 41613 19261 41647 19295
rect 14289 19193 14323 19227
rect 31861 19193 31895 19227
rect 34529 19193 34563 19227
rect 40049 19193 40083 19227
rect 5089 19125 5123 19159
rect 8309 19125 8343 19159
rect 8953 19125 8987 19159
rect 15485 19125 15519 19159
rect 18061 19125 18095 19159
rect 19441 19125 19475 19159
rect 23029 19125 23063 19159
rect 23489 19125 23523 19159
rect 26525 19125 26559 19159
rect 31769 19125 31803 19159
rect 32965 19125 32999 19159
rect 34345 19125 34379 19159
rect 37013 19125 37047 19159
rect 39497 19125 39531 19159
rect 40785 19125 40819 19159
rect 10425 18921 10459 18955
rect 12633 18921 12667 18955
rect 13737 18921 13771 18955
rect 17601 18921 17635 18955
rect 23305 18921 23339 18955
rect 25776 18921 25810 18955
rect 28457 18921 28491 18955
rect 32045 18921 32079 18955
rect 33425 18921 33459 18955
rect 36829 18921 36863 18955
rect 24869 18853 24903 18887
rect 39313 18853 39347 18887
rect 40049 18853 40083 18887
rect 40233 18853 40267 18887
rect 2053 18785 2087 18819
rect 3433 18785 3467 18819
rect 4445 18785 4479 18819
rect 6285 18785 6319 18819
rect 8217 18785 8251 18819
rect 9597 18785 9631 18819
rect 9689 18785 9723 18819
rect 10885 18785 10919 18819
rect 14473 18785 14507 18819
rect 14749 18785 14783 18819
rect 16865 18785 16899 18819
rect 18061 18785 18095 18819
rect 18153 18785 18187 18819
rect 18613 18785 18647 18819
rect 20361 18785 20395 18819
rect 21097 18785 21131 18819
rect 23121 18785 23155 18819
rect 23949 18785 23983 18819
rect 25513 18785 25547 18819
rect 27721 18785 27755 18819
rect 29101 18785 29135 18819
rect 1777 18717 1811 18751
rect 4169 18717 4203 18751
rect 6009 18717 6043 18751
rect 13093 18717 13127 18751
rect 16957 18717 16991 18751
rect 19625 18717 19659 18751
rect 23673 18717 23707 18751
rect 28917 18717 28951 18751
rect 29745 18717 29779 18751
rect 30849 18717 30883 18751
rect 32321 18717 32355 18751
rect 33609 18717 33643 18751
rect 34897 18717 34931 18751
rect 35173 18717 35207 18751
rect 36185 18717 36219 18751
rect 37105 18717 37139 18751
rect 37473 18717 37507 18751
rect 39497 18717 39531 18751
rect 8033 18649 8067 18683
rect 9505 18649 9539 18683
rect 10609 18649 10643 18683
rect 11161 18649 11195 18683
rect 15025 18649 15059 18683
rect 17969 18649 18003 18683
rect 21373 18649 21407 18683
rect 24685 18649 24719 18683
rect 31493 18649 31527 18683
rect 31769 18649 31803 18683
rect 34161 18649 34195 18683
rect 38669 18649 38703 18683
rect 39865 18649 39899 18683
rect 3617 18581 3651 18615
rect 7665 18581 7699 18615
rect 8125 18581 8159 18615
rect 8769 18581 8803 18615
rect 9137 18581 9171 18615
rect 10241 18581 10275 18615
rect 14289 18581 14323 18615
rect 16497 18581 16531 18615
rect 18797 18581 18831 18615
rect 19073 18581 19107 18615
rect 19349 18581 19383 18615
rect 22845 18581 22879 18615
rect 23765 18581 23799 18615
rect 25237 18581 25271 18615
rect 27261 18581 27295 18615
rect 28825 18581 28859 18615
rect 30389 18581 30423 18615
rect 32965 18581 32999 18615
rect 34253 18581 34287 18615
rect 34805 18581 34839 18615
rect 38117 18581 38151 18615
rect 38761 18581 38795 18615
rect 10333 18377 10367 18411
rect 12265 18377 12299 18411
rect 12633 18377 12667 18411
rect 14841 18377 14875 18411
rect 15301 18377 15335 18411
rect 19165 18377 19199 18411
rect 21465 18377 21499 18411
rect 24869 18377 24903 18411
rect 32137 18377 32171 18411
rect 32781 18377 32815 18411
rect 39405 18377 39439 18411
rect 5641 18309 5675 18343
rect 7481 18309 7515 18343
rect 9689 18309 9723 18343
rect 11713 18309 11747 18343
rect 11989 18309 12023 18343
rect 13461 18309 13495 18343
rect 14289 18309 14323 18343
rect 17233 18309 17267 18343
rect 22661 18309 22695 18343
rect 23397 18309 23431 18343
rect 26065 18309 26099 18343
rect 30941 18309 30975 18343
rect 31769 18309 31803 18343
rect 1777 18241 1811 18275
rect 3617 18241 3651 18275
rect 6745 18241 6779 18275
rect 8953 18241 8987 18275
rect 10701 18241 10735 18275
rect 12725 18241 12759 18275
rect 15209 18241 15243 18275
rect 16129 18241 16163 18275
rect 17325 18241 17359 18275
rect 18061 18241 18095 18275
rect 19533 18241 19567 18275
rect 20821 18241 20855 18275
rect 22017 18241 22051 18275
rect 23121 18241 23155 18275
rect 25329 18241 25363 18275
rect 28089 18241 28123 18275
rect 30297 18241 30331 18275
rect 31585 18241 31619 18275
rect 33241 18241 33275 18275
rect 34805 18241 34839 18275
rect 35817 18241 35851 18275
rect 36737 18241 36771 18275
rect 37565 18241 37599 18275
rect 38209 18241 38243 18275
rect 39129 18241 39163 18275
rect 2053 18173 2087 18207
rect 3893 18173 3927 18207
rect 5733 18173 5767 18207
rect 5917 18173 5951 18207
rect 8401 18173 8435 18207
rect 10793 18173 10827 18207
rect 10977 18173 11011 18207
rect 12909 18173 12943 18207
rect 15393 18173 15427 18207
rect 17509 18173 17543 18207
rect 19625 18173 19659 18207
rect 19717 18173 19751 18207
rect 27169 18173 27203 18207
rect 28365 18173 28399 18207
rect 33517 18173 33551 18207
rect 34529 18173 34563 18207
rect 5273 18105 5307 18139
rect 16313 18105 16347 18139
rect 16865 18105 16899 18139
rect 32413 18105 32447 18139
rect 8217 18037 8251 18071
rect 8677 18037 8711 18071
rect 11529 18037 11563 18071
rect 18705 18037 18739 18071
rect 20177 18037 20211 18071
rect 20453 18037 20487 18071
rect 26617 18037 26651 18071
rect 26801 18037 26835 18071
rect 27721 18037 27755 18071
rect 29837 18037 29871 18071
rect 32505 18037 32539 18071
rect 36461 18037 36495 18071
rect 37013 18037 37047 18071
rect 37657 18037 37691 18071
rect 38393 18037 38427 18071
rect 38945 18037 38979 18071
rect 7297 17833 7331 17867
rect 11805 17833 11839 17867
rect 12909 17833 12943 17867
rect 14289 17833 14323 17867
rect 15393 17833 15427 17867
rect 25132 17833 25166 17867
rect 35541 17833 35575 17867
rect 4169 17765 4203 17799
rect 20269 17765 20303 17799
rect 26617 17765 26651 17799
rect 28825 17765 28859 17799
rect 36921 17765 36955 17799
rect 2053 17697 2087 17731
rect 3617 17697 3651 17731
rect 4813 17697 4847 17731
rect 8401 17697 8435 17731
rect 10977 17697 11011 17731
rect 11161 17697 11195 17731
rect 12357 17697 12391 17731
rect 13553 17697 13587 17731
rect 14473 17697 14507 17731
rect 15853 17697 15887 17731
rect 18889 17697 18923 17731
rect 20913 17697 20947 17731
rect 22385 17697 22419 17731
rect 24869 17697 24903 17731
rect 27077 17697 27111 17731
rect 29193 17697 29227 17731
rect 30297 17697 30331 17731
rect 33793 17697 33827 17731
rect 1777 17629 1811 17663
rect 3893 17629 3927 17663
rect 4353 17629 4387 17663
rect 9873 17629 9907 17663
rect 14749 17629 14783 17663
rect 18245 17629 18279 17663
rect 22109 17629 22143 17663
rect 24409 17629 24443 17663
rect 30941 17629 30975 17663
rect 32045 17629 32079 17663
rect 33149 17629 33183 17663
rect 34253 17629 34287 17663
rect 34897 17629 34931 17663
rect 36185 17629 36219 17663
rect 37565 17629 37599 17663
rect 37841 17629 37875 17663
rect 5089 17561 5123 17595
rect 7205 17561 7239 17595
rect 8217 17561 8251 17595
rect 9137 17561 9171 17595
rect 11621 17561 11655 17595
rect 12081 17561 12115 17595
rect 13369 17561 13403 17595
rect 16129 17561 16163 17595
rect 19533 17561 19567 17595
rect 27353 17561 27387 17595
rect 29285 17561 29319 17595
rect 36737 17561 36771 17595
rect 3341 17493 3375 17527
rect 6561 17493 6595 17527
rect 7849 17493 7883 17527
rect 8309 17493 8343 17527
rect 10517 17493 10551 17527
rect 10885 17493 10919 17527
rect 12265 17493 12299 17527
rect 12633 17493 12667 17527
rect 13277 17493 13311 17527
rect 17601 17493 17635 17527
rect 19625 17493 19659 17527
rect 20637 17493 20671 17527
rect 20729 17493 20763 17527
rect 21465 17493 21499 17527
rect 23857 17493 23891 17527
rect 24225 17493 24259 17527
rect 29745 17493 29779 17527
rect 30113 17493 30147 17527
rect 30205 17493 30239 17527
rect 31585 17493 31619 17527
rect 32689 17493 32723 17527
rect 34069 17493 34103 17527
rect 34529 17493 34563 17527
rect 36001 17493 36035 17527
rect 37381 17493 37415 17527
rect 5273 17289 5307 17323
rect 5733 17289 5767 17323
rect 8033 17289 8067 17323
rect 9965 17289 9999 17323
rect 10793 17289 10827 17323
rect 14197 17289 14231 17323
rect 14749 17289 14783 17323
rect 17049 17289 17083 17323
rect 21281 17289 21315 17323
rect 22477 17289 22511 17323
rect 22569 17289 22603 17323
rect 23857 17289 23891 17323
rect 29653 17289 29687 17323
rect 30757 17289 30791 17323
rect 34069 17289 34103 17323
rect 35909 17289 35943 17323
rect 15485 17221 15519 17255
rect 15945 17221 15979 17255
rect 18153 17221 18187 17255
rect 23949 17221 23983 17255
rect 31585 17221 31619 17255
rect 1777 17153 1811 17187
rect 3617 17153 3651 17187
rect 5641 17153 5675 17187
rect 6561 17153 6595 17187
rect 7205 17153 7239 17187
rect 9229 17153 9263 17187
rect 10885 17153 10919 17187
rect 11713 17153 11747 17187
rect 16957 17153 16991 17187
rect 17417 17153 17451 17187
rect 20453 17153 20487 17187
rect 21465 17153 21499 17187
rect 24685 17153 24719 17187
rect 26801 17153 26835 17187
rect 27905 17153 27939 17187
rect 30113 17153 30147 17187
rect 32321 17153 32355 17187
rect 33425 17153 33459 17187
rect 34621 17153 34655 17187
rect 2053 17085 2087 17119
rect 4169 17085 4203 17119
rect 5917 17085 5951 17119
rect 8125 17085 8159 17119
rect 8217 17085 8251 17119
rect 9321 17085 9355 17119
rect 9505 17085 9539 17119
rect 10977 17085 11011 17119
rect 11989 17085 12023 17119
rect 14841 17085 14875 17119
rect 15025 17085 15059 17119
rect 16037 17085 16071 17119
rect 16221 17085 16255 17119
rect 17877 17085 17911 17119
rect 20545 17085 20579 17119
rect 20637 17085 20671 17119
rect 22753 17085 22787 17119
rect 24133 17085 24167 17119
rect 24961 17085 24995 17119
rect 27261 17085 27295 17119
rect 28181 17085 28215 17119
rect 35265 17085 35299 17119
rect 8861 17017 8895 17051
rect 13921 17017 13955 17051
rect 14381 17017 14415 17051
rect 19625 17017 19659 17051
rect 20085 17017 20119 17051
rect 22109 17017 22143 17051
rect 23213 17017 23247 17051
rect 26433 17017 26467 17051
rect 31769 17017 31803 17051
rect 7665 16949 7699 16983
rect 10057 16949 10091 16983
rect 10425 16949 10459 16983
rect 13461 16949 13495 16983
rect 14105 16949 14139 16983
rect 15577 16949 15611 16983
rect 23489 16949 23523 16983
rect 31033 16949 31067 16983
rect 32965 16949 32999 16983
rect 34713 16949 34747 16983
rect 6101 16745 6135 16779
rect 9229 16745 9263 16779
rect 15393 16745 15427 16779
rect 15761 16745 15795 16779
rect 16681 16745 16715 16779
rect 19698 16745 19732 16779
rect 27445 16745 27479 16779
rect 29377 16745 29411 16779
rect 29653 16745 29687 16779
rect 3433 16677 3467 16711
rect 17141 16677 17175 16711
rect 21833 16677 21867 16711
rect 3525 16609 3559 16643
rect 7205 16609 7239 16643
rect 8493 16609 8527 16643
rect 9689 16609 9723 16643
rect 9873 16609 9907 16643
rect 10885 16609 10919 16643
rect 11069 16609 11103 16643
rect 12449 16609 12483 16643
rect 13645 16609 13679 16643
rect 14841 16609 14875 16643
rect 17601 16609 17635 16643
rect 17785 16609 17819 16643
rect 18981 16609 19015 16643
rect 19441 16609 19475 16643
rect 23765 16609 23799 16643
rect 23949 16609 23983 16643
rect 24501 16609 24535 16643
rect 25329 16609 25363 16643
rect 26525 16609 26559 16643
rect 27905 16609 27939 16643
rect 28089 16609 28123 16643
rect 30665 16609 30699 16643
rect 30941 16609 30975 16643
rect 32229 16609 32263 16643
rect 33241 16609 33275 16643
rect 33517 16609 33551 16643
rect 1777 16541 1811 16575
rect 4169 16541 4203 16575
rect 4997 16541 5031 16575
rect 7113 16541 7147 16575
rect 11529 16541 11563 16575
rect 12265 16541 12299 16575
rect 13369 16541 13403 16575
rect 15577 16541 15611 16575
rect 16037 16541 16071 16575
rect 18429 16541 18463 16575
rect 21465 16541 21499 16575
rect 22201 16541 22235 16575
rect 22845 16541 22879 16575
rect 26341 16541 26375 16575
rect 27813 16541 27847 16575
rect 28825 16541 28859 16575
rect 30205 16541 30239 16575
rect 31953 16541 31987 16575
rect 2513 16473 2547 16507
rect 6009 16473 6043 16507
rect 7021 16473 7055 16507
rect 8217 16473 8251 16507
rect 14657 16473 14691 16507
rect 14749 16473 14783 16507
rect 17509 16473 17543 16507
rect 23673 16473 23707 16507
rect 34989 16473 35023 16507
rect 35449 16473 35483 16507
rect 6653 16405 6687 16439
rect 7849 16405 7883 16439
rect 8309 16405 8343 16439
rect 9597 16405 9631 16439
rect 10425 16405 10459 16439
rect 10793 16405 10827 16439
rect 11805 16405 11839 16439
rect 12173 16405 12207 16439
rect 13001 16405 13035 16439
rect 13461 16405 13495 16439
rect 14105 16405 14139 16439
rect 14289 16405 14323 16439
rect 18521 16405 18555 16439
rect 23305 16405 23339 16439
rect 24777 16405 24811 16439
rect 25145 16405 25179 16439
rect 25237 16405 25271 16439
rect 25973 16405 26007 16439
rect 26433 16405 26467 16439
rect 27077 16405 27111 16439
rect 28641 16405 28675 16439
rect 29101 16405 29135 16439
rect 30021 16405 30055 16439
rect 35081 16405 35115 16439
rect 5641 16201 5675 16235
rect 9137 16201 9171 16235
rect 9229 16201 9263 16235
rect 10425 16201 10459 16235
rect 11345 16201 11379 16235
rect 11713 16201 11747 16235
rect 19349 16201 19383 16235
rect 19809 16201 19843 16235
rect 22017 16201 22051 16235
rect 22385 16201 22419 16235
rect 26617 16201 26651 16235
rect 4629 16133 4663 16167
rect 5733 16133 5767 16167
rect 11069 16133 11103 16167
rect 12449 16133 12483 16167
rect 21005 16133 21039 16167
rect 22477 16133 22511 16167
rect 31125 16133 31159 16167
rect 1777 16065 1811 16099
rect 3617 16065 3651 16099
rect 6929 16065 6963 16099
rect 7941 16065 7975 16099
rect 12357 16065 12391 16099
rect 13369 16065 13403 16099
rect 14841 16065 14875 16099
rect 14933 16065 14967 16099
rect 15669 16065 15703 16099
rect 19717 16065 19751 16099
rect 20913 16065 20947 16099
rect 23213 16065 23247 16099
rect 23489 16065 23523 16099
rect 23765 16065 23799 16099
rect 24869 16065 24903 16099
rect 27169 16065 27203 16099
rect 28273 16065 28307 16099
rect 30481 16065 30515 16099
rect 31769 16065 31803 16099
rect 32597 16065 32631 16099
rect 33793 16065 33827 16099
rect 34069 16065 34103 16099
rect 2053 15997 2087 16031
rect 5825 15997 5859 16031
rect 8033 15997 8067 16031
rect 8125 15997 8159 16031
rect 9321 15997 9355 16031
rect 10517 15997 10551 16031
rect 10609 15997 10643 16031
rect 11805 15997 11839 16031
rect 12633 15997 12667 16031
rect 15117 15997 15151 16031
rect 16865 15997 16899 16031
rect 17141 15997 17175 16031
rect 19901 15997 19935 16031
rect 21189 15997 21223 16031
rect 22569 15997 22603 16031
rect 25145 15997 25179 16031
rect 27813 15997 27847 16031
rect 29469 15997 29503 16031
rect 32321 15997 32355 16031
rect 7113 15929 7147 15963
rect 7573 15929 7607 15963
rect 11989 15929 12023 15963
rect 14473 15929 14507 15963
rect 19073 15929 19107 15963
rect 20545 15929 20579 15963
rect 21649 15929 21683 15963
rect 28917 15929 28951 15963
rect 5273 15861 5307 15895
rect 6561 15861 6595 15895
rect 8769 15861 8803 15895
rect 10057 15861 10091 15895
rect 13093 15861 13127 15895
rect 14013 15861 14047 15895
rect 14289 15861 14323 15895
rect 16313 15861 16347 15895
rect 18613 15861 18647 15895
rect 23029 15861 23063 15895
rect 24409 15861 24443 15895
rect 30021 15861 30055 15895
rect 31585 15861 31619 15895
rect 33609 15861 33643 15895
rect 7573 15657 7607 15691
rect 14473 15657 14507 15691
rect 16497 15657 16531 15691
rect 19533 15657 19567 15691
rect 27813 15657 27847 15691
rect 27997 15657 28031 15691
rect 32413 15657 32447 15691
rect 3617 15589 3651 15623
rect 20545 15589 20579 15623
rect 31953 15589 31987 15623
rect 2053 15521 2087 15555
rect 4997 15521 5031 15555
rect 5273 15521 5307 15555
rect 8033 15521 8067 15555
rect 8125 15521 8159 15555
rect 9689 15521 9723 15555
rect 10977 15521 11011 15555
rect 14749 15521 14783 15555
rect 19073 15521 19107 15555
rect 20177 15521 20211 15555
rect 23949 15521 23983 15555
rect 24593 15521 24627 15555
rect 24869 15521 24903 15555
rect 25973 15521 26007 15555
rect 26985 15521 27019 15555
rect 27537 15521 27571 15555
rect 1777 15453 1811 15487
rect 4353 15453 4387 15487
rect 8677 15453 8711 15487
rect 9505 15453 9539 15487
rect 11621 15453 11655 15487
rect 13921 15453 13955 15487
rect 16957 15453 16991 15487
rect 21005 15453 21039 15487
rect 25881 15453 25915 15487
rect 26893 15453 26927 15487
rect 27721 15453 27755 15487
rect 28365 15453 28399 15487
rect 28641 15453 28675 15487
rect 29745 15453 29779 15487
rect 30021 15453 30055 15487
rect 31493 15453 31527 15487
rect 32137 15453 32171 15487
rect 32781 15453 32815 15487
rect 3433 15385 3467 15419
rect 7021 15385 7055 15419
rect 7941 15385 7975 15419
rect 10885 15385 10919 15419
rect 11897 15385 11931 15419
rect 13737 15385 13771 15419
rect 15025 15385 15059 15419
rect 17220 15385 17254 15419
rect 19993 15385 20027 15419
rect 21281 15385 21315 15419
rect 23673 15385 23707 15419
rect 30849 15385 30883 15419
rect 3985 15317 4019 15351
rect 4445 15317 4479 15351
rect 9137 15317 9171 15351
rect 9597 15317 9631 15351
rect 10425 15317 10459 15351
rect 10793 15317 10827 15351
rect 13369 15317 13403 15351
rect 14105 15317 14139 15351
rect 18705 15317 18739 15351
rect 19901 15317 19935 15351
rect 22753 15317 22787 15351
rect 23305 15317 23339 15351
rect 23765 15317 23799 15351
rect 26433 15317 26467 15351
rect 26801 15317 26835 15351
rect 31309 15317 31343 15351
rect 32597 15317 32631 15351
rect 4537 15113 4571 15147
rect 5733 15113 5767 15147
rect 8033 15113 8067 15147
rect 9689 15113 9723 15147
rect 11621 15113 11655 15147
rect 12265 15113 12299 15147
rect 12725 15113 12759 15147
rect 14381 15113 14415 15147
rect 15577 15113 15611 15147
rect 21465 15113 21499 15147
rect 5641 15045 5675 15079
rect 9597 15045 9631 15079
rect 12633 15045 12667 15079
rect 13737 15045 13771 15079
rect 19993 15045 20027 15079
rect 24593 15045 24627 15079
rect 1777 14977 1811 15011
rect 3617 14977 3651 15011
rect 4445 14977 4479 15011
rect 6653 14977 6687 15011
rect 7941 14977 7975 15011
rect 10793 14977 10827 15011
rect 13553 14977 13587 15011
rect 14749 14977 14783 15011
rect 15945 14977 15979 15011
rect 16037 14977 16071 15011
rect 16681 14977 16715 15011
rect 17233 14977 17267 15011
rect 22293 14977 22327 15011
rect 24409 14977 24443 15011
rect 27629 14977 27663 15011
rect 28733 14977 28767 15011
rect 29837 14977 29871 15011
rect 30941 14977 30975 15011
rect 2053 14909 2087 14943
rect 4721 14909 4755 14943
rect 5825 14909 5859 14943
rect 8125 14909 8159 14943
rect 8953 14909 8987 14943
rect 9781 14909 9815 14943
rect 10885 14909 10919 14943
rect 11069 14909 11103 14943
rect 12817 14909 12851 14943
rect 14105 14909 14139 14943
rect 14841 14909 14875 14943
rect 15025 14909 15059 14943
rect 16221 14909 16255 14943
rect 18981 14909 19015 14943
rect 19717 14909 19751 14943
rect 22569 14909 22603 14943
rect 24869 14909 24903 14943
rect 25145 14909 25179 14943
rect 28273 14909 28307 14943
rect 6837 14841 6871 14875
rect 16865 14841 16899 14875
rect 24041 14841 24075 14875
rect 27169 14841 27203 14875
rect 3433 14773 3467 14807
rect 4077 14773 4111 14807
rect 5273 14773 5307 14807
rect 7205 14773 7239 14807
rect 7573 14773 7607 14807
rect 8769 14773 8803 14807
rect 9229 14773 9263 14807
rect 10425 14773 10459 14807
rect 11805 14773 11839 14807
rect 11989 14773 12023 14807
rect 19349 14773 19383 14807
rect 21833 14773 21867 14807
rect 26617 14773 26651 14807
rect 27077 14773 27111 14807
rect 29377 14773 29411 14807
rect 30481 14773 30515 14807
rect 31585 14773 31619 14807
rect 31861 14773 31895 14807
rect 3433 14569 3467 14603
rect 3893 14569 3927 14603
rect 13553 14569 13587 14603
rect 13921 14569 13955 14603
rect 18889 14569 18923 14603
rect 28917 14569 28951 14603
rect 30389 14569 30423 14603
rect 8585 14501 8619 14535
rect 10425 14501 10459 14535
rect 24409 14501 24443 14535
rect 26249 14501 26283 14535
rect 26433 14501 26467 14535
rect 2053 14433 2087 14467
rect 3985 14433 4019 14467
rect 5089 14433 5123 14467
rect 5273 14433 5307 14467
rect 10885 14433 10919 14467
rect 10977 14433 11011 14467
rect 14197 14433 14231 14467
rect 17141 14433 17175 14467
rect 20177 14433 20211 14467
rect 20913 14433 20947 14467
rect 21925 14433 21959 14467
rect 23305 14433 23339 14467
rect 24041 14433 24075 14467
rect 25881 14433 25915 14467
rect 31125 14433 31159 14467
rect 1777 14365 1811 14399
rect 5825 14365 5859 14399
rect 8401 14365 8435 14399
rect 8953 14365 8987 14399
rect 9137 14365 9171 14399
rect 9413 14365 9447 14399
rect 10793 14365 10827 14399
rect 11805 14365 11839 14399
rect 14657 14365 14691 14399
rect 20637 14365 20671 14399
rect 21741 14365 21775 14399
rect 25605 14365 25639 14399
rect 27169 14365 27203 14399
rect 28273 14365 28307 14399
rect 29745 14365 29779 14399
rect 30849 14365 30883 14399
rect 4997 14297 5031 14331
rect 6101 14297 6135 14331
rect 7849 14297 7883 14331
rect 11437 14297 11471 14331
rect 12081 14297 12115 14331
rect 14933 14297 14967 14331
rect 17417 14297 17451 14331
rect 19441 14297 19475 14331
rect 21097 14297 21131 14331
rect 22569 14297 22603 14331
rect 23857 14297 23891 14331
rect 24869 14297 24903 14331
rect 3617 14229 3651 14263
rect 4629 14229 4663 14263
rect 16405 14229 16439 14263
rect 16773 14229 16807 14263
rect 21373 14229 21407 14263
rect 21833 14229 21867 14263
rect 24133 14229 24167 14263
rect 24777 14229 24811 14263
rect 25237 14229 25271 14263
rect 25697 14229 25731 14263
rect 26617 14229 26651 14263
rect 27813 14229 27847 14263
rect 29377 14229 29411 14263
rect 7389 14025 7423 14059
rect 8125 14025 8159 14059
rect 8585 14025 8619 14059
rect 12173 14025 12207 14059
rect 15577 14025 15611 14059
rect 16405 14025 16439 14059
rect 16681 14025 16715 14059
rect 19533 14025 19567 14059
rect 19901 14025 19935 14059
rect 19993 14025 20027 14059
rect 20729 14025 20763 14059
rect 22201 14025 22235 14059
rect 23029 14025 23063 14059
rect 23857 14025 23891 14059
rect 24225 14025 24259 14059
rect 25513 14025 25547 14059
rect 25605 14025 25639 14059
rect 26249 14025 26283 14059
rect 26341 14025 26375 14059
rect 29653 14025 29687 14059
rect 30297 14025 30331 14059
rect 3709 13957 3743 13991
rect 6009 13957 6043 13991
rect 6561 13957 6595 13991
rect 7297 13957 7331 13991
rect 13553 13957 13587 13991
rect 14381 13957 14415 13991
rect 17417 13957 17451 13991
rect 29193 13957 29227 13991
rect 1593 13889 1627 13923
rect 3985 13889 4019 13923
rect 8493 13889 8527 13923
rect 11805 13889 11839 13923
rect 12541 13889 12575 13923
rect 13277 13889 13311 13923
rect 14289 13889 14323 13923
rect 15669 13889 15703 13923
rect 16221 13889 16255 13923
rect 17141 13889 17175 13923
rect 21097 13889 21131 13923
rect 21189 13889 21223 13923
rect 21925 13889 21959 13923
rect 24317 13889 24351 13923
rect 27169 13889 27203 13923
rect 28549 13889 28583 13923
rect 29837 13889 29871 13923
rect 30481 13889 30515 13923
rect 30757 13889 30791 13923
rect 2053 13821 2087 13855
rect 3525 13821 3559 13855
rect 6377 13821 6411 13855
rect 7481 13821 7515 13855
rect 8677 13821 8711 13855
rect 9321 13821 9355 13855
rect 12633 13821 12667 13855
rect 12817 13821 12851 13855
rect 13369 13821 13403 13855
rect 14565 13821 14599 13855
rect 15761 13821 15795 13855
rect 18889 13821 18923 13855
rect 20085 13821 20119 13855
rect 21281 13821 21315 13855
rect 22293 13821 22327 13855
rect 23121 13821 23155 13855
rect 23213 13821 23247 13855
rect 24409 13821 24443 13855
rect 25789 13821 25823 13855
rect 3341 13753 3375 13787
rect 11529 13753 11563 13787
rect 13921 13753 13955 13787
rect 15209 13753 15243 13787
rect 4242 13685 4276 13719
rect 6929 13685 6963 13719
rect 9584 13685 9618 13719
rect 11069 13685 11103 13719
rect 13737 13685 13771 13719
rect 19257 13685 19291 13719
rect 22661 13685 22695 13719
rect 25145 13685 25179 13719
rect 27813 13685 27847 13719
rect 3617 13481 3651 13515
rect 3985 13481 4019 13515
rect 8585 13481 8619 13515
rect 16313 13481 16347 13515
rect 16497 13481 16531 13515
rect 16957 13481 16991 13515
rect 23857 13481 23891 13515
rect 4445 13413 4479 13447
rect 9137 13413 9171 13447
rect 18153 13413 18187 13447
rect 19349 13413 19383 13447
rect 29653 13413 29687 13447
rect 2053 13345 2087 13379
rect 4905 13345 4939 13379
rect 4997 13345 5031 13379
rect 6101 13345 6135 13379
rect 6285 13345 6319 13379
rect 9781 13345 9815 13379
rect 10885 13345 10919 13379
rect 11897 13345 11931 13379
rect 14289 13345 14323 13379
rect 17417 13345 17451 13379
rect 17601 13345 17635 13379
rect 18613 13345 18647 13379
rect 18797 13345 18831 13379
rect 19625 13345 19659 13379
rect 22017 13345 22051 13379
rect 25145 13345 25179 13379
rect 1593 13277 1627 13311
rect 4077 13277 4111 13311
rect 6837 13277 6871 13311
rect 9597 13277 9631 13311
rect 10701 13277 10735 13311
rect 18521 13277 18555 13311
rect 20269 13277 20303 13311
rect 22477 13277 22511 13311
rect 24041 13277 24075 13311
rect 24961 13277 24995 13311
rect 25789 13277 25823 13311
rect 27169 13277 27203 13311
rect 28273 13277 28307 13311
rect 4813 13209 4847 13243
rect 6009 13209 6043 13243
rect 7113 13209 7147 13243
rect 10793 13209 10827 13243
rect 11621 13209 11655 13243
rect 12173 13209 12207 13243
rect 14565 13209 14599 13243
rect 20545 13209 20579 13243
rect 23213 13209 23247 13243
rect 27813 13209 27847 13243
rect 28917 13209 28951 13243
rect 3433 13141 3467 13175
rect 5641 13141 5675 13175
rect 9505 13141 9539 13175
rect 10333 13141 10367 13175
rect 11345 13141 11379 13175
rect 13645 13141 13679 13175
rect 16037 13141 16071 13175
rect 17325 13141 17359 13175
rect 24593 13141 24627 13175
rect 25053 13141 25087 13175
rect 26433 13141 26467 13175
rect 26709 13141 26743 13175
rect 2973 12937 3007 12971
rect 5917 12937 5951 12971
rect 10885 12937 10919 12971
rect 11989 12937 12023 12971
rect 12449 12937 12483 12971
rect 13645 12937 13679 12971
rect 16957 12937 16991 12971
rect 17693 12937 17727 12971
rect 22569 12937 22603 12971
rect 4445 12869 4479 12903
rect 10057 12869 10091 12903
rect 10793 12869 10827 12903
rect 14841 12869 14875 12903
rect 16681 12869 16715 12903
rect 23213 12869 23247 12903
rect 25145 12869 25179 12903
rect 25881 12869 25915 12903
rect 1869 12801 1903 12835
rect 3341 12801 3375 12835
rect 4169 12801 4203 12835
rect 6469 12801 6503 12835
rect 6561 12801 6595 12835
rect 7205 12801 7239 12835
rect 11621 12801 11655 12835
rect 12357 12801 12391 12835
rect 13553 12801 13587 12835
rect 14289 12801 14323 12835
rect 14749 12801 14783 12835
rect 15945 12801 15979 12835
rect 16037 12801 16071 12835
rect 17601 12801 17635 12835
rect 18429 12801 18463 12835
rect 18705 12801 18739 12835
rect 19717 12801 19751 12835
rect 22109 12801 22143 12835
rect 26341 12801 26375 12835
rect 27169 12801 27203 12835
rect 28365 12801 28399 12835
rect 1593 12733 1627 12767
rect 3433 12733 3467 12767
rect 3525 12733 3559 12767
rect 7665 12733 7699 12767
rect 7941 12733 7975 12767
rect 9689 12733 9723 12767
rect 11069 12733 11103 12767
rect 12541 12733 12575 12767
rect 13829 12733 13863 12767
rect 15025 12733 15059 12767
rect 16221 12733 16255 12767
rect 17877 12733 17911 12767
rect 19993 12733 20027 12767
rect 22937 12733 22971 12767
rect 24685 12733 24719 12767
rect 28917 12733 28951 12767
rect 13185 12665 13219 12699
rect 22293 12665 22327 12699
rect 10425 12597 10459 12631
rect 14381 12597 14415 12631
rect 15577 12597 15611 12631
rect 17233 12597 17267 12631
rect 21465 12597 21499 12631
rect 26525 12597 26559 12631
rect 27813 12597 27847 12631
rect 2237 12393 2271 12427
rect 4077 12393 4111 12427
rect 9045 12393 9079 12427
rect 9413 12393 9447 12427
rect 13001 12393 13035 12427
rect 18889 12393 18923 12427
rect 25697 12393 25731 12427
rect 28457 12393 28491 12427
rect 4997 12325 5031 12359
rect 11805 12325 11839 12359
rect 14105 12325 14139 12359
rect 18981 12325 19015 12359
rect 8585 12257 8619 12291
rect 9965 12257 9999 12291
rect 11161 12257 11195 12291
rect 12357 12257 12391 12291
rect 13553 12257 13587 12291
rect 15485 12257 15519 12291
rect 16129 12257 16163 12291
rect 18337 12257 18371 12291
rect 19441 12257 19475 12291
rect 20085 12257 20119 12291
rect 22293 12257 22327 12291
rect 2789 12189 2823 12223
rect 4353 12189 4387 12223
rect 5457 12189 5491 12223
rect 7481 12189 7515 12223
rect 7941 12189 7975 12223
rect 12265 12189 12299 12223
rect 13461 12189 13495 12223
rect 25053 12189 25087 12223
rect 27169 12189 27203 12223
rect 2145 12121 2179 12155
rect 3433 12121 3467 12155
rect 5733 12121 5767 12155
rect 10977 12121 11011 12155
rect 12173 12121 12207 12155
rect 14473 12121 14507 12155
rect 14749 12121 14783 12155
rect 16405 12121 16439 12155
rect 20361 12121 20395 12155
rect 22569 12121 22603 12155
rect 28365 12121 28399 12155
rect 28825 12121 28859 12155
rect 1593 12053 1627 12087
rect 1777 12053 1811 12087
rect 3801 12053 3835 12087
rect 9781 12053 9815 12087
rect 9873 12053 9907 12087
rect 10609 12053 10643 12087
rect 11069 12053 11103 12087
rect 13369 12053 13403 12087
rect 17877 12053 17911 12087
rect 21833 12053 21867 12087
rect 24041 12053 24075 12087
rect 24501 12053 24535 12087
rect 27813 12053 27847 12087
rect 1409 11849 1443 11883
rect 2605 11849 2639 11883
rect 11989 11849 12023 11883
rect 15485 11849 15519 11883
rect 17325 11849 17359 11883
rect 17417 11849 17451 11883
rect 21649 11849 21683 11883
rect 24593 11849 24627 11883
rect 28273 11849 28307 11883
rect 5641 11781 5675 11815
rect 6469 11781 6503 11815
rect 6561 11781 6595 11815
rect 7481 11781 7515 11815
rect 10149 11781 10183 11815
rect 10977 11781 11011 11815
rect 11713 11781 11747 11815
rect 13461 11781 13495 11815
rect 21833 11781 21867 11815
rect 1961 11713 1995 11747
rect 3065 11713 3099 11747
rect 4169 11713 4203 11747
rect 7205 11713 7239 11747
rect 9413 11713 9447 11747
rect 11161 11713 11195 11747
rect 12357 11713 12391 11747
rect 12449 11713 12483 11747
rect 13185 11713 13219 11747
rect 15853 11713 15887 11747
rect 20453 11713 20487 11747
rect 20729 11713 20763 11747
rect 22477 11713 22511 11747
rect 25697 11713 25731 11747
rect 27169 11713 27203 11747
rect 5733 11645 5767 11679
rect 5825 11645 5859 11679
rect 12633 11645 12667 11679
rect 15945 11645 15979 11679
rect 16129 11645 16163 11679
rect 17601 11645 17635 11679
rect 18245 11645 18279 11679
rect 18521 11645 18555 11679
rect 22753 11645 22787 11679
rect 26341 11645 26375 11679
rect 4813 11577 4847 11611
rect 14933 11577 14967 11611
rect 22109 11577 22143 11611
rect 1593 11509 1627 11543
rect 3709 11509 3743 11543
rect 5273 11509 5307 11543
rect 8953 11509 8987 11543
rect 16957 11509 16991 11543
rect 19993 11509 20027 11543
rect 24225 11509 24259 11543
rect 27813 11509 27847 11543
rect 2329 11305 2363 11339
rect 3433 11305 3467 11339
rect 7205 11305 7239 11339
rect 13829 11305 13863 11339
rect 17398 11305 17432 11339
rect 23213 11305 23247 11339
rect 26341 11305 26375 11339
rect 32137 11305 32171 11339
rect 4261 11237 4295 11271
rect 11069 11237 11103 11271
rect 14381 11237 14415 11271
rect 18889 11237 18923 11271
rect 20637 11237 20671 11271
rect 25237 11237 25271 11271
rect 27445 11237 27479 11271
rect 4813 11169 4847 11203
rect 6561 11169 6595 11203
rect 8309 11169 8343 11203
rect 8401 11169 8435 11203
rect 9137 11169 9171 11203
rect 9965 11169 9999 11203
rect 10149 11169 10183 11203
rect 13277 11169 13311 11203
rect 13645 11169 13679 11203
rect 16405 11169 16439 11203
rect 17141 11169 17175 11203
rect 20177 11169 20211 11203
rect 21005 11169 21039 11203
rect 22753 11169 22787 11203
rect 23673 11169 23707 11203
rect 23765 11169 23799 11203
rect 29745 11169 29779 11203
rect 1685 11101 1719 11135
rect 2789 11101 2823 11135
rect 4077 11101 4111 11135
rect 8953 11101 8987 11135
rect 9873 11101 9907 11135
rect 11529 11101 11563 11135
rect 14657 11101 14691 11135
rect 19441 11101 19475 11135
rect 23581 11101 23615 11135
rect 24593 11101 24627 11135
rect 25697 11101 25731 11135
rect 26801 11101 26835 11135
rect 28917 11101 28951 11135
rect 5089 11033 5123 11067
rect 7113 11033 7147 11067
rect 8217 11033 8251 11067
rect 10885 11033 10919 11067
rect 11805 11033 11839 11067
rect 14197 11033 14231 11067
rect 14933 11033 14967 11067
rect 16773 11033 16807 11067
rect 21281 11033 21315 11067
rect 27997 11033 28031 11067
rect 28181 11033 28215 11067
rect 28733 11033 28767 11067
rect 29193 11033 29227 11067
rect 30021 11033 30055 11067
rect 31769 11033 31803 11067
rect 7849 10965 7883 10999
rect 9505 10965 9539 10999
rect 1593 10761 1627 10795
rect 6929 10761 6963 10795
rect 11713 10761 11747 10795
rect 14565 10761 14599 10795
rect 16313 10761 16347 10795
rect 22385 10761 22419 10795
rect 22477 10761 22511 10795
rect 29469 10761 29503 10795
rect 6009 10693 6043 10727
rect 10241 10693 10275 10727
rect 14933 10693 14967 10727
rect 15761 10693 15795 10727
rect 17785 10693 17819 10727
rect 27261 10693 27295 10727
rect 1961 10625 1995 10659
rect 3065 10625 3099 10659
rect 4169 10625 4203 10659
rect 5365 10625 5399 10659
rect 7021 10625 7055 10659
rect 12265 10625 12299 10659
rect 16129 10625 16163 10659
rect 17509 10625 17543 10659
rect 19717 10625 19751 10659
rect 23121 10625 23155 10659
rect 23489 10625 23523 10659
rect 24593 10625 24627 10659
rect 25237 10625 25271 10659
rect 25697 10625 25731 10659
rect 27445 10625 27479 10659
rect 28825 10625 28859 10659
rect 7205 10557 7239 10591
rect 7757 10557 7791 10591
rect 8033 10557 8067 10591
rect 9781 10557 9815 10591
rect 10977 10557 11011 10591
rect 12541 10557 12575 10591
rect 16865 10557 16899 10591
rect 19993 10557 20027 10591
rect 22569 10557 22603 10591
rect 24133 10557 24167 10591
rect 1501 10489 1535 10523
rect 22017 10489 22051 10523
rect 26341 10489 26375 10523
rect 2605 10421 2639 10455
rect 3709 10421 3743 10455
rect 4813 10421 4847 10455
rect 6561 10421 6595 10455
rect 11621 10421 11655 10455
rect 11989 10421 12023 10455
rect 14013 10421 14047 10455
rect 14381 10421 14415 10455
rect 19257 10421 19291 10455
rect 21465 10421 21499 10455
rect 27721 10421 27755 10455
rect 3433 10217 3467 10251
rect 11253 10217 11287 10251
rect 19073 10217 19107 10251
rect 3985 10149 4019 10183
rect 7205 10149 7239 10183
rect 10885 10149 10919 10183
rect 13829 10149 13863 10183
rect 16221 10149 16255 10183
rect 18705 10149 18739 10183
rect 23857 10149 23891 10183
rect 27215 10149 27249 10183
rect 6101 10081 6135 10115
rect 8309 10081 8343 10115
rect 8401 10081 8435 10115
rect 11529 10081 11563 10115
rect 13553 10081 13587 10115
rect 16681 10081 16715 10115
rect 18429 10081 18463 10115
rect 19809 10081 19843 10115
rect 1685 10013 1719 10047
rect 2789 10013 2823 10047
rect 4261 10013 4295 10047
rect 5457 10013 5491 10047
rect 6561 10013 6595 10047
rect 9137 10013 9171 10047
rect 14473 10013 14507 10047
rect 19533 10013 19567 10047
rect 22109 10013 22143 10047
rect 23213 10013 23247 10047
rect 24961 10013 24995 10047
rect 25421 10013 25455 10047
rect 26985 10013 27019 10047
rect 9413 9945 9447 9979
rect 11805 9945 11839 9979
rect 14749 9945 14783 9979
rect 16957 9945 16991 9979
rect 2329 9877 2363 9911
rect 4905 9877 4939 9911
rect 7481 9877 7515 9911
rect 7849 9877 7883 9911
rect 8217 9877 8251 9911
rect 13277 9877 13311 9911
rect 14197 9877 14231 9911
rect 21281 9877 21315 9911
rect 22753 9877 22787 9911
rect 24777 9877 24811 9911
rect 26065 9877 26099 9911
rect 26617 9877 26651 9911
rect 28273 9877 28307 9911
rect 6561 9673 6595 9707
rect 27813 9673 27847 9707
rect 11253 9605 11287 9639
rect 14749 9605 14783 9639
rect 19901 9605 19935 9639
rect 23857 9605 23891 9639
rect 2053 9537 2087 9571
rect 3157 9537 3191 9571
rect 4261 9537 4295 9571
rect 5365 9537 5399 9571
rect 6009 9537 6043 9571
rect 6745 9537 6779 9571
rect 7573 9537 7607 9571
rect 7665 9537 7699 9571
rect 10793 9537 10827 9571
rect 11713 9537 11747 9571
rect 14473 9537 14507 9571
rect 19809 9537 19843 9571
rect 20637 9537 20671 9571
rect 22017 9537 22051 9571
rect 23213 9537 23247 9571
rect 24593 9537 24627 9571
rect 25697 9537 25731 9571
rect 27169 9537 27203 9571
rect 3801 9469 3835 9503
rect 4905 9469 4939 9503
rect 7757 9469 7791 9503
rect 8493 9469 8527 9503
rect 8769 9469 8803 9503
rect 10977 9469 11011 9503
rect 16221 9469 16255 9503
rect 16865 9469 16899 9503
rect 17141 9469 17175 9503
rect 20085 9469 20119 9503
rect 1593 9401 1627 9435
rect 13737 9401 13771 9435
rect 19441 9401 19475 9435
rect 25237 9401 25271 9435
rect 26341 9401 26375 9435
rect 1685 9333 1719 9367
rect 2697 9333 2731 9367
rect 7205 9333 7239 9367
rect 10241 9333 10275 9367
rect 11970 9333 12004 9367
rect 13461 9333 13495 9367
rect 13921 9333 13955 9367
rect 14197 9333 14231 9367
rect 18613 9333 18647 9367
rect 21281 9333 21315 9367
rect 22661 9333 22695 9367
rect 3801 9129 3835 9163
rect 13737 9129 13771 9163
rect 14289 9129 14323 9163
rect 20085 9129 20119 9163
rect 23765 9129 23799 9163
rect 26341 9129 26375 9163
rect 27445 9129 27479 9163
rect 28273 9129 28307 9163
rect 2329 9061 2363 9095
rect 6285 9061 6319 9095
rect 12725 9061 12759 9095
rect 22661 9061 22695 9095
rect 12173 8993 12207 9027
rect 14933 8993 14967 9027
rect 16221 8993 16255 9027
rect 21557 8993 21591 9027
rect 1685 8925 1719 8959
rect 2789 8925 2823 8959
rect 4261 8925 4295 8959
rect 5641 8925 5675 8959
rect 6745 8925 6779 8959
rect 7941 8925 7975 8959
rect 9137 8925 9171 8959
rect 11989 8925 12023 8959
rect 13093 8925 13127 8959
rect 17141 8925 17175 8959
rect 18245 8925 18279 8959
rect 18889 8925 18923 8959
rect 19441 8925 19475 8959
rect 20913 8925 20947 8959
rect 22028 8925 22062 8959
rect 23121 8925 23155 8959
rect 24593 8925 24627 8959
rect 25697 8925 25731 8959
rect 27169 8925 27203 8959
rect 9781 8857 9815 8891
rect 10241 8857 10275 8891
rect 10977 8857 11011 8891
rect 14657 8857 14691 8891
rect 17785 8857 17819 8891
rect 3433 8789 3467 8823
rect 4905 8789 4939 8823
rect 5273 8789 5307 8823
rect 7389 8789 7423 8823
rect 8585 8789 8619 8823
rect 11621 8789 11655 8823
rect 12081 8789 12115 8823
rect 14749 8789 14783 8823
rect 15577 8789 15611 8823
rect 15945 8789 15979 8823
rect 16037 8789 16071 8823
rect 16589 8789 16623 8823
rect 16865 8789 16899 8823
rect 25237 8789 25271 8823
rect 27629 8789 27663 8823
rect 28089 8789 28123 8823
rect 1593 8585 1627 8619
rect 1685 8585 1719 8619
rect 3801 8585 3835 8619
rect 4905 8585 4939 8619
rect 6009 8585 6043 8619
rect 13185 8585 13219 8619
rect 19533 8585 19567 8619
rect 20637 8585 20671 8619
rect 22661 8585 22695 8619
rect 23765 8585 23799 8619
rect 24225 8585 24259 8619
rect 26065 8585 26099 8619
rect 7205 8517 7239 8551
rect 9781 8517 9815 8551
rect 16773 8517 16807 8551
rect 24685 8517 24719 8551
rect 25605 8517 25639 8551
rect 2053 8449 2087 8483
rect 3157 8449 3191 8483
rect 4261 8449 4295 8483
rect 5365 8449 5399 8483
rect 6561 8449 6595 8483
rect 7665 8449 7699 8483
rect 8309 8449 8343 8483
rect 8769 8449 8803 8483
rect 10793 8449 10827 8483
rect 11529 8449 11563 8483
rect 12357 8449 12391 8483
rect 13553 8449 13587 8483
rect 14657 8449 14691 8483
rect 15669 8449 15703 8483
rect 17417 8449 17451 8483
rect 18889 8449 18923 8483
rect 19993 8449 20027 8483
rect 22017 8449 22051 8483
rect 23121 8449 23155 8483
rect 24869 8449 24903 8483
rect 25421 8449 25455 8483
rect 10057 8381 10091 8415
rect 10885 8381 10919 8415
rect 10977 8381 11011 8415
rect 12449 8381 12483 8415
rect 12633 8381 12667 8415
rect 13645 8381 13679 8415
rect 13737 8381 13771 8415
rect 14381 8381 14415 8415
rect 18061 8381 18095 8415
rect 21097 8381 21131 8415
rect 10425 8313 10459 8347
rect 11989 8313 12023 8347
rect 2697 8245 2731 8279
rect 9413 8245 9447 8279
rect 9965 8245 9999 8279
rect 16313 8245 16347 8279
rect 2329 8041 2363 8075
rect 3433 8041 3467 8075
rect 4721 8041 4755 8075
rect 6193 8041 6227 8075
rect 7481 8041 7515 8075
rect 8585 8041 8619 8075
rect 9873 8041 9907 8075
rect 13737 8041 13771 8075
rect 17049 8041 17083 8075
rect 18153 8041 18187 8075
rect 22661 8041 22695 8075
rect 23765 8041 23799 8075
rect 14105 7973 14139 8007
rect 21557 7973 21591 8007
rect 5825 7905 5859 7939
rect 9229 7905 9263 7939
rect 10425 7905 10459 7939
rect 14657 7905 14691 7939
rect 18613 7905 18647 7939
rect 19441 7905 19475 7939
rect 24869 7905 24903 7939
rect 25237 7905 25271 7939
rect 1685 7837 1719 7871
rect 2789 7837 2823 7871
rect 4077 7837 4111 7871
rect 5181 7837 5215 7871
rect 6561 7837 6595 7871
rect 7941 7837 7975 7871
rect 10241 7837 10275 7871
rect 11529 7837 11563 7871
rect 11989 7837 12023 7871
rect 12633 7837 12667 7871
rect 13093 7837 13127 7871
rect 15301 7837 15335 7871
rect 16405 7837 16439 7871
rect 17509 7837 17543 7871
rect 19717 7837 19751 7871
rect 20913 7837 20947 7871
rect 22017 7837 22051 7871
rect 23121 7837 23155 7871
rect 11345 7769 11379 7803
rect 24685 7769 24719 7803
rect 7205 7701 7239 7735
rect 10333 7701 10367 7735
rect 10885 7701 10919 7735
rect 14289 7701 14323 7735
rect 15945 7701 15979 7735
rect 1501 7497 1535 7531
rect 2513 7497 2547 7531
rect 3617 7497 3651 7531
rect 4721 7497 4755 7531
rect 4997 7497 5031 7531
rect 9597 7497 9631 7531
rect 10057 7497 10091 7531
rect 11529 7497 11563 7531
rect 15209 7497 15243 7531
rect 16865 7497 16899 7531
rect 18337 7497 18371 7531
rect 20085 7497 20119 7531
rect 21465 7497 21499 7531
rect 23765 7497 23799 7531
rect 7389 7429 7423 7463
rect 11161 7429 11195 7463
rect 14013 7429 14047 7463
rect 18797 7429 18831 7463
rect 21189 7429 21223 7463
rect 22293 7429 22327 7463
rect 24869 7429 24903 7463
rect 1869 7361 1903 7395
rect 2973 7361 3007 7395
rect 4077 7361 4111 7395
rect 5365 7361 5399 7395
rect 6745 7361 6779 7395
rect 7849 7361 7883 7395
rect 8953 7361 8987 7395
rect 10425 7361 10459 7395
rect 12265 7361 12299 7395
rect 13369 7361 13403 7395
rect 14565 7361 14599 7395
rect 15669 7361 15703 7395
rect 17049 7361 17083 7395
rect 17693 7361 17727 7395
rect 19441 7361 19475 7395
rect 20545 7361 20579 7395
rect 22017 7361 22051 7395
rect 24225 7361 24259 7395
rect 6009 7293 6043 7327
rect 10517 7293 10551 7327
rect 10701 7293 10735 7327
rect 12909 7293 12943 7327
rect 11345 7225 11379 7259
rect 11897 7225 11931 7259
rect 24409 7225 24443 7259
rect 6469 7157 6503 7191
rect 8493 7157 8527 7191
rect 11713 7157 11747 7191
rect 16313 7157 16347 7191
rect 17325 7157 17359 7191
rect 6377 6953 6411 6987
rect 9873 6953 9907 6987
rect 20177 6953 20211 6987
rect 22477 6953 22511 6987
rect 23857 6953 23891 6987
rect 8585 6817 8619 6851
rect 10793 6817 10827 6851
rect 12633 6817 12667 6851
rect 13737 6817 13771 6851
rect 14565 6817 14599 6851
rect 16405 6817 16439 6851
rect 17417 6817 17451 6851
rect 18521 6817 18555 6851
rect 1685 6749 1719 6783
rect 2513 6749 2547 6783
rect 3433 6749 3467 6783
rect 3893 6749 3927 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 5273 6749 5307 6783
rect 5733 6749 5767 6783
rect 6837 6749 6871 6783
rect 7481 6749 7515 6783
rect 7941 6749 7975 6783
rect 9045 6749 9079 6783
rect 9137 6749 9171 6783
rect 11529 6749 11563 6783
rect 11989 6749 12023 6783
rect 13093 6749 13127 6783
rect 15209 6749 15243 6783
rect 15485 6749 15519 6783
rect 16773 6749 16807 6783
rect 17877 6749 17911 6783
rect 19533 6749 19567 6783
rect 20637 6749 20671 6783
rect 21281 6749 21315 6783
rect 21833 6749 21867 6783
rect 3249 6681 3283 6715
rect 9689 6681 9723 6715
rect 23029 6681 23063 6715
rect 23213 6681 23247 6715
rect 1777 6613 1811 6647
rect 2605 6613 2639 6647
rect 3985 6613 4019 6647
rect 10149 6613 10183 6647
rect 10517 6613 10551 6647
rect 10609 6613 10643 6647
rect 11345 6613 11379 6647
rect 4905 6409 4939 6443
rect 10057 6409 10091 6443
rect 12633 6409 12667 6443
rect 15209 6409 15243 6443
rect 17509 6409 17543 6443
rect 19717 6409 19751 6443
rect 20821 6409 20855 6443
rect 21281 6409 21315 6443
rect 23765 6409 23799 6443
rect 7849 6341 7883 6375
rect 8953 6341 8987 6375
rect 16313 6341 16347 6375
rect 1593 6273 1627 6307
rect 3065 6273 3099 6307
rect 3617 6273 3651 6307
rect 4261 6273 4295 6307
rect 5365 6273 5399 6307
rect 7205 6273 7239 6307
rect 8309 6273 8343 6307
rect 9413 6273 9447 6307
rect 10517 6273 10551 6307
rect 11989 6273 12023 6307
rect 13461 6273 13495 6307
rect 14565 6273 14599 6307
rect 15669 6273 15703 6307
rect 16865 6273 16899 6307
rect 17969 6273 18003 6307
rect 19073 6273 19107 6307
rect 20177 6273 20211 6307
rect 21465 6273 21499 6307
rect 22201 6273 22235 6307
rect 22477 6273 22511 6307
rect 22845 6273 22879 6307
rect 1869 6205 1903 6239
rect 6009 6205 6043 6239
rect 6561 6205 6595 6239
rect 18613 6205 18647 6239
rect 2881 6137 2915 6171
rect 13093 6137 13127 6171
rect 3709 6069 3743 6103
rect 6469 6069 6503 6103
rect 11161 6069 11195 6103
rect 11713 6069 11747 6103
rect 12909 6069 12943 6103
rect 14105 6069 14139 6103
rect 22017 6069 22051 6103
rect 23121 6069 23155 6103
rect 23305 6069 23339 6103
rect 2789 5865 2823 5899
rect 5457 5865 5491 5899
rect 7481 5865 7515 5899
rect 10425 5865 10459 5899
rect 11529 5865 11563 5899
rect 12633 5865 12667 5899
rect 13737 5865 13771 5899
rect 19349 5865 19383 5899
rect 20729 5865 20763 5899
rect 3433 5797 3467 5831
rect 18889 5797 18923 5831
rect 21189 5797 21223 5831
rect 1869 5729 1903 5763
rect 4905 5729 4939 5763
rect 6377 5729 6411 5763
rect 9137 5729 9171 5763
rect 15301 5729 15335 5763
rect 17141 5729 17175 5763
rect 17417 5729 17451 5763
rect 19441 5729 19475 5763
rect 19717 5729 19751 5763
rect 21649 5729 21683 5763
rect 23305 5729 23339 5763
rect 23857 5729 23891 5763
rect 1593 5661 1627 5695
rect 3249 5661 3283 5695
rect 4261 5661 4295 5695
rect 5733 5661 5767 5695
rect 6837 5661 6871 5695
rect 7941 5661 7975 5695
rect 9781 5661 9815 5695
rect 10885 5661 10919 5695
rect 11989 5661 12023 5695
rect 13093 5661 13127 5695
rect 14289 5661 14323 5695
rect 20913 5661 20947 5695
rect 21373 5661 21407 5695
rect 22712 5661 22746 5695
rect 3893 5593 3927 5627
rect 14473 5593 14507 5627
rect 22799 5593 22833 5627
rect 5181 5525 5215 5559
rect 8585 5525 8619 5559
rect 16497 5525 16531 5559
rect 3893 5321 3927 5355
rect 4169 5321 4203 5355
rect 6561 5321 6595 5355
rect 7849 5321 7883 5355
rect 8953 5321 8987 5355
rect 11621 5321 11655 5355
rect 12817 5321 12851 5355
rect 15209 5321 15243 5355
rect 17509 5321 17543 5355
rect 21557 5321 21591 5355
rect 5273 5253 5307 5287
rect 5825 5253 5859 5287
rect 14013 5253 14047 5287
rect 22753 5253 22787 5287
rect 22845 5253 22879 5287
rect 24961 5253 24995 5287
rect 26617 5253 26651 5287
rect 31309 5253 31343 5287
rect 1685 5185 1719 5219
rect 4629 5185 4663 5219
rect 7205 5185 7239 5219
rect 8309 5185 8343 5219
rect 9413 5185 9447 5219
rect 10517 5185 10551 5219
rect 11161 5185 11195 5219
rect 12173 5185 12207 5219
rect 13369 5185 13403 5219
rect 14565 5185 14599 5219
rect 15669 5185 15703 5219
rect 16865 5185 16899 5219
rect 18705 5185 18739 5219
rect 19993 5185 20027 5219
rect 21097 5185 21131 5219
rect 21833 5185 21867 5219
rect 22236 5184 22270 5218
rect 2789 5117 2823 5151
rect 3065 5117 3099 5151
rect 11713 5117 11747 5151
rect 18061 5117 18095 5151
rect 18429 5117 18463 5151
rect 19717 5117 19751 5151
rect 24777 5117 24811 5151
rect 27169 5117 27203 5151
rect 27353 5117 27387 5151
rect 28917 5117 28951 5151
rect 29469 5117 29503 5151
rect 29653 5117 29687 5151
rect 6009 5049 6043 5083
rect 2329 4981 2363 5015
rect 4353 4981 4387 5015
rect 10057 4981 10091 5015
rect 16313 4981 16347 5015
rect 21189 4981 21223 5015
rect 22339 4981 22373 5015
rect 3433 4777 3467 4811
rect 4629 4777 4663 4811
rect 5273 4777 5307 4811
rect 6561 4777 6595 4811
rect 7481 4777 7515 4811
rect 8585 4777 8619 4811
rect 9965 4777 9999 4811
rect 11805 4777 11839 4811
rect 12081 4777 12115 4811
rect 13093 4777 13127 4811
rect 14933 4777 14967 4811
rect 18613 4777 18647 4811
rect 18981 4777 19015 4811
rect 21005 4777 21039 4811
rect 22477 4777 22511 4811
rect 23075 4777 23109 4811
rect 10241 4709 10275 4743
rect 24731 4709 24765 4743
rect 1869 4641 1903 4675
rect 10701 4641 10735 4675
rect 10977 4641 11011 4675
rect 15669 4641 15703 4675
rect 19441 4641 19475 4675
rect 19717 4641 19751 4675
rect 21925 4641 21959 4675
rect 25881 4641 25915 4675
rect 27077 4641 27111 4675
rect 1593 4573 1627 4607
rect 2973 4573 3007 4607
rect 3157 4573 3191 4607
rect 3985 4573 4019 4607
rect 5181 4573 5215 4607
rect 6837 4573 6871 4607
rect 7941 4573 7975 4607
rect 9321 4573 9355 4607
rect 12449 4573 12483 4607
rect 14289 4573 14323 4607
rect 17969 4573 18003 4607
rect 20913 4573 20947 4607
rect 22972 4573 23006 4607
rect 24628 4573 24662 4607
rect 25697 4573 25731 4607
rect 5917 4505 5951 4539
rect 6101 4505 6135 4539
rect 15853 4505 15887 4539
rect 17509 4505 17543 4539
rect 8953 4437 8987 4471
rect 13461 4437 13495 4471
rect 13553 4437 13587 4471
rect 20545 4437 20579 4471
rect 21373 4437 21407 4471
rect 5825 4233 5859 4267
rect 14197 4233 14231 4267
rect 19165 4233 19199 4267
rect 20453 4233 20487 4267
rect 21097 4233 21131 4267
rect 5181 4165 5215 4199
rect 7573 4165 7607 4199
rect 7665 4165 7699 4199
rect 10977 4165 11011 4199
rect 12357 4165 12391 4199
rect 1593 4097 1627 4131
rect 2881 4097 2915 4131
rect 3985 4097 4019 4131
rect 4629 4097 4663 4131
rect 5365 4097 5399 4131
rect 6009 4097 6043 4131
rect 6561 4097 6595 4131
rect 7205 4097 7239 4131
rect 8401 4097 8435 4131
rect 8861 4097 8895 4131
rect 9597 4097 9631 4131
rect 11713 4097 11747 4131
rect 13093 4097 13127 4131
rect 13553 4097 13587 4131
rect 14657 4097 14691 4131
rect 16129 4097 16163 4131
rect 19441 4097 19475 4131
rect 20637 4097 20671 4131
rect 21557 4097 21591 4131
rect 1869 4029 1903 4063
rect 9321 4029 9355 4063
rect 10517 4029 10551 4063
rect 11161 4029 11195 4063
rect 16865 4029 16899 4063
rect 17049 4029 17083 4063
rect 18705 4029 18739 4063
rect 21833 4029 21867 4063
rect 3525 3893 3559 3927
rect 8493 3893 8527 3927
rect 9137 3893 9171 3927
rect 10241 3893 10275 3927
rect 12909 3893 12943 3927
rect 15301 3893 15335 3927
rect 15669 3893 15703 3927
rect 16221 3893 16255 3927
rect 19533 3893 19567 3927
rect 19901 3893 19935 3927
rect 2329 3689 2363 3723
rect 5273 3689 5307 3723
rect 9045 3689 9079 3723
rect 11253 3689 11287 3723
rect 13001 3689 13035 3723
rect 7021 3621 7055 3655
rect 11713 3621 11747 3655
rect 14565 3621 14599 3655
rect 15301 3621 15335 3655
rect 15761 3621 15795 3655
rect 15945 3621 15979 3655
rect 3985 3553 4019 3587
rect 5733 3553 5767 3587
rect 9137 3553 9171 3587
rect 20729 3553 20763 3587
rect 1685 3485 1719 3519
rect 2789 3485 2823 3519
rect 4629 3485 4663 3519
rect 6009 3485 6043 3519
rect 7205 3485 7239 3519
rect 8401 3485 8435 3519
rect 9505 3485 9539 3519
rect 10149 3485 10183 3519
rect 10609 3485 10643 3519
rect 11897 3485 11931 3519
rect 12357 3485 12391 3519
rect 16313 3485 16347 3519
rect 16589 3485 16623 3519
rect 17601 3485 17635 3519
rect 17877 3485 17911 3519
rect 19625 3485 19659 3519
rect 20269 3485 20303 3519
rect 8585 3417 8619 3451
rect 13553 3417 13587 3451
rect 14381 3417 14415 3451
rect 15117 3417 15151 3451
rect 15669 3417 15703 3451
rect 19073 3417 19107 3451
rect 3433 3349 3467 3383
rect 7665 3349 7699 3383
rect 18797 3349 18831 3383
rect 19441 3349 19475 3383
rect 20085 3349 20119 3383
rect 2881 3145 2915 3179
rect 10609 3145 10643 3179
rect 18061 3145 18095 3179
rect 20821 3145 20855 3179
rect 5825 3077 5859 3111
rect 14841 3077 14875 3111
rect 15025 3077 15059 3111
rect 15853 3077 15887 3111
rect 18705 3077 18739 3111
rect 20361 3077 20395 3111
rect 3065 3009 3099 3043
rect 3525 3009 3559 3043
rect 4629 3009 4663 3043
rect 5273 3009 5307 3043
rect 6561 3009 6595 3043
rect 7205 3009 7239 3043
rect 7757 3009 7791 3043
rect 8861 3009 8895 3043
rect 10885 3009 10919 3043
rect 11345 3009 11379 3043
rect 11805 3009 11839 3043
rect 12541 3009 12575 3043
rect 13093 3009 13127 3043
rect 13553 3009 13587 3043
rect 14105 3009 14139 3043
rect 17233 3009 17267 3043
rect 18521 3009 18555 3043
rect 22201 3009 22235 3043
rect 22477 3009 22511 3043
rect 1593 2941 1627 2975
rect 1869 2941 1903 2975
rect 8401 2941 8435 2975
rect 9137 2941 9171 2975
rect 16957 2941 16991 2975
rect 16405 2873 16439 2907
rect 4169 2805 4203 2839
rect 11897 2805 11931 2839
rect 12633 2805 12667 2839
rect 13369 2805 13403 2839
rect 14197 2805 14231 2839
rect 15393 2805 15427 2839
rect 15945 2805 15979 2839
rect 22017 2805 22051 2839
rect 2881 2601 2915 2635
rect 6377 2601 6411 2635
rect 9137 2601 9171 2635
rect 13829 2601 13863 2635
rect 14933 2601 14967 2635
rect 16957 2601 16991 2635
rect 17601 2601 17635 2635
rect 20085 2601 20119 2635
rect 22017 2601 22051 2635
rect 22569 2601 22603 2635
rect 25513 2601 25547 2635
rect 28181 2601 28215 2635
rect 30849 2601 30883 2635
rect 33517 2601 33551 2635
rect 3801 2533 3835 2567
rect 8677 2533 8711 2567
rect 18245 2533 18279 2567
rect 19441 2533 19475 2567
rect 1869 2465 1903 2499
rect 3249 2465 3283 2499
rect 4629 2465 4663 2499
rect 5825 2465 5859 2499
rect 6101 2465 6135 2499
rect 7297 2465 7331 2499
rect 9965 2465 9999 2499
rect 12633 2465 12667 2499
rect 36369 2465 36403 2499
rect 1593 2397 1627 2431
rect 4353 2397 4387 2431
rect 7021 2397 7055 2431
rect 9597 2397 9631 2431
rect 12357 2397 12391 2431
rect 15485 2397 15519 2431
rect 15761 2397 15795 2431
rect 17141 2397 17175 2431
rect 17785 2397 17819 2431
rect 18429 2397 18463 2431
rect 19625 2397 19659 2431
rect 20269 2397 20303 2431
rect 22201 2397 22235 2431
rect 25697 2397 25731 2431
rect 25973 2397 26007 2431
rect 28365 2397 28399 2431
rect 28641 2397 28675 2431
rect 31033 2397 31067 2431
rect 31309 2397 31343 2431
rect 33701 2397 33735 2431
rect 33977 2397 34011 2431
rect 36093 2397 36127 2431
rect 37289 2397 37323 2431
rect 14841 2329 14875 2363
rect 20729 2329 20763 2363
rect 2789 2261 2823 2295
rect 8493 2261 8527 2295
rect 9045 2261 9079 2295
rect 11161 2261 11195 2295
rect 11529 2261 11563 2295
rect 14197 2261 14231 2295
rect 14381 2261 14415 2295
rect 18797 2261 18831 2295
rect 18981 2261 19015 2295
<< metal1 >>
rect 7742 26936 7748 26988
rect 7800 26976 7806 26988
rect 21726 26976 21732 26988
rect 7800 26948 21732 26976
rect 7800 26936 7806 26948
rect 21726 26936 21732 26948
rect 21784 26936 21790 26988
rect 10226 26868 10232 26920
rect 10284 26908 10290 26920
rect 19702 26908 19708 26920
rect 10284 26880 19708 26908
rect 10284 26868 10290 26880
rect 19702 26868 19708 26880
rect 19760 26868 19766 26920
rect 22922 26840 22928 26852
rect 17236 26812 22928 26840
rect 9490 26596 9496 26648
rect 9548 26636 9554 26648
rect 17236 26636 17264 26812
rect 22922 26800 22928 26812
rect 22980 26800 22986 26852
rect 23382 26800 23388 26852
rect 23440 26840 23446 26852
rect 33686 26840 33692 26852
rect 23440 26812 33692 26840
rect 23440 26800 23446 26812
rect 33686 26800 33692 26812
rect 33744 26800 33750 26852
rect 29822 26772 29828 26784
rect 9548 26608 17264 26636
rect 17328 26744 29828 26772
rect 9548 26596 9554 26608
rect 16850 26528 16856 26580
rect 16908 26568 16914 26580
rect 17328 26568 17356 26744
rect 29822 26732 29828 26744
rect 29880 26732 29886 26784
rect 36538 26704 36544 26716
rect 22066 26676 36544 26704
rect 20530 26596 20536 26648
rect 20588 26636 20594 26648
rect 22066 26636 22094 26676
rect 36538 26664 36544 26676
rect 36596 26664 36602 26716
rect 20588 26608 22094 26636
rect 20588 26596 20594 26608
rect 25958 26596 25964 26648
rect 26016 26636 26022 26648
rect 34606 26636 34612 26648
rect 26016 26608 34612 26636
rect 26016 26596 26022 26608
rect 34606 26596 34612 26608
rect 34664 26596 34670 26648
rect 16908 26540 17356 26568
rect 16908 26528 16914 26540
rect 17770 26528 17776 26580
rect 17828 26568 17834 26580
rect 42886 26568 42892 26580
rect 17828 26540 42892 26568
rect 17828 26528 17834 26540
rect 42886 26528 42892 26540
rect 42944 26528 42950 26580
rect 17218 26460 17224 26512
rect 17276 26500 17282 26512
rect 41598 26500 41604 26512
rect 17276 26472 41604 26500
rect 17276 26460 17282 26472
rect 41598 26460 41604 26472
rect 41656 26460 41662 26512
rect 18874 26432 18880 26444
rect 2746 26404 18880 26432
rect 1302 26324 1308 26376
rect 1360 26364 1366 26376
rect 2746 26364 2774 26404
rect 18874 26392 18880 26404
rect 18932 26392 18938 26444
rect 19058 26392 19064 26444
rect 19116 26432 19122 26444
rect 40954 26432 40960 26444
rect 19116 26404 40960 26432
rect 19116 26392 19122 26404
rect 40954 26392 40960 26404
rect 41012 26392 41018 26444
rect 1360 26336 2774 26364
rect 1360 26324 1366 26336
rect 14734 26324 14740 26376
rect 14792 26364 14798 26376
rect 14792 26336 24164 26364
rect 14792 26324 14798 26336
rect 566 26256 572 26308
rect 624 26296 630 26308
rect 22094 26296 22100 26308
rect 624 26268 22100 26296
rect 624 26256 630 26268
rect 22094 26256 22100 26268
rect 22152 26256 22158 26308
rect 5258 26188 5264 26240
rect 5316 26228 5322 26240
rect 20070 26228 20076 26240
rect 5316 26200 20076 26228
rect 5316 26188 5322 26200
rect 20070 26188 20076 26200
rect 20128 26188 20134 26240
rect 22370 26188 22376 26240
rect 22428 26228 22434 26240
rect 23382 26228 23388 26240
rect 22428 26200 23388 26228
rect 22428 26188 22434 26200
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 14182 26120 14188 26172
rect 14240 26160 14246 26172
rect 19058 26160 19064 26172
rect 14240 26132 19064 26160
rect 14240 26120 14246 26132
rect 19058 26120 19064 26132
rect 19116 26120 19122 26172
rect 24136 26160 24164 26336
rect 28258 26324 28264 26376
rect 28316 26364 28322 26376
rect 45922 26364 45928 26376
rect 28316 26336 45928 26364
rect 28316 26324 28322 26336
rect 45922 26324 45928 26336
rect 45980 26324 45986 26376
rect 26970 26256 26976 26308
rect 27028 26296 27034 26308
rect 36814 26296 36820 26308
rect 27028 26268 36820 26296
rect 27028 26256 27034 26268
rect 36814 26256 36820 26268
rect 36872 26256 36878 26308
rect 26878 26188 26884 26240
rect 26936 26228 26942 26240
rect 37274 26228 37280 26240
rect 26936 26200 37280 26228
rect 26936 26188 26942 26200
rect 37274 26188 37280 26200
rect 37332 26188 37338 26240
rect 33870 26160 33876 26172
rect 24136 26132 33876 26160
rect 33870 26120 33876 26132
rect 33928 26120 33934 26172
rect 17586 26052 17592 26104
rect 17644 26092 17650 26104
rect 39114 26092 39120 26104
rect 17644 26064 39120 26092
rect 17644 26052 17650 26064
rect 39114 26052 39120 26064
rect 39172 26052 39178 26104
rect 12618 25984 12624 26036
rect 12676 26024 12682 26036
rect 39758 26024 39764 26036
rect 12676 25996 39764 26024
rect 12676 25984 12682 25996
rect 39758 25984 39764 25996
rect 39816 25984 39822 26036
rect 8938 25916 8944 25968
rect 8996 25956 9002 25968
rect 34698 25956 34704 25968
rect 8996 25928 34704 25956
rect 8996 25916 9002 25928
rect 34698 25916 34704 25928
rect 34756 25916 34762 25968
rect 7558 25848 7564 25900
rect 7616 25888 7622 25900
rect 17862 25888 17868 25900
rect 7616 25860 17868 25888
rect 7616 25848 7622 25860
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 21266 25848 21272 25900
rect 21324 25888 21330 25900
rect 41874 25888 41880 25900
rect 21324 25860 41880 25888
rect 21324 25848 21330 25860
rect 41874 25848 41880 25860
rect 41932 25848 41938 25900
rect 6638 25780 6644 25832
rect 6696 25820 6702 25832
rect 36998 25820 37004 25832
rect 6696 25792 37004 25820
rect 6696 25780 6702 25792
rect 36998 25780 37004 25792
rect 37056 25780 37062 25832
rect 3878 25712 3884 25764
rect 3936 25752 3942 25764
rect 41138 25752 41144 25764
rect 3936 25724 41144 25752
rect 3936 25712 3942 25724
rect 41138 25712 41144 25724
rect 41196 25712 41202 25764
rect 8294 25644 8300 25696
rect 8352 25684 8358 25696
rect 22094 25684 22100 25696
rect 8352 25656 22100 25684
rect 8352 25644 8358 25656
rect 22094 25644 22100 25656
rect 22152 25644 22158 25696
rect 22278 25644 22284 25696
rect 22336 25684 22342 25696
rect 29546 25684 29552 25696
rect 22336 25656 29552 25684
rect 22336 25644 22342 25656
rect 29546 25644 29552 25656
rect 29604 25644 29610 25696
rect 2038 25576 2044 25628
rect 2096 25616 2102 25628
rect 16206 25616 16212 25628
rect 2096 25588 16212 25616
rect 2096 25576 2102 25588
rect 16206 25576 16212 25588
rect 16264 25576 16270 25628
rect 17034 25576 17040 25628
rect 17092 25616 17098 25628
rect 31938 25616 31944 25628
rect 17092 25588 31944 25616
rect 17092 25576 17098 25588
rect 31938 25576 31944 25588
rect 31996 25576 32002 25628
rect 2130 25508 2136 25560
rect 2188 25548 2194 25560
rect 14550 25548 14556 25560
rect 2188 25520 14556 25548
rect 2188 25508 2194 25520
rect 14550 25508 14556 25520
rect 14608 25508 14614 25560
rect 14826 25508 14832 25560
rect 14884 25548 14890 25560
rect 33778 25548 33784 25560
rect 14884 25520 33784 25548
rect 14884 25508 14890 25520
rect 33778 25508 33784 25520
rect 33836 25508 33842 25560
rect 9214 25440 9220 25492
rect 9272 25480 9278 25492
rect 20806 25480 20812 25492
rect 9272 25452 20812 25480
rect 9272 25440 9278 25452
rect 20806 25440 20812 25452
rect 20864 25440 20870 25492
rect 21082 25440 21088 25492
rect 21140 25480 21146 25492
rect 40310 25480 40316 25492
rect 21140 25452 40316 25480
rect 21140 25440 21146 25452
rect 40310 25440 40316 25452
rect 40368 25440 40374 25492
rect 17494 25372 17500 25424
rect 17552 25412 17558 25424
rect 40402 25412 40408 25424
rect 17552 25384 40408 25412
rect 17552 25372 17558 25384
rect 40402 25372 40408 25384
rect 40460 25372 40466 25424
rect 15010 25304 15016 25356
rect 15068 25344 15074 25356
rect 15068 25316 17172 25344
rect 15068 25304 15074 25316
rect 7098 25236 7104 25288
rect 7156 25276 7162 25288
rect 16942 25276 16948 25288
rect 7156 25248 16948 25276
rect 7156 25236 7162 25248
rect 16942 25236 16948 25248
rect 17000 25236 17006 25288
rect 17144 25276 17172 25316
rect 18690 25304 18696 25356
rect 18748 25344 18754 25356
rect 43622 25344 43628 25356
rect 18748 25316 43628 25344
rect 18748 25304 18754 25316
rect 43622 25304 43628 25316
rect 43680 25304 43686 25356
rect 17144 25248 22048 25276
rect 1854 25168 1860 25220
rect 1912 25208 1918 25220
rect 1912 25180 16528 25208
rect 1912 25168 1918 25180
rect 6730 25100 6736 25152
rect 6788 25140 6794 25152
rect 16390 25140 16396 25152
rect 6788 25112 16396 25140
rect 6788 25100 6794 25112
rect 16390 25100 16396 25112
rect 16448 25100 16454 25152
rect 16500 25140 16528 25180
rect 17512 25180 17954 25208
rect 17512 25140 17540 25180
rect 16500 25112 17540 25140
rect 17926 25140 17954 25180
rect 20806 25168 20812 25220
rect 20864 25208 20870 25220
rect 21910 25208 21916 25220
rect 20864 25180 21916 25208
rect 20864 25168 20870 25180
rect 21910 25168 21916 25180
rect 21968 25168 21974 25220
rect 22020 25208 22048 25248
rect 22094 25236 22100 25288
rect 22152 25276 22158 25288
rect 22554 25276 22560 25288
rect 22152 25248 22560 25276
rect 22152 25236 22158 25248
rect 22554 25236 22560 25248
rect 22612 25236 22618 25288
rect 22646 25236 22652 25288
rect 22704 25276 22710 25288
rect 22704 25248 27200 25276
rect 22704 25236 22710 25248
rect 23934 25208 23940 25220
rect 22020 25180 23940 25208
rect 23934 25168 23940 25180
rect 23992 25168 23998 25220
rect 27172 25208 27200 25248
rect 30374 25236 30380 25288
rect 30432 25276 30438 25288
rect 44358 25276 44364 25288
rect 30432 25248 44364 25276
rect 30432 25236 30438 25248
rect 44358 25236 44364 25248
rect 44416 25236 44422 25288
rect 36630 25208 36636 25220
rect 27172 25180 36636 25208
rect 36630 25168 36636 25180
rect 36688 25168 36694 25220
rect 19886 25140 19892 25152
rect 17926 25112 19892 25140
rect 19886 25100 19892 25112
rect 19944 25100 19950 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 36170 25140 36176 25152
rect 20036 25112 36176 25140
rect 20036 25100 20042 25112
rect 36170 25100 36176 25112
rect 36228 25100 36234 25152
rect 4062 25032 4068 25084
rect 4120 25072 4126 25084
rect 10042 25072 10048 25084
rect 4120 25044 10048 25072
rect 4120 25032 4126 25044
rect 10042 25032 10048 25044
rect 10100 25032 10106 25084
rect 12066 25032 12072 25084
rect 12124 25072 12130 25084
rect 12124 25044 16436 25072
rect 12124 25032 12130 25044
rect 4522 24964 4528 25016
rect 4580 25004 4586 25016
rect 15838 25004 15844 25016
rect 4580 24976 15844 25004
rect 4580 24964 4586 24976
rect 15838 24964 15844 24976
rect 15896 24964 15902 25016
rect 5718 24896 5724 24948
rect 5776 24936 5782 24948
rect 13722 24936 13728 24948
rect 5776 24908 13728 24936
rect 5776 24896 5782 24908
rect 13722 24896 13728 24908
rect 13780 24896 13786 24948
rect 16408 24936 16436 25044
rect 16942 25032 16948 25084
rect 17000 25072 17006 25084
rect 23382 25072 23388 25084
rect 17000 25044 23388 25072
rect 17000 25032 17006 25044
rect 23382 25032 23388 25044
rect 23440 25032 23446 25084
rect 24578 25032 24584 25084
rect 24636 25072 24642 25084
rect 26234 25072 26240 25084
rect 24636 25044 26240 25072
rect 24636 25032 24642 25044
rect 26234 25032 26240 25044
rect 26292 25032 26298 25084
rect 28718 25032 28724 25084
rect 28776 25072 28782 25084
rect 39206 25072 39212 25084
rect 28776 25044 39212 25072
rect 28776 25032 28782 25044
rect 39206 25032 39212 25044
rect 39264 25032 39270 25084
rect 16482 24964 16488 25016
rect 16540 25004 16546 25016
rect 16540 24976 22094 25004
rect 16540 24964 16546 24976
rect 18138 24936 18144 24948
rect 16408 24908 18144 24936
rect 18138 24896 18144 24908
rect 18196 24896 18202 24948
rect 20254 24896 20260 24948
rect 20312 24936 20318 24948
rect 20714 24936 20720 24948
rect 20312 24908 20720 24936
rect 20312 24896 20318 24908
rect 20714 24896 20720 24908
rect 20772 24896 20778 24948
rect 3326 24828 3332 24880
rect 3384 24868 3390 24880
rect 4890 24868 4896 24880
rect 3384 24840 4896 24868
rect 3384 24828 3390 24840
rect 4890 24828 4896 24840
rect 4948 24828 4954 24880
rect 8386 24828 8392 24880
rect 8444 24868 8450 24880
rect 11054 24868 11060 24880
rect 8444 24840 11060 24868
rect 8444 24828 8450 24840
rect 11054 24828 11060 24840
rect 11112 24828 11118 24880
rect 13630 24828 13636 24880
rect 13688 24868 13694 24880
rect 17954 24868 17960 24880
rect 13688 24840 17960 24868
rect 13688 24828 13694 24840
rect 17954 24828 17960 24840
rect 18012 24828 18018 24880
rect 18506 24828 18512 24880
rect 18564 24868 18570 24880
rect 20806 24868 20812 24880
rect 18564 24840 20812 24868
rect 18564 24828 18570 24840
rect 20806 24828 20812 24840
rect 20864 24828 20870 24880
rect 6546 24760 6552 24812
rect 6604 24800 6610 24812
rect 21358 24800 21364 24812
rect 6604 24772 21364 24800
rect 6604 24760 6610 24772
rect 21358 24760 21364 24772
rect 21416 24760 21422 24812
rect 22066 24800 22094 24976
rect 23474 24964 23480 25016
rect 23532 25004 23538 25016
rect 35802 25004 35808 25016
rect 23532 24976 35808 25004
rect 23532 24964 23538 24976
rect 35802 24964 35808 24976
rect 35860 24964 35866 25016
rect 22830 24896 22836 24948
rect 22888 24936 22894 24948
rect 26970 24936 26976 24948
rect 22888 24908 26976 24936
rect 22888 24896 22894 24908
rect 26970 24896 26976 24908
rect 27028 24896 27034 24948
rect 28810 24896 28816 24948
rect 28868 24936 28874 24948
rect 31110 24936 31116 24948
rect 28868 24908 31116 24936
rect 28868 24896 28874 24908
rect 31110 24896 31116 24908
rect 31168 24896 31174 24948
rect 32674 24896 32680 24948
rect 32732 24936 32738 24948
rect 42058 24936 42064 24948
rect 32732 24908 42064 24936
rect 32732 24896 32738 24908
rect 42058 24896 42064 24908
rect 42116 24896 42122 24948
rect 22554 24828 22560 24880
rect 22612 24868 22618 24880
rect 24578 24868 24584 24880
rect 22612 24840 24584 24868
rect 22612 24828 22618 24840
rect 24578 24828 24584 24840
rect 24636 24828 24642 24880
rect 24670 24828 24676 24880
rect 24728 24868 24734 24880
rect 29178 24868 29184 24880
rect 24728 24840 29184 24868
rect 24728 24828 24734 24840
rect 29178 24828 29184 24840
rect 29236 24828 29242 24880
rect 30650 24868 30656 24880
rect 29288 24840 30656 24868
rect 25958 24800 25964 24812
rect 22066 24772 25964 24800
rect 25958 24760 25964 24772
rect 26016 24760 26022 24812
rect 26234 24760 26240 24812
rect 26292 24800 26298 24812
rect 29288 24800 29316 24840
rect 30650 24828 30656 24840
rect 30708 24828 30714 24880
rect 26292 24772 29316 24800
rect 26292 24760 26298 24772
rect 13722 24692 13728 24744
rect 13780 24732 13786 24744
rect 16298 24732 16304 24744
rect 13780 24704 16304 24732
rect 13780 24692 13786 24704
rect 16298 24692 16304 24704
rect 16356 24692 16362 24744
rect 17862 24692 17868 24744
rect 17920 24732 17926 24744
rect 22554 24732 22560 24744
rect 17920 24704 22560 24732
rect 17920 24692 17926 24704
rect 22554 24692 22560 24704
rect 22612 24692 22618 24744
rect 22830 24692 22836 24744
rect 22888 24732 22894 24744
rect 28350 24732 28356 24744
rect 22888 24704 28356 24732
rect 22888 24692 22894 24704
rect 28350 24692 28356 24704
rect 28408 24692 28414 24744
rect 12342 24624 12348 24676
rect 12400 24664 12406 24676
rect 25774 24664 25780 24676
rect 12400 24636 25780 24664
rect 12400 24624 12406 24636
rect 25774 24624 25780 24636
rect 25832 24624 25838 24676
rect 26602 24624 26608 24676
rect 26660 24664 26666 24676
rect 29914 24664 29920 24676
rect 26660 24636 29920 24664
rect 26660 24624 26666 24636
rect 29914 24624 29920 24636
rect 29972 24624 29978 24676
rect 13998 24556 14004 24608
rect 14056 24596 14062 24608
rect 16850 24596 16856 24608
rect 14056 24568 16856 24596
rect 14056 24556 14062 24568
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 16942 24556 16948 24608
rect 17000 24596 17006 24608
rect 17126 24596 17132 24608
rect 17000 24568 17132 24596
rect 17000 24556 17006 24568
rect 17126 24556 17132 24568
rect 17184 24556 17190 24608
rect 17954 24556 17960 24608
rect 18012 24596 18018 24608
rect 19794 24596 19800 24608
rect 18012 24568 19800 24596
rect 18012 24556 18018 24568
rect 19794 24556 19800 24568
rect 19852 24556 19858 24608
rect 20346 24556 20352 24608
rect 20404 24596 20410 24608
rect 26050 24596 26056 24608
rect 20404 24568 26056 24596
rect 20404 24556 20410 24568
rect 26050 24556 26056 24568
rect 26108 24556 26114 24608
rect 29454 24556 29460 24608
rect 29512 24596 29518 24608
rect 37458 24596 37464 24608
rect 29512 24568 37464 24596
rect 29512 24556 29518 24568
rect 37458 24556 37464 24568
rect 37516 24556 37522 24608
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 842 24352 848 24404
rect 900 24392 906 24404
rect 900 24364 3924 24392
rect 900 24352 906 24364
rect 3237 24259 3295 24265
rect 3237 24225 3249 24259
rect 3283 24256 3295 24259
rect 3510 24256 3516 24268
rect 3283 24228 3516 24256
rect 3283 24225 3295 24228
rect 3237 24219 3295 24225
rect 3510 24216 3516 24228
rect 3568 24216 3574 24268
rect 3896 24256 3924 24364
rect 3970 24352 3976 24404
rect 4028 24392 4034 24404
rect 7466 24392 7472 24404
rect 4028 24364 7472 24392
rect 4028 24352 4034 24364
rect 7466 24352 7472 24364
rect 7524 24352 7530 24404
rect 11422 24392 11428 24404
rect 7576 24364 11428 24392
rect 7576 24324 7604 24364
rect 11422 24352 11428 24364
rect 11480 24352 11486 24404
rect 12406 24364 14872 24392
rect 5092 24296 7604 24324
rect 5092 24256 5120 24296
rect 9306 24284 9312 24336
rect 9364 24284 9370 24336
rect 3896 24228 5120 24256
rect 5813 24259 5871 24265
rect 5813 24225 5825 24259
rect 5859 24256 5871 24259
rect 7374 24256 7380 24268
rect 5859 24228 7380 24256
rect 5859 24225 5871 24228
rect 5813 24219 5871 24225
rect 7374 24216 7380 24228
rect 7432 24216 7438 24268
rect 8205 24259 8263 24265
rect 8205 24225 8217 24259
rect 8251 24256 8263 24259
rect 9324 24256 9352 24284
rect 11514 24256 11520 24268
rect 8251 24228 9352 24256
rect 9692 24228 11520 24256
rect 8251 24225 8263 24228
rect 8205 24219 8263 24225
rect 2222 24148 2228 24200
rect 2280 24148 2286 24200
rect 4157 24191 4215 24197
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4706 24188 4712 24200
rect 4203 24160 4712 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4706 24148 4712 24160
rect 4764 24148 4770 24200
rect 4798 24148 4804 24200
rect 4856 24148 4862 24200
rect 6546 24148 6552 24200
rect 6604 24148 6610 24200
rect 7285 24191 7343 24197
rect 7285 24157 7297 24191
rect 7331 24157 7343 24191
rect 7285 24151 7343 24157
rect 9033 24191 9091 24197
rect 9033 24157 9045 24191
rect 9079 24188 9091 24191
rect 9309 24191 9367 24197
rect 9309 24188 9321 24191
rect 9079 24160 9321 24188
rect 9079 24157 9091 24160
rect 9033 24151 9091 24157
rect 9309 24157 9321 24160
rect 9355 24188 9367 24191
rect 9692 24188 9720 24228
rect 11514 24216 11520 24228
rect 11572 24216 11578 24268
rect 9355 24160 9720 24188
rect 9355 24157 9367 24160
rect 9309 24151 9367 24157
rect 1581 24123 1639 24129
rect 1581 24089 1593 24123
rect 1627 24120 1639 24123
rect 7300 24120 7328 24151
rect 9766 24148 9772 24200
rect 9824 24148 9830 24200
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24188 11667 24191
rect 11885 24191 11943 24197
rect 11885 24188 11897 24191
rect 11655 24160 11897 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 11885 24157 11897 24160
rect 11931 24188 11943 24191
rect 12406 24188 12434 24364
rect 14458 24324 14464 24336
rect 13556 24296 14464 24324
rect 13556 24265 13584 24296
rect 14458 24284 14464 24296
rect 14516 24284 14522 24336
rect 14844 24324 14872 24364
rect 16666 24352 16672 24404
rect 16724 24392 16730 24404
rect 24762 24392 24768 24404
rect 16724 24364 24768 24392
rect 16724 24352 16730 24364
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 25774 24352 25780 24404
rect 25832 24352 25838 24404
rect 25958 24392 25964 24404
rect 25884 24364 25964 24392
rect 16850 24324 16856 24336
rect 14844 24296 16856 24324
rect 16850 24284 16856 24296
rect 16908 24284 16914 24336
rect 18138 24284 18144 24336
rect 18196 24324 18202 24336
rect 21450 24324 21456 24336
rect 18196 24296 21456 24324
rect 18196 24284 18202 24296
rect 21450 24284 21456 24296
rect 21508 24284 21514 24336
rect 24854 24284 24860 24336
rect 24912 24324 24918 24336
rect 25884 24324 25912 24364
rect 25958 24352 25964 24364
rect 26016 24392 26022 24404
rect 26016 24364 38608 24392
rect 26016 24352 26022 24364
rect 24912 24296 25912 24324
rect 25976 24296 27108 24324
rect 24912 24284 24918 24296
rect 13541 24259 13599 24265
rect 13541 24225 13553 24259
rect 13587 24225 13599 24259
rect 13541 24219 13599 24225
rect 14366 24216 14372 24268
rect 14424 24256 14430 24268
rect 16117 24259 16175 24265
rect 14424 24228 14964 24256
rect 14424 24216 14430 24228
rect 11931 24160 12434 24188
rect 11931 24157 11943 24160
rect 11885 24151 11943 24157
rect 12526 24148 12532 24200
rect 12584 24148 12590 24200
rect 14458 24148 14464 24200
rect 14516 24188 14522 24200
rect 14936 24197 14964 24228
rect 16117 24225 16129 24259
rect 16163 24256 16175 24259
rect 18966 24256 18972 24268
rect 16163 24228 18972 24256
rect 16163 24225 16175 24228
rect 16117 24219 16175 24225
rect 18966 24216 18972 24228
rect 19024 24216 19030 24268
rect 20622 24256 20628 24268
rect 19720 24228 20628 24256
rect 14921 24191 14979 24197
rect 14516 24160 14872 24188
rect 14516 24148 14522 24160
rect 10134 24120 10140 24132
rect 1627 24092 5120 24120
rect 7300 24092 10140 24120
rect 1627 24089 1639 24092
rect 1581 24083 1639 24089
rect 1762 24012 1768 24064
rect 1820 24012 1826 24064
rect 3510 24012 3516 24064
rect 3568 24052 3574 24064
rect 3973 24055 4031 24061
rect 3973 24052 3985 24055
rect 3568 24024 3985 24052
rect 3568 24012 3574 24024
rect 3973 24021 3985 24024
rect 4019 24021 4031 24055
rect 5092 24052 5120 24092
rect 10134 24080 10140 24092
rect 10192 24080 10198 24132
rect 10965 24123 11023 24129
rect 10965 24089 10977 24123
rect 11011 24120 11023 24123
rect 13814 24120 13820 24132
rect 11011 24092 13820 24120
rect 11011 24089 11023 24092
rect 10965 24083 11023 24089
rect 13814 24080 13820 24092
rect 13872 24080 13878 24132
rect 7374 24052 7380 24064
rect 5092 24024 7380 24052
rect 3973 24015 4031 24021
rect 7374 24012 7380 24024
rect 7432 24012 7438 24064
rect 9122 24012 9128 24064
rect 9180 24012 9186 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 11790 24012 11796 24064
rect 11848 24052 11854 24064
rect 12434 24052 12440 24064
rect 11848 24024 12440 24052
rect 11848 24012 11854 24024
rect 12434 24012 12440 24024
rect 12492 24012 12498 24064
rect 12526 24012 12532 24064
rect 12584 24052 12590 24064
rect 14182 24052 14188 24064
rect 12584 24024 14188 24052
rect 12584 24012 12590 24024
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 14274 24012 14280 24064
rect 14332 24012 14338 24064
rect 14844 24052 14872 24160
rect 14921 24157 14933 24191
rect 14967 24157 14979 24191
rect 14921 24151 14979 24157
rect 16850 24148 16856 24200
rect 16908 24148 16914 24200
rect 19610 24148 19616 24200
rect 19668 24148 19674 24200
rect 16758 24080 16764 24132
rect 16816 24120 16822 24132
rect 17129 24123 17187 24129
rect 17129 24120 17141 24123
rect 16816 24092 17141 24120
rect 16816 24080 16822 24092
rect 17129 24089 17141 24092
rect 17175 24089 17187 24123
rect 18414 24120 18420 24132
rect 18354 24092 18420 24120
rect 17129 24083 17187 24089
rect 18414 24080 18420 24092
rect 18472 24120 18478 24132
rect 19518 24120 19524 24132
rect 18472 24092 19524 24120
rect 18472 24080 18478 24092
rect 19518 24080 19524 24092
rect 19576 24120 19582 24132
rect 19720 24120 19748 24228
rect 20622 24216 20628 24228
rect 20680 24216 20686 24268
rect 20898 24216 20904 24268
rect 20956 24216 20962 24268
rect 21542 24216 21548 24268
rect 21600 24256 21606 24268
rect 22465 24259 22523 24265
rect 22465 24256 22477 24259
rect 21600 24228 22477 24256
rect 21600 24216 21606 24228
rect 22465 24225 22477 24228
rect 22511 24225 22523 24259
rect 22465 24219 22523 24225
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 25130 24256 25136 24268
rect 22612 24228 25136 24256
rect 22612 24216 22618 24228
rect 25130 24216 25136 24228
rect 25188 24216 25194 24268
rect 25225 24259 25283 24265
rect 25225 24225 25237 24259
rect 25271 24256 25283 24259
rect 25976 24256 26004 24296
rect 25271 24228 26004 24256
rect 25271 24225 25283 24228
rect 25225 24219 25283 24225
rect 26050 24216 26056 24268
rect 26108 24256 26114 24268
rect 26329 24259 26387 24265
rect 26329 24256 26341 24259
rect 26108 24228 26341 24256
rect 26108 24216 26114 24228
rect 26329 24225 26341 24228
rect 26375 24225 26387 24259
rect 26329 24219 26387 24225
rect 26418 24216 26424 24268
rect 26476 24216 26482 24268
rect 27080 24256 27108 24296
rect 27154 24284 27160 24336
rect 27212 24284 27218 24336
rect 29086 24324 29092 24336
rect 27632 24296 29092 24324
rect 27632 24256 27660 24296
rect 29086 24284 29092 24296
rect 29144 24324 29150 24336
rect 29144 24296 29868 24324
rect 29144 24284 29150 24296
rect 27080 24228 27660 24256
rect 27706 24216 27712 24268
rect 27764 24216 27770 24268
rect 27798 24216 27804 24268
rect 27856 24256 27862 24268
rect 28997 24259 29055 24265
rect 27856 24228 28488 24256
rect 27856 24216 27862 24228
rect 20070 24148 20076 24200
rect 20128 24148 20134 24200
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 22189 24191 22247 24197
rect 20220 24160 22140 24188
rect 20220 24148 20226 24160
rect 19576 24092 19748 24120
rect 22112 24120 22140 24160
rect 22189 24157 22201 24191
rect 22235 24188 22247 24191
rect 22278 24188 22284 24200
rect 22235 24160 22284 24188
rect 22235 24157 22247 24160
rect 22189 24151 22247 24157
rect 22278 24148 22284 24160
rect 22336 24148 22342 24200
rect 24762 24188 24768 24200
rect 23768 24160 24768 24188
rect 23768 24120 23796 24160
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 25041 24191 25099 24197
rect 25041 24157 25053 24191
rect 25087 24157 25099 24191
rect 26436 24188 26464 24216
rect 27617 24191 27675 24197
rect 27617 24188 27629 24191
rect 26436 24160 27629 24188
rect 25041 24151 25099 24157
rect 27617 24157 27629 24160
rect 27663 24157 27675 24191
rect 27617 24151 27675 24157
rect 22112 24092 23796 24120
rect 23845 24123 23903 24129
rect 19576 24080 19582 24092
rect 23845 24089 23857 24123
rect 23891 24120 23903 24123
rect 24949 24123 25007 24129
rect 24949 24120 24961 24123
rect 23891 24092 24961 24120
rect 23891 24089 23903 24092
rect 23845 24083 23903 24089
rect 24949 24089 24961 24092
rect 24995 24089 25007 24123
rect 25056 24120 25084 24151
rect 28350 24148 28356 24200
rect 28408 24148 28414 24200
rect 28460 24188 28488 24228
rect 28997 24225 29009 24259
rect 29043 24256 29055 24259
rect 29178 24256 29184 24268
rect 29043 24228 29184 24256
rect 29043 24225 29055 24228
rect 28997 24219 29055 24225
rect 29178 24216 29184 24228
rect 29236 24216 29242 24268
rect 29270 24216 29276 24268
rect 29328 24256 29334 24268
rect 29730 24256 29736 24268
rect 29328 24228 29736 24256
rect 29328 24216 29334 24228
rect 29730 24216 29736 24228
rect 29788 24216 29794 24268
rect 29840 24256 29868 24296
rect 29914 24284 29920 24336
rect 29972 24324 29978 24336
rect 29972 24296 34928 24324
rect 29972 24284 29978 24296
rect 32214 24256 32220 24268
rect 29840 24228 32220 24256
rect 32214 24216 32220 24228
rect 32272 24216 32278 24268
rect 32324 24228 34192 24256
rect 30009 24191 30067 24197
rect 30009 24188 30021 24191
rect 28460 24160 30021 24188
rect 30009 24157 30021 24160
rect 30055 24157 30067 24191
rect 30009 24151 30067 24157
rect 31018 24148 31024 24200
rect 31076 24148 31082 24200
rect 32324 24197 32352 24228
rect 32309 24191 32367 24197
rect 32309 24157 32321 24191
rect 32355 24157 32367 24191
rect 32309 24151 32367 24157
rect 32953 24191 33011 24197
rect 32953 24157 32965 24191
rect 32999 24188 33011 24191
rect 33413 24191 33471 24197
rect 33413 24188 33425 24191
rect 32999 24160 33425 24188
rect 32999 24157 33011 24160
rect 32953 24151 33011 24157
rect 33413 24157 33425 24160
rect 33459 24157 33471 24191
rect 33413 24151 33471 24157
rect 27246 24120 27252 24132
rect 25056 24092 27252 24120
rect 24949 24083 25007 24089
rect 27246 24080 27252 24092
rect 27304 24080 27310 24132
rect 27430 24080 27436 24132
rect 27488 24120 27494 24132
rect 34057 24123 34115 24129
rect 34057 24120 34069 24123
rect 27488 24092 34069 24120
rect 27488 24080 27494 24092
rect 34057 24089 34069 24092
rect 34103 24089 34115 24123
rect 34164 24120 34192 24228
rect 34330 24148 34336 24200
rect 34388 24148 34394 24200
rect 34900 24197 34928 24296
rect 36630 24284 36636 24336
rect 36688 24284 36694 24336
rect 36998 24284 37004 24336
rect 37056 24324 37062 24336
rect 37056 24296 38516 24324
rect 37056 24284 37062 24296
rect 34885 24191 34943 24197
rect 34885 24157 34897 24191
rect 34931 24157 34943 24191
rect 34885 24151 34943 24157
rect 35989 24191 36047 24197
rect 35989 24157 36001 24191
rect 36035 24188 36047 24191
rect 37366 24188 37372 24200
rect 36035 24160 37372 24188
rect 36035 24157 36047 24160
rect 35989 24151 36047 24157
rect 37366 24148 37372 24160
rect 37424 24148 37430 24200
rect 37458 24148 37464 24200
rect 37516 24148 37522 24200
rect 35529 24123 35587 24129
rect 35529 24120 35541 24123
rect 34164 24092 35541 24120
rect 34057 24083 34115 24089
rect 35529 24089 35541 24092
rect 35575 24089 35587 24123
rect 35529 24083 35587 24089
rect 35618 24080 35624 24132
rect 35676 24120 35682 24132
rect 38105 24123 38163 24129
rect 38105 24120 38117 24123
rect 35676 24092 38117 24120
rect 35676 24080 35682 24092
rect 38105 24089 38117 24092
rect 38151 24089 38163 24123
rect 38488 24120 38516 24296
rect 38580 24197 38608 24364
rect 45922 24352 45928 24404
rect 45980 24392 45986 24404
rect 49421 24395 49479 24401
rect 49421 24392 49433 24395
rect 45980 24364 49433 24392
rect 45980 24352 45986 24364
rect 49421 24361 49433 24364
rect 49467 24361 49479 24395
rect 49421 24355 49479 24361
rect 39390 24284 39396 24336
rect 39448 24324 39454 24336
rect 44910 24324 44916 24336
rect 39448 24296 44916 24324
rect 39448 24284 39454 24296
rect 44910 24284 44916 24296
rect 44968 24284 44974 24336
rect 42613 24259 42671 24265
rect 42613 24225 42625 24259
rect 42659 24256 42671 24259
rect 45833 24259 45891 24265
rect 45833 24256 45845 24259
rect 42659 24228 45845 24256
rect 42659 24225 42671 24228
rect 42613 24219 42671 24225
rect 45833 24225 45845 24228
rect 45879 24225 45891 24259
rect 45833 24219 45891 24225
rect 38565 24191 38623 24197
rect 38565 24157 38577 24191
rect 38611 24157 38623 24191
rect 38565 24151 38623 24157
rect 40037 24191 40095 24197
rect 40037 24157 40049 24191
rect 40083 24157 40095 24191
rect 40037 24151 40095 24157
rect 41233 24191 41291 24197
rect 41233 24157 41245 24191
rect 41279 24188 41291 24191
rect 41414 24188 41420 24200
rect 41279 24160 41420 24188
rect 41279 24157 41291 24160
rect 41233 24151 41291 24157
rect 40052 24120 40080 24151
rect 41414 24148 41420 24160
rect 41472 24148 41478 24200
rect 41506 24148 41512 24200
rect 41564 24148 41570 24200
rect 42794 24148 42800 24200
rect 42852 24188 42858 24200
rect 42889 24191 42947 24197
rect 42889 24188 42901 24191
rect 42852 24160 42901 24188
rect 42852 24148 42858 24160
rect 42889 24157 42901 24160
rect 42935 24157 42947 24191
rect 42889 24151 42947 24157
rect 43898 24148 43904 24200
rect 43956 24148 43962 24200
rect 44450 24148 44456 24200
rect 44508 24188 44514 24200
rect 45189 24191 45247 24197
rect 45189 24188 45201 24191
rect 44508 24160 45201 24188
rect 44508 24148 44514 24160
rect 45189 24157 45201 24160
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 46569 24191 46627 24197
rect 46569 24157 46581 24191
rect 46615 24157 46627 24191
rect 46569 24151 46627 24157
rect 47765 24191 47823 24197
rect 47765 24157 47777 24191
rect 47811 24188 47823 24191
rect 48406 24188 48412 24200
rect 47811 24160 48412 24188
rect 47811 24157 47823 24160
rect 47765 24151 47823 24157
rect 38488 24092 40080 24120
rect 38105 24083 38163 24089
rect 42702 24080 42708 24132
rect 42760 24120 42766 24132
rect 46109 24123 46167 24129
rect 46109 24120 46121 24123
rect 42760 24092 46121 24120
rect 42760 24080 42766 24092
rect 46109 24089 46121 24092
rect 46155 24089 46167 24123
rect 46584 24120 46612 24151
rect 48406 24148 48412 24160
rect 48464 24148 48470 24200
rect 48869 24191 48927 24197
rect 48869 24157 48881 24191
rect 48915 24188 48927 24191
rect 49234 24188 49240 24200
rect 48915 24160 49240 24188
rect 48915 24157 48927 24160
rect 48869 24151 48927 24157
rect 49234 24148 49240 24160
rect 49292 24148 49298 24200
rect 49326 24120 49332 24132
rect 46584 24092 49332 24120
rect 46109 24083 46167 24089
rect 49326 24080 49332 24092
rect 49384 24080 49390 24132
rect 17862 24052 17868 24064
rect 14844 24024 17868 24052
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 18601 24055 18659 24061
rect 18601 24021 18613 24055
rect 18647 24052 18659 24055
rect 18782 24052 18788 24064
rect 18647 24024 18788 24052
rect 18647 24021 18659 24024
rect 18601 24015 18659 24021
rect 18782 24012 18788 24024
rect 18840 24012 18846 24064
rect 19058 24012 19064 24064
rect 19116 24012 19122 24064
rect 19429 24055 19487 24061
rect 19429 24021 19441 24055
rect 19475 24052 19487 24055
rect 24486 24052 24492 24064
rect 19475 24024 24492 24052
rect 19475 24021 19487 24024
rect 19429 24015 19487 24021
rect 24486 24012 24492 24024
rect 24544 24012 24550 24064
rect 24578 24012 24584 24064
rect 24636 24012 24642 24064
rect 25866 24012 25872 24064
rect 25924 24052 25930 24064
rect 26145 24055 26203 24061
rect 26145 24052 26157 24055
rect 25924 24024 26157 24052
rect 25924 24012 25930 24024
rect 26145 24021 26157 24024
rect 26191 24021 26203 24055
rect 26145 24015 26203 24021
rect 26237 24055 26295 24061
rect 26237 24021 26249 24055
rect 26283 24052 26295 24055
rect 26326 24052 26332 24064
rect 26283 24024 26332 24052
rect 26283 24021 26295 24024
rect 26237 24015 26295 24021
rect 26326 24012 26332 24024
rect 26384 24012 26390 24064
rect 26510 24012 26516 24064
rect 26568 24052 26574 24064
rect 27525 24055 27583 24061
rect 27525 24052 27537 24055
rect 26568 24024 27537 24052
rect 26568 24012 26574 24024
rect 27525 24021 27537 24024
rect 27571 24021 27583 24055
rect 27525 24015 27583 24021
rect 29270 24012 29276 24064
rect 29328 24012 29334 24064
rect 29362 24012 29368 24064
rect 29420 24052 29426 24064
rect 31665 24055 31723 24061
rect 31665 24052 31677 24055
rect 29420 24024 31677 24052
rect 29420 24012 29426 24024
rect 31665 24021 31677 24024
rect 31711 24021 31723 24055
rect 31665 24015 31723 24021
rect 32030 24012 32036 24064
rect 32088 24052 32094 24064
rect 35434 24052 35440 24064
rect 32088 24024 35440 24052
rect 32088 24012 32094 24024
rect 35434 24012 35440 24024
rect 35492 24012 35498 24064
rect 37458 24012 37464 24064
rect 37516 24052 37522 24064
rect 39209 24055 39267 24061
rect 39209 24052 39221 24055
rect 37516 24024 39221 24052
rect 37516 24012 37522 24024
rect 39209 24021 39221 24024
rect 39255 24021 39267 24055
rect 39209 24015 39267 24021
rect 39482 24012 39488 24064
rect 39540 24012 39546 24064
rect 39666 24012 39672 24064
rect 39724 24052 39730 24064
rect 40681 24055 40739 24061
rect 40681 24052 40693 24055
rect 39724 24024 40693 24052
rect 39724 24012 39730 24024
rect 40681 24021 40693 24024
rect 40727 24021 40739 24055
rect 40681 24015 40739 24021
rect 42886 24012 42892 24064
rect 42944 24052 42950 24064
rect 43806 24052 43812 24064
rect 42944 24024 43812 24052
rect 42944 24012 42950 24024
rect 43806 24012 43812 24024
rect 43864 24012 43870 24064
rect 44542 24012 44548 24064
rect 44600 24012 44606 24064
rect 47213 24055 47271 24061
rect 47213 24021 47225 24055
rect 47259 24052 47271 24055
rect 48314 24052 48320 24064
rect 47259 24024 48320 24052
rect 47259 24021 47271 24024
rect 47213 24015 47271 24021
rect 48314 24012 48320 24024
rect 48372 24012 48378 24064
rect 48409 24055 48467 24061
rect 48409 24021 48421 24055
rect 48455 24052 48467 24055
rect 48498 24052 48504 24064
rect 48455 24024 48504 24052
rect 48455 24021 48467 24024
rect 48409 24015 48467 24021
rect 48498 24012 48504 24024
rect 48556 24012 48562 24064
rect 48958 24012 48964 24064
rect 49016 24052 49022 24064
rect 49053 24055 49111 24061
rect 49053 24052 49065 24055
rect 49016 24024 49065 24052
rect 49016 24012 49022 24024
rect 49053 24021 49065 24024
rect 49099 24021 49111 24055
rect 49053 24015 49111 24021
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 1762 23808 1768 23860
rect 1820 23848 1826 23860
rect 14458 23848 14464 23860
rect 1820 23820 14464 23848
rect 1820 23808 1826 23820
rect 14458 23808 14464 23820
rect 14516 23808 14522 23860
rect 16298 23808 16304 23860
rect 16356 23848 16362 23860
rect 18966 23848 18972 23860
rect 16356 23820 18972 23848
rect 16356 23808 16362 23820
rect 18966 23808 18972 23820
rect 19024 23808 19030 23860
rect 19058 23808 19064 23860
rect 19116 23848 19122 23860
rect 21545 23851 21603 23857
rect 21545 23848 21557 23851
rect 19116 23820 21557 23848
rect 19116 23808 19122 23820
rect 21545 23817 21557 23820
rect 21591 23848 21603 23851
rect 22278 23848 22284 23860
rect 21591 23820 22284 23848
rect 21591 23817 21603 23820
rect 21545 23811 21603 23817
rect 22278 23808 22284 23820
rect 22336 23808 22342 23860
rect 23753 23851 23811 23857
rect 23753 23817 23765 23851
rect 23799 23848 23811 23851
rect 24854 23848 24860 23860
rect 23799 23820 24860 23848
rect 23799 23817 23811 23820
rect 23753 23811 23811 23817
rect 24854 23808 24860 23820
rect 24912 23808 24918 23860
rect 29362 23848 29368 23860
rect 25148 23820 29368 23848
rect 750 23740 756 23792
rect 808 23780 814 23792
rect 9122 23780 9128 23792
rect 808 23752 4660 23780
rect 808 23740 814 23752
rect 1949 23715 2007 23721
rect 1949 23681 1961 23715
rect 1995 23712 2007 23715
rect 2961 23715 3019 23721
rect 1995 23684 2728 23712
rect 1995 23681 2007 23684
rect 1949 23675 2007 23681
rect 2041 23647 2099 23653
rect 2041 23644 2053 23647
rect 1964 23616 2053 23644
rect 1964 23588 1992 23616
rect 2041 23613 2053 23616
rect 2087 23613 2099 23647
rect 2041 23607 2099 23613
rect 2225 23647 2283 23653
rect 2225 23613 2237 23647
rect 2271 23644 2283 23647
rect 2406 23644 2412 23656
rect 2271 23616 2412 23644
rect 2271 23613 2283 23616
rect 2225 23607 2283 23613
rect 2406 23604 2412 23616
rect 2464 23604 2470 23656
rect 1946 23536 1952 23588
rect 2004 23536 2010 23588
rect 2700 23576 2728 23684
rect 2961 23681 2973 23715
rect 3007 23681 3019 23715
rect 2961 23675 3019 23681
rect 3973 23715 4031 23721
rect 3973 23681 3985 23715
rect 4019 23712 4031 23715
rect 4154 23712 4160 23724
rect 4019 23684 4160 23712
rect 4019 23681 4031 23684
rect 3973 23675 4031 23681
rect 2774 23604 2780 23656
rect 2832 23644 2838 23656
rect 2976 23644 3004 23675
rect 4154 23672 4160 23684
rect 4212 23672 4218 23724
rect 4632 23721 4660 23752
rect 6564 23752 9128 23780
rect 6564 23721 6592 23752
rect 9122 23740 9128 23752
rect 9180 23740 9186 23792
rect 10965 23783 11023 23789
rect 10965 23749 10977 23783
rect 11011 23780 11023 23783
rect 11790 23780 11796 23792
rect 11011 23752 11796 23780
rect 11011 23749 11023 23752
rect 10965 23743 11023 23749
rect 11790 23740 11796 23752
rect 11848 23740 11854 23792
rect 12250 23740 12256 23792
rect 12308 23740 12314 23792
rect 12342 23740 12348 23792
rect 12400 23740 12406 23792
rect 13906 23780 13912 23792
rect 12636 23752 13912 23780
rect 4617 23715 4675 23721
rect 4617 23681 4629 23715
rect 4663 23681 4675 23715
rect 6549 23715 6607 23721
rect 4617 23675 4675 23681
rect 4724 23684 6500 23712
rect 4724 23644 4752 23684
rect 2832 23616 2912 23644
rect 2976 23616 4752 23644
rect 2832 23604 2838 23616
rect 2884 23576 2912 23616
rect 5442 23604 5448 23656
rect 5500 23604 5506 23656
rect 6472 23644 6500 23684
rect 6549 23681 6561 23715
rect 6595 23681 6607 23715
rect 6549 23675 6607 23681
rect 6730 23672 6736 23724
rect 6788 23712 6794 23724
rect 6825 23715 6883 23721
rect 6825 23712 6837 23715
rect 6788 23684 6837 23712
rect 6788 23672 6794 23684
rect 6825 23681 6837 23684
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 8021 23715 8079 23721
rect 8021 23681 8033 23715
rect 8067 23681 8079 23715
rect 8021 23675 8079 23681
rect 7926 23644 7932 23656
rect 6472 23616 7932 23644
rect 7926 23604 7932 23616
rect 7984 23604 7990 23656
rect 4982 23576 4988 23588
rect 2700 23548 2774 23576
rect 2884 23548 4988 23576
rect 1581 23511 1639 23517
rect 1581 23477 1593 23511
rect 1627 23508 1639 23511
rect 2590 23508 2596 23520
rect 1627 23480 2596 23508
rect 1627 23477 1639 23480
rect 1581 23471 1639 23477
rect 2590 23468 2596 23480
rect 2648 23468 2654 23520
rect 2746 23508 2774 23548
rect 4982 23536 4988 23548
rect 5040 23536 5046 23588
rect 5350 23536 5356 23588
rect 5408 23576 5414 23588
rect 8036 23576 8064 23675
rect 9858 23672 9864 23724
rect 9916 23672 9922 23724
rect 11701 23715 11759 23721
rect 11701 23681 11713 23715
rect 11747 23712 11759 23715
rect 12268 23712 12296 23740
rect 12636 23712 12664 23752
rect 13906 23740 13912 23752
rect 13964 23740 13970 23792
rect 14277 23783 14335 23789
rect 14277 23749 14289 23783
rect 14323 23780 14335 23783
rect 15746 23780 15752 23792
rect 14323 23752 15752 23780
rect 14323 23749 14335 23752
rect 14277 23743 14335 23749
rect 15746 23740 15752 23752
rect 15804 23740 15810 23792
rect 15930 23740 15936 23792
rect 15988 23780 15994 23792
rect 17586 23780 17592 23792
rect 15988 23752 17592 23780
rect 15988 23740 15994 23752
rect 17586 23740 17592 23752
rect 17644 23740 17650 23792
rect 18141 23783 18199 23789
rect 18141 23749 18153 23783
rect 18187 23780 18199 23783
rect 19150 23780 19156 23792
rect 18187 23752 19156 23780
rect 18187 23749 18199 23752
rect 18141 23743 18199 23749
rect 19150 23740 19156 23752
rect 19208 23740 19214 23792
rect 19518 23740 19524 23792
rect 19576 23740 19582 23792
rect 21358 23740 21364 23792
rect 21416 23780 21422 23792
rect 22554 23780 22560 23792
rect 21416 23752 22560 23780
rect 21416 23740 21422 23752
rect 22554 23740 22560 23752
rect 22612 23740 22618 23792
rect 23290 23740 23296 23792
rect 23348 23740 23354 23792
rect 24213 23783 24271 23789
rect 24213 23749 24225 23783
rect 24259 23780 24271 23783
rect 25038 23780 25044 23792
rect 24259 23752 25044 23780
rect 24259 23749 24271 23752
rect 24213 23743 24271 23749
rect 25038 23740 25044 23752
rect 25096 23740 25102 23792
rect 25148 23789 25176 23820
rect 29362 23808 29368 23820
rect 29420 23808 29426 23860
rect 31018 23808 31024 23860
rect 31076 23848 31082 23860
rect 32953 23851 33011 23857
rect 32953 23848 32965 23851
rect 31076 23820 32965 23848
rect 31076 23808 31082 23820
rect 32953 23817 32965 23820
rect 32999 23817 33011 23851
rect 32953 23811 33011 23817
rect 33686 23808 33692 23860
rect 33744 23848 33750 23860
rect 34425 23851 34483 23857
rect 34425 23848 34437 23851
rect 33744 23820 34437 23848
rect 33744 23808 33750 23820
rect 34425 23817 34437 23820
rect 34471 23848 34483 23851
rect 34471 23820 36124 23848
rect 34471 23817 34483 23820
rect 34425 23811 34483 23817
rect 25133 23783 25191 23789
rect 25133 23749 25145 23783
rect 25179 23749 25191 23783
rect 27062 23780 27068 23792
rect 26358 23752 27068 23780
rect 25133 23743 25191 23749
rect 27062 23740 27068 23752
rect 27120 23780 27126 23792
rect 27706 23780 27712 23792
rect 27120 23752 27712 23780
rect 27120 23740 27126 23752
rect 27706 23740 27712 23752
rect 27764 23740 27770 23792
rect 28810 23780 28816 23792
rect 28658 23766 28816 23780
rect 28644 23752 28816 23766
rect 11747 23684 12296 23712
rect 12544 23684 12664 23712
rect 13265 23715 13323 23721
rect 11747 23681 11759 23684
rect 11701 23675 11759 23681
rect 9125 23647 9183 23653
rect 9125 23613 9137 23647
rect 9171 23644 9183 23647
rect 9950 23644 9956 23656
rect 9171 23616 9956 23644
rect 9171 23613 9183 23616
rect 9125 23607 9183 23613
rect 9950 23604 9956 23616
rect 10008 23604 10014 23656
rect 12342 23644 12348 23656
rect 10060 23616 12348 23644
rect 5408 23548 8064 23576
rect 5408 23536 5414 23548
rect 8110 23536 8116 23588
rect 8168 23576 8174 23588
rect 10060 23576 10088 23616
rect 12342 23604 12348 23616
rect 12400 23604 12406 23656
rect 12544 23653 12572 23684
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13354 23712 13360 23724
rect 13311 23684 13360 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13354 23672 13360 23684
rect 13412 23672 13418 23724
rect 14918 23672 14924 23724
rect 14976 23672 14982 23724
rect 17129 23715 17187 23721
rect 17129 23681 17141 23715
rect 17175 23712 17187 23715
rect 18506 23712 18512 23724
rect 17175 23684 18512 23712
rect 17175 23681 17187 23684
rect 17129 23675 17187 23681
rect 18506 23672 18512 23684
rect 18564 23672 18570 23724
rect 20990 23672 20996 23724
rect 21048 23672 21054 23724
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 16117 23647 16175 23653
rect 16117 23613 16129 23647
rect 16163 23644 16175 23647
rect 18322 23644 18328 23656
rect 16163 23616 18328 23644
rect 16163 23613 16175 23616
rect 16117 23607 16175 23613
rect 18322 23604 18328 23616
rect 18380 23604 18386 23656
rect 18782 23604 18788 23656
rect 18840 23604 18846 23656
rect 19061 23647 19119 23653
rect 19061 23644 19073 23647
rect 18892 23616 19073 23644
rect 8168 23548 10088 23576
rect 11609 23579 11667 23585
rect 8168 23536 8174 23548
rect 11609 23545 11621 23579
rect 11655 23576 11667 23579
rect 15194 23576 15200 23588
rect 11655 23548 12572 23576
rect 11655 23545 11667 23548
rect 11609 23539 11667 23545
rect 7650 23508 7656 23520
rect 2746 23480 7656 23508
rect 7650 23468 7656 23480
rect 7708 23468 7714 23520
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 9674 23508 9680 23520
rect 7984 23480 9680 23508
rect 7984 23468 7990 23480
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 11885 23511 11943 23517
rect 11885 23477 11897 23511
rect 11931 23508 11943 23511
rect 12158 23508 12164 23520
rect 11931 23480 12164 23508
rect 11931 23477 11943 23480
rect 11885 23471 11943 23477
rect 12158 23468 12164 23480
rect 12216 23468 12222 23520
rect 12544 23508 12572 23548
rect 13832 23548 15200 23576
rect 13832 23508 13860 23548
rect 15194 23536 15200 23548
rect 15252 23536 15258 23588
rect 15286 23536 15292 23588
rect 15344 23576 15350 23588
rect 18230 23576 18236 23588
rect 15344 23548 18236 23576
rect 15344 23536 15350 23548
rect 18230 23536 18236 23548
rect 18288 23536 18294 23588
rect 18690 23536 18696 23588
rect 18748 23576 18754 23588
rect 18892 23576 18920 23616
rect 19061 23613 19073 23616
rect 19107 23613 19119 23647
rect 19061 23607 19119 23613
rect 19150 23604 19156 23656
rect 19208 23644 19214 23656
rect 19208 23616 20116 23644
rect 19208 23604 19214 23616
rect 18748 23548 18920 23576
rect 20088 23576 20116 23616
rect 20898 23604 20904 23656
rect 20956 23644 20962 23656
rect 22005 23647 22063 23653
rect 22005 23644 22017 23647
rect 20956 23616 22017 23644
rect 20956 23604 20962 23616
rect 22005 23613 22017 23616
rect 22051 23613 22063 23647
rect 22005 23607 22063 23613
rect 22281 23647 22339 23653
rect 22281 23613 22293 23647
rect 22327 23644 22339 23647
rect 22370 23644 22376 23656
rect 22327 23616 22376 23644
rect 22327 23613 22339 23616
rect 22281 23607 22339 23613
rect 22370 23604 22376 23616
rect 22428 23604 22434 23656
rect 22738 23604 22744 23656
rect 22796 23644 22802 23656
rect 22922 23644 22928 23656
rect 22796 23616 22928 23644
rect 22796 23604 22802 23616
rect 22922 23604 22928 23616
rect 22980 23604 22986 23656
rect 24854 23644 24860 23656
rect 23400 23616 24860 23644
rect 23400 23588 23428 23616
rect 24854 23604 24860 23616
rect 24912 23604 24918 23656
rect 26418 23644 26424 23656
rect 24964 23616 26424 23644
rect 20088 23548 20208 23576
rect 18748 23536 18754 23548
rect 12544 23480 13860 23508
rect 13906 23468 13912 23520
rect 13964 23508 13970 23520
rect 18708 23508 18736 23536
rect 13964 23480 18736 23508
rect 13964 23468 13970 23480
rect 18782 23468 18788 23520
rect 18840 23508 18846 23520
rect 20070 23508 20076 23520
rect 18840 23480 20076 23508
rect 18840 23468 18846 23480
rect 20070 23468 20076 23480
rect 20128 23468 20134 23520
rect 20180 23508 20208 23548
rect 20346 23536 20352 23588
rect 20404 23576 20410 23588
rect 21177 23579 21235 23585
rect 21177 23576 21189 23579
rect 20404 23548 21189 23576
rect 20404 23536 20410 23548
rect 21177 23545 21189 23548
rect 21223 23545 21235 23579
rect 21177 23539 21235 23545
rect 23382 23536 23388 23588
rect 23440 23536 23446 23588
rect 24964 23576 24992 23616
rect 26418 23604 26424 23616
rect 26476 23604 26482 23656
rect 27157 23647 27215 23653
rect 27157 23644 27169 23647
rect 27080 23616 27169 23644
rect 24780 23548 24992 23576
rect 20533 23511 20591 23517
rect 20533 23508 20545 23511
rect 20180 23480 20545 23508
rect 20533 23477 20545 23480
rect 20579 23508 20591 23511
rect 24780 23508 24808 23548
rect 26602 23536 26608 23588
rect 26660 23536 26666 23588
rect 20579 23480 24808 23508
rect 20579 23477 20591 23480
rect 20533 23471 20591 23477
rect 24854 23468 24860 23520
rect 24912 23508 24918 23520
rect 27080 23508 27108 23616
rect 27157 23613 27169 23616
rect 27203 23613 27215 23647
rect 27157 23607 27215 23613
rect 27430 23604 27436 23656
rect 27488 23604 27494 23656
rect 27798 23604 27804 23656
rect 27856 23644 27862 23656
rect 28644 23644 28672 23752
rect 28810 23740 28816 23752
rect 28868 23740 28874 23792
rect 28902 23740 28908 23792
rect 28960 23780 28966 23792
rect 31386 23780 31392 23792
rect 28960 23752 31392 23780
rect 28960 23740 28966 23752
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 32030 23780 32036 23792
rect 31680 23752 32036 23780
rect 28994 23672 29000 23724
rect 29052 23712 29058 23724
rect 29365 23715 29423 23721
rect 29365 23712 29377 23715
rect 29052 23684 29377 23712
rect 29052 23672 29058 23684
rect 29365 23681 29377 23684
rect 29411 23681 29423 23715
rect 29365 23675 29423 23681
rect 29472 23684 29776 23712
rect 27856 23616 28672 23644
rect 27856 23604 27862 23616
rect 28810 23604 28816 23656
rect 28868 23644 28874 23656
rect 29472 23644 29500 23684
rect 28868 23616 29500 23644
rect 28868 23604 28874 23616
rect 29638 23604 29644 23656
rect 29696 23604 29702 23656
rect 29748 23644 29776 23684
rect 30742 23672 30748 23724
rect 30800 23712 30806 23724
rect 30837 23715 30895 23721
rect 30837 23712 30849 23715
rect 30800 23684 30849 23712
rect 30800 23672 30806 23684
rect 30837 23681 30849 23684
rect 30883 23681 30895 23715
rect 31680 23712 31708 23752
rect 32030 23740 32036 23752
rect 32088 23740 32094 23792
rect 32214 23740 32220 23792
rect 32272 23780 32278 23792
rect 34057 23783 34115 23789
rect 32272 23752 33456 23780
rect 32272 23740 32278 23752
rect 30837 23675 30895 23681
rect 30944 23684 31708 23712
rect 30944 23644 30972 23684
rect 32306 23672 32312 23724
rect 32364 23672 32370 23724
rect 33428 23721 33456 23752
rect 34057 23749 34069 23783
rect 34103 23780 34115 23783
rect 36096 23780 36124 23820
rect 40310 23808 40316 23860
rect 40368 23808 40374 23860
rect 41414 23808 41420 23860
rect 41472 23848 41478 23860
rect 47029 23851 47087 23857
rect 47029 23848 47041 23851
rect 41472 23820 47041 23848
rect 41472 23808 41478 23820
rect 47029 23817 47041 23820
rect 47075 23817 47087 23851
rect 47029 23811 47087 23817
rect 48406 23808 48412 23860
rect 48464 23808 48470 23860
rect 34103 23752 36032 23780
rect 36096 23752 40632 23780
rect 34103 23749 34115 23752
rect 34057 23743 34115 23749
rect 33413 23715 33471 23721
rect 33413 23681 33425 23715
rect 33459 23681 33471 23715
rect 33413 23675 33471 23681
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23712 34943 23715
rect 35618 23712 35624 23724
rect 34931 23684 35624 23712
rect 34931 23681 34943 23684
rect 34885 23675 34943 23681
rect 35618 23672 35624 23684
rect 35676 23672 35682 23724
rect 36004 23721 36032 23752
rect 35989 23715 36047 23721
rect 35989 23681 36001 23715
rect 36035 23681 36047 23715
rect 35989 23675 36047 23681
rect 37461 23715 37519 23721
rect 37461 23681 37473 23715
rect 37507 23681 37519 23715
rect 37461 23675 37519 23681
rect 38565 23715 38623 23721
rect 38565 23681 38577 23715
rect 38611 23681 38623 23715
rect 38565 23675 38623 23681
rect 29748 23616 30972 23644
rect 31110 23604 31116 23656
rect 31168 23644 31174 23656
rect 31573 23647 31631 23653
rect 31573 23644 31585 23647
rect 31168 23616 31585 23644
rect 31168 23604 31174 23616
rect 31573 23613 31585 23616
rect 31619 23613 31631 23647
rect 31573 23607 31631 23613
rect 31662 23604 31668 23656
rect 31720 23644 31726 23656
rect 35529 23647 35587 23653
rect 31720 23616 34928 23644
rect 31720 23604 31726 23616
rect 28905 23579 28963 23585
rect 28905 23545 28917 23579
rect 28951 23576 28963 23579
rect 29454 23576 29460 23588
rect 28951 23548 29460 23576
rect 28951 23545 28963 23548
rect 28905 23539 28963 23545
rect 29454 23536 29460 23548
rect 29512 23536 29518 23588
rect 29730 23536 29736 23588
rect 29788 23576 29794 23588
rect 34517 23579 34575 23585
rect 34517 23576 34529 23579
rect 29788 23548 34529 23576
rect 29788 23536 29794 23548
rect 34517 23545 34529 23548
rect 34563 23545 34575 23579
rect 34900 23576 34928 23616
rect 35529 23613 35541 23647
rect 35575 23644 35587 23647
rect 37476 23644 37504 23675
rect 35575 23616 37504 23644
rect 38580 23644 38608 23675
rect 39666 23672 39672 23724
rect 39724 23672 39730 23724
rect 40494 23644 40500 23656
rect 38580 23616 40500 23644
rect 35575 23613 35587 23616
rect 35529 23607 35587 23613
rect 40494 23604 40500 23616
rect 40552 23604 40558 23656
rect 38105 23579 38163 23585
rect 38105 23576 38117 23579
rect 34900 23548 38117 23576
rect 34517 23539 34575 23545
rect 38105 23545 38117 23548
rect 38151 23545 38163 23579
rect 38105 23539 38163 23545
rect 39942 23536 39948 23588
rect 40000 23576 40006 23588
rect 40604 23576 40632 23752
rect 42702 23740 42708 23792
rect 42760 23740 42766 23792
rect 42886 23740 42892 23792
rect 42944 23740 42950 23792
rect 47213 23783 47271 23789
rect 47213 23780 47225 23783
rect 43548 23752 47225 23780
rect 40773 23715 40831 23721
rect 40773 23681 40785 23715
rect 40819 23712 40831 23715
rect 41782 23712 41788 23724
rect 40819 23684 41788 23712
rect 40819 23681 40831 23684
rect 40773 23675 40831 23681
rect 41782 23672 41788 23684
rect 41840 23672 41846 23724
rect 42061 23715 42119 23721
rect 42061 23681 42073 23715
rect 42107 23681 42119 23715
rect 42061 23675 42119 23681
rect 42076 23644 42104 23675
rect 42794 23672 42800 23724
rect 42852 23712 42858 23724
rect 43165 23715 43223 23721
rect 43165 23712 43177 23715
rect 42852 23684 43177 23712
rect 42852 23672 42858 23684
rect 43165 23681 43177 23684
rect 43211 23681 43223 23715
rect 43165 23675 43223 23681
rect 43346 23672 43352 23724
rect 43404 23712 43410 23724
rect 43548 23721 43576 23752
rect 47213 23749 47225 23752
rect 47259 23749 47271 23783
rect 47213 23743 47271 23749
rect 47302 23740 47308 23792
rect 47360 23780 47366 23792
rect 49421 23783 49479 23789
rect 49421 23780 49433 23783
rect 47360 23752 49433 23780
rect 47360 23740 47366 23752
rect 49421 23749 49433 23752
rect 49467 23749 49479 23783
rect 49421 23743 49479 23749
rect 43533 23715 43591 23721
rect 43533 23712 43545 23715
rect 43404 23684 43545 23712
rect 43404 23672 43410 23684
rect 43533 23681 43545 23684
rect 43579 23681 43591 23715
rect 43533 23675 43591 23681
rect 44818 23672 44824 23724
rect 44876 23672 44882 23724
rect 46201 23715 46259 23721
rect 46201 23712 46213 23715
rect 45526 23684 46213 23712
rect 43438 23644 43444 23656
rect 42076 23616 43444 23644
rect 43438 23604 43444 23616
rect 43496 23604 43502 23656
rect 43809 23647 43867 23653
rect 43809 23613 43821 23647
rect 43855 23613 43867 23647
rect 43809 23607 43867 23613
rect 41417 23579 41475 23585
rect 41417 23576 41429 23579
rect 40000 23548 40540 23576
rect 40604 23548 41429 23576
rect 40000 23536 40006 23548
rect 27154 23508 27160 23520
rect 24912 23480 27160 23508
rect 24912 23468 24918 23480
rect 27154 23468 27160 23480
rect 27212 23468 27218 23520
rect 27246 23468 27252 23520
rect 27304 23508 27310 23520
rect 28994 23508 29000 23520
rect 27304 23480 29000 23508
rect 27304 23468 27310 23480
rect 28994 23468 29000 23480
rect 29052 23468 29058 23520
rect 29270 23468 29276 23520
rect 29328 23508 29334 23520
rect 30469 23511 30527 23517
rect 30469 23508 30481 23511
rect 29328 23480 30481 23508
rect 29328 23468 29334 23480
rect 30469 23477 30481 23480
rect 30515 23508 30527 23511
rect 31754 23508 31760 23520
rect 30515 23480 31760 23508
rect 30515 23477 30527 23480
rect 30469 23471 30527 23477
rect 31754 23468 31760 23480
rect 31812 23468 31818 23520
rect 35986 23468 35992 23520
rect 36044 23508 36050 23520
rect 36633 23511 36691 23517
rect 36633 23508 36645 23511
rect 36044 23480 36645 23508
rect 36044 23468 36050 23480
rect 36633 23477 36645 23480
rect 36679 23477 36691 23511
rect 36633 23471 36691 23477
rect 37090 23468 37096 23520
rect 37148 23468 37154 23520
rect 38562 23468 38568 23520
rect 38620 23508 38626 23520
rect 39209 23511 39267 23517
rect 39209 23508 39221 23511
rect 38620 23480 39221 23508
rect 38620 23468 38626 23480
rect 39209 23477 39221 23480
rect 39255 23477 39267 23511
rect 40512 23508 40540 23548
rect 41417 23545 41429 23548
rect 41463 23545 41475 23579
rect 41417 23539 41475 23545
rect 41874 23536 41880 23588
rect 41932 23536 41938 23588
rect 43824 23508 43852 23607
rect 44836 23576 44864 23672
rect 44910 23604 44916 23656
rect 44968 23644 44974 23656
rect 45526 23644 45554 23684
rect 46201 23681 46213 23684
rect 46247 23681 46259 23715
rect 46201 23675 46259 23681
rect 47026 23672 47032 23724
rect 47084 23712 47090 23724
rect 47765 23715 47823 23721
rect 47765 23712 47777 23715
rect 47084 23684 47777 23712
rect 47084 23672 47090 23684
rect 47765 23681 47777 23684
rect 47811 23681 47823 23715
rect 47765 23675 47823 23681
rect 48866 23672 48872 23724
rect 48924 23672 48930 23724
rect 44968 23616 45554 23644
rect 44968 23604 44974 23616
rect 45922 23604 45928 23656
rect 45980 23604 45986 23656
rect 46934 23576 46940 23588
rect 44836 23548 46940 23576
rect 46934 23536 46940 23548
rect 46992 23536 46998 23588
rect 40512 23480 43852 23508
rect 39209 23471 39267 23477
rect 44174 23468 44180 23520
rect 44232 23508 44238 23520
rect 45465 23511 45523 23517
rect 45465 23508 45477 23511
rect 44232 23480 45477 23508
rect 44232 23468 44238 23480
rect 45465 23477 45477 23480
rect 45511 23477 45523 23511
rect 45465 23471 45523 23477
rect 49050 23468 49056 23520
rect 49108 23468 49114 23520
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 2866 23264 2872 23316
rect 2924 23304 2930 23316
rect 4154 23304 4160 23316
rect 2924 23276 4160 23304
rect 2924 23264 2930 23276
rect 4154 23264 4160 23276
rect 4212 23264 4218 23316
rect 8018 23264 8024 23316
rect 8076 23304 8082 23316
rect 12618 23304 12624 23316
rect 8076 23276 12624 23304
rect 8076 23264 8082 23276
rect 12618 23264 12624 23276
rect 12676 23264 12682 23316
rect 13538 23264 13544 23316
rect 13596 23304 13602 23316
rect 14182 23304 14188 23316
rect 13596 23276 14188 23304
rect 13596 23264 13602 23276
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 18877 23307 18935 23313
rect 18877 23273 18889 23307
rect 18923 23304 18935 23307
rect 18923 23276 23796 23304
rect 18923 23273 18935 23276
rect 18877 23267 18935 23273
rect 3602 23196 3608 23248
rect 3660 23196 3666 23248
rect 7282 23236 7288 23248
rect 4172 23208 7288 23236
rect 3421 23171 3479 23177
rect 3421 23137 3433 23171
rect 3467 23168 3479 23171
rect 4172 23168 4200 23208
rect 7282 23196 7288 23208
rect 7340 23236 7346 23248
rect 7340 23208 9076 23236
rect 7340 23196 7346 23208
rect 3467 23140 4200 23168
rect 4249 23171 4307 23177
rect 3467 23137 3479 23140
rect 3421 23131 3479 23137
rect 4249 23137 4261 23171
rect 4295 23168 4307 23171
rect 5258 23168 5264 23180
rect 4295 23140 5264 23168
rect 4295 23137 4307 23140
rect 4249 23131 4307 23137
rect 5258 23128 5264 23140
rect 5316 23128 5322 23180
rect 6086 23128 6092 23180
rect 6144 23128 6150 23180
rect 7834 23128 7840 23180
rect 7892 23128 7898 23180
rect 9048 23168 9076 23208
rect 9646 23208 10640 23236
rect 9646 23168 9674 23208
rect 9048 23140 9674 23168
rect 10502 23128 10508 23180
rect 10560 23128 10566 23180
rect 10612 23168 10640 23208
rect 13906 23196 13912 23248
rect 13964 23196 13970 23248
rect 14090 23196 14096 23248
rect 14148 23236 14154 23248
rect 14148 23208 17264 23236
rect 14148 23196 14154 23208
rect 11790 23168 11796 23180
rect 10612 23140 11796 23168
rect 11790 23128 11796 23140
rect 11848 23128 11854 23180
rect 11882 23128 11888 23180
rect 11940 23168 11946 23180
rect 12802 23168 12808 23180
rect 11940 23140 12808 23168
rect 11940 23128 11946 23140
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 13538 23128 13544 23180
rect 13596 23168 13602 23180
rect 14734 23168 14740 23180
rect 13596 23140 14740 23168
rect 13596 23128 13602 23140
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 16850 23128 16856 23180
rect 16908 23168 16914 23180
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 16908 23140 17141 23168
rect 16908 23128 16914 23140
rect 17129 23137 17141 23140
rect 17175 23137 17187 23171
rect 17236 23168 17264 23208
rect 17405 23171 17463 23177
rect 17405 23168 17417 23171
rect 17236 23140 17417 23168
rect 17129 23131 17187 23137
rect 17405 23137 17417 23140
rect 17451 23168 17463 23171
rect 17770 23168 17776 23180
rect 17451 23140 17776 23168
rect 17451 23137 17463 23140
rect 17405 23131 17463 23137
rect 17770 23128 17776 23140
rect 17828 23128 17834 23180
rect 20070 23128 20076 23180
rect 20128 23168 20134 23180
rect 20898 23168 20904 23180
rect 20128 23140 20904 23168
rect 20128 23128 20134 23140
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 22278 23128 22284 23180
rect 22336 23128 22342 23180
rect 22557 23171 22615 23177
rect 22557 23137 22569 23171
rect 22603 23168 22615 23171
rect 22646 23168 22652 23180
rect 22603 23140 22652 23168
rect 22603 23137 22615 23140
rect 22557 23131 22615 23137
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 23290 23128 23296 23180
rect 23348 23168 23354 23180
rect 23348 23140 23704 23168
rect 23348 23128 23354 23140
rect 23676 23112 23704 23140
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 1854 23100 1860 23112
rect 1811 23072 1860 23100
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23069 4031 23103
rect 3973 23063 4031 23069
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23100 5503 23103
rect 6178 23100 6184 23112
rect 5491 23072 6184 23100
rect 5491 23069 5503 23072
rect 5445 23063 5503 23069
rect 2774 22992 2780 23044
rect 2832 22992 2838 23044
rect 3988 23032 4016 23063
rect 6178 23060 6184 23072
rect 6236 23060 6242 23112
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 8018 23100 8024 23112
rect 7423 23072 8024 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 9490 23060 9496 23112
rect 9548 23060 9554 23112
rect 11146 23060 11152 23112
rect 11204 23060 11210 23112
rect 14642 23060 14648 23112
rect 14700 23060 14706 23112
rect 15470 23060 15476 23112
rect 15528 23060 15534 23112
rect 16393 23103 16451 23109
rect 16393 23069 16405 23103
rect 16439 23100 16451 23103
rect 16439 23072 16988 23100
rect 16439 23069 16451 23072
rect 16393 23063 16451 23069
rect 11054 23032 11060 23044
rect 3988 23004 11060 23032
rect 11054 22992 11060 23004
rect 11112 22992 11118 23044
rect 11422 22992 11428 23044
rect 11480 22992 11486 23044
rect 12986 23032 12992 23044
rect 12650 23004 12992 23032
rect 9030 22924 9036 22976
rect 9088 22924 9094 22976
rect 9398 22924 9404 22976
rect 9456 22964 9462 22976
rect 10778 22964 10784 22976
rect 9456 22936 10784 22964
rect 9456 22924 9462 22936
rect 10778 22924 10784 22936
rect 10836 22964 10842 22976
rect 12728 22964 12756 23004
rect 12986 22992 12992 23004
rect 13044 22992 13050 23044
rect 13173 23035 13231 23041
rect 13173 23001 13185 23035
rect 13219 23032 13231 23035
rect 13354 23032 13360 23044
rect 13219 23004 13360 23032
rect 13219 23001 13231 23004
rect 13173 22995 13231 23001
rect 13354 22992 13360 23004
rect 13412 22992 13418 23044
rect 13541 23035 13599 23041
rect 13541 23001 13553 23035
rect 13587 23032 13599 23035
rect 16960 23032 16988 23072
rect 23658 23060 23664 23112
rect 23716 23060 23722 23112
rect 23768 23100 23796 23276
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 24854 23304 24860 23316
rect 23900 23276 24860 23304
rect 23900 23264 23906 23276
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 26050 23264 26056 23316
rect 26108 23304 26114 23316
rect 29638 23304 29644 23316
rect 26108 23276 29644 23304
rect 26108 23264 26114 23276
rect 29638 23264 29644 23276
rect 29696 23264 29702 23316
rect 30190 23264 30196 23316
rect 30248 23304 30254 23316
rect 32214 23304 32220 23316
rect 30248 23276 32220 23304
rect 30248 23264 30254 23276
rect 32214 23264 32220 23276
rect 32272 23264 32278 23316
rect 32306 23264 32312 23316
rect 32364 23304 32370 23316
rect 32953 23307 33011 23313
rect 32953 23304 32965 23307
rect 32364 23276 32965 23304
rect 32364 23264 32370 23276
rect 32953 23273 32965 23276
rect 32999 23273 33011 23307
rect 36633 23307 36691 23313
rect 36633 23304 36645 23307
rect 32953 23267 33011 23273
rect 33060 23276 36645 23304
rect 24118 23196 24124 23248
rect 24176 23236 24182 23248
rect 24762 23236 24768 23248
rect 24176 23208 24768 23236
rect 24176 23196 24182 23208
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 25314 23196 25320 23248
rect 25372 23236 25378 23248
rect 25372 23208 26648 23236
rect 25372 23196 25378 23208
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23168 25283 23171
rect 25774 23168 25780 23180
rect 25271 23140 25780 23168
rect 25271 23137 25283 23140
rect 25225 23131 25283 23137
rect 25774 23128 25780 23140
rect 25832 23128 25838 23180
rect 25958 23128 25964 23180
rect 26016 23168 26022 23180
rect 26329 23171 26387 23177
rect 26329 23168 26341 23171
rect 26016 23140 26341 23168
rect 26016 23128 26022 23140
rect 26329 23137 26341 23140
rect 26375 23137 26387 23171
rect 26329 23131 26387 23137
rect 23768 23072 26096 23100
rect 17678 23032 17684 23044
rect 13587 23004 16160 23032
rect 16960 23004 17684 23032
rect 13587 23001 13599 23004
rect 13541 22995 13599 23001
rect 10836 22936 12756 22964
rect 10836 22924 10842 22936
rect 13722 22924 13728 22976
rect 13780 22924 13786 22976
rect 14274 22924 14280 22976
rect 14332 22924 14338 22976
rect 14734 22924 14740 22976
rect 14792 22924 14798 22976
rect 16132 22964 16160 23004
rect 17678 22992 17684 23004
rect 17736 22992 17742 23044
rect 18414 22992 18420 23044
rect 18472 22992 18478 23044
rect 20254 22992 20260 23044
rect 20312 23032 20318 23044
rect 20349 23035 20407 23041
rect 20349 23032 20361 23035
rect 20312 23004 20361 23032
rect 20312 22992 20318 23004
rect 20349 23001 20361 23004
rect 20395 23001 20407 23035
rect 20349 22995 20407 23001
rect 17218 22964 17224 22976
rect 16132 22936 17224 22964
rect 17218 22924 17224 22936
rect 17276 22924 17282 22976
rect 18966 22924 18972 22976
rect 19024 22964 19030 22976
rect 19429 22967 19487 22973
rect 19429 22964 19441 22967
rect 19024 22936 19441 22964
rect 19024 22924 19030 22936
rect 19429 22933 19441 22936
rect 19475 22933 19487 22967
rect 20364 22964 20392 22995
rect 20622 22992 20628 23044
rect 20680 23032 20686 23044
rect 20680 23004 20838 23032
rect 21652 23004 22094 23032
rect 20680 22992 20686 23004
rect 21082 22964 21088 22976
rect 20364 22936 21088 22964
rect 19429 22927 19487 22933
rect 21082 22924 21088 22936
rect 21140 22924 21146 22976
rect 21174 22924 21180 22976
rect 21232 22964 21238 22976
rect 21652 22964 21680 23004
rect 21232 22936 21680 22964
rect 21232 22924 21238 22936
rect 21818 22924 21824 22976
rect 21876 22924 21882 22976
rect 22066 22964 22094 23004
rect 23290 22992 23296 23044
rect 23348 22992 23354 23044
rect 23860 23004 24624 23032
rect 23860 22964 23888 23004
rect 22066 22936 23888 22964
rect 24029 22967 24087 22973
rect 24029 22933 24041 22967
rect 24075 22964 24087 22967
rect 24118 22964 24124 22976
rect 24075 22936 24124 22964
rect 24075 22933 24087 22936
rect 24029 22927 24087 22933
rect 24118 22924 24124 22936
rect 24176 22924 24182 22976
rect 24596 22973 24624 23004
rect 24946 22992 24952 23044
rect 25004 22992 25010 23044
rect 26068 23032 26096 23072
rect 26142 23060 26148 23112
rect 26200 23100 26206 23112
rect 26237 23103 26295 23109
rect 26237 23100 26249 23103
rect 26200 23072 26249 23100
rect 26200 23060 26206 23072
rect 26237 23069 26249 23072
rect 26283 23069 26295 23103
rect 26620 23100 26648 23208
rect 26694 23196 26700 23248
rect 26752 23236 26758 23248
rect 27246 23236 27252 23248
rect 26752 23208 27252 23236
rect 26752 23196 26758 23208
rect 27246 23196 27252 23208
rect 27304 23196 27310 23248
rect 29086 23196 29092 23248
rect 29144 23196 29150 23248
rect 31754 23196 31760 23248
rect 31812 23236 31818 23248
rect 31941 23239 31999 23245
rect 31941 23236 31953 23239
rect 31812 23208 31953 23236
rect 31812 23196 31818 23208
rect 31941 23205 31953 23208
rect 31987 23205 31999 23239
rect 33060 23236 33088 23276
rect 36633 23273 36645 23276
rect 36679 23273 36691 23307
rect 36633 23267 36691 23273
rect 40494 23264 40500 23316
rect 40552 23304 40558 23316
rect 40681 23307 40739 23313
rect 40681 23304 40693 23307
rect 40552 23276 40693 23304
rect 40552 23264 40558 23276
rect 40681 23273 40693 23276
rect 40727 23273 40739 23307
rect 40681 23267 40739 23273
rect 41782 23264 41788 23316
rect 41840 23264 41846 23316
rect 43162 23304 43168 23316
rect 42812 23276 43168 23304
rect 31941 23199 31999 23205
rect 32324 23208 33088 23236
rect 27154 23128 27160 23180
rect 27212 23168 27218 23180
rect 27341 23171 27399 23177
rect 27341 23168 27353 23171
rect 27212 23140 27353 23168
rect 27212 23128 27218 23140
rect 27341 23137 27353 23140
rect 27387 23137 27399 23171
rect 27341 23131 27399 23137
rect 27617 23171 27675 23177
rect 27617 23137 27629 23171
rect 27663 23168 27675 23171
rect 28902 23168 28908 23180
rect 27663 23140 28908 23168
rect 27663 23137 27675 23140
rect 27617 23131 27675 23137
rect 28902 23128 28908 23140
rect 28960 23128 28966 23180
rect 30009 23171 30067 23177
rect 30009 23137 30021 23171
rect 30055 23168 30067 23171
rect 32324 23168 32352 23208
rect 33410 23196 33416 23248
rect 33468 23236 33474 23248
rect 34057 23239 34115 23245
rect 34057 23236 34069 23239
rect 33468 23208 34069 23236
rect 33468 23196 33474 23208
rect 34057 23205 34069 23208
rect 34103 23205 34115 23239
rect 34057 23199 34115 23205
rect 36354 23196 36360 23248
rect 36412 23236 36418 23248
rect 36412 23208 37872 23236
rect 36412 23196 36418 23208
rect 30055 23140 32352 23168
rect 30055 23137 30067 23140
rect 30009 23131 30067 23137
rect 32490 23128 32496 23180
rect 32548 23168 32554 23180
rect 37090 23168 37096 23180
rect 32548 23140 37096 23168
rect 32548 23128 32554 23140
rect 37090 23128 37096 23140
rect 37148 23168 37154 23180
rect 37737 23171 37795 23177
rect 37737 23168 37749 23171
rect 37148 23140 37749 23168
rect 37148 23128 37154 23140
rect 37737 23137 37749 23140
rect 37783 23137 37795 23171
rect 37844 23168 37872 23208
rect 39574 23196 39580 23248
rect 39632 23236 39638 23248
rect 41230 23236 41236 23248
rect 39632 23208 41236 23236
rect 39632 23196 39638 23208
rect 41230 23196 41236 23208
rect 41288 23196 41294 23248
rect 42812 23236 42840 23276
rect 43162 23264 43168 23276
rect 43220 23264 43226 23316
rect 43438 23264 43444 23316
rect 43496 23304 43502 23316
rect 43993 23307 44051 23313
rect 43993 23304 44005 23307
rect 43496 23276 44005 23304
rect 43496 23264 43502 23276
rect 43993 23273 44005 23276
rect 44039 23273 44051 23307
rect 43993 23267 44051 23273
rect 44358 23264 44364 23316
rect 44416 23304 44422 23316
rect 44453 23307 44511 23313
rect 44453 23304 44465 23307
rect 44416 23276 44465 23304
rect 44416 23264 44422 23276
rect 44453 23273 44465 23276
rect 44499 23273 44511 23307
rect 44453 23267 44511 23273
rect 46658 23264 46664 23316
rect 46716 23304 46722 23316
rect 48866 23304 48872 23316
rect 46716 23276 48872 23304
rect 46716 23264 46722 23276
rect 48866 23264 48872 23276
rect 48924 23264 48930 23316
rect 49326 23264 49332 23316
rect 49384 23264 49390 23316
rect 41386 23208 42840 23236
rect 42889 23239 42947 23245
rect 41386 23168 41414 23208
rect 42889 23205 42901 23239
rect 42935 23236 42947 23239
rect 43622 23236 43628 23248
rect 42935 23208 43628 23236
rect 42935 23205 42947 23208
rect 42889 23199 42947 23205
rect 43622 23196 43628 23208
rect 43680 23196 43686 23248
rect 46106 23196 46112 23248
rect 46164 23196 46170 23248
rect 48498 23236 48504 23248
rect 46400 23208 48504 23236
rect 44542 23168 44548 23180
rect 37844 23140 41414 23168
rect 42260 23140 44548 23168
rect 37737 23131 37795 23137
rect 26620 23072 27108 23100
rect 26237 23063 26295 23069
rect 26694 23032 26700 23044
rect 26068 23004 26700 23032
rect 26694 22992 26700 23004
rect 26752 22992 26758 23044
rect 24581 22967 24639 22973
rect 24581 22933 24593 22967
rect 24627 22933 24639 22967
rect 24581 22927 24639 22933
rect 25041 22967 25099 22973
rect 25041 22933 25053 22967
rect 25087 22964 25099 22967
rect 25498 22964 25504 22976
rect 25087 22936 25504 22964
rect 25087 22933 25099 22936
rect 25041 22927 25099 22933
rect 25498 22924 25504 22936
rect 25556 22924 25562 22976
rect 25590 22924 25596 22976
rect 25648 22964 25654 22976
rect 25777 22967 25835 22973
rect 25777 22964 25789 22967
rect 25648 22936 25789 22964
rect 25648 22924 25654 22936
rect 25777 22933 25789 22936
rect 25823 22933 25835 22967
rect 25777 22927 25835 22933
rect 25866 22924 25872 22976
rect 25924 22964 25930 22976
rect 26050 22964 26056 22976
rect 25924 22936 26056 22964
rect 25924 22924 25930 22936
rect 26050 22924 26056 22936
rect 26108 22964 26114 22976
rect 26145 22967 26203 22973
rect 26145 22964 26157 22967
rect 26108 22936 26157 22964
rect 26108 22924 26114 22936
rect 26145 22933 26157 22936
rect 26191 22964 26203 22967
rect 26878 22964 26884 22976
rect 26191 22936 26884 22964
rect 26191 22933 26203 22936
rect 26145 22927 26203 22933
rect 26878 22924 26884 22936
rect 26936 22964 26942 22976
rect 26973 22967 27031 22973
rect 26973 22964 26985 22967
rect 26936 22936 26985 22964
rect 26936 22924 26942 22936
rect 26973 22933 26985 22936
rect 27019 22933 27031 22967
rect 27080 22964 27108 23072
rect 29270 23060 29276 23112
rect 29328 23100 29334 23112
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29328 23072 29745 23100
rect 29328 23060 29334 23072
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 31386 23060 31392 23112
rect 31444 23100 31450 23112
rect 32309 23103 32367 23109
rect 32309 23100 32321 23103
rect 31444 23072 32321 23100
rect 31444 23060 31450 23072
rect 32309 23069 32321 23072
rect 32355 23069 32367 23103
rect 32309 23063 32367 23069
rect 33134 23060 33140 23112
rect 33192 23100 33198 23112
rect 33413 23103 33471 23109
rect 33413 23100 33425 23103
rect 33192 23072 33425 23100
rect 33192 23060 33198 23072
rect 33413 23069 33425 23072
rect 33459 23069 33471 23103
rect 34885 23103 34943 23109
rect 34885 23100 34897 23103
rect 33413 23063 33471 23069
rect 33520 23072 34897 23100
rect 27706 22992 27712 23044
rect 27764 23032 27770 23044
rect 27764 23004 28106 23032
rect 27764 22992 27770 23004
rect 28994 22992 29000 23044
rect 29052 23032 29058 23044
rect 29638 23032 29644 23044
rect 29052 23004 29644 23032
rect 29052 22992 29058 23004
rect 29638 22992 29644 23004
rect 29696 22992 29702 23044
rect 30098 22992 30104 23044
rect 30156 23032 30162 23044
rect 33520 23032 33548 23072
rect 34885 23069 34897 23072
rect 34931 23069 34943 23103
rect 34885 23063 34943 23069
rect 35986 23060 35992 23112
rect 36044 23060 36050 23112
rect 36814 23060 36820 23112
rect 36872 23100 36878 23112
rect 37277 23103 37335 23109
rect 37277 23100 37289 23103
rect 36872 23072 37289 23100
rect 36872 23060 36878 23072
rect 37277 23069 37289 23072
rect 37323 23069 37335 23103
rect 37277 23063 37335 23069
rect 40034 23060 40040 23112
rect 40092 23060 40098 23112
rect 41138 23060 41144 23112
rect 41196 23060 41202 23112
rect 42260 23109 42288 23140
rect 44542 23128 44548 23140
rect 44600 23128 44606 23180
rect 42245 23103 42303 23109
rect 42245 23069 42257 23103
rect 42291 23069 42303 23103
rect 42245 23063 42303 23069
rect 43349 23103 43407 23109
rect 43349 23069 43361 23103
rect 43395 23100 43407 23103
rect 44174 23100 44180 23112
rect 43395 23072 44180 23100
rect 43395 23069 43407 23072
rect 43349 23063 43407 23069
rect 44174 23060 44180 23072
rect 44232 23060 44238 23112
rect 44634 23060 44640 23112
rect 44692 23060 44698 23112
rect 45189 23103 45247 23109
rect 45189 23069 45201 23103
rect 45235 23100 45247 23103
rect 46400 23100 46428 23208
rect 48498 23196 48504 23208
rect 48556 23196 48562 23248
rect 48225 23171 48283 23177
rect 48225 23168 48237 23171
rect 46492 23140 48237 23168
rect 46492 23109 46520 23140
rect 48225 23137 48237 23140
rect 48271 23137 48283 23171
rect 48225 23131 48283 23137
rect 45235 23072 46428 23100
rect 46477 23103 46535 23109
rect 45235 23069 45247 23072
rect 45189 23063 45247 23069
rect 46477 23069 46489 23103
rect 46523 23069 46535 23103
rect 46477 23063 46535 23069
rect 47581 23103 47639 23109
rect 47581 23069 47593 23103
rect 47627 23100 47639 23103
rect 48498 23100 48504 23112
rect 47627 23072 48504 23100
rect 47627 23069 47639 23072
rect 47581 23063 47639 23069
rect 48498 23060 48504 23072
rect 48556 23060 48562 23112
rect 48685 23103 48743 23109
rect 48685 23069 48697 23103
rect 48731 23100 48743 23103
rect 49326 23100 49332 23112
rect 48731 23072 49332 23100
rect 48731 23069 48743 23072
rect 48685 23063 48743 23069
rect 49326 23060 49332 23072
rect 49384 23060 49390 23112
rect 30156 23004 30498 23032
rect 31312 23004 33548 23032
rect 30156 22992 30162 23004
rect 29730 22964 29736 22976
rect 27080 22936 29736 22964
rect 26973 22927 27031 22933
rect 29730 22924 29736 22936
rect 29788 22924 29794 22976
rect 30190 22924 30196 22976
rect 30248 22964 30254 22976
rect 31312 22964 31340 23004
rect 33962 22992 33968 23044
rect 34020 23032 34026 23044
rect 35529 23035 35587 23041
rect 35529 23032 35541 23035
rect 34020 23004 35541 23032
rect 34020 22992 34026 23004
rect 35529 23001 35541 23004
rect 35575 23001 35587 23035
rect 38013 23035 38071 23041
rect 35529 22995 35587 23001
rect 35636 23004 37228 23032
rect 30248 22936 31340 22964
rect 31481 22967 31539 22973
rect 30248 22924 30254 22936
rect 31481 22933 31493 22967
rect 31527 22964 31539 22967
rect 31570 22964 31576 22976
rect 31527 22936 31576 22964
rect 31527 22933 31539 22936
rect 31481 22927 31539 22933
rect 31570 22924 31576 22936
rect 31628 22924 31634 22976
rect 31849 22967 31907 22973
rect 31849 22933 31861 22967
rect 31895 22964 31907 22967
rect 31938 22964 31944 22976
rect 31895 22936 31944 22964
rect 31895 22933 31907 22936
rect 31849 22927 31907 22933
rect 31938 22924 31944 22936
rect 31996 22964 32002 22976
rect 33042 22964 33048 22976
rect 31996 22936 33048 22964
rect 31996 22924 32002 22936
rect 33042 22924 33048 22936
rect 33100 22924 33106 22976
rect 33502 22924 33508 22976
rect 33560 22964 33566 22976
rect 34333 22967 34391 22973
rect 34333 22964 34345 22967
rect 33560 22936 34345 22964
rect 33560 22924 33566 22936
rect 34333 22933 34345 22936
rect 34379 22933 34391 22967
rect 34333 22927 34391 22933
rect 34790 22924 34796 22976
rect 34848 22964 34854 22976
rect 35636 22964 35664 23004
rect 34848 22936 35664 22964
rect 34848 22924 34854 22936
rect 37090 22924 37096 22976
rect 37148 22924 37154 22976
rect 37200 22964 37228 23004
rect 38013 23001 38025 23035
rect 38059 23032 38071 23035
rect 38286 23032 38292 23044
rect 38059 23004 38292 23032
rect 38059 23001 38071 23004
rect 38013 22995 38071 23001
rect 38286 22992 38292 23004
rect 38344 22992 38350 23044
rect 40310 23032 40316 23044
rect 39238 23004 40316 23032
rect 39316 22964 39344 23004
rect 40310 22992 40316 23004
rect 40368 23032 40374 23044
rect 42794 23032 42800 23044
rect 40368 23004 42800 23032
rect 40368 22992 40374 23004
rect 42794 22992 42800 23004
rect 42852 22992 42858 23044
rect 37200 22936 39344 22964
rect 39482 22924 39488 22976
rect 39540 22924 39546 22976
rect 39758 22924 39764 22976
rect 39816 22964 39822 22976
rect 41046 22964 41052 22976
rect 39816 22936 41052 22964
rect 39816 22924 39822 22936
rect 41046 22924 41052 22936
rect 41104 22924 41110 22976
rect 45830 22924 45836 22976
rect 45888 22924 45894 22976
rect 47121 22967 47179 22973
rect 47121 22933 47133 22967
rect 47167 22964 47179 22967
rect 47210 22964 47216 22976
rect 47167 22936 47216 22964
rect 47167 22933 47179 22936
rect 47121 22927 47179 22933
rect 47210 22924 47216 22936
rect 47268 22924 47274 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 3881 22763 3939 22769
rect 3881 22729 3893 22763
rect 3927 22760 3939 22763
rect 4341 22763 4399 22769
rect 4341 22760 4353 22763
rect 3927 22732 4353 22760
rect 3927 22729 3939 22732
rect 3881 22723 3939 22729
rect 4341 22729 4353 22732
rect 4387 22760 4399 22763
rect 4522 22760 4528 22772
rect 4387 22732 4528 22760
rect 4387 22729 4399 22732
rect 4341 22723 4399 22729
rect 4522 22720 4528 22732
rect 4580 22720 4586 22772
rect 6656 22732 18552 22760
rect 6656 22701 6684 22732
rect 6641 22695 6699 22701
rect 2746 22664 4660 22692
rect 1765 22627 1823 22633
rect 1765 22593 1777 22627
rect 1811 22624 1823 22627
rect 2038 22624 2044 22636
rect 1811 22596 2044 22624
rect 1811 22593 1823 22596
rect 1765 22587 1823 22593
rect 2038 22584 2044 22596
rect 2096 22584 2102 22636
rect 2746 22624 2774 22664
rect 4632 22633 4660 22664
rect 6641 22661 6653 22695
rect 6687 22661 6699 22695
rect 6641 22655 6699 22661
rect 8570 22652 8576 22704
rect 8628 22652 8634 22704
rect 9493 22695 9551 22701
rect 9493 22692 9505 22695
rect 8772 22664 9505 22692
rect 2148 22596 2774 22624
rect 3329 22627 3387 22633
rect 382 22516 388 22568
rect 440 22556 446 22568
rect 2148 22556 2176 22596
rect 3329 22593 3341 22627
rect 3375 22624 3387 22627
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3375 22596 3801 22624
rect 3375 22593 3387 22596
rect 3329 22587 3387 22593
rect 3789 22593 3801 22596
rect 3835 22624 3847 22627
rect 4617 22627 4675 22633
rect 3835 22596 4568 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 440 22528 2176 22556
rect 440 22516 446 22528
rect 2222 22516 2228 22568
rect 2280 22516 2286 22568
rect 4062 22516 4068 22568
rect 4120 22516 4126 22568
rect 3418 22380 3424 22432
rect 3476 22380 3482 22432
rect 4540 22420 4568 22596
rect 4617 22593 4629 22627
rect 4663 22593 4675 22627
rect 4617 22587 4675 22593
rect 7558 22584 7564 22636
rect 7616 22584 7622 22636
rect 7742 22584 7748 22636
rect 7800 22624 7806 22636
rect 8772 22624 8800 22664
rect 9493 22661 9505 22664
rect 9539 22661 9551 22695
rect 10778 22692 10784 22704
rect 10718 22664 10784 22692
rect 9493 22655 9551 22661
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 11974 22652 11980 22704
rect 12032 22652 12038 22704
rect 12526 22652 12532 22704
rect 12584 22652 12590 22704
rect 12986 22652 12992 22704
rect 13044 22652 13050 22704
rect 14461 22695 14519 22701
rect 14461 22661 14473 22695
rect 14507 22692 14519 22695
rect 14507 22664 16068 22692
rect 14507 22661 14519 22664
rect 14461 22655 14519 22661
rect 7800 22596 8800 22624
rect 7800 22584 7806 22596
rect 11146 22584 11152 22636
rect 11204 22624 11210 22636
rect 12250 22624 12256 22636
rect 11204 22596 12256 22624
rect 11204 22584 11210 22596
rect 12250 22584 12256 22596
rect 12308 22584 12314 22636
rect 14550 22584 14556 22636
rect 14608 22624 14614 22636
rect 14826 22624 14832 22636
rect 14608 22596 14832 22624
rect 14608 22584 14614 22596
rect 14826 22584 14832 22596
rect 14884 22584 14890 22636
rect 14918 22584 14924 22636
rect 14976 22584 14982 22636
rect 16040 22624 16068 22664
rect 16114 22652 16120 22704
rect 16172 22652 16178 22704
rect 17129 22695 17187 22701
rect 17129 22661 17141 22695
rect 17175 22692 17187 22695
rect 17218 22692 17224 22704
rect 17175 22664 17224 22692
rect 17175 22661 17187 22664
rect 17129 22655 17187 22661
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 18414 22692 18420 22704
rect 18354 22664 18420 22692
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 16574 22624 16580 22636
rect 16040 22596 16580 22624
rect 16574 22584 16580 22596
rect 16632 22584 16638 22636
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 6638 22516 6644 22568
rect 6696 22556 6702 22568
rect 6825 22559 6883 22565
rect 6825 22556 6837 22559
rect 6696 22528 6837 22556
rect 6696 22516 6702 22528
rect 6825 22525 6837 22528
rect 6871 22525 6883 22559
rect 6825 22519 6883 22525
rect 8662 22516 8668 22568
rect 8720 22556 8726 22568
rect 9217 22559 9275 22565
rect 9217 22556 9229 22559
rect 8720 22528 9229 22556
rect 8720 22516 8726 22528
rect 9217 22525 9229 22528
rect 9263 22525 9275 22559
rect 15470 22556 15476 22568
rect 9217 22519 9275 22525
rect 9324 22528 15476 22556
rect 5994 22448 6000 22500
rect 6052 22488 6058 22500
rect 9324 22488 9352 22528
rect 15470 22516 15476 22528
rect 15528 22516 15534 22568
rect 16850 22516 16856 22568
rect 16908 22516 16914 22568
rect 6052 22460 9352 22488
rect 11609 22491 11667 22497
rect 6052 22448 6058 22460
rect 11609 22457 11621 22491
rect 11655 22488 11667 22491
rect 16114 22488 16120 22500
rect 11655 22460 12020 22488
rect 11655 22457 11667 22460
rect 11609 22451 11667 22457
rect 8386 22420 8392 22432
rect 4540 22392 8392 22420
rect 8386 22380 8392 22392
rect 8444 22380 8450 22432
rect 9950 22380 9956 22432
rect 10008 22420 10014 22432
rect 10965 22423 11023 22429
rect 10965 22420 10977 22423
rect 10008 22392 10977 22420
rect 10008 22380 10014 22392
rect 10965 22389 10977 22392
rect 11011 22389 11023 22423
rect 10965 22383 11023 22389
rect 11330 22380 11336 22432
rect 11388 22380 11394 22432
rect 11422 22380 11428 22432
rect 11480 22420 11486 22432
rect 11701 22423 11759 22429
rect 11701 22420 11713 22423
rect 11480 22392 11713 22420
rect 11480 22380 11486 22392
rect 11701 22389 11713 22392
rect 11747 22389 11759 22423
rect 11992 22420 12020 22460
rect 13924 22460 16120 22488
rect 13924 22420 13952 22460
rect 16114 22448 16120 22460
rect 16172 22448 16178 22500
rect 18524 22488 18552 22732
rect 18598 22720 18604 22772
rect 18656 22760 18662 22772
rect 25317 22763 25375 22769
rect 25317 22760 25329 22763
rect 18656 22732 25329 22760
rect 18656 22720 18662 22732
rect 25317 22729 25329 22732
rect 25363 22729 25375 22763
rect 29362 22760 29368 22772
rect 25317 22723 25375 22729
rect 25424 22732 29368 22760
rect 19981 22695 20039 22701
rect 19981 22661 19993 22695
rect 20027 22692 20039 22695
rect 20070 22692 20076 22704
rect 20027 22664 20076 22692
rect 20027 22661 20039 22664
rect 19981 22655 20039 22661
rect 20070 22652 20076 22664
rect 20128 22652 20134 22704
rect 20622 22652 20628 22704
rect 20680 22652 20686 22704
rect 23382 22692 23388 22704
rect 23124 22664 23388 22692
rect 22005 22627 22063 22633
rect 22005 22593 22017 22627
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 19061 22559 19119 22565
rect 19061 22525 19073 22559
rect 19107 22556 19119 22559
rect 19610 22556 19616 22568
rect 19107 22528 19616 22556
rect 19107 22525 19119 22528
rect 19061 22519 19119 22525
rect 19610 22516 19616 22528
rect 19668 22516 19674 22568
rect 19702 22516 19708 22568
rect 19760 22516 19766 22568
rect 20990 22556 20996 22568
rect 19812 22528 20996 22556
rect 19812 22488 19840 22528
rect 20990 22516 20996 22528
rect 21048 22556 21054 22568
rect 21453 22559 21511 22565
rect 21453 22556 21465 22559
rect 21048 22528 21465 22556
rect 21048 22516 21054 22528
rect 21453 22525 21465 22528
rect 21499 22525 21511 22559
rect 22020 22556 22048 22587
rect 22278 22584 22284 22636
rect 22336 22624 22342 22636
rect 23124 22633 23152 22664
rect 23382 22652 23388 22664
rect 23440 22652 23446 22704
rect 23658 22652 23664 22704
rect 23716 22692 23722 22704
rect 23716 22664 23874 22692
rect 23716 22652 23722 22664
rect 25222 22652 25228 22704
rect 25280 22692 25286 22704
rect 25424 22692 25452 22732
rect 29362 22720 29368 22732
rect 29420 22720 29426 22772
rect 29454 22720 29460 22772
rect 29512 22760 29518 22772
rect 30006 22760 30012 22772
rect 29512 22732 30012 22760
rect 29512 22720 29518 22732
rect 30006 22720 30012 22732
rect 30064 22720 30070 22772
rect 31386 22760 31392 22772
rect 30208 22732 31392 22760
rect 25280 22664 25452 22692
rect 25516 22664 26464 22692
rect 25280 22652 25286 22664
rect 23109 22627 23167 22633
rect 23109 22624 23121 22627
rect 22336 22596 23121 22624
rect 22336 22584 22342 22596
rect 23109 22593 23121 22596
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 24762 22584 24768 22636
rect 24820 22584 24826 22636
rect 25130 22584 25136 22636
rect 25188 22624 25194 22636
rect 25516 22624 25544 22664
rect 25188 22596 25544 22624
rect 25685 22627 25743 22633
rect 25188 22584 25194 22596
rect 25685 22593 25697 22627
rect 25731 22624 25743 22627
rect 26436 22624 26464 22664
rect 27154 22652 27160 22704
rect 27212 22692 27218 22704
rect 27212 22664 28488 22692
rect 27212 22652 27218 22664
rect 28460 22636 28488 22664
rect 28718 22652 28724 22704
rect 28776 22652 28782 22704
rect 30098 22692 30104 22704
rect 29946 22664 30104 22692
rect 30098 22652 30104 22664
rect 30156 22652 30162 22704
rect 25731 22596 26372 22624
rect 26436 22596 27384 22624
rect 25731 22593 25743 22596
rect 25685 22587 25743 22593
rect 23385 22559 23443 22565
rect 22020 22528 23244 22556
rect 21453 22519 21511 22525
rect 18524 22460 19840 22488
rect 11992 22392 13952 22420
rect 11701 22383 11759 22389
rect 13998 22380 14004 22432
rect 14056 22380 14062 22432
rect 14645 22423 14703 22429
rect 14645 22389 14657 22423
rect 14691 22420 14703 22423
rect 14826 22420 14832 22432
rect 14691 22392 14832 22420
rect 14691 22389 14703 22392
rect 14645 22383 14703 22389
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 18601 22423 18659 22429
rect 18601 22389 18613 22423
rect 18647 22420 18659 22423
rect 20346 22420 20352 22432
rect 18647 22392 20352 22420
rect 18647 22389 18659 22392
rect 18601 22383 18659 22389
rect 20346 22380 20352 22392
rect 20404 22380 20410 22432
rect 22646 22380 22652 22432
rect 22704 22380 22710 22432
rect 23216 22420 23244 22528
rect 23385 22525 23397 22559
rect 23431 22556 23443 22559
rect 23474 22556 23480 22568
rect 23431 22528 23480 22556
rect 23431 22525 23443 22528
rect 23385 22519 23443 22525
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 23934 22516 23940 22568
rect 23992 22556 23998 22568
rect 24118 22556 24124 22568
rect 23992 22528 24124 22556
rect 23992 22516 23998 22528
rect 24118 22516 24124 22528
rect 24176 22516 24182 22568
rect 24670 22420 24676 22432
rect 23216 22392 24676 22420
rect 24670 22380 24676 22392
rect 24728 22380 24734 22432
rect 24780 22420 24808 22584
rect 25774 22516 25780 22568
rect 25832 22516 25838 22568
rect 25958 22516 25964 22568
rect 26016 22516 26022 22568
rect 26344 22565 26372 22596
rect 26329 22559 26387 22565
rect 26329 22525 26341 22559
rect 26375 22556 26387 22559
rect 27154 22556 27160 22568
rect 26375 22528 27160 22556
rect 26375 22525 26387 22528
rect 26329 22519 26387 22525
rect 27154 22516 27160 22528
rect 27212 22516 27218 22568
rect 24857 22491 24915 22497
rect 24857 22457 24869 22491
rect 24903 22488 24915 22491
rect 25976 22488 26004 22516
rect 27249 22491 27307 22497
rect 27249 22488 27261 22491
rect 24903 22460 26004 22488
rect 26344 22460 27261 22488
rect 24903 22457 24915 22460
rect 24857 22451 24915 22457
rect 26344 22432 26372 22460
rect 27249 22457 27261 22460
rect 27295 22457 27307 22491
rect 27249 22451 27307 22457
rect 25866 22420 25872 22432
rect 24780 22392 25872 22420
rect 25866 22380 25872 22392
rect 25924 22380 25930 22432
rect 26326 22380 26332 22432
rect 26384 22380 26390 22432
rect 26605 22423 26663 22429
rect 26605 22389 26617 22423
rect 26651 22420 26663 22423
rect 26789 22423 26847 22429
rect 26789 22420 26801 22423
rect 26651 22392 26801 22420
rect 26651 22389 26663 22392
rect 26605 22383 26663 22389
rect 26789 22389 26801 22392
rect 26835 22420 26847 22423
rect 26878 22420 26884 22432
rect 26835 22392 26884 22420
rect 26835 22389 26847 22392
rect 26789 22383 26847 22389
rect 26878 22380 26884 22392
rect 26936 22380 26942 22432
rect 27356 22420 27384 22596
rect 27614 22584 27620 22636
rect 27672 22584 27678 22636
rect 28442 22584 28448 22636
rect 28500 22584 28506 22636
rect 27706 22516 27712 22568
rect 27764 22516 27770 22568
rect 27893 22559 27951 22565
rect 27893 22525 27905 22559
rect 27939 22556 27951 22559
rect 30208 22556 30236 22732
rect 31386 22720 31392 22732
rect 31444 22720 31450 22772
rect 31754 22720 31760 22772
rect 31812 22760 31818 22772
rect 31941 22763 31999 22769
rect 31941 22760 31953 22763
rect 31812 22732 31953 22760
rect 31812 22720 31818 22732
rect 31941 22729 31953 22732
rect 31987 22760 31999 22763
rect 32490 22760 32496 22772
rect 31987 22732 32496 22760
rect 31987 22729 31999 22732
rect 31941 22723 31999 22729
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 34330 22720 34336 22772
rect 34388 22720 34394 22772
rect 35434 22720 35440 22772
rect 35492 22760 35498 22772
rect 35529 22763 35587 22769
rect 35529 22760 35541 22763
rect 35492 22732 35541 22760
rect 35492 22720 35498 22732
rect 35529 22729 35541 22732
rect 35575 22729 35587 22763
rect 35529 22723 35587 22729
rect 35894 22720 35900 22772
rect 35952 22760 35958 22772
rect 36633 22763 36691 22769
rect 36633 22760 36645 22763
rect 35952 22732 36645 22760
rect 35952 22720 35958 22732
rect 36633 22729 36645 22732
rect 36679 22729 36691 22763
rect 36633 22723 36691 22729
rect 36814 22720 36820 22772
rect 36872 22760 36878 22772
rect 36909 22763 36967 22769
rect 36909 22760 36921 22763
rect 36872 22732 36921 22760
rect 36872 22720 36878 22732
rect 36909 22729 36921 22732
rect 36955 22729 36967 22763
rect 36909 22723 36967 22729
rect 37366 22720 37372 22772
rect 37424 22760 37430 22772
rect 38105 22763 38163 22769
rect 38105 22760 38117 22763
rect 37424 22732 38117 22760
rect 37424 22720 37430 22732
rect 38105 22729 38117 22732
rect 38151 22729 38163 22763
rect 38105 22723 38163 22729
rect 38930 22720 38936 22772
rect 38988 22760 38994 22772
rect 40494 22760 40500 22772
rect 38988 22732 40500 22760
rect 38988 22720 38994 22732
rect 40494 22720 40500 22732
rect 40552 22720 40558 22772
rect 41417 22763 41475 22769
rect 41417 22729 41429 22763
rect 41463 22760 41475 22763
rect 43898 22760 43904 22772
rect 41463 22732 43904 22760
rect 41463 22729 41475 22732
rect 41417 22723 41475 22729
rect 43898 22720 43904 22732
rect 43956 22720 43962 22772
rect 47213 22763 47271 22769
rect 47213 22760 47225 22763
rect 44652 22732 47225 22760
rect 44652 22704 44680 22732
rect 47213 22729 47225 22732
rect 47259 22729 47271 22763
rect 47213 22723 47271 22729
rect 31113 22695 31171 22701
rect 31113 22661 31125 22695
rect 31159 22692 31171 22695
rect 31202 22692 31208 22704
rect 31159 22664 31208 22692
rect 31159 22661 31171 22664
rect 31113 22655 31171 22661
rect 31202 22652 31208 22664
rect 31260 22652 31266 22704
rect 31294 22652 31300 22704
rect 31352 22692 31358 22704
rect 44634 22692 44640 22704
rect 31352 22664 44640 22692
rect 31352 22652 31358 22664
rect 44634 22652 44640 22664
rect 44692 22652 44698 22704
rect 45370 22652 45376 22704
rect 45428 22692 45434 22704
rect 45428 22664 46520 22692
rect 45428 22652 45434 22664
rect 46492 22636 46520 22664
rect 46934 22652 46940 22704
rect 46992 22692 46998 22704
rect 47029 22695 47087 22701
rect 47029 22692 47041 22695
rect 46992 22664 47041 22692
rect 46992 22652 46998 22664
rect 47029 22661 47041 22664
rect 47075 22661 47087 22695
rect 47029 22655 47087 22661
rect 47302 22652 47308 22704
rect 47360 22692 47366 22704
rect 47857 22695 47915 22701
rect 47857 22692 47869 22695
rect 47360 22664 47869 22692
rect 47360 22652 47366 22664
rect 47857 22661 47869 22664
rect 47903 22661 47915 22695
rect 47857 22655 47915 22661
rect 31021 22627 31079 22633
rect 31021 22593 31033 22627
rect 31067 22624 31079 22627
rect 31478 22624 31484 22636
rect 31067 22596 31484 22624
rect 31067 22593 31079 22596
rect 31021 22587 31079 22593
rect 31478 22584 31484 22596
rect 31536 22584 31542 22636
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 33318 22624 33324 22636
rect 32355 22596 33324 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 33318 22584 33324 22596
rect 33376 22584 33382 22636
rect 33413 22627 33471 22633
rect 33413 22593 33425 22627
rect 33459 22624 33471 22627
rect 33962 22624 33968 22636
rect 33459 22596 33968 22624
rect 33459 22593 33471 22596
rect 33413 22587 33471 22593
rect 33962 22584 33968 22596
rect 34020 22584 34026 22636
rect 34057 22627 34115 22633
rect 34057 22593 34069 22627
rect 34103 22624 34115 22627
rect 34885 22627 34943 22633
rect 34885 22624 34897 22627
rect 34103 22596 34897 22624
rect 34103 22593 34115 22596
rect 34057 22587 34115 22593
rect 34885 22593 34897 22596
rect 34931 22593 34943 22627
rect 34885 22587 34943 22593
rect 35989 22627 36047 22633
rect 35989 22593 36001 22627
rect 36035 22624 36047 22627
rect 37182 22624 37188 22636
rect 36035 22596 37188 22624
rect 36035 22593 36047 22596
rect 35989 22587 36047 22593
rect 37182 22584 37188 22596
rect 37240 22584 37246 22636
rect 37458 22584 37464 22636
rect 37516 22584 37522 22636
rect 38562 22584 38568 22636
rect 38620 22584 38626 22636
rect 39206 22584 39212 22636
rect 39264 22584 39270 22636
rect 39666 22584 39672 22636
rect 39724 22584 39730 22636
rect 40773 22627 40831 22633
rect 40773 22624 40785 22627
rect 40144 22596 40785 22624
rect 27939 22528 30236 22556
rect 31297 22559 31355 22565
rect 27939 22525 27951 22528
rect 27893 22519 27951 22525
rect 31297 22525 31309 22559
rect 31343 22556 31355 22559
rect 31570 22556 31576 22568
rect 31343 22528 31576 22556
rect 31343 22525 31355 22528
rect 31297 22519 31355 22525
rect 27522 22448 27528 22500
rect 27580 22488 27586 22500
rect 27908 22488 27936 22519
rect 31570 22516 31576 22528
rect 31628 22556 31634 22568
rect 40034 22556 40040 22568
rect 31628 22528 40040 22556
rect 31628 22516 31634 22528
rect 40034 22516 40040 22528
rect 40092 22516 40098 22568
rect 27580 22460 27936 22488
rect 27580 22448 27586 22460
rect 29730 22448 29736 22500
rect 29788 22488 29794 22500
rect 32953 22491 33011 22497
rect 32953 22488 32965 22491
rect 29788 22460 32965 22488
rect 29788 22448 29794 22460
rect 32953 22457 32965 22460
rect 32999 22457 33011 22491
rect 32953 22451 33011 22457
rect 33042 22448 33048 22500
rect 33100 22488 33106 22500
rect 34609 22491 34667 22497
rect 33100 22460 34468 22488
rect 33100 22448 33106 22460
rect 28902 22420 28908 22432
rect 27356 22392 28908 22420
rect 28902 22380 28908 22392
rect 28960 22380 28966 22432
rect 29914 22380 29920 22432
rect 29972 22420 29978 22432
rect 30190 22420 30196 22432
rect 29972 22392 30196 22420
rect 29972 22380 29978 22392
rect 30190 22380 30196 22392
rect 30248 22380 30254 22432
rect 30282 22380 30288 22432
rect 30340 22420 30346 22432
rect 30653 22423 30711 22429
rect 30653 22420 30665 22423
rect 30340 22392 30665 22420
rect 30340 22380 30346 22392
rect 30653 22389 30665 22392
rect 30699 22389 30711 22423
rect 30653 22383 30711 22389
rect 31754 22380 31760 22432
rect 31812 22420 31818 22432
rect 32490 22420 32496 22432
rect 31812 22392 32496 22420
rect 31812 22380 31818 22392
rect 32490 22380 32496 22392
rect 32548 22380 32554 22432
rect 34440 22420 34468 22460
rect 34609 22457 34621 22491
rect 34655 22488 34667 22491
rect 34790 22488 34796 22500
rect 34655 22460 34796 22488
rect 34655 22457 34667 22460
rect 34609 22451 34667 22457
rect 34790 22448 34796 22460
rect 34848 22448 34854 22500
rect 36998 22448 37004 22500
rect 37056 22488 37062 22500
rect 40144 22488 40172 22596
rect 40773 22593 40785 22596
rect 40819 22593 40831 22627
rect 40773 22587 40831 22593
rect 41046 22584 41052 22636
rect 41104 22624 41110 22636
rect 42889 22627 42947 22633
rect 42889 22624 42901 22627
rect 41104 22596 42901 22624
rect 41104 22584 41110 22596
rect 42889 22593 42901 22596
rect 42935 22593 42947 22627
rect 42889 22587 42947 22593
rect 43714 22584 43720 22636
rect 43772 22624 43778 22636
rect 43901 22627 43959 22633
rect 43901 22624 43913 22627
rect 43772 22596 43913 22624
rect 43772 22584 43778 22596
rect 43901 22593 43913 22596
rect 43947 22624 43959 22627
rect 44910 22624 44916 22636
rect 43947 22596 44916 22624
rect 43947 22593 43959 22596
rect 43901 22587 43959 22593
rect 44910 22584 44916 22596
rect 44968 22584 44974 22636
rect 45002 22584 45008 22636
rect 45060 22584 45066 22636
rect 45094 22584 45100 22636
rect 45152 22624 45158 22636
rect 45741 22627 45799 22633
rect 45741 22624 45753 22627
rect 45152 22596 45753 22624
rect 45152 22584 45158 22596
rect 45741 22593 45753 22596
rect 45787 22593 45799 22627
rect 45741 22587 45799 22593
rect 41874 22516 41880 22568
rect 41932 22516 41938 22568
rect 42613 22559 42671 22565
rect 42613 22525 42625 22559
rect 42659 22525 42671 22559
rect 42613 22519 42671 22525
rect 37056 22460 40172 22488
rect 42628 22488 42656 22519
rect 43162 22516 43168 22568
rect 43220 22556 43226 22568
rect 43990 22556 43996 22568
rect 43220 22528 43996 22556
rect 43220 22516 43226 22528
rect 43990 22516 43996 22528
rect 44048 22516 44054 22568
rect 45020 22556 45048 22584
rect 45646 22556 45652 22568
rect 45020 22528 45652 22556
rect 45646 22516 45652 22528
rect 45704 22516 45710 22568
rect 45756 22556 45784 22587
rect 46474 22584 46480 22636
rect 46532 22584 46538 22636
rect 48314 22584 48320 22636
rect 48372 22624 48378 22636
rect 48685 22627 48743 22633
rect 48685 22624 48697 22627
rect 48372 22596 48697 22624
rect 48372 22584 48378 22596
rect 48685 22593 48697 22596
rect 48731 22593 48743 22627
rect 48685 22587 48743 22593
rect 48409 22559 48467 22565
rect 48409 22556 48421 22559
rect 45756 22528 48421 22556
rect 48409 22525 48421 22528
rect 48455 22525 48467 22559
rect 48409 22519 48467 22525
rect 44358 22488 44364 22500
rect 42628 22460 44364 22488
rect 37056 22448 37062 22460
rect 44358 22448 44364 22460
rect 44416 22448 44422 22500
rect 44818 22448 44824 22500
rect 44876 22488 44882 22500
rect 45925 22491 45983 22497
rect 45925 22488 45937 22491
rect 44876 22460 45937 22488
rect 44876 22448 44882 22460
rect 45925 22457 45937 22460
rect 45971 22457 45983 22491
rect 45925 22451 45983 22457
rect 37016 22420 37044 22448
rect 34440 22392 37044 22420
rect 40126 22380 40132 22432
rect 40184 22420 40190 22432
rect 40313 22423 40371 22429
rect 40313 22420 40325 22423
rect 40184 22392 40325 22420
rect 40184 22380 40190 22392
rect 40313 22389 40325 22392
rect 40359 22389 40371 22423
rect 40313 22383 40371 22389
rect 40862 22380 40868 22432
rect 40920 22420 40926 22432
rect 43438 22420 43444 22432
rect 40920 22392 43444 22420
rect 40920 22380 40926 22392
rect 43438 22380 43444 22392
rect 43496 22380 43502 22432
rect 44542 22380 44548 22432
rect 44600 22380 44606 22432
rect 45186 22380 45192 22432
rect 45244 22380 45250 22432
rect 46658 22380 46664 22432
rect 46716 22380 46722 22432
rect 46934 22380 46940 22432
rect 46992 22420 46998 22432
rect 47949 22423 48007 22429
rect 47949 22420 47961 22423
rect 46992 22392 47961 22420
rect 46992 22380 46998 22392
rect 47949 22389 47961 22392
rect 47995 22389 48007 22423
rect 47949 22383 48007 22389
rect 48682 22380 48688 22432
rect 48740 22420 48746 22432
rect 49329 22423 49387 22429
rect 49329 22420 49341 22423
rect 48740 22392 49341 22420
rect 48740 22380 48746 22392
rect 49329 22389 49341 22392
rect 49375 22389 49387 22423
rect 49329 22383 49387 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 3326 22176 3332 22228
rect 3384 22216 3390 22228
rect 4338 22216 4344 22228
rect 3384 22188 4344 22216
rect 3384 22176 3390 22188
rect 4338 22176 4344 22188
rect 4396 22176 4402 22228
rect 4614 22176 4620 22228
rect 4672 22216 4678 22228
rect 14734 22216 14740 22228
rect 4672 22188 14740 22216
rect 4672 22176 4678 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 16298 22216 16304 22228
rect 14884 22188 16304 22216
rect 14884 22176 14890 22188
rect 16298 22176 16304 22188
rect 16356 22176 16362 22228
rect 16574 22176 16580 22228
rect 16632 22216 16638 22228
rect 17392 22219 17450 22225
rect 17392 22216 17404 22219
rect 16632 22188 17404 22216
rect 16632 22176 16638 22188
rect 17392 22185 17404 22188
rect 17438 22216 17450 22219
rect 17494 22216 17500 22228
rect 17438 22188 17500 22216
rect 17438 22185 17450 22188
rect 17392 22179 17450 22185
rect 17494 22176 17500 22188
rect 17552 22176 17558 22228
rect 17954 22176 17960 22228
rect 18012 22216 18018 22228
rect 19426 22216 19432 22228
rect 18012 22188 19432 22216
rect 18012 22176 18018 22188
rect 19426 22176 19432 22188
rect 19484 22176 19490 22228
rect 21266 22216 21272 22228
rect 19536 22188 21272 22216
rect 3970 22108 3976 22160
rect 4028 22148 4034 22160
rect 4246 22148 4252 22160
rect 4028 22120 4252 22148
rect 4028 22108 4034 22120
rect 4246 22108 4252 22120
rect 4304 22108 4310 22160
rect 11882 22148 11888 22160
rect 9784 22120 11888 22148
rect 1486 22040 1492 22092
rect 1544 22080 1550 22092
rect 2041 22083 2099 22089
rect 2041 22080 2053 22083
rect 1544 22052 2053 22080
rect 1544 22040 1550 22052
rect 2041 22049 2053 22052
rect 2087 22049 2099 22083
rect 2041 22043 2099 22049
rect 3326 22040 3332 22092
rect 3384 22080 3390 22092
rect 4433 22083 4491 22089
rect 4433 22080 4445 22083
rect 3384 22052 4445 22080
rect 3384 22040 3390 22052
rect 4433 22049 4445 22052
rect 4479 22049 4491 22083
rect 4433 22043 4491 22049
rect 7006 22040 7012 22092
rect 7064 22080 7070 22092
rect 9784 22089 9812 22120
rect 11882 22108 11888 22120
rect 11940 22108 11946 22160
rect 12710 22108 12716 22160
rect 12768 22148 12774 22160
rect 16758 22148 16764 22160
rect 12768 22120 16764 22148
rect 12768 22108 12774 22120
rect 16758 22108 16764 22120
rect 16816 22108 16822 22160
rect 19536 22148 19564 22188
rect 21266 22176 21272 22188
rect 21324 22176 21330 22228
rect 22646 22176 22652 22228
rect 22704 22216 22710 22228
rect 26034 22219 26092 22225
rect 26034 22216 26046 22219
rect 22704 22188 26046 22216
rect 22704 22176 22710 22188
rect 26034 22185 26046 22188
rect 26080 22185 26092 22219
rect 26034 22179 26092 22185
rect 26142 22176 26148 22228
rect 26200 22216 26206 22228
rect 26200 22188 27108 22216
rect 26200 22176 26206 22188
rect 18524 22120 19564 22148
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 7064 22052 7297 22080
rect 7064 22040 7070 22052
rect 7285 22049 7297 22052
rect 7331 22049 7343 22083
rect 7285 22043 7343 22049
rect 9769 22083 9827 22089
rect 9769 22049 9781 22083
rect 9815 22080 9827 22083
rect 9953 22083 10011 22089
rect 9815 22052 9849 22080
rect 9815 22049 9827 22052
rect 9769 22043 9827 22049
rect 9953 22049 9965 22083
rect 9999 22080 10011 22083
rect 10410 22080 10416 22092
rect 9999 22052 10416 22080
rect 9999 22049 10011 22052
rect 9953 22043 10011 22049
rect 10410 22040 10416 22052
rect 10468 22040 10474 22092
rect 11238 22040 11244 22092
rect 11296 22040 11302 22092
rect 13446 22040 13452 22092
rect 13504 22040 13510 22092
rect 13648 22052 14872 22080
rect 1578 21972 1584 22024
rect 1636 21972 1642 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 6089 22015 6147 22021
rect 6089 21981 6101 22015
rect 6135 21981 6147 22015
rect 6089 21975 6147 21981
rect 3421 21947 3479 21953
rect 3421 21913 3433 21947
rect 3467 21944 3479 21947
rect 5534 21944 5540 21956
rect 3467 21916 5540 21944
rect 3467 21913 3479 21916
rect 3421 21907 3479 21913
rect 5534 21904 5540 21916
rect 5592 21904 5598 21956
rect 6104 21944 6132 21975
rect 6914 21972 6920 22024
rect 6972 21972 6978 22024
rect 8573 22015 8631 22021
rect 8573 21981 8585 22015
rect 8619 22012 8631 22015
rect 8619 21984 10640 22012
rect 8619 21981 8631 21984
rect 8573 21975 8631 21981
rect 8386 21944 8392 21956
rect 6104 21916 8392 21944
rect 8386 21904 8392 21916
rect 8444 21904 8450 21956
rect 8680 21916 8984 21944
rect 3326 21836 3332 21888
rect 3384 21876 3390 21888
rect 3513 21879 3571 21885
rect 3513 21876 3525 21879
rect 3384 21848 3525 21876
rect 3384 21836 3390 21848
rect 3513 21845 3525 21848
rect 3559 21845 3571 21879
rect 3513 21839 3571 21845
rect 5810 21836 5816 21888
rect 5868 21836 5874 21888
rect 6273 21879 6331 21885
rect 6273 21845 6285 21879
rect 6319 21876 6331 21879
rect 6822 21876 6828 21888
rect 6319 21848 6828 21876
rect 6319 21845 6331 21848
rect 6273 21839 6331 21845
rect 6822 21836 6828 21848
rect 6880 21836 6886 21888
rect 7374 21836 7380 21888
rect 7432 21876 7438 21888
rect 8680 21876 8708 21916
rect 7432 21848 8708 21876
rect 7432 21836 7438 21848
rect 8754 21836 8760 21888
rect 8812 21836 8818 21888
rect 8956 21876 8984 21916
rect 9030 21904 9036 21956
rect 9088 21904 9094 21956
rect 10318 21944 10324 21956
rect 9232 21916 10324 21944
rect 9232 21876 9260 21916
rect 10318 21904 10324 21916
rect 10376 21904 10382 21956
rect 10612 21944 10640 21984
rect 10686 21972 10692 22024
rect 10744 21972 10750 22024
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 13538 21944 13544 21956
rect 10612 21916 13544 21944
rect 13538 21904 13544 21916
rect 13596 21904 13602 21956
rect 8956 21848 9260 21876
rect 9306 21836 9312 21888
rect 9364 21836 9370 21888
rect 9674 21836 9680 21888
rect 9732 21836 9738 21888
rect 11146 21836 11152 21888
rect 11204 21876 11210 21888
rect 13648 21876 13676 22052
rect 14274 21972 14280 22024
rect 14332 22012 14338 22024
rect 14553 22015 14611 22021
rect 14553 22012 14565 22015
rect 14332 21984 14565 22012
rect 14332 21972 14338 21984
rect 14553 21981 14565 21984
rect 14599 21981 14611 22015
rect 14553 21975 14611 21981
rect 14642 21972 14648 22024
rect 14700 22012 14706 22024
rect 14737 22015 14795 22021
rect 14737 22012 14749 22015
rect 14700 21984 14749 22012
rect 14700 21972 14706 21984
rect 14737 21981 14749 21984
rect 14783 21981 14795 22015
rect 14737 21975 14795 21981
rect 14844 21944 14872 22052
rect 15102 22040 15108 22092
rect 15160 22080 15166 22092
rect 15657 22083 15715 22089
rect 15657 22080 15669 22083
rect 15160 22052 15669 22080
rect 15160 22040 15166 22052
rect 15657 22049 15669 22052
rect 15703 22049 15715 22083
rect 15657 22043 15715 22049
rect 16850 22040 16856 22092
rect 16908 22080 16914 22092
rect 17129 22083 17187 22089
rect 17129 22080 17141 22083
rect 16908 22052 17141 22080
rect 16908 22040 16914 22052
rect 17129 22049 17141 22052
rect 17175 22080 17187 22083
rect 17494 22080 17500 22092
rect 17175 22052 17500 22080
rect 17175 22049 17187 22052
rect 17129 22043 17187 22049
rect 17494 22040 17500 22052
rect 17552 22040 17558 22092
rect 18046 22040 18052 22092
rect 18104 22080 18110 22092
rect 18524 22080 18552 22120
rect 19794 22108 19800 22160
rect 19852 22148 19858 22160
rect 22094 22148 22100 22160
rect 19852 22120 22100 22148
rect 19852 22108 19858 22120
rect 22094 22108 22100 22120
rect 22152 22108 22158 22160
rect 23106 22108 23112 22160
rect 23164 22148 23170 22160
rect 23293 22151 23351 22157
rect 23293 22148 23305 22151
rect 23164 22120 23305 22148
rect 23164 22108 23170 22120
rect 23293 22117 23305 22120
rect 23339 22117 23351 22151
rect 25682 22148 25688 22160
rect 23293 22111 23351 22117
rect 24044 22120 25688 22148
rect 18104 22052 18552 22080
rect 18104 22040 18110 22052
rect 15194 21972 15200 22024
rect 15252 21972 15258 22024
rect 18524 21998 18552 22052
rect 19610 22040 19616 22092
rect 19668 22080 19674 22092
rect 20070 22080 20076 22092
rect 19668 22052 20076 22080
rect 19668 22040 19674 22052
rect 20070 22040 20076 22052
rect 20128 22040 20134 22092
rect 20714 22040 20720 22092
rect 20772 22080 20778 22092
rect 20809 22083 20867 22089
rect 20809 22080 20821 22083
rect 20772 22052 20821 22080
rect 20772 22040 20778 22052
rect 20809 22049 20821 22052
rect 20855 22049 20867 22083
rect 20809 22043 20867 22049
rect 21450 22040 21456 22092
rect 21508 22080 21514 22092
rect 22646 22080 22652 22092
rect 21508 22052 22652 22080
rect 21508 22040 21514 22052
rect 22646 22040 22652 22052
rect 22704 22040 22710 22092
rect 22738 22040 22744 22092
rect 22796 22080 22802 22092
rect 22833 22083 22891 22089
rect 22833 22080 22845 22083
rect 22796 22052 22845 22080
rect 22796 22040 22802 22052
rect 22833 22049 22845 22052
rect 22879 22049 22891 22083
rect 22833 22043 22891 22049
rect 23934 22040 23940 22092
rect 23992 22040 23998 22092
rect 19460 22015 19518 22021
rect 19460 21981 19472 22015
rect 19506 22012 19518 22015
rect 20254 22012 20260 22024
rect 19506 21984 20260 22012
rect 19506 21981 19518 21984
rect 19460 21975 19518 21981
rect 20254 21972 20260 21984
rect 20312 21972 20318 22024
rect 20346 21972 20352 22024
rect 20404 21972 20410 22024
rect 22189 22015 22247 22021
rect 22189 21981 22201 22015
rect 22235 22012 22247 22015
rect 23566 22012 23572 22024
rect 22235 21984 23572 22012
rect 22235 21981 22247 21984
rect 22189 21975 22247 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 23753 22015 23811 22021
rect 23753 21981 23765 22015
rect 23799 22012 23811 22015
rect 24044 22012 24072 22120
rect 25682 22108 25688 22120
rect 25740 22108 25746 22160
rect 27080 22148 27108 22188
rect 27246 22176 27252 22228
rect 27304 22216 27310 22228
rect 27890 22216 27896 22228
rect 27304 22188 27896 22216
rect 27304 22176 27310 22188
rect 27890 22176 27896 22188
rect 27948 22176 27954 22228
rect 28442 22176 28448 22228
rect 28500 22216 28506 22228
rect 29089 22219 29147 22225
rect 29089 22216 29101 22219
rect 28500 22188 29101 22216
rect 28500 22176 28506 22188
rect 29089 22185 29101 22188
rect 29135 22216 29147 22219
rect 29270 22216 29276 22228
rect 29135 22188 29276 22216
rect 29135 22185 29147 22188
rect 29089 22179 29147 22185
rect 29270 22176 29276 22188
rect 29328 22176 29334 22228
rect 29638 22176 29644 22228
rect 29696 22216 29702 22228
rect 29733 22219 29791 22225
rect 29733 22216 29745 22219
rect 29696 22188 29745 22216
rect 29696 22176 29702 22188
rect 29733 22185 29745 22188
rect 29779 22185 29791 22219
rect 29733 22179 29791 22185
rect 30006 22176 30012 22228
rect 30064 22216 30070 22228
rect 30064 22188 30420 22216
rect 30064 22176 30070 22188
rect 30282 22148 30288 22160
rect 27080 22120 30288 22148
rect 30282 22108 30288 22120
rect 30340 22108 30346 22160
rect 25130 22040 25136 22092
rect 25188 22040 25194 22092
rect 26050 22080 26056 22092
rect 25700 22052 26056 22080
rect 23799 21984 24072 22012
rect 23799 21981 23811 21984
rect 23753 21975 23811 21981
rect 17678 21944 17684 21956
rect 14844 21916 17684 21944
rect 17678 21904 17684 21916
rect 17736 21904 17742 21956
rect 19705 21947 19763 21953
rect 18708 21916 19334 21944
rect 11204 21848 13676 21876
rect 14185 21879 14243 21885
rect 11204 21836 11210 21848
rect 14185 21845 14197 21879
rect 14231 21876 14243 21879
rect 16206 21876 16212 21888
rect 14231 21848 16212 21876
rect 14231 21845 14243 21848
rect 14185 21839 14243 21845
rect 16206 21836 16212 21848
rect 16264 21836 16270 21888
rect 17586 21836 17592 21888
rect 17644 21876 17650 21888
rect 18708 21876 18736 21916
rect 17644 21848 18736 21876
rect 18877 21879 18935 21885
rect 17644 21836 17650 21848
rect 18877 21845 18889 21879
rect 18923 21876 18935 21879
rect 19150 21876 19156 21888
rect 18923 21848 19156 21876
rect 18923 21845 18935 21848
rect 18877 21839 18935 21845
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 19306 21876 19334 21916
rect 19705 21913 19717 21947
rect 19751 21944 19763 21947
rect 20622 21944 20628 21956
rect 19751 21916 20628 21944
rect 19751 21913 19763 21916
rect 19705 21907 19763 21913
rect 20622 21904 20628 21916
rect 20680 21904 20686 21956
rect 24949 21947 25007 21953
rect 20732 21916 24624 21944
rect 19426 21876 19432 21888
rect 19306 21848 19432 21876
rect 19426 21836 19432 21848
rect 19484 21836 19490 21888
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 20732 21876 20760 21916
rect 19668 21848 20760 21876
rect 19668 21836 19674 21848
rect 22738 21836 22744 21888
rect 22796 21876 22802 21888
rect 23661 21879 23719 21885
rect 23661 21876 23673 21879
rect 22796 21848 23673 21876
rect 22796 21836 22802 21848
rect 23661 21845 23673 21848
rect 23707 21876 23719 21879
rect 24394 21876 24400 21888
rect 23707 21848 24400 21876
rect 23707 21845 23719 21848
rect 23661 21839 23719 21845
rect 24394 21836 24400 21848
rect 24452 21836 24458 21888
rect 24596 21885 24624 21916
rect 24949 21913 24961 21947
rect 24995 21944 25007 21947
rect 25700 21944 25728 22052
rect 26050 22040 26056 22052
rect 26108 22040 26114 22092
rect 27522 22040 27528 22092
rect 27580 22040 27586 22092
rect 30392 22089 30420 22188
rect 30558 22176 30564 22228
rect 30616 22216 30622 22228
rect 39666 22216 39672 22228
rect 30616 22188 39672 22216
rect 30616 22176 30622 22188
rect 39666 22176 39672 22188
rect 39724 22176 39730 22228
rect 40218 22176 40224 22228
rect 40276 22216 40282 22228
rect 41690 22216 41696 22228
rect 40276 22188 41696 22216
rect 40276 22176 40282 22188
rect 41690 22176 41696 22188
rect 41748 22176 41754 22228
rect 43530 22176 43536 22228
rect 43588 22216 43594 22228
rect 43588 22188 45968 22216
rect 43588 22176 43594 22188
rect 35066 22108 35072 22160
rect 35124 22148 35130 22160
rect 45002 22148 45008 22160
rect 35124 22120 45008 22148
rect 35124 22108 35130 22120
rect 45002 22108 45008 22120
rect 45060 22108 45066 22160
rect 30377 22083 30435 22089
rect 27632 22052 29868 22080
rect 25777 22015 25835 22021
rect 25777 21981 25789 22015
rect 25823 21981 25835 22015
rect 25777 21975 25835 21981
rect 24995 21916 25728 21944
rect 25792 21944 25820 21975
rect 27338 21972 27344 22024
rect 27396 22012 27402 22024
rect 27632 22012 27660 22052
rect 29840 22024 29868 22052
rect 30377 22049 30389 22083
rect 30423 22080 30435 22083
rect 31849 22083 31907 22089
rect 31849 22080 31861 22083
rect 30423 22052 30457 22080
rect 30852 22052 31861 22080
rect 30423 22049 30435 22052
rect 30377 22043 30435 22049
rect 27396 21984 27660 22012
rect 27985 22015 28043 22021
rect 27396 21972 27402 21984
rect 27985 21981 27997 22015
rect 28031 22012 28043 22015
rect 28810 22012 28816 22024
rect 28031 21984 28816 22012
rect 28031 21981 28043 21984
rect 27985 21975 28043 21981
rect 28810 21972 28816 21984
rect 28868 21972 28874 22024
rect 29822 21972 29828 22024
rect 29880 22012 29886 22024
rect 30101 22015 30159 22021
rect 30101 22012 30113 22015
rect 29880 21984 30113 22012
rect 29880 21972 29886 21984
rect 30101 21981 30113 21984
rect 30147 22012 30159 22015
rect 30852 22012 30880 22052
rect 31849 22049 31861 22052
rect 31895 22049 31907 22083
rect 31849 22043 31907 22049
rect 33318 22040 33324 22092
rect 33376 22080 33382 22092
rect 34057 22083 34115 22089
rect 34057 22080 34069 22083
rect 33376 22052 34069 22080
rect 33376 22040 33382 22052
rect 34057 22049 34069 22052
rect 34103 22049 34115 22083
rect 34057 22043 34115 22049
rect 36998 22040 37004 22092
rect 37056 22040 37062 22092
rect 37182 22040 37188 22092
rect 37240 22080 37246 22092
rect 39209 22083 39267 22089
rect 39209 22080 39221 22083
rect 37240 22052 39221 22080
rect 37240 22040 37246 22052
rect 39209 22049 39221 22052
rect 39255 22049 39267 22083
rect 39209 22043 39267 22049
rect 40313 22083 40371 22089
rect 40313 22049 40325 22083
rect 40359 22080 40371 22083
rect 40402 22080 40408 22092
rect 40359 22052 40408 22080
rect 40359 22049 40371 22052
rect 40313 22043 40371 22049
rect 40402 22040 40408 22052
rect 40460 22040 40466 22092
rect 41598 22040 41604 22092
rect 41656 22040 41662 22092
rect 45830 22080 45836 22092
rect 42628 22052 45836 22080
rect 30147 21984 30880 22012
rect 30147 21981 30159 21984
rect 30101 21975 30159 21981
rect 30926 21972 30932 22024
rect 30984 21972 30990 22024
rect 31573 22015 31631 22021
rect 31573 21981 31585 22015
rect 31619 22012 31631 22015
rect 32309 22015 32367 22021
rect 32309 22012 32321 22015
rect 31619 21984 32321 22012
rect 31619 21981 31631 21984
rect 31573 21975 31631 21981
rect 32309 21981 32321 21984
rect 32355 21981 32367 22015
rect 32309 21975 32367 21981
rect 33042 21972 33048 22024
rect 33100 21972 33106 22024
rect 33410 21972 33416 22024
rect 33468 21972 33474 22024
rect 34514 21972 34520 22024
rect 34572 22012 34578 22024
rect 34885 22015 34943 22021
rect 34885 22012 34897 22015
rect 34572 21984 34897 22012
rect 34572 21972 34578 21984
rect 34885 21981 34897 21984
rect 34931 21981 34943 22015
rect 34885 21975 34943 21981
rect 34974 21972 34980 22024
rect 35032 22012 35038 22024
rect 35989 22015 36047 22021
rect 35989 22012 36001 22015
rect 35032 21984 36001 22012
rect 35032 21972 35038 21984
rect 35989 21981 36001 21984
rect 36035 21981 36047 22015
rect 35989 21975 36047 21981
rect 37461 22015 37519 22021
rect 37461 21981 37473 22015
rect 37507 22012 37519 22015
rect 37507 21984 37688 22012
rect 37507 21981 37519 21984
rect 37461 21975 37519 21981
rect 25958 21944 25964 21956
rect 25792 21916 25964 21944
rect 24995 21913 25007 21916
rect 24949 21907 25007 21913
rect 25958 21904 25964 21916
rect 26016 21904 26022 21956
rect 26326 21944 26332 21956
rect 26068 21916 26332 21944
rect 24581 21879 24639 21885
rect 24581 21845 24593 21879
rect 24627 21845 24639 21879
rect 24581 21839 24639 21845
rect 25041 21879 25099 21885
rect 25041 21845 25053 21879
rect 25087 21876 25099 21879
rect 25314 21876 25320 21888
rect 25087 21848 25320 21876
rect 25087 21845 25099 21848
rect 25041 21839 25099 21845
rect 25314 21836 25320 21848
rect 25372 21836 25378 21888
rect 25406 21836 25412 21888
rect 25464 21876 25470 21888
rect 26068 21876 26096 21916
rect 26326 21904 26332 21916
rect 26384 21904 26390 21956
rect 27062 21904 27068 21956
rect 27120 21904 27126 21956
rect 32953 21947 33011 21953
rect 32953 21944 32965 21947
rect 27540 21916 32965 21944
rect 25464 21848 26096 21876
rect 25464 21836 25470 21848
rect 26234 21836 26240 21888
rect 26292 21876 26298 21888
rect 27540 21876 27568 21916
rect 32953 21913 32965 21916
rect 32999 21913 33011 21947
rect 33060 21944 33088 21972
rect 34790 21944 34796 21956
rect 33060 21916 34796 21944
rect 32953 21907 33011 21913
rect 34790 21904 34796 21916
rect 34848 21904 34854 21956
rect 36078 21904 36084 21956
rect 36136 21944 36142 21956
rect 37090 21944 37096 21956
rect 36136 21916 37096 21944
rect 36136 21904 36142 21916
rect 37090 21904 37096 21916
rect 37148 21904 37154 21956
rect 37660 21944 37688 21984
rect 37826 21972 37832 22024
rect 37884 22012 37890 22024
rect 38565 22015 38623 22021
rect 38565 22012 38577 22015
rect 37884 21984 38577 22012
rect 37884 21972 37890 21984
rect 38565 21981 38577 21984
rect 38611 21981 38623 22015
rect 38565 21975 38623 21981
rect 38838 21972 38844 22024
rect 38896 22012 38902 22024
rect 40037 22015 40095 22021
rect 40037 22012 40049 22015
rect 38896 21984 40049 22012
rect 38896 21972 38902 21984
rect 40037 21981 40049 21984
rect 40083 21981 40095 22015
rect 40037 21975 40095 21981
rect 40678 21972 40684 22024
rect 40736 22012 40742 22024
rect 42628 22021 42656 22052
rect 45830 22040 45836 22052
rect 45888 22040 45894 22092
rect 41325 22015 41383 22021
rect 41325 22012 41337 22015
rect 40736 21984 41337 22012
rect 40736 21972 40742 21984
rect 41325 21981 41337 21984
rect 41371 21981 41383 22015
rect 41325 21975 41383 21981
rect 42613 22015 42671 22021
rect 42613 21981 42625 22015
rect 42659 21981 42671 22015
rect 42613 21975 42671 21981
rect 43717 22015 43775 22021
rect 43717 21981 43729 22015
rect 43763 21981 43775 22015
rect 43717 21975 43775 21981
rect 40126 21944 40132 21956
rect 37660 21916 40132 21944
rect 40126 21904 40132 21916
rect 40184 21904 40190 21956
rect 40402 21904 40408 21956
rect 40460 21944 40466 21956
rect 43732 21944 43760 21975
rect 44358 21972 44364 22024
rect 44416 21972 44422 22024
rect 45940 22021 45968 22188
rect 46474 22176 46480 22228
rect 46532 22216 46538 22228
rect 46661 22219 46719 22225
rect 46661 22216 46673 22219
rect 46532 22188 46673 22216
rect 46532 22176 46538 22188
rect 46661 22185 46673 22188
rect 46707 22185 46719 22219
rect 46661 22179 46719 22185
rect 46014 22108 46020 22160
rect 46072 22148 46078 22160
rect 46845 22151 46903 22157
rect 46845 22148 46857 22151
rect 46072 22120 46857 22148
rect 46072 22108 46078 22120
rect 46845 22117 46857 22120
rect 46891 22148 46903 22151
rect 46891 22120 47256 22148
rect 46891 22117 46903 22120
rect 46845 22111 46903 22117
rect 47228 22021 47256 22120
rect 48498 22040 48504 22092
rect 48556 22080 48562 22092
rect 49329 22083 49387 22089
rect 49329 22080 49341 22083
rect 48556 22052 49341 22080
rect 48556 22040 48562 22052
rect 49329 22049 49341 22052
rect 49375 22049 49387 22083
rect 49329 22043 49387 22049
rect 45189 22015 45247 22021
rect 45189 21981 45201 22015
rect 45235 21981 45247 22015
rect 45189 21975 45247 21981
rect 45925 22015 45983 22021
rect 45925 21981 45937 22015
rect 45971 22012 45983 22015
rect 46477 22015 46535 22021
rect 46477 22012 46489 22015
rect 45971 21984 46489 22012
rect 45971 21981 45983 21984
rect 45925 21975 45983 21981
rect 46477 21981 46489 21984
rect 46523 21981 46535 22015
rect 46477 21975 46535 21981
rect 47213 22015 47271 22021
rect 47213 21981 47225 22015
rect 47259 21981 47271 22015
rect 47213 21975 47271 21981
rect 40460 21916 43760 21944
rect 40460 21904 40466 21916
rect 26292 21848 27568 21876
rect 26292 21836 26298 21848
rect 27614 21836 27620 21888
rect 27672 21876 27678 21888
rect 28629 21879 28687 21885
rect 28629 21876 28641 21879
rect 27672 21848 28641 21876
rect 27672 21836 27678 21848
rect 28629 21845 28641 21848
rect 28675 21845 28687 21879
rect 28629 21839 28687 21845
rect 28902 21836 28908 21888
rect 28960 21876 28966 21888
rect 30006 21876 30012 21888
rect 28960 21848 30012 21876
rect 28960 21836 28966 21848
rect 30006 21836 30012 21848
rect 30064 21836 30070 21888
rect 30193 21879 30251 21885
rect 30193 21845 30205 21879
rect 30239 21876 30251 21879
rect 30282 21876 30288 21888
rect 30239 21848 30288 21876
rect 30239 21845 30251 21848
rect 30193 21839 30251 21845
rect 30282 21836 30288 21848
rect 30340 21836 30346 21888
rect 30742 21836 30748 21888
rect 30800 21876 30806 21888
rect 33042 21876 33048 21888
rect 30800 21848 33048 21876
rect 30800 21836 30806 21848
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 34330 21836 34336 21888
rect 34388 21836 34394 21888
rect 34422 21836 34428 21888
rect 34480 21876 34486 21888
rect 35529 21879 35587 21885
rect 35529 21876 35541 21879
rect 34480 21848 35541 21876
rect 34480 21836 34486 21848
rect 35529 21845 35541 21848
rect 35575 21845 35587 21879
rect 35529 21839 35587 21845
rect 35618 21836 35624 21888
rect 35676 21876 35682 21888
rect 36633 21879 36691 21885
rect 36633 21876 36645 21879
rect 35676 21848 36645 21876
rect 35676 21836 35682 21848
rect 36633 21845 36645 21848
rect 36679 21845 36691 21879
rect 36633 21839 36691 21845
rect 37182 21836 37188 21888
rect 37240 21876 37246 21888
rect 38105 21879 38163 21885
rect 38105 21876 38117 21879
rect 37240 21848 38117 21876
rect 37240 21836 37246 21848
rect 38105 21845 38117 21848
rect 38151 21845 38163 21879
rect 38105 21839 38163 21845
rect 38746 21836 38752 21888
rect 38804 21876 38810 21888
rect 39485 21879 39543 21885
rect 39485 21876 39497 21879
rect 38804 21848 39497 21876
rect 38804 21836 38810 21848
rect 39485 21845 39497 21848
rect 39531 21845 39543 21879
rect 39485 21839 39543 21845
rect 43254 21836 43260 21888
rect 43312 21836 43318 21888
rect 43732 21876 43760 21916
rect 44174 21904 44180 21956
rect 44232 21944 44238 21956
rect 45204 21944 45232 21975
rect 47854 21972 47860 22024
rect 47912 22012 47918 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 47912 21984 47961 22012
rect 47912 21972 47918 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 48682 21972 48688 22024
rect 48740 21972 48746 22024
rect 45278 21944 45284 21956
rect 44232 21916 45284 21944
rect 44232 21904 44238 21916
rect 45278 21904 45284 21916
rect 45336 21904 45342 21956
rect 45462 21904 45468 21956
rect 45520 21944 45526 21956
rect 45520 21904 45554 21944
rect 44637 21879 44695 21885
rect 44637 21876 44649 21879
rect 43732 21848 44649 21876
rect 44637 21845 44649 21848
rect 44683 21845 44695 21879
rect 44637 21839 44695 21845
rect 45370 21836 45376 21888
rect 45428 21836 45434 21888
rect 45526 21876 45554 21904
rect 46109 21879 46167 21885
rect 46109 21876 46121 21879
rect 45526 21848 46121 21876
rect 46109 21845 46121 21848
rect 46155 21845 46167 21879
rect 46109 21839 46167 21845
rect 47394 21836 47400 21888
rect 47452 21836 47458 21888
rect 47854 21836 47860 21888
rect 47912 21876 47918 21888
rect 48133 21879 48191 21885
rect 48133 21876 48145 21879
rect 47912 21848 48145 21876
rect 47912 21836 47918 21848
rect 48133 21845 48145 21848
rect 48179 21845 48191 21879
rect 48133 21839 48191 21845
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 5169 21675 5227 21681
rect 5169 21641 5181 21675
rect 5215 21672 5227 21675
rect 5718 21672 5724 21684
rect 5215 21644 5724 21672
rect 5215 21641 5227 21644
rect 5169 21635 5227 21641
rect 5718 21632 5724 21644
rect 5776 21632 5782 21684
rect 6457 21675 6515 21681
rect 6457 21641 6469 21675
rect 6503 21672 6515 21675
rect 6917 21675 6975 21681
rect 6917 21672 6929 21675
rect 6503 21644 6929 21672
rect 6503 21641 6515 21644
rect 6457 21635 6515 21641
rect 6917 21641 6929 21644
rect 6963 21672 6975 21675
rect 7098 21672 7104 21684
rect 6963 21644 7104 21672
rect 6963 21641 6975 21644
rect 6917 21635 6975 21641
rect 7098 21632 7104 21644
rect 7156 21632 7162 21684
rect 11701 21675 11759 21681
rect 11701 21672 11713 21675
rect 8404 21644 11713 21672
rect 4430 21564 4436 21616
rect 4488 21604 4494 21616
rect 6270 21604 6276 21616
rect 4488 21576 6276 21604
rect 4488 21564 4494 21576
rect 6270 21564 6276 21576
rect 6328 21564 6334 21616
rect 7009 21607 7067 21613
rect 7009 21573 7021 21607
rect 7055 21604 7067 21607
rect 8404 21604 8432 21644
rect 11701 21641 11713 21644
rect 11747 21641 11759 21675
rect 11701 21635 11759 21641
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12161 21675 12219 21681
rect 12161 21672 12173 21675
rect 12124 21644 12173 21672
rect 12124 21632 12130 21644
rect 12161 21641 12173 21644
rect 12207 21641 12219 21675
rect 12161 21635 12219 21641
rect 15289 21675 15347 21681
rect 15289 21641 15301 21675
rect 15335 21672 15347 21675
rect 15335 21644 21128 21672
rect 15335 21641 15347 21644
rect 15289 21635 15347 21641
rect 21100 21616 21128 21644
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 23934 21672 23940 21684
rect 23348 21644 23940 21672
rect 23348 21632 23354 21644
rect 23934 21632 23940 21644
rect 23992 21672 23998 21684
rect 23992 21644 24072 21672
rect 23992 21632 23998 21644
rect 9398 21604 9404 21616
rect 7055 21576 8432 21604
rect 9246 21576 9404 21604
rect 7055 21573 7067 21576
rect 7009 21567 7067 21573
rect 9398 21564 9404 21576
rect 9456 21564 9462 21616
rect 9953 21607 10011 21613
rect 9953 21573 9965 21607
rect 9999 21604 10011 21607
rect 9999 21576 12204 21604
rect 9999 21573 10011 21576
rect 9953 21567 10011 21573
rect 1670 21496 1676 21548
rect 1728 21496 1734 21548
rect 3602 21496 3608 21548
rect 3660 21496 3666 21548
rect 5626 21496 5632 21548
rect 5684 21496 5690 21548
rect 10229 21539 10287 21545
rect 10229 21505 10241 21539
rect 10275 21505 10287 21539
rect 10229 21499 10287 21505
rect 2774 21428 2780 21480
rect 2832 21428 2838 21480
rect 4154 21428 4160 21480
rect 4212 21428 4218 21480
rect 5905 21471 5963 21477
rect 5905 21437 5917 21471
rect 5951 21468 5963 21471
rect 7098 21468 7104 21480
rect 5951 21440 7104 21468
rect 5951 21437 5963 21440
rect 5905 21431 5963 21437
rect 7098 21428 7104 21440
rect 7156 21428 7162 21480
rect 7193 21471 7251 21477
rect 7193 21437 7205 21471
rect 7239 21468 7251 21471
rect 7558 21468 7564 21480
rect 7239 21440 7564 21468
rect 7239 21437 7251 21440
rect 7193 21431 7251 21437
rect 7558 21428 7564 21440
rect 7616 21428 7622 21480
rect 7745 21471 7803 21477
rect 7745 21437 7757 21471
rect 7791 21437 7803 21471
rect 7745 21431 7803 21437
rect 2498 21360 2504 21412
rect 2556 21400 2562 21412
rect 7006 21400 7012 21412
rect 2556 21372 7012 21400
rect 2556 21360 2562 21372
rect 7006 21360 7012 21372
rect 7064 21360 7070 21412
rect 5261 21335 5319 21341
rect 5261 21301 5273 21335
rect 5307 21332 5319 21335
rect 5442 21332 5448 21344
rect 5307 21304 5448 21332
rect 5307 21301 5319 21304
rect 5261 21295 5319 21301
rect 5442 21292 5448 21304
rect 5500 21292 5506 21344
rect 6546 21292 6552 21344
rect 6604 21292 6610 21344
rect 7760 21332 7788 21431
rect 8018 21428 8024 21480
rect 8076 21428 8082 21480
rect 8386 21428 8392 21480
rect 8444 21468 8450 21480
rect 10244 21468 10272 21499
rect 10318 21496 10324 21548
rect 10376 21536 10382 21548
rect 12069 21539 12127 21545
rect 12069 21536 12081 21539
rect 10376 21508 12081 21536
rect 10376 21496 10382 21508
rect 12069 21505 12081 21508
rect 12115 21505 12127 21539
rect 12176 21536 12204 21576
rect 12250 21564 12256 21616
rect 12308 21604 12314 21616
rect 12308 21576 12940 21604
rect 12308 21564 12314 21576
rect 12710 21536 12716 21548
rect 12176 21508 12716 21536
rect 12069 21499 12127 21505
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 10502 21468 10508 21480
rect 8444 21440 10508 21468
rect 8444 21428 8450 21440
rect 10502 21428 10508 21440
rect 10560 21428 10566 21480
rect 10962 21428 10968 21480
rect 11020 21428 11026 21480
rect 12250 21428 12256 21480
rect 12308 21428 12314 21480
rect 12912 21477 12940 21576
rect 15102 21564 15108 21616
rect 15160 21564 15166 21616
rect 18414 21604 18420 21616
rect 15672 21576 18420 21604
rect 14458 21536 14464 21548
rect 14306 21508 14464 21536
rect 14458 21496 14464 21508
rect 14516 21536 14522 21548
rect 15672 21536 15700 21576
rect 18414 21564 18420 21576
rect 18472 21564 18478 21616
rect 18874 21564 18880 21616
rect 18932 21604 18938 21616
rect 18969 21607 19027 21613
rect 18969 21604 18981 21607
rect 18932 21576 18981 21604
rect 18932 21564 18938 21576
rect 18969 21573 18981 21576
rect 19015 21604 19027 21607
rect 19058 21604 19064 21616
rect 19015 21576 19064 21604
rect 19015 21573 19027 21576
rect 18969 21567 19027 21573
rect 19058 21564 19064 21576
rect 19116 21564 19122 21616
rect 20622 21604 20628 21616
rect 20194 21576 20628 21604
rect 20622 21564 20628 21576
rect 20680 21604 20686 21616
rect 20990 21604 20996 21616
rect 20680 21576 20996 21604
rect 20680 21564 20686 21576
rect 20990 21564 20996 21576
rect 21048 21564 21054 21616
rect 21082 21564 21088 21616
rect 21140 21564 21146 21616
rect 23658 21564 23664 21616
rect 23716 21564 23722 21616
rect 24044 21604 24072 21644
rect 25038 21632 25044 21684
rect 25096 21672 25102 21684
rect 26605 21675 26663 21681
rect 26605 21672 26617 21675
rect 25096 21644 26617 21672
rect 25096 21632 25102 21644
rect 26605 21641 26617 21644
rect 26651 21672 26663 21675
rect 27522 21672 27528 21684
rect 26651 21644 27528 21672
rect 26651 21641 26663 21644
rect 26605 21635 26663 21641
rect 27522 21632 27528 21644
rect 27580 21672 27586 21684
rect 27617 21675 27675 21681
rect 27617 21672 27629 21675
rect 27580 21644 27629 21672
rect 27580 21632 27586 21644
rect 27617 21641 27629 21644
rect 27663 21641 27675 21675
rect 27617 21635 27675 21641
rect 27709 21675 27767 21681
rect 27709 21641 27721 21675
rect 27755 21672 27767 21675
rect 28350 21672 28356 21684
rect 27755 21644 28356 21672
rect 27755 21641 27767 21644
rect 27709 21635 27767 21641
rect 28350 21632 28356 21644
rect 28408 21632 28414 21684
rect 28644 21644 28856 21672
rect 25961 21607 26019 21613
rect 24044 21576 24150 21604
rect 25961 21573 25973 21607
rect 26007 21604 26019 21607
rect 26050 21604 26056 21616
rect 26007 21576 26056 21604
rect 26007 21573 26019 21576
rect 25961 21567 26019 21573
rect 26050 21564 26056 21576
rect 26108 21564 26114 21616
rect 26142 21564 26148 21616
rect 26200 21564 26206 21616
rect 26237 21607 26295 21613
rect 26237 21573 26249 21607
rect 26283 21604 26295 21607
rect 27890 21604 27896 21616
rect 26283 21576 27896 21604
rect 26283 21573 26295 21576
rect 26237 21567 26295 21573
rect 27890 21564 27896 21576
rect 27948 21564 27954 21616
rect 27982 21564 27988 21616
rect 28040 21604 28046 21616
rect 28644 21604 28672 21644
rect 28040 21576 28672 21604
rect 28040 21564 28046 21576
rect 28718 21564 28724 21616
rect 28776 21564 28782 21616
rect 28828 21604 28856 21644
rect 29012 21644 30052 21672
rect 29012 21604 29040 21644
rect 28828 21576 29040 21604
rect 30024 21604 30052 21644
rect 30926 21632 30932 21684
rect 30984 21672 30990 21684
rect 32953 21675 33011 21681
rect 32953 21672 32965 21675
rect 30984 21644 32965 21672
rect 30984 21632 30990 21644
rect 32953 21641 32965 21644
rect 32999 21641 33011 21675
rect 32953 21635 33011 21641
rect 33042 21632 33048 21684
rect 33100 21672 33106 21684
rect 34333 21675 34391 21681
rect 34333 21672 34345 21675
rect 33100 21644 34345 21672
rect 33100 21632 33106 21644
rect 34333 21641 34345 21644
rect 34379 21641 34391 21675
rect 34333 21635 34391 21641
rect 36538 21632 36544 21684
rect 36596 21672 36602 21684
rect 36633 21675 36691 21681
rect 36633 21672 36645 21675
rect 36596 21644 36645 21672
rect 36596 21632 36602 21644
rect 36633 21641 36645 21644
rect 36679 21641 36691 21675
rect 36633 21635 36691 21641
rect 37090 21632 37096 21684
rect 37148 21672 37154 21684
rect 37826 21672 37832 21684
rect 37148 21644 37832 21672
rect 37148 21632 37154 21644
rect 37826 21632 37832 21644
rect 37884 21632 37890 21684
rect 38286 21632 38292 21684
rect 38344 21672 38350 21684
rect 43254 21672 43260 21684
rect 38344 21644 43260 21672
rect 38344 21632 38350 21644
rect 43254 21632 43260 21644
rect 43312 21632 43318 21684
rect 44082 21632 44088 21684
rect 44140 21632 44146 21684
rect 44910 21632 44916 21684
rect 44968 21672 44974 21684
rect 45189 21675 45247 21681
rect 45189 21672 45201 21675
rect 44968 21644 45201 21672
rect 44968 21632 44974 21644
rect 45189 21641 45201 21644
rect 45235 21641 45247 21675
rect 45189 21635 45247 21641
rect 45278 21632 45284 21684
rect 45336 21672 45342 21684
rect 45557 21675 45615 21681
rect 45557 21672 45569 21675
rect 45336 21644 45569 21672
rect 45336 21632 45342 21644
rect 45557 21641 45569 21644
rect 45603 21641 45615 21675
rect 45557 21635 45615 21641
rect 45646 21632 45652 21684
rect 45704 21672 45710 21684
rect 45741 21675 45799 21681
rect 45741 21672 45753 21675
rect 45704 21644 45753 21672
rect 45704 21632 45710 21644
rect 45741 21641 45753 21644
rect 45787 21641 45799 21675
rect 45741 21635 45799 21641
rect 47026 21632 47032 21684
rect 47084 21632 47090 21684
rect 47673 21675 47731 21681
rect 47673 21641 47685 21675
rect 47719 21672 47731 21675
rect 47762 21672 47768 21684
rect 47719 21644 47768 21672
rect 47719 21641 47731 21644
rect 47673 21635 47731 21641
rect 47762 21632 47768 21644
rect 47820 21632 47826 21684
rect 30024 21576 31248 21604
rect 14516 21508 15700 21536
rect 14516 21496 14522 21508
rect 15930 21496 15936 21548
rect 15988 21536 15994 21548
rect 16482 21536 16488 21548
rect 15988 21508 16488 21536
rect 15988 21496 15994 21508
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 17037 21539 17095 21545
rect 17037 21505 17049 21539
rect 17083 21536 17095 21539
rect 17126 21536 17132 21548
rect 17083 21508 17132 21536
rect 17083 21505 17095 21508
rect 17037 21499 17095 21505
rect 17126 21496 17132 21508
rect 17184 21496 17190 21548
rect 17770 21536 17776 21548
rect 17236 21508 17776 21536
rect 12897 21471 12955 21477
rect 12897 21437 12909 21471
rect 12943 21468 12955 21471
rect 13173 21471 13231 21477
rect 12943 21440 13032 21468
rect 12943 21437 12955 21440
rect 12897 21431 12955 21437
rect 9493 21403 9551 21409
rect 9493 21369 9505 21403
rect 9539 21400 9551 21403
rect 9582 21400 9588 21412
rect 9539 21372 9588 21400
rect 9539 21369 9551 21372
rect 9493 21363 9551 21369
rect 9582 21360 9588 21372
rect 9640 21360 9646 21412
rect 8662 21332 8668 21344
rect 7760 21304 8668 21332
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 13004 21332 13032 21440
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 13538 21468 13544 21480
rect 13219 21440 13544 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 14826 21468 14832 21480
rect 13780 21440 14832 21468
rect 13780 21428 13786 21440
rect 14826 21428 14832 21440
rect 14884 21468 14890 21480
rect 15102 21468 15108 21480
rect 14884 21440 15108 21468
rect 14884 21428 14890 21440
rect 15102 21428 15108 21440
rect 15160 21428 15166 21480
rect 15746 21428 15752 21480
rect 15804 21468 15810 21480
rect 16025 21471 16083 21477
rect 16025 21468 16037 21471
rect 15804 21440 16037 21468
rect 15804 21428 15810 21440
rect 16025 21437 16037 21440
rect 16071 21437 16083 21471
rect 16025 21431 16083 21437
rect 16114 21428 16120 21480
rect 16172 21468 16178 21480
rect 16209 21471 16267 21477
rect 16209 21468 16221 21471
rect 16172 21440 16221 21468
rect 16172 21428 16178 21440
rect 16209 21437 16221 21440
rect 16255 21437 16267 21471
rect 16209 21431 16267 21437
rect 14366 21360 14372 21412
rect 14424 21400 14430 21412
rect 16224 21400 16252 21431
rect 16758 21428 16764 21480
rect 16816 21468 16822 21480
rect 17236 21468 17264 21508
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 20254 21496 20260 21548
rect 20312 21536 20318 21548
rect 20312 21508 21772 21536
rect 20312 21496 20318 21508
rect 16816 21440 17264 21468
rect 16816 21428 16822 21440
rect 17310 21428 17316 21480
rect 17368 21428 17374 21480
rect 17494 21428 17500 21480
rect 17552 21468 17558 21480
rect 18693 21471 18751 21477
rect 18693 21468 18705 21471
rect 17552 21440 18705 21468
rect 17552 21428 17558 21440
rect 18693 21437 18705 21440
rect 18739 21437 18751 21471
rect 18693 21431 18751 21437
rect 17954 21400 17960 21412
rect 14424 21372 16160 21400
rect 16224 21372 17960 21400
rect 14424 21360 14430 21372
rect 13538 21332 13544 21344
rect 13004 21304 13544 21332
rect 13538 21292 13544 21304
rect 13596 21292 13602 21344
rect 14645 21335 14703 21341
rect 14645 21301 14657 21335
rect 14691 21332 14703 21335
rect 14918 21332 14924 21344
rect 14691 21304 14924 21332
rect 14691 21301 14703 21304
rect 14645 21295 14703 21301
rect 14918 21292 14924 21304
rect 14976 21292 14982 21344
rect 15378 21292 15384 21344
rect 15436 21332 15442 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15436 21304 15577 21332
rect 15436 21292 15442 21304
rect 15565 21301 15577 21304
rect 15611 21301 15623 21335
rect 16132 21332 16160 21372
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 16298 21332 16304 21344
rect 16132 21304 16304 21332
rect 15565 21295 15623 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 18708 21332 18736 21431
rect 19058 21428 19064 21480
rect 19116 21468 19122 21480
rect 21634 21468 21640 21480
rect 19116 21440 21640 21468
rect 19116 21428 19122 21440
rect 21634 21428 21640 21440
rect 21692 21428 21698 21480
rect 21744 21468 21772 21508
rect 22002 21496 22008 21548
rect 22060 21496 22066 21548
rect 25314 21496 25320 21548
rect 25372 21536 25378 21548
rect 27430 21536 27436 21548
rect 25372 21508 27436 21536
rect 25372 21496 25378 21508
rect 27430 21496 27436 21508
rect 27488 21496 27494 21548
rect 27522 21496 27528 21548
rect 27580 21536 27586 21548
rect 28074 21536 28080 21548
rect 27580 21508 28080 21536
rect 27580 21496 27586 21508
rect 28074 21496 28080 21508
rect 28132 21496 28138 21548
rect 28442 21496 28448 21548
rect 28500 21496 28506 21548
rect 29730 21496 29736 21548
rect 29788 21536 29794 21548
rect 30650 21536 30656 21548
rect 29788 21508 30656 21536
rect 29788 21496 29794 21508
rect 30650 21496 30656 21508
rect 30708 21496 30714 21548
rect 30742 21496 30748 21548
rect 30800 21536 30806 21548
rect 31021 21539 31079 21545
rect 31021 21536 31033 21539
rect 30800 21508 31033 21536
rect 30800 21496 30806 21508
rect 31021 21505 31033 21508
rect 31067 21505 31079 21539
rect 31021 21499 31079 21505
rect 31110 21496 31116 21548
rect 31168 21496 31174 21548
rect 31220 21536 31248 21576
rect 31754 21564 31760 21616
rect 31812 21604 31818 21616
rect 31812 21576 32444 21604
rect 31812 21564 31818 21576
rect 32309 21539 32367 21545
rect 32309 21536 32321 21539
rect 31220 21508 32321 21536
rect 32309 21505 32321 21508
rect 32355 21505 32367 21539
rect 32416 21536 32444 21576
rect 32582 21564 32588 21616
rect 32640 21604 32646 21616
rect 32766 21604 32772 21616
rect 32640 21576 32772 21604
rect 32640 21564 32646 21576
rect 32766 21564 32772 21576
rect 32824 21564 32830 21616
rect 32858 21564 32864 21616
rect 32916 21604 32922 21616
rect 32916 21576 44956 21604
rect 32916 21564 32922 21576
rect 33318 21536 33324 21548
rect 32416 21508 33324 21536
rect 32309 21499 32367 21505
rect 33318 21496 33324 21508
rect 33376 21496 33382 21548
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21536 33471 21539
rect 34422 21536 34428 21548
rect 33459 21508 34428 21536
rect 33459 21505 33471 21508
rect 33413 21499 33471 21505
rect 34422 21496 34428 21508
rect 34480 21496 34486 21548
rect 34885 21539 34943 21545
rect 34885 21505 34897 21539
rect 34931 21536 34943 21539
rect 35618 21536 35624 21548
rect 34931 21508 35624 21536
rect 34931 21505 34943 21508
rect 34885 21499 34943 21505
rect 35618 21496 35624 21508
rect 35676 21496 35682 21548
rect 35894 21496 35900 21548
rect 35952 21536 35958 21548
rect 35989 21539 36047 21545
rect 35989 21536 36001 21539
rect 35952 21508 36001 21536
rect 35952 21496 35958 21508
rect 35989 21505 36001 21508
rect 36035 21505 36047 21539
rect 35989 21499 36047 21505
rect 37734 21496 37740 21548
rect 37792 21496 37798 21548
rect 38746 21496 38752 21548
rect 38804 21496 38810 21548
rect 39482 21496 39488 21548
rect 39540 21536 39546 21548
rect 39850 21536 39856 21548
rect 39540 21508 39856 21536
rect 39540 21496 39546 21508
rect 39850 21496 39856 21508
rect 39908 21496 39914 21548
rect 40957 21539 41015 21545
rect 40957 21536 40969 21539
rect 40052 21508 40969 21536
rect 22370 21468 22376 21480
rect 21744 21440 22376 21468
rect 22370 21428 22376 21440
rect 22428 21468 22434 21480
rect 22741 21471 22799 21477
rect 22741 21468 22753 21471
rect 22428 21440 22753 21468
rect 22428 21428 22434 21440
rect 22741 21437 22753 21440
rect 22787 21437 22799 21471
rect 22741 21431 22799 21437
rect 23382 21428 23388 21480
rect 23440 21428 23446 21480
rect 23658 21428 23664 21480
rect 23716 21468 23722 21480
rect 27706 21468 27712 21480
rect 23716 21440 27712 21468
rect 23716 21428 23722 21440
rect 27706 21428 27712 21440
rect 27764 21428 27770 21480
rect 27801 21471 27859 21477
rect 27801 21437 27813 21471
rect 27847 21437 27859 21471
rect 27801 21431 27859 21437
rect 20441 21403 20499 21409
rect 20441 21369 20453 21403
rect 20487 21400 20499 21403
rect 22278 21400 22284 21412
rect 20487 21372 22284 21400
rect 20487 21369 20499 21372
rect 20441 21363 20499 21369
rect 22278 21360 22284 21372
rect 22336 21360 22342 21412
rect 23106 21360 23112 21412
rect 23164 21400 23170 21412
rect 23290 21400 23296 21412
rect 23164 21372 23296 21400
rect 23164 21360 23170 21372
rect 23290 21360 23296 21372
rect 23348 21360 23354 21412
rect 19702 21332 19708 21344
rect 18708 21304 19708 21332
rect 19702 21292 19708 21304
rect 19760 21332 19766 21344
rect 20254 21332 20260 21344
rect 19760 21304 20260 21332
rect 19760 21292 19766 21304
rect 20254 21292 20260 21304
rect 20312 21292 20318 21344
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 21361 21335 21419 21341
rect 21361 21332 21373 21335
rect 21324 21304 21373 21332
rect 21324 21292 21330 21304
rect 21361 21301 21373 21304
rect 21407 21332 21419 21335
rect 21634 21332 21640 21344
rect 21407 21304 21640 21332
rect 21407 21301 21419 21304
rect 21361 21295 21419 21301
rect 21634 21292 21640 21304
rect 21692 21332 21698 21344
rect 22002 21332 22008 21344
rect 21692 21304 22008 21332
rect 21692 21292 21698 21304
rect 22002 21292 22008 21304
rect 22060 21292 22066 21344
rect 23400 21332 23428 21428
rect 24670 21360 24676 21412
rect 24728 21400 24734 21412
rect 25130 21400 25136 21412
rect 24728 21372 25136 21400
rect 24728 21360 24734 21372
rect 25130 21360 25136 21372
rect 25188 21360 25194 21412
rect 26510 21400 26516 21412
rect 25608 21372 26516 21400
rect 24118 21332 24124 21344
rect 23400 21304 24124 21332
rect 24118 21292 24124 21304
rect 24176 21292 24182 21344
rect 24394 21292 24400 21344
rect 24452 21332 24458 21344
rect 25608 21332 25636 21372
rect 26510 21360 26516 21372
rect 26568 21360 26574 21412
rect 26602 21360 26608 21412
rect 26660 21400 26666 21412
rect 27062 21400 27068 21412
rect 26660 21372 27068 21400
rect 26660 21360 26666 21372
rect 27062 21360 27068 21372
rect 27120 21400 27126 21412
rect 27338 21400 27344 21412
rect 27120 21372 27344 21400
rect 27120 21360 27126 21372
rect 27338 21360 27344 21372
rect 27396 21360 27402 21412
rect 27816 21400 27844 21431
rect 27890 21428 27896 21480
rect 27948 21468 27954 21480
rect 29914 21468 29920 21480
rect 27948 21440 29920 21468
rect 27948 21428 27954 21440
rect 29914 21428 29920 21440
rect 29972 21428 29978 21480
rect 30193 21471 30251 21477
rect 30193 21437 30205 21471
rect 30239 21468 30251 21471
rect 31205 21471 31263 21477
rect 31205 21468 31217 21471
rect 30239 21440 31217 21468
rect 30239 21437 30251 21440
rect 30193 21431 30251 21437
rect 31205 21437 31217 21440
rect 31251 21468 31263 21471
rect 34974 21468 34980 21480
rect 31251 21440 34980 21468
rect 31251 21437 31263 21440
rect 31205 21431 31263 21437
rect 34974 21428 34980 21440
rect 35032 21428 35038 21480
rect 36998 21428 37004 21480
rect 37056 21468 37062 21480
rect 37461 21471 37519 21477
rect 37461 21468 37473 21471
rect 37056 21440 37473 21468
rect 37056 21428 37062 21440
rect 37461 21437 37473 21440
rect 37507 21437 37519 21471
rect 37461 21431 37519 21437
rect 27982 21400 27988 21412
rect 27816 21372 27988 21400
rect 27982 21360 27988 21372
rect 28040 21360 28046 21412
rect 30098 21360 30104 21412
rect 30156 21400 30162 21412
rect 30156 21372 31754 21400
rect 30156 21360 30162 21372
rect 24452 21304 25636 21332
rect 24452 21292 24458 21304
rect 25682 21292 25688 21344
rect 25740 21292 25746 21344
rect 27246 21292 27252 21344
rect 27304 21292 27310 21344
rect 27522 21292 27528 21344
rect 27580 21332 27586 21344
rect 30653 21335 30711 21341
rect 30653 21332 30665 21335
rect 27580 21304 30665 21332
rect 27580 21292 27586 21304
rect 30653 21301 30665 21304
rect 30699 21301 30711 21335
rect 31726 21332 31754 21372
rect 31938 21360 31944 21412
rect 31996 21400 32002 21412
rect 40052 21400 40080 21508
rect 40957 21505 40969 21508
rect 41003 21536 41015 21539
rect 41782 21536 41788 21548
rect 41003 21508 41788 21536
rect 41003 21505 41015 21508
rect 40957 21499 41015 21505
rect 41782 21496 41788 21508
rect 41840 21496 41846 21548
rect 42518 21496 42524 21548
rect 42576 21536 42582 21548
rect 42705 21539 42763 21545
rect 42705 21536 42717 21539
rect 42576 21508 42717 21536
rect 42576 21496 42582 21508
rect 42705 21505 42717 21508
rect 42751 21505 42763 21539
rect 42705 21499 42763 21505
rect 43441 21539 43499 21545
rect 43441 21505 43453 21539
rect 43487 21536 43499 21539
rect 43622 21536 43628 21548
rect 43487 21508 43628 21536
rect 43487 21505 43499 21508
rect 43441 21499 43499 21505
rect 43622 21496 43628 21508
rect 43680 21496 43686 21548
rect 43990 21496 43996 21548
rect 44048 21536 44054 21548
rect 44928 21545 44956 21576
rect 44269 21539 44327 21545
rect 44269 21536 44281 21539
rect 44048 21508 44281 21536
rect 44048 21496 44054 21508
rect 44269 21505 44281 21508
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 44913 21539 44971 21545
rect 44913 21505 44925 21539
rect 44959 21536 44971 21539
rect 45373 21539 45431 21545
rect 45373 21536 45385 21539
rect 44959 21508 45385 21536
rect 44959 21505 44971 21508
rect 44913 21499 44971 21505
rect 45373 21505 45385 21508
rect 45419 21505 45431 21539
rect 45373 21499 45431 21505
rect 47210 21496 47216 21548
rect 47268 21496 47274 21548
rect 47762 21496 47768 21548
rect 47820 21536 47826 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 47820 21508 47961 21536
rect 47820 21496 47826 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 41601 21471 41659 21477
rect 41601 21437 41613 21471
rect 41647 21468 41659 21471
rect 44450 21468 44456 21480
rect 41647 21440 44456 21468
rect 41647 21437 41659 21440
rect 41601 21431 41659 21437
rect 44450 21428 44456 21440
rect 44508 21428 44514 21480
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 31996 21372 40080 21400
rect 40144 21372 40632 21400
rect 31996 21360 32002 21372
rect 31846 21332 31852 21344
rect 31726 21304 31852 21332
rect 30653 21295 30711 21301
rect 31846 21292 31852 21304
rect 31904 21292 31910 21344
rect 32122 21292 32128 21344
rect 32180 21332 32186 21344
rect 32582 21332 32588 21344
rect 32180 21304 32588 21332
rect 32180 21292 32186 21304
rect 32582 21292 32588 21304
rect 32640 21292 32646 21344
rect 33502 21292 33508 21344
rect 33560 21332 33566 21344
rect 34057 21335 34115 21341
rect 34057 21332 34069 21335
rect 33560 21304 34069 21332
rect 33560 21292 33566 21304
rect 34057 21301 34069 21304
rect 34103 21301 34115 21335
rect 34057 21295 34115 21301
rect 34609 21335 34667 21341
rect 34609 21301 34621 21335
rect 34655 21332 34667 21335
rect 35250 21332 35256 21344
rect 34655 21304 35256 21332
rect 34655 21301 34667 21304
rect 34609 21295 34667 21301
rect 35250 21292 35256 21304
rect 35308 21292 35314 21344
rect 35529 21335 35587 21341
rect 35529 21301 35541 21335
rect 35575 21332 35587 21335
rect 35986 21332 35992 21344
rect 35575 21304 35992 21332
rect 35575 21301 35587 21304
rect 35529 21295 35587 21301
rect 35986 21292 35992 21304
rect 36044 21292 36050 21344
rect 36538 21292 36544 21344
rect 36596 21332 36602 21344
rect 36998 21332 37004 21344
rect 36596 21304 37004 21332
rect 36596 21292 36602 21304
rect 36998 21292 37004 21304
rect 37056 21292 37062 21344
rect 38194 21292 38200 21344
rect 38252 21332 38258 21344
rect 39393 21335 39451 21341
rect 39393 21332 39405 21335
rect 38252 21304 39405 21332
rect 38252 21292 38258 21304
rect 39393 21301 39405 21304
rect 39439 21301 39451 21335
rect 39393 21295 39451 21301
rect 39482 21292 39488 21344
rect 39540 21332 39546 21344
rect 40144 21332 40172 21372
rect 39540 21304 40172 21332
rect 39540 21292 39546 21304
rect 40218 21292 40224 21344
rect 40276 21332 40282 21344
rect 40497 21335 40555 21341
rect 40497 21332 40509 21335
rect 40276 21304 40509 21332
rect 40276 21292 40282 21304
rect 40497 21301 40509 21304
rect 40543 21301 40555 21335
rect 40604 21332 40632 21372
rect 41322 21360 41328 21412
rect 41380 21400 41386 21412
rect 42061 21403 42119 21409
rect 42061 21400 42073 21403
rect 41380 21372 42073 21400
rect 41380 21360 41386 21372
rect 42061 21369 42073 21372
rect 42107 21369 42119 21403
rect 42061 21363 42119 21369
rect 41877 21335 41935 21341
rect 41877 21332 41889 21335
rect 40604 21304 41889 21332
rect 40497 21295 40555 21301
rect 41877 21301 41889 21304
rect 41923 21301 41935 21335
rect 41877 21295 41935 21301
rect 42794 21292 42800 21344
rect 42852 21292 42858 21344
rect 43530 21292 43536 21344
rect 43588 21292 43594 21344
rect 44726 21292 44732 21344
rect 44784 21292 44790 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 3602 21088 3608 21140
rect 3660 21128 3666 21140
rect 3786 21128 3792 21140
rect 3660 21100 3792 21128
rect 3660 21088 3666 21100
rect 3786 21088 3792 21100
rect 3844 21088 3850 21140
rect 10965 21131 11023 21137
rect 6288 21100 10456 21128
rect 3513 21063 3571 21069
rect 3513 21029 3525 21063
rect 3559 21060 3571 21063
rect 6288 21060 6316 21100
rect 3559 21032 6316 21060
rect 3559 21029 3571 21032
rect 3513 21023 3571 21029
rect 7558 21020 7564 21072
rect 7616 21060 7622 21072
rect 9950 21060 9956 21072
rect 7616 21032 9956 21060
rect 7616 21020 7622 21032
rect 9950 21020 9956 21032
rect 10008 21020 10014 21072
rect 2038 20952 2044 21004
rect 2096 20952 2102 21004
rect 3786 20952 3792 21004
rect 3844 20992 3850 21004
rect 4433 20995 4491 21001
rect 4433 20992 4445 20995
rect 3844 20964 4445 20992
rect 3844 20952 3850 20964
rect 4433 20961 4445 20964
rect 4479 20961 4491 20995
rect 4433 20955 4491 20961
rect 6822 20952 6828 21004
rect 6880 20992 6886 21004
rect 6880 20964 7788 20992
rect 6880 20952 6886 20964
rect 7576 20936 7604 20964
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 2222 20924 2228 20936
rect 1811 20896 2228 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 4062 20884 4068 20936
rect 4120 20884 4126 20936
rect 6178 20884 6184 20936
rect 6236 20884 6242 20936
rect 7558 20884 7564 20936
rect 7616 20884 7622 20936
rect 7760 20924 7788 20964
rect 7834 20952 7840 21004
rect 7892 20992 7898 21004
rect 8389 20995 8447 21001
rect 8389 20992 8401 20995
rect 7892 20964 8401 20992
rect 7892 20952 7898 20964
rect 8389 20961 8401 20964
rect 8435 20961 8447 20995
rect 9398 20992 9404 21004
rect 8389 20955 8447 20961
rect 8496 20964 9404 20992
rect 8496 20924 8524 20964
rect 9398 20952 9404 20964
rect 9456 20952 9462 21004
rect 10042 20952 10048 21004
rect 10100 20952 10106 21004
rect 7760 20896 8524 20924
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 10428 20924 10456 21100
rect 10965 21097 10977 21131
rect 11011 21128 11023 21131
rect 14366 21128 14372 21140
rect 11011 21100 14372 21128
rect 11011 21097 11023 21100
rect 10965 21091 11023 21097
rect 14366 21088 14372 21100
rect 14424 21088 14430 21140
rect 14553 21131 14611 21137
rect 14553 21097 14565 21131
rect 14599 21128 14611 21131
rect 15102 21128 15108 21140
rect 14599 21100 15108 21128
rect 14599 21097 14611 21100
rect 14553 21091 14611 21097
rect 15102 21088 15108 21100
rect 15160 21088 15166 21140
rect 15746 21088 15752 21140
rect 15804 21088 15810 21140
rect 16574 21128 16580 21140
rect 16132 21100 16580 21128
rect 10502 21020 10508 21072
rect 10560 21060 10566 21072
rect 14277 21063 14335 21069
rect 10560 21032 12940 21060
rect 10560 21020 10566 21032
rect 11517 20995 11575 21001
rect 11517 20961 11529 20995
rect 11563 20992 11575 20995
rect 11563 20964 12756 20992
rect 11563 20961 11575 20964
rect 11517 20955 11575 20961
rect 11974 20924 11980 20936
rect 10428 20896 11980 20924
rect 9309 20887 9367 20893
rect 2590 20816 2596 20868
rect 2648 20856 2654 20868
rect 5810 20856 5816 20868
rect 2648 20828 5816 20856
rect 2648 20816 2654 20828
rect 5810 20816 5816 20828
rect 5868 20816 5874 20868
rect 6454 20816 6460 20868
rect 6512 20816 6518 20868
rect 9324 20856 9352 20887
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12728 20924 12756 20964
rect 12802 20952 12808 21004
rect 12860 20952 12866 21004
rect 12912 20992 12940 21032
rect 14277 21029 14289 21063
rect 14323 21060 14335 21063
rect 16132 21060 16160 21100
rect 16574 21088 16580 21100
rect 16632 21088 16638 21140
rect 20162 21128 20168 21140
rect 17236 21100 20168 21128
rect 16390 21060 16396 21072
rect 14323 21032 16160 21060
rect 16224 21032 16396 21060
rect 14323 21029 14335 21032
rect 14277 21023 14335 21029
rect 14642 20992 14648 21004
rect 12912 20964 14648 20992
rect 14642 20952 14648 20964
rect 14700 20952 14706 21004
rect 15105 20995 15163 21001
rect 14752 20964 15056 20992
rect 13817 20927 13875 20933
rect 13817 20924 13829 20927
rect 12728 20896 13829 20924
rect 13817 20893 13829 20896
rect 13863 20924 13875 20927
rect 14366 20924 14372 20936
rect 13863 20896 14372 20924
rect 13863 20893 13875 20896
rect 13817 20887 13875 20893
rect 14366 20884 14372 20896
rect 14424 20884 14430 20936
rect 10502 20856 10508 20868
rect 9324 20828 10508 20856
rect 10502 20816 10508 20828
rect 10560 20816 10566 20868
rect 11149 20859 11207 20865
rect 11149 20825 11161 20859
rect 11195 20856 11207 20859
rect 13725 20859 13783 20865
rect 11195 20828 13676 20856
rect 11195 20825 11207 20828
rect 11149 20819 11207 20825
rect 3421 20791 3479 20797
rect 3421 20757 3433 20791
rect 3467 20788 3479 20791
rect 5534 20788 5540 20800
rect 3467 20760 5540 20788
rect 3467 20757 3479 20760
rect 3421 20751 3479 20757
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 5718 20748 5724 20800
rect 5776 20748 5782 20800
rect 5902 20748 5908 20800
rect 5960 20748 5966 20800
rect 7834 20748 7840 20800
rect 7892 20788 7898 20800
rect 7929 20791 7987 20797
rect 7929 20788 7941 20791
rect 7892 20760 7941 20788
rect 7892 20748 7898 20760
rect 7929 20757 7941 20760
rect 7975 20757 7987 20791
rect 7929 20751 7987 20757
rect 10134 20748 10140 20800
rect 10192 20788 10198 20800
rect 11238 20788 11244 20800
rect 10192 20760 11244 20788
rect 10192 20748 10198 20760
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 11330 20748 11336 20800
rect 11388 20788 11394 20800
rect 11514 20788 11520 20800
rect 11388 20760 11520 20788
rect 11388 20748 11394 20760
rect 11514 20748 11520 20760
rect 11572 20748 11578 20800
rect 11698 20748 11704 20800
rect 11756 20748 11762 20800
rect 13648 20788 13676 20828
rect 13725 20825 13737 20859
rect 13771 20856 13783 20859
rect 14642 20856 14648 20868
rect 13771 20828 14648 20856
rect 13771 20825 13783 20828
rect 13725 20819 13783 20825
rect 14642 20816 14648 20828
rect 14700 20816 14706 20868
rect 14752 20788 14780 20964
rect 15028 20924 15056 20964
rect 15105 20961 15117 20995
rect 15151 20992 15163 20995
rect 15194 20992 15200 21004
rect 15151 20964 15200 20992
rect 15151 20961 15163 20964
rect 15105 20955 15163 20961
rect 15194 20952 15200 20964
rect 15252 20952 15258 21004
rect 16224 21001 16252 21032
rect 16390 21020 16396 21032
rect 16448 21020 16454 21072
rect 16209 20995 16267 21001
rect 16209 20992 16221 20995
rect 15304 20964 16221 20992
rect 15304 20924 15332 20964
rect 16209 20961 16221 20964
rect 16255 20961 16267 20995
rect 16209 20955 16267 20961
rect 16298 20952 16304 21004
rect 16356 20952 16362 21004
rect 17236 20992 17264 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 23474 21128 23480 21140
rect 21928 21100 23480 21128
rect 17310 21020 17316 21072
rect 17368 21060 17374 21072
rect 17862 21060 17868 21072
rect 17368 21032 17868 21060
rect 17368 21020 17374 21032
rect 17862 21020 17868 21032
rect 17920 21020 17926 21072
rect 18800 21032 19564 21060
rect 16500 20964 17356 20992
rect 15028 20896 15332 20924
rect 16114 20884 16120 20936
rect 16172 20924 16178 20936
rect 16500 20924 16528 20964
rect 16172 20896 16528 20924
rect 16172 20884 16178 20896
rect 16574 20884 16580 20936
rect 16632 20924 16638 20936
rect 17328 20933 17356 20964
rect 17494 20952 17500 21004
rect 17552 20952 17558 21004
rect 18598 20952 18604 21004
rect 18656 20952 18662 21004
rect 18800 21001 18828 21032
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20961 18843 20995
rect 19536 20992 19564 21032
rect 21082 21020 21088 21072
rect 21140 21060 21146 21072
rect 21453 21063 21511 21069
rect 21453 21060 21465 21063
rect 21140 21032 21465 21060
rect 21140 21020 21146 21032
rect 21453 21029 21465 21032
rect 21499 21029 21511 21063
rect 21453 21023 21511 21029
rect 21928 20992 21956 21100
rect 23474 21088 23480 21100
rect 23532 21088 23538 21140
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 27246 21128 27252 21140
rect 23624 21100 27252 21128
rect 23624 21088 23630 21100
rect 27246 21088 27252 21100
rect 27304 21088 27310 21140
rect 27706 21088 27712 21140
rect 27764 21088 27770 21140
rect 28442 21088 28448 21140
rect 28500 21128 28506 21140
rect 29089 21131 29147 21137
rect 29089 21128 29101 21131
rect 28500 21100 29101 21128
rect 28500 21088 28506 21100
rect 29089 21097 29101 21100
rect 29135 21097 29147 21131
rect 29089 21091 29147 21097
rect 29270 21088 29276 21140
rect 29328 21128 29334 21140
rect 30742 21128 30748 21140
rect 29328 21100 30748 21128
rect 29328 21088 29334 21100
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 31478 21088 31484 21140
rect 31536 21128 31542 21140
rect 31536 21100 31616 21128
rect 31536 21088 31542 21100
rect 25406 21060 25412 21072
rect 22388 21032 25412 21060
rect 19536 20964 21956 20992
rect 22281 20995 22339 21001
rect 18785 20955 18843 20961
rect 22281 20961 22293 20995
rect 22327 20992 22339 20995
rect 22388 20992 22416 21032
rect 25406 21020 25412 21032
rect 25464 21020 25470 21072
rect 27430 21020 27436 21072
rect 27488 21060 27494 21072
rect 28718 21060 28724 21072
rect 27488 21032 28724 21060
rect 27488 21020 27494 21032
rect 28718 21020 28724 21032
rect 28776 21020 28782 21072
rect 28810 21020 28816 21072
rect 28868 21020 28874 21072
rect 31205 21063 31263 21069
rect 31205 21029 31217 21063
rect 31251 21029 31263 21063
rect 31205 21023 31263 21029
rect 22327 20964 22416 20992
rect 22465 20995 22523 21001
rect 22327 20961 22339 20964
rect 22281 20955 22339 20961
rect 22465 20961 22477 20995
rect 22511 20961 22523 20995
rect 22465 20955 22523 20961
rect 17313 20927 17371 20933
rect 16632 20896 16988 20924
rect 16632 20884 16638 20896
rect 14826 20816 14832 20868
rect 14884 20816 14890 20868
rect 15013 20859 15071 20865
rect 15013 20825 15025 20859
rect 15059 20856 15071 20859
rect 15654 20856 15660 20868
rect 15059 20828 15660 20856
rect 15059 20825 15071 20828
rect 15013 20819 15071 20825
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 15838 20816 15844 20868
rect 15896 20856 15902 20868
rect 16850 20856 16856 20868
rect 15896 20828 16856 20856
rect 15896 20816 15902 20828
rect 16850 20816 16856 20828
rect 16908 20816 16914 20868
rect 16960 20856 16988 20896
rect 17313 20893 17325 20927
rect 17359 20893 17371 20927
rect 17313 20887 17371 20893
rect 17402 20884 17408 20936
rect 17460 20924 17466 20936
rect 18414 20924 18420 20936
rect 17460 20896 18420 20924
rect 17460 20884 17466 20896
rect 18414 20884 18420 20896
rect 18472 20884 18478 20936
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20924 18567 20927
rect 18966 20924 18972 20936
rect 18555 20896 18972 20924
rect 18555 20893 18567 20896
rect 18509 20887 18567 20893
rect 18966 20884 18972 20896
rect 19024 20884 19030 20936
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 22189 20927 22247 20933
rect 22189 20924 22201 20927
rect 21284 20896 22201 20924
rect 19058 20856 19064 20868
rect 16960 20828 19064 20856
rect 19058 20816 19064 20828
rect 19116 20816 19122 20868
rect 19705 20859 19763 20865
rect 19705 20825 19717 20859
rect 19751 20856 19763 20859
rect 19978 20856 19984 20868
rect 19751 20828 19984 20856
rect 19751 20825 19763 20828
rect 19705 20819 19763 20825
rect 19978 20816 19984 20828
rect 20036 20816 20042 20868
rect 20990 20856 20996 20868
rect 20930 20828 20996 20856
rect 20990 20816 20996 20828
rect 21048 20816 21054 20868
rect 13648 20760 14780 20788
rect 14844 20788 14872 20816
rect 21284 20800 21312 20896
rect 22189 20893 22201 20896
rect 22235 20893 22247 20927
rect 22189 20887 22247 20893
rect 21358 20816 21364 20868
rect 21416 20856 21422 20868
rect 22480 20856 22508 20955
rect 23566 20952 23572 21004
rect 23624 20952 23630 21004
rect 23661 20995 23719 21001
rect 23661 20961 23673 20995
rect 23707 20961 23719 20995
rect 23661 20955 23719 20961
rect 22554 20884 22560 20936
rect 22612 20924 22618 20936
rect 23198 20924 23204 20936
rect 22612 20896 23204 20924
rect 22612 20884 22618 20896
rect 23198 20884 23204 20896
rect 23256 20884 23262 20936
rect 23477 20927 23535 20933
rect 23477 20893 23489 20927
rect 23523 20924 23535 20927
rect 23584 20924 23612 20952
rect 23523 20896 23612 20924
rect 23523 20893 23535 20896
rect 23477 20887 23535 20893
rect 23566 20856 23572 20868
rect 21416 20828 21956 20856
rect 22480 20828 23572 20856
rect 21416 20816 21422 20828
rect 14921 20791 14979 20797
rect 14921 20788 14933 20791
rect 14844 20760 14933 20788
rect 14921 20757 14933 20760
rect 14967 20757 14979 20791
rect 14921 20751 14979 20757
rect 16114 20748 16120 20800
rect 16172 20748 16178 20800
rect 16942 20748 16948 20800
rect 17000 20748 17006 20800
rect 17402 20748 17408 20800
rect 17460 20748 17466 20800
rect 18141 20791 18199 20797
rect 18141 20757 18153 20791
rect 18187 20788 18199 20791
rect 18874 20788 18880 20800
rect 18187 20760 18880 20788
rect 18187 20757 18199 20760
rect 18141 20751 18199 20757
rect 18874 20748 18880 20760
rect 18932 20748 18938 20800
rect 20714 20748 20720 20800
rect 20772 20788 20778 20800
rect 21177 20791 21235 20797
rect 21177 20788 21189 20791
rect 20772 20760 21189 20788
rect 20772 20748 20778 20760
rect 21177 20757 21189 20760
rect 21223 20757 21235 20791
rect 21177 20751 21235 20757
rect 21266 20748 21272 20800
rect 21324 20788 21330 20800
rect 21729 20791 21787 20797
rect 21729 20788 21741 20791
rect 21324 20760 21741 20788
rect 21324 20748 21330 20760
rect 21729 20757 21741 20760
rect 21775 20757 21787 20791
rect 21729 20751 21787 20757
rect 21818 20748 21824 20800
rect 21876 20748 21882 20800
rect 21928 20788 21956 20828
rect 23566 20816 23572 20828
rect 23624 20816 23630 20868
rect 22554 20788 22560 20800
rect 21928 20760 22560 20788
rect 22554 20748 22560 20760
rect 22612 20748 22618 20800
rect 22738 20748 22744 20800
rect 22796 20788 22802 20800
rect 23017 20791 23075 20797
rect 23017 20788 23029 20791
rect 22796 20760 23029 20788
rect 22796 20748 22802 20760
rect 23017 20757 23029 20760
rect 23063 20757 23075 20791
rect 23017 20751 23075 20757
rect 23198 20748 23204 20800
rect 23256 20788 23262 20800
rect 23385 20791 23443 20797
rect 23385 20788 23397 20791
rect 23256 20760 23397 20788
rect 23256 20748 23262 20760
rect 23385 20757 23397 20760
rect 23431 20757 23443 20791
rect 23385 20751 23443 20757
rect 23474 20748 23480 20800
rect 23532 20788 23538 20800
rect 23676 20788 23704 20955
rect 23934 20952 23940 21004
rect 23992 20992 23998 21004
rect 25130 20992 25136 21004
rect 23992 20964 25136 20992
rect 23992 20952 23998 20964
rect 25130 20952 25136 20964
rect 25188 20952 25194 21004
rect 25222 20952 25228 21004
rect 25280 20952 25286 21004
rect 25314 20952 25320 21004
rect 25372 20992 25378 21004
rect 31220 20992 31248 21023
rect 25372 20964 31248 20992
rect 25372 20952 25378 20964
rect 24118 20884 24124 20936
rect 24176 20924 24182 20936
rect 24213 20927 24271 20933
rect 24213 20924 24225 20927
rect 24176 20896 24225 20924
rect 24176 20884 24182 20896
rect 24213 20893 24225 20896
rect 24259 20924 24271 20927
rect 25958 20924 25964 20936
rect 24259 20896 25964 20924
rect 24259 20893 24271 20896
rect 24213 20887 24271 20893
rect 25958 20884 25964 20896
rect 26016 20884 26022 20936
rect 27338 20884 27344 20936
rect 27396 20884 27402 20936
rect 27706 20884 27712 20936
rect 27764 20924 27770 20936
rect 27982 20924 27988 20936
rect 27764 20896 27988 20924
rect 27764 20884 27770 20896
rect 27982 20884 27988 20896
rect 28040 20884 28046 20936
rect 31588 20933 31616 21100
rect 31846 21088 31852 21140
rect 31904 21128 31910 21140
rect 32858 21128 32864 21140
rect 31904 21100 32864 21128
rect 31904 21088 31910 21100
rect 32858 21088 32864 21100
rect 32916 21088 32922 21140
rect 34698 21088 34704 21140
rect 34756 21128 34762 21140
rect 35069 21131 35127 21137
rect 35069 21128 35081 21131
rect 34756 21100 35081 21128
rect 34756 21088 34762 21100
rect 35069 21097 35081 21100
rect 35115 21097 35127 21131
rect 35069 21091 35127 21097
rect 35176 21100 37320 21128
rect 32490 21020 32496 21072
rect 32548 21060 32554 21072
rect 35176 21060 35204 21100
rect 37182 21060 37188 21072
rect 32548 21032 35204 21060
rect 35820 21032 37188 21060
rect 32548 21020 32554 21032
rect 31849 20995 31907 21001
rect 31849 20961 31861 20995
rect 31895 20992 31907 20995
rect 32122 20992 32128 21004
rect 31895 20964 32128 20992
rect 31895 20961 31907 20964
rect 31849 20955 31907 20961
rect 32122 20952 32128 20964
rect 32180 20952 32186 21004
rect 32582 20952 32588 21004
rect 32640 20992 32646 21004
rect 35820 21001 35848 21032
rect 37182 21020 37188 21032
rect 37240 21020 37246 21072
rect 37292 21060 37320 21100
rect 38838 21088 38844 21140
rect 38896 21088 38902 21140
rect 40678 21088 40684 21140
rect 40736 21088 40742 21140
rect 41325 21131 41383 21137
rect 41325 21097 41337 21131
rect 41371 21128 41383 21131
rect 41966 21128 41972 21140
rect 41371 21100 41972 21128
rect 41371 21097 41383 21100
rect 41325 21091 41383 21097
rect 41966 21088 41972 21100
rect 42024 21088 42030 21140
rect 44082 21088 44088 21140
rect 44140 21128 44146 21140
rect 44637 21131 44695 21137
rect 44637 21128 44649 21131
rect 44140 21100 44649 21128
rect 44140 21088 44146 21100
rect 44637 21097 44649 21100
rect 44683 21097 44695 21131
rect 44637 21091 44695 21097
rect 48409 21131 48467 21137
rect 48409 21097 48421 21131
rect 48455 21128 48467 21131
rect 48590 21128 48596 21140
rect 48455 21100 48596 21128
rect 48455 21097 48467 21100
rect 48409 21091 48467 21097
rect 48590 21088 48596 21100
rect 48648 21088 48654 21140
rect 49326 21088 49332 21140
rect 49384 21088 49390 21140
rect 43993 21063 44051 21069
rect 43993 21060 44005 21063
rect 37292 21032 44005 21060
rect 43993 21029 44005 21032
rect 44039 21029 44051 21063
rect 43993 21023 44051 21029
rect 35805 20995 35863 21001
rect 32640 20964 35664 20992
rect 32640 20952 32646 20964
rect 28169 20927 28227 20933
rect 28169 20893 28181 20927
rect 28215 20924 28227 20927
rect 31573 20927 31631 20933
rect 28215 20896 31524 20924
rect 28215 20893 28227 20896
rect 28169 20887 28227 20893
rect 25041 20859 25099 20865
rect 25041 20825 25053 20859
rect 25087 20856 25099 20859
rect 26142 20856 26148 20868
rect 25087 20828 26148 20856
rect 25087 20825 25099 20828
rect 25041 20819 25099 20825
rect 26142 20816 26148 20828
rect 26200 20816 26206 20868
rect 26234 20816 26240 20868
rect 26292 20816 26298 20868
rect 27798 20816 27804 20868
rect 27856 20856 27862 20868
rect 29825 20859 29883 20865
rect 27856 20828 29776 20856
rect 27856 20816 27862 20828
rect 23532 20760 23704 20788
rect 23532 20748 23538 20760
rect 24670 20748 24676 20800
rect 24728 20748 24734 20800
rect 25133 20791 25191 20797
rect 25133 20757 25145 20791
rect 25179 20788 25191 20791
rect 27522 20788 27528 20800
rect 25179 20760 27528 20788
rect 25179 20757 25191 20760
rect 25133 20751 25191 20757
rect 27522 20748 27528 20760
rect 27580 20748 27586 20800
rect 28074 20748 28080 20800
rect 28132 20788 28138 20800
rect 28810 20788 28816 20800
rect 28132 20760 28816 20788
rect 28132 20748 28138 20760
rect 28810 20748 28816 20760
rect 28868 20788 28874 20800
rect 29270 20788 29276 20800
rect 28868 20760 29276 20788
rect 28868 20748 28874 20760
rect 29270 20748 29276 20760
rect 29328 20748 29334 20800
rect 29748 20788 29776 20828
rect 29825 20825 29837 20859
rect 29871 20856 29883 20859
rect 30098 20856 30104 20868
rect 29871 20828 30104 20856
rect 29871 20825 29883 20828
rect 29825 20819 29883 20825
rect 30098 20816 30104 20828
rect 30156 20816 30162 20868
rect 30650 20816 30656 20868
rect 30708 20856 30714 20868
rect 31496 20856 31524 20896
rect 31573 20893 31585 20927
rect 31619 20893 31631 20927
rect 31573 20887 31631 20893
rect 31662 20884 31668 20936
rect 31720 20884 31726 20936
rect 31938 20884 31944 20936
rect 31996 20924 32002 20936
rect 32401 20927 32459 20933
rect 32401 20924 32413 20927
rect 31996 20896 32413 20924
rect 31996 20884 32002 20896
rect 32401 20893 32413 20896
rect 32447 20893 32459 20927
rect 32401 20887 32459 20893
rect 33502 20884 33508 20936
rect 33560 20884 33566 20936
rect 34517 20927 34575 20933
rect 34517 20893 34529 20927
rect 34563 20924 34575 20927
rect 35434 20924 35440 20936
rect 34563 20896 35440 20924
rect 34563 20893 34575 20896
rect 34517 20887 34575 20893
rect 35434 20884 35440 20896
rect 35492 20884 35498 20936
rect 33045 20859 33103 20865
rect 33045 20856 33057 20859
rect 30708 20828 31248 20856
rect 31496 20828 33057 20856
rect 30708 20816 30714 20828
rect 31110 20788 31116 20800
rect 29748 20760 31116 20788
rect 31110 20748 31116 20760
rect 31168 20748 31174 20800
rect 31220 20788 31248 20828
rect 33045 20825 33057 20828
rect 33091 20825 33103 20859
rect 34977 20859 35035 20865
rect 34977 20856 34989 20859
rect 33045 20819 33103 20825
rect 34072 20828 34989 20856
rect 31754 20788 31760 20800
rect 31220 20760 31760 20788
rect 31754 20748 31760 20760
rect 31812 20748 31818 20800
rect 32214 20748 32220 20800
rect 32272 20788 32278 20800
rect 34072 20788 34100 20828
rect 34977 20825 34989 20828
rect 35023 20856 35035 20859
rect 35529 20859 35587 20865
rect 35529 20856 35541 20859
rect 35023 20828 35541 20856
rect 35023 20825 35035 20828
rect 34977 20819 35035 20825
rect 35529 20825 35541 20828
rect 35575 20825 35587 20859
rect 35636 20856 35664 20964
rect 35805 20961 35817 20995
rect 35851 20961 35863 20995
rect 35805 20955 35863 20961
rect 36081 20995 36139 21001
rect 36081 20961 36093 20995
rect 36127 20992 36139 20995
rect 36170 20992 36176 21004
rect 36127 20964 36176 20992
rect 36127 20961 36139 20964
rect 36081 20955 36139 20961
rect 36170 20952 36176 20964
rect 36228 20952 36234 21004
rect 37200 20964 44220 20992
rect 36262 20884 36268 20936
rect 36320 20924 36326 20936
rect 37093 20927 37151 20933
rect 37093 20924 37105 20927
rect 36320 20896 37105 20924
rect 36320 20884 36326 20896
rect 37093 20893 37105 20896
rect 37139 20893 37151 20927
rect 37093 20887 37151 20893
rect 37200 20856 37228 20964
rect 38194 20884 38200 20936
rect 38252 20884 38258 20936
rect 39206 20884 39212 20936
rect 39264 20924 39270 20936
rect 39482 20924 39488 20936
rect 39264 20896 39488 20924
rect 39264 20884 39270 20896
rect 39482 20884 39488 20896
rect 39540 20884 39546 20936
rect 40034 20884 40040 20936
rect 40092 20884 40098 20936
rect 41969 20927 42027 20933
rect 41969 20893 41981 20927
rect 42015 20924 42027 20927
rect 42058 20924 42064 20936
rect 42015 20896 42064 20924
rect 42015 20893 42027 20896
rect 41969 20887 42027 20893
rect 42058 20884 42064 20896
rect 42116 20884 42122 20936
rect 43438 20884 43444 20936
rect 43496 20924 43502 20936
rect 44192 20933 44220 20964
rect 43533 20927 43591 20933
rect 43533 20924 43545 20927
rect 43496 20896 43545 20924
rect 43496 20884 43502 20896
rect 43533 20893 43545 20896
rect 43579 20893 43591 20927
rect 43533 20887 43591 20893
rect 44177 20927 44235 20933
rect 44177 20893 44189 20927
rect 44223 20924 44235 20927
rect 44453 20927 44511 20933
rect 44453 20924 44465 20927
rect 44223 20896 44465 20924
rect 44223 20893 44235 20896
rect 44177 20887 44235 20893
rect 44453 20893 44465 20896
rect 44499 20893 44511 20927
rect 44453 20887 44511 20893
rect 48590 20884 48596 20936
rect 48648 20924 48654 20936
rect 48685 20927 48743 20933
rect 48685 20924 48697 20927
rect 48648 20896 48697 20924
rect 48648 20884 48654 20896
rect 48685 20893 48697 20896
rect 48731 20893 48743 20927
rect 48685 20887 48743 20893
rect 35636 20828 37228 20856
rect 41233 20859 41291 20865
rect 35529 20819 35587 20825
rect 41233 20825 41245 20859
rect 41279 20856 41291 20859
rect 41322 20856 41328 20868
rect 41279 20828 41328 20856
rect 41279 20825 41291 20828
rect 41233 20819 41291 20825
rect 41322 20816 41328 20828
rect 41380 20816 41386 20868
rect 42702 20816 42708 20868
rect 42760 20816 42766 20868
rect 42889 20859 42947 20865
rect 42889 20825 42901 20859
rect 42935 20856 42947 20859
rect 43898 20856 43904 20868
rect 42935 20828 43904 20856
rect 42935 20825 42947 20828
rect 42889 20819 42947 20825
rect 43898 20816 43904 20828
rect 43956 20816 43962 20868
rect 32272 20760 34100 20788
rect 32272 20748 32278 20760
rect 34146 20748 34152 20800
rect 34204 20748 34210 20800
rect 37734 20748 37740 20800
rect 37792 20748 37798 20800
rect 39298 20748 39304 20800
rect 39356 20748 39362 20800
rect 42058 20748 42064 20800
rect 42116 20748 42122 20800
rect 43346 20748 43352 20800
rect 43404 20748 43410 20800
rect 47762 20748 47768 20800
rect 47820 20748 47826 20800
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 3786 20544 3792 20596
rect 3844 20584 3850 20596
rect 10686 20584 10692 20596
rect 3844 20556 10692 20584
rect 3844 20544 3850 20556
rect 10686 20544 10692 20556
rect 10744 20544 10750 20596
rect 11054 20544 11060 20596
rect 11112 20584 11118 20596
rect 11701 20587 11759 20593
rect 11701 20584 11713 20587
rect 11112 20556 11713 20584
rect 11112 20544 11118 20556
rect 11701 20553 11713 20556
rect 11747 20553 11759 20587
rect 11701 20547 11759 20553
rect 12342 20544 12348 20596
rect 12400 20544 12406 20596
rect 12820 20556 16068 20584
rect 3697 20519 3755 20525
rect 3697 20485 3709 20519
rect 3743 20516 3755 20519
rect 4246 20516 4252 20528
rect 3743 20488 4252 20516
rect 3743 20485 3755 20488
rect 3697 20479 3755 20485
rect 4246 20476 4252 20488
rect 4304 20476 4310 20528
rect 8481 20519 8539 20525
rect 8481 20516 8493 20519
rect 5920 20488 8493 20516
rect 1118 20408 1124 20460
rect 1176 20448 1182 20460
rect 1581 20451 1639 20457
rect 1581 20448 1593 20451
rect 1176 20420 1593 20448
rect 1176 20408 1182 20420
rect 1581 20417 1593 20420
rect 1627 20417 1639 20451
rect 1581 20411 1639 20417
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 3970 20448 3976 20460
rect 3559 20420 3976 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 5626 20408 5632 20460
rect 5684 20408 5690 20460
rect 1394 20340 1400 20392
rect 1452 20380 1458 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1452 20352 2053 20380
rect 1452 20340 1458 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 4249 20383 4307 20389
rect 4249 20349 4261 20383
rect 4295 20380 4307 20383
rect 4295 20352 4384 20380
rect 4295 20349 4307 20352
rect 4249 20343 4307 20349
rect 4356 20244 4384 20352
rect 4522 20340 4528 20392
rect 4580 20340 4586 20392
rect 5258 20340 5264 20392
rect 5316 20380 5322 20392
rect 5920 20380 5948 20488
rect 8481 20485 8493 20488
rect 8527 20516 8539 20519
rect 8941 20519 8999 20525
rect 8941 20516 8953 20519
rect 8527 20488 8953 20516
rect 8527 20485 8539 20488
rect 8481 20479 8539 20485
rect 8941 20485 8953 20488
rect 8987 20485 8999 20519
rect 8941 20479 8999 20485
rect 10870 20476 10876 20528
rect 10928 20516 10934 20528
rect 12713 20519 12771 20525
rect 12713 20516 12725 20519
rect 10928 20488 12725 20516
rect 10928 20476 10934 20488
rect 12713 20485 12725 20488
rect 12759 20485 12771 20519
rect 12713 20479 12771 20485
rect 6733 20451 6791 20457
rect 6733 20448 6745 20451
rect 6012 20420 6745 20448
rect 6012 20389 6040 20420
rect 6733 20417 6745 20420
rect 6779 20448 6791 20451
rect 6914 20448 6920 20460
rect 6779 20420 6920 20448
rect 6779 20417 6791 20420
rect 6733 20411 6791 20417
rect 6914 20408 6920 20420
rect 6972 20408 6978 20460
rect 5316 20352 5948 20380
rect 5997 20383 6055 20389
rect 5316 20340 5322 20352
rect 5997 20349 6009 20383
rect 6043 20349 6055 20383
rect 5997 20343 6055 20349
rect 7006 20340 7012 20392
rect 7064 20340 7070 20392
rect 8662 20340 8668 20392
rect 8720 20340 8726 20392
rect 10060 20380 10088 20434
rect 10502 20408 10508 20460
rect 10560 20448 10566 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10560 20420 10977 20448
rect 10560 20408 10566 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 11790 20408 11796 20460
rect 11848 20448 11854 20460
rect 11885 20451 11943 20457
rect 11885 20448 11897 20451
rect 11848 20420 11897 20448
rect 11848 20408 11854 20420
rect 11885 20417 11897 20420
rect 11931 20417 11943 20451
rect 12820 20448 12848 20556
rect 12894 20476 12900 20528
rect 12952 20516 12958 20528
rect 13817 20519 13875 20525
rect 13817 20516 13829 20519
rect 12952 20488 13829 20516
rect 12952 20476 12958 20488
rect 13817 20485 13829 20488
rect 13863 20516 13875 20519
rect 14090 20516 14096 20528
rect 13863 20488 14096 20516
rect 13863 20485 13875 20488
rect 13817 20479 13875 20485
rect 14090 20476 14096 20488
rect 14148 20476 14154 20528
rect 14458 20476 14464 20528
rect 14516 20476 14522 20528
rect 16040 20525 16068 20556
rect 16850 20544 16856 20596
rect 16908 20584 16914 20596
rect 17310 20584 17316 20596
rect 16908 20556 17316 20584
rect 16908 20544 16914 20556
rect 17310 20544 17316 20556
rect 17368 20544 17374 20596
rect 17586 20544 17592 20596
rect 17644 20544 17650 20596
rect 18233 20587 18291 20593
rect 18233 20553 18245 20587
rect 18279 20584 18291 20587
rect 18279 20556 19380 20584
rect 18279 20553 18291 20556
rect 18233 20547 18291 20553
rect 16025 20519 16083 20525
rect 16025 20485 16037 20519
rect 16071 20485 16083 20519
rect 16025 20479 16083 20485
rect 16390 20476 16396 20528
rect 16448 20516 16454 20528
rect 18138 20516 18144 20528
rect 16448 20488 18144 20516
rect 16448 20476 16454 20488
rect 18138 20476 18144 20488
rect 18196 20476 18202 20528
rect 18322 20476 18328 20528
rect 18380 20516 18386 20528
rect 18877 20519 18935 20525
rect 18877 20516 18889 20519
rect 18380 20488 18889 20516
rect 18380 20476 18386 20488
rect 18877 20485 18889 20488
rect 18923 20485 18935 20519
rect 19352 20516 19380 20556
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 20898 20584 20904 20596
rect 19484 20556 20904 20584
rect 19484 20544 19490 20556
rect 19352 20488 19472 20516
rect 18877 20479 18935 20485
rect 19444 20460 19472 20488
rect 11885 20411 11943 20417
rect 12406 20420 12848 20448
rect 10778 20380 10784 20392
rect 8772 20352 10784 20380
rect 6546 20312 6552 20324
rect 5552 20284 6552 20312
rect 5552 20244 5580 20284
rect 6546 20272 6552 20284
rect 6604 20272 6610 20324
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 8772 20312 8800 20352
rect 10778 20340 10784 20352
rect 10836 20380 10842 20392
rect 11054 20380 11060 20392
rect 10836 20352 11060 20380
rect 10836 20340 10842 20352
rect 11054 20340 11060 20352
rect 11112 20340 11118 20392
rect 11422 20340 11428 20392
rect 11480 20380 11486 20392
rect 12406 20380 12434 20420
rect 15470 20408 15476 20460
rect 15528 20448 15534 20460
rect 16209 20451 16267 20457
rect 16209 20448 16221 20451
rect 15528 20420 16221 20448
rect 15528 20408 15534 20420
rect 16209 20417 16221 20420
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 16298 20408 16304 20460
rect 16356 20448 16362 20460
rect 17218 20448 17224 20460
rect 16356 20420 17224 20448
rect 16356 20408 16362 20420
rect 17218 20408 17224 20420
rect 17276 20448 17282 20460
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 17276 20420 17509 20448
rect 17276 20408 17282 20420
rect 17497 20417 17509 20420
rect 17543 20417 17555 20451
rect 17497 20411 17555 20417
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 18598 20448 18604 20460
rect 17644 20420 18604 20448
rect 17644 20408 17650 20420
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 18966 20408 18972 20460
rect 19024 20408 19030 20460
rect 19426 20408 19432 20460
rect 19484 20408 19490 20460
rect 19720 20457 19748 20556
rect 20898 20544 20904 20556
rect 20956 20584 20962 20596
rect 22186 20584 22192 20596
rect 20956 20556 22192 20584
rect 20956 20544 20962 20556
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 23566 20544 23572 20596
rect 23624 20544 23630 20596
rect 24118 20544 24124 20596
rect 24176 20544 24182 20596
rect 26145 20587 26203 20593
rect 25135 20556 26004 20584
rect 25135 20528 25163 20556
rect 21634 20516 21640 20528
rect 21206 20488 21640 20516
rect 21634 20476 21640 20488
rect 21692 20516 21698 20528
rect 21818 20516 21824 20528
rect 21692 20488 21824 20516
rect 21692 20476 21698 20488
rect 21818 20476 21824 20488
rect 21876 20476 21882 20528
rect 23934 20516 23940 20528
rect 21928 20488 23940 20516
rect 19705 20451 19763 20457
rect 19705 20417 19717 20451
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 21266 20408 21272 20460
rect 21324 20448 21330 20460
rect 21928 20448 21956 20488
rect 23934 20476 23940 20488
rect 23992 20476 23998 20528
rect 25130 20476 25136 20528
rect 25188 20476 25194 20528
rect 25976 20516 26004 20556
rect 26145 20553 26157 20587
rect 26191 20584 26203 20587
rect 26191 20556 26740 20584
rect 26191 20553 26203 20556
rect 26145 20547 26203 20553
rect 26602 20516 26608 20528
rect 25976 20488 26608 20516
rect 26602 20476 26608 20488
rect 26660 20476 26666 20528
rect 26712 20516 26740 20556
rect 26786 20544 26792 20596
rect 26844 20544 26850 20596
rect 26896 20556 27384 20584
rect 26896 20516 26924 20556
rect 26712 20488 26924 20516
rect 26970 20476 26976 20528
rect 27028 20516 27034 20528
rect 27154 20516 27160 20528
rect 27028 20488 27160 20516
rect 27028 20476 27034 20488
rect 27154 20476 27160 20488
rect 27212 20476 27218 20528
rect 27356 20516 27384 20556
rect 27430 20544 27436 20596
rect 27488 20584 27494 20596
rect 34146 20584 34152 20596
rect 27488 20556 34152 20584
rect 27488 20544 27494 20556
rect 34146 20544 34152 20556
rect 34204 20544 34210 20596
rect 34606 20544 34612 20596
rect 34664 20544 34670 20596
rect 35529 20587 35587 20593
rect 35529 20553 35541 20587
rect 35575 20584 35587 20587
rect 35894 20584 35900 20596
rect 35575 20556 35900 20584
rect 35575 20553 35587 20556
rect 35529 20547 35587 20553
rect 35894 20544 35900 20556
rect 35952 20544 35958 20596
rect 36722 20544 36728 20596
rect 36780 20584 36786 20596
rect 36780 20556 38700 20584
rect 36780 20544 36786 20556
rect 27798 20516 27804 20528
rect 27356 20488 27804 20516
rect 27798 20476 27804 20488
rect 27856 20476 27862 20528
rect 29730 20476 29736 20528
rect 29788 20476 29794 20528
rect 31754 20476 31760 20528
rect 31812 20476 31818 20528
rect 36633 20519 36691 20525
rect 36633 20516 36645 20519
rect 32232 20488 36645 20516
rect 21324 20420 21956 20448
rect 21324 20408 21330 20420
rect 22002 20408 22008 20460
rect 22060 20408 22066 20460
rect 22186 20408 22192 20460
rect 22244 20448 22250 20460
rect 23477 20451 23535 20457
rect 22244 20420 22876 20448
rect 22244 20408 22250 20420
rect 11480 20352 12434 20380
rect 12805 20383 12863 20389
rect 11480 20340 11486 20352
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 12805 20343 12863 20349
rect 6788 20284 8800 20312
rect 6788 20272 6794 20284
rect 9950 20272 9956 20324
rect 10008 20312 10014 20324
rect 11149 20315 11207 20321
rect 11149 20312 11161 20315
rect 10008 20284 11161 20312
rect 10008 20272 10014 20284
rect 11149 20281 11161 20284
rect 11195 20281 11207 20315
rect 11149 20275 11207 20281
rect 4356 20216 5580 20244
rect 5718 20204 5724 20256
rect 5776 20244 5782 20256
rect 5902 20244 5908 20256
rect 5776 20216 5908 20244
rect 5776 20204 5782 20216
rect 5902 20204 5908 20216
rect 5960 20244 5966 20256
rect 8110 20244 8116 20256
rect 5960 20216 8116 20244
rect 5960 20204 5966 20216
rect 8110 20204 8116 20216
rect 8168 20204 8174 20256
rect 8386 20204 8392 20256
rect 8444 20204 8450 20256
rect 8570 20204 8576 20256
rect 8628 20244 8634 20256
rect 9306 20244 9312 20256
rect 8628 20216 9312 20244
rect 8628 20204 8634 20216
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9674 20204 9680 20256
rect 9732 20244 9738 20256
rect 10410 20244 10416 20256
rect 9732 20216 10416 20244
rect 9732 20204 9738 20216
rect 10410 20204 10416 20216
rect 10468 20204 10474 20256
rect 12820 20244 12848 20343
rect 12986 20340 12992 20392
rect 13044 20340 13050 20392
rect 13538 20340 13544 20392
rect 13596 20340 13602 20392
rect 15289 20383 15347 20389
rect 15289 20380 15301 20383
rect 13648 20352 15301 20380
rect 13004 20312 13032 20340
rect 13648 20312 13676 20352
rect 15289 20349 15301 20352
rect 15335 20380 15347 20383
rect 16482 20380 16488 20392
rect 15335 20352 16488 20380
rect 15335 20349 15347 20352
rect 15289 20343 15347 20349
rect 16482 20340 16488 20352
rect 16540 20340 16546 20392
rect 17681 20383 17739 20389
rect 17681 20380 17693 20383
rect 16592 20352 17693 20380
rect 16390 20312 16396 20324
rect 13004 20284 13676 20312
rect 15580 20284 16396 20312
rect 15580 20244 15608 20284
rect 16390 20272 16396 20284
rect 16448 20272 16454 20324
rect 16592 20312 16620 20352
rect 17681 20349 17693 20352
rect 17727 20349 17739 20383
rect 17681 20343 17739 20349
rect 16500 20284 16620 20312
rect 16500 20256 16528 20284
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17402 20312 17408 20324
rect 17000 20284 17408 20312
rect 17000 20272 17006 20284
rect 17402 20272 17408 20284
rect 17460 20272 17466 20324
rect 17696 20312 17724 20343
rect 17954 20340 17960 20392
rect 18012 20380 18018 20392
rect 18782 20380 18788 20392
rect 18012 20352 18788 20380
rect 18012 20340 18018 20352
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 19058 20340 19064 20392
rect 19116 20340 19122 20392
rect 19981 20383 20039 20389
rect 19981 20349 19993 20383
rect 20027 20380 20039 20383
rect 20530 20380 20536 20392
rect 20027 20352 20536 20380
rect 20027 20349 20039 20352
rect 19981 20343 20039 20349
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 21450 20340 21456 20392
rect 21508 20340 21514 20392
rect 22462 20340 22468 20392
rect 22520 20380 22526 20392
rect 22738 20380 22744 20392
rect 22520 20352 22744 20380
rect 22520 20340 22526 20352
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 22848 20389 22876 20420
rect 23477 20417 23489 20451
rect 23523 20448 23535 20451
rect 23566 20448 23572 20460
rect 23523 20420 23572 20448
rect 23523 20417 23535 20420
rect 23477 20411 23535 20417
rect 23566 20408 23572 20420
rect 23624 20408 23630 20460
rect 26510 20408 26516 20460
rect 26568 20448 26574 20460
rect 27525 20451 27583 20457
rect 27525 20448 27537 20451
rect 26568 20420 27537 20448
rect 26568 20408 26574 20420
rect 27525 20417 27537 20420
rect 27571 20448 27583 20451
rect 27571 20420 27752 20448
rect 27571 20417 27583 20420
rect 27525 20411 27583 20417
rect 22833 20383 22891 20389
rect 22833 20349 22845 20383
rect 22879 20380 22891 20383
rect 24397 20383 24455 20389
rect 24397 20380 24409 20383
rect 22879 20352 24409 20380
rect 22879 20349 22891 20352
rect 22833 20343 22891 20349
rect 24397 20349 24409 20352
rect 24443 20349 24455 20383
rect 24397 20343 24455 20349
rect 24673 20383 24731 20389
rect 24673 20349 24685 20383
rect 24719 20380 24731 20383
rect 27430 20380 27436 20392
rect 24719 20352 27436 20380
rect 24719 20349 24731 20352
rect 24673 20343 24731 20349
rect 27430 20340 27436 20352
rect 27488 20340 27494 20392
rect 27617 20383 27675 20389
rect 27617 20380 27629 20383
rect 27540 20352 27629 20380
rect 17862 20312 17868 20324
rect 17696 20284 17868 20312
rect 17862 20272 17868 20284
rect 17920 20272 17926 20324
rect 18138 20272 18144 20324
rect 18196 20312 18202 20324
rect 18966 20312 18972 20324
rect 18196 20284 18972 20312
rect 18196 20272 18202 20284
rect 18966 20272 18972 20284
rect 19024 20272 19030 20324
rect 21008 20284 21588 20312
rect 12820 20216 15608 20244
rect 15654 20204 15660 20256
rect 15712 20204 15718 20256
rect 16482 20204 16488 20256
rect 16540 20204 16546 20256
rect 17129 20247 17187 20253
rect 17129 20213 17141 20247
rect 17175 20244 17187 20247
rect 17678 20244 17684 20256
rect 17175 20216 17684 20244
rect 17175 20213 17187 20216
rect 17129 20207 17187 20213
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 18506 20204 18512 20256
rect 18564 20204 18570 20256
rect 19150 20204 19156 20256
rect 19208 20244 19214 20256
rect 21008 20244 21036 20284
rect 19208 20216 21036 20244
rect 21560 20244 21588 20284
rect 21634 20272 21640 20324
rect 21692 20312 21698 20324
rect 23382 20312 23388 20324
rect 21692 20284 23388 20312
rect 21692 20272 21698 20284
rect 23382 20272 23388 20284
rect 23440 20272 23446 20324
rect 27246 20272 27252 20324
rect 27304 20312 27310 20324
rect 27540 20312 27568 20352
rect 27617 20349 27629 20352
rect 27663 20349 27675 20383
rect 27617 20343 27675 20349
rect 27304 20284 27568 20312
rect 27304 20272 27310 20284
rect 22830 20244 22836 20256
rect 21560 20216 22836 20244
rect 19208 20204 19214 20216
rect 22830 20204 22836 20216
rect 22888 20204 22894 20256
rect 22922 20204 22928 20256
rect 22980 20244 22986 20256
rect 23658 20244 23664 20256
rect 22980 20216 23664 20244
rect 22980 20204 22986 20216
rect 23658 20204 23664 20216
rect 23716 20204 23722 20256
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 25406 20244 25412 20256
rect 24912 20216 25412 20244
rect 24912 20204 24918 20216
rect 25406 20204 25412 20216
rect 25464 20204 25470 20256
rect 27154 20204 27160 20256
rect 27212 20204 27218 20256
rect 27724 20244 27752 20420
rect 28442 20408 28448 20460
rect 28500 20408 28506 20460
rect 31018 20408 31024 20460
rect 31076 20408 31082 20460
rect 32232 20448 32260 20488
rect 36633 20485 36645 20488
rect 36679 20485 36691 20519
rect 36633 20479 36691 20485
rect 31220 20420 32260 20448
rect 27798 20340 27804 20392
rect 27856 20340 27862 20392
rect 28721 20383 28779 20389
rect 28721 20349 28733 20383
rect 28767 20380 28779 20383
rect 28767 20352 31064 20380
rect 28767 20349 28779 20352
rect 28721 20343 28779 20349
rect 30650 20272 30656 20324
rect 30708 20272 30714 20324
rect 31036 20312 31064 20352
rect 31110 20340 31116 20392
rect 31168 20340 31174 20392
rect 31220 20312 31248 20420
rect 32306 20408 32312 20460
rect 32364 20408 32370 20460
rect 33410 20408 33416 20460
rect 33468 20408 33474 20460
rect 34885 20451 34943 20457
rect 34885 20417 34897 20451
rect 34931 20448 34943 20451
rect 35526 20448 35532 20460
rect 34931 20420 35532 20448
rect 34931 20417 34943 20420
rect 34885 20411 34943 20417
rect 35526 20408 35532 20420
rect 35584 20408 35590 20460
rect 35986 20408 35992 20460
rect 36044 20408 36050 20460
rect 37366 20408 37372 20460
rect 37424 20448 37430 20460
rect 37737 20451 37795 20457
rect 37737 20448 37749 20451
rect 37424 20420 37749 20448
rect 37424 20408 37430 20420
rect 37737 20417 37749 20420
rect 37783 20417 37795 20451
rect 37737 20411 37795 20417
rect 31294 20340 31300 20392
rect 31352 20340 31358 20392
rect 34054 20340 34060 20392
rect 34112 20340 34118 20392
rect 34330 20340 34336 20392
rect 34388 20340 34394 20392
rect 36630 20340 36636 20392
rect 36688 20380 36694 20392
rect 37461 20383 37519 20389
rect 37461 20380 37473 20383
rect 36688 20352 37473 20380
rect 36688 20340 36694 20352
rect 37461 20349 37473 20352
rect 37507 20349 37519 20383
rect 38672 20380 38700 20556
rect 38764 20556 41644 20584
rect 38764 20457 38792 20556
rect 41506 20516 41512 20528
rect 40052 20488 41512 20516
rect 38749 20451 38807 20457
rect 38749 20417 38761 20451
rect 38795 20417 38807 20451
rect 38749 20411 38807 20417
rect 39022 20408 39028 20460
rect 39080 20408 39086 20460
rect 40052 20457 40080 20488
rect 41506 20476 41512 20488
rect 41564 20476 41570 20528
rect 41616 20516 41644 20556
rect 43438 20544 43444 20596
rect 43496 20544 43502 20596
rect 48866 20544 48872 20596
rect 48924 20584 48930 20596
rect 49421 20587 49479 20593
rect 49421 20584 49433 20587
rect 48924 20556 49433 20584
rect 48924 20544 48930 20556
rect 49421 20553 49433 20556
rect 49467 20553 49479 20587
rect 49421 20547 49479 20553
rect 44542 20516 44548 20528
rect 41616 20488 44548 20516
rect 44542 20476 44548 20488
rect 44600 20476 44606 20528
rect 49234 20476 49240 20528
rect 49292 20476 49298 20528
rect 40037 20451 40095 20457
rect 40037 20417 40049 20451
rect 40083 20417 40095 20451
rect 40037 20411 40095 20417
rect 40310 20408 40316 20460
rect 40368 20408 40374 20460
rect 41230 20408 41236 20460
rect 41288 20408 41294 20460
rect 42797 20451 42855 20457
rect 42797 20448 42809 20451
rect 41340 20420 42809 20448
rect 39482 20380 39488 20392
rect 38672 20352 39488 20380
rect 37461 20343 37519 20349
rect 39482 20340 39488 20352
rect 39540 20340 39546 20392
rect 41340 20312 41368 20420
rect 42797 20417 42809 20420
rect 42843 20448 42855 20451
rect 43073 20451 43131 20457
rect 43073 20448 43085 20451
rect 42843 20420 43085 20448
rect 42843 20417 42855 20420
rect 42797 20411 42855 20417
rect 43073 20417 43085 20420
rect 43119 20417 43131 20451
rect 43073 20411 43131 20417
rect 41414 20340 41420 20392
rect 41472 20380 41478 20392
rect 41509 20383 41567 20389
rect 41509 20380 41521 20383
rect 41472 20352 41521 20380
rect 41472 20340 41478 20352
rect 41509 20349 41521 20352
rect 41555 20349 41567 20383
rect 41509 20343 41567 20349
rect 31036 20284 31248 20312
rect 36832 20284 41368 20312
rect 29270 20244 29276 20256
rect 27724 20216 29276 20244
rect 29270 20204 29276 20216
rect 29328 20204 29334 20256
rect 29362 20204 29368 20256
rect 29420 20244 29426 20256
rect 30193 20247 30251 20253
rect 30193 20244 30205 20247
rect 29420 20216 30205 20244
rect 29420 20204 29426 20216
rect 30193 20213 30205 20216
rect 30239 20244 30251 20247
rect 31386 20244 31392 20256
rect 30239 20216 31392 20244
rect 30239 20213 30251 20216
rect 30193 20207 30251 20213
rect 31386 20204 31392 20216
rect 31444 20204 31450 20256
rect 31938 20204 31944 20256
rect 31996 20204 32002 20256
rect 32214 20204 32220 20256
rect 32272 20244 32278 20256
rect 32953 20247 33011 20253
rect 32953 20244 32965 20247
rect 32272 20216 32965 20244
rect 32272 20204 32278 20216
rect 32953 20213 32965 20216
rect 32999 20213 33011 20247
rect 32953 20207 33011 20213
rect 33042 20204 33048 20256
rect 33100 20244 33106 20256
rect 36832 20244 36860 20284
rect 42702 20272 42708 20324
rect 42760 20312 42766 20324
rect 43257 20315 43315 20321
rect 43257 20312 43269 20315
rect 42760 20284 43269 20312
rect 42760 20272 42766 20284
rect 43257 20281 43269 20284
rect 43303 20281 43315 20315
rect 43257 20275 43315 20281
rect 33100 20216 36860 20244
rect 33100 20204 33106 20216
rect 36998 20204 37004 20256
rect 37056 20204 37062 20256
rect 40586 20204 40592 20256
rect 40644 20244 40650 20256
rect 40773 20247 40831 20253
rect 40773 20244 40785 20247
rect 40644 20216 40785 20244
rect 40644 20204 40650 20216
rect 40773 20213 40785 20216
rect 40819 20213 40831 20247
rect 40773 20207 40831 20213
rect 40862 20204 40868 20256
rect 40920 20244 40926 20256
rect 42613 20247 42671 20253
rect 42613 20244 42625 20247
rect 40920 20216 42625 20244
rect 40920 20204 40926 20216
rect 42613 20213 42625 20216
rect 42659 20213 42671 20247
rect 42613 20207 42671 20213
rect 43622 20204 43628 20256
rect 43680 20204 43686 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 3605 20043 3663 20049
rect 3605 20009 3617 20043
rect 3651 20040 3663 20043
rect 3786 20040 3792 20052
rect 3651 20012 3792 20040
rect 3651 20009 3663 20012
rect 3605 20003 3663 20009
rect 3786 20000 3792 20012
rect 3844 20000 3850 20052
rect 3881 20043 3939 20049
rect 3881 20009 3893 20043
rect 3927 20040 3939 20043
rect 8570 20040 8576 20052
rect 3927 20012 8576 20040
rect 3927 20009 3939 20012
rect 3881 20003 3939 20009
rect 1486 19864 1492 19916
rect 1544 19904 1550 19916
rect 3988 19913 4016 20012
rect 8570 20000 8576 20012
rect 8628 20000 8634 20052
rect 9030 20000 9036 20052
rect 9088 20000 9094 20052
rect 9398 20000 9404 20052
rect 9456 20040 9462 20052
rect 12437 20043 12495 20049
rect 9456 20012 11376 20040
rect 9456 20000 9462 20012
rect 8110 19932 8116 19984
rect 8168 19972 8174 19984
rect 11348 19972 11376 20012
rect 12437 20009 12449 20043
rect 12483 20040 12495 20043
rect 12483 20012 16712 20040
rect 12483 20009 12495 20012
rect 12437 20003 12495 20009
rect 12713 19975 12771 19981
rect 12713 19972 12725 19975
rect 8168 19944 10180 19972
rect 11348 19944 12725 19972
rect 8168 19932 8174 19944
rect 2041 19907 2099 19913
rect 2041 19904 2053 19907
rect 1544 19876 2053 19904
rect 1544 19864 1550 19876
rect 2041 19873 2053 19876
rect 2087 19873 2099 19907
rect 2041 19867 2099 19873
rect 3973 19907 4031 19913
rect 3973 19873 3985 19907
rect 4019 19873 4031 19907
rect 6178 19904 6184 19916
rect 3973 19867 4031 19873
rect 4632 19876 6184 19904
rect 1026 19796 1032 19848
rect 1084 19836 1090 19848
rect 1581 19839 1639 19845
rect 1581 19836 1593 19839
rect 1084 19808 1593 19836
rect 1084 19796 1090 19808
rect 1581 19805 1593 19808
rect 1627 19805 1639 19839
rect 1581 19799 1639 19805
rect 3418 19796 3424 19848
rect 3476 19836 3482 19848
rect 4430 19836 4436 19848
rect 3476 19808 4436 19836
rect 3476 19796 3482 19808
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 4632 19845 4660 19876
rect 6178 19864 6184 19876
rect 6236 19864 6242 19916
rect 6546 19864 6552 19916
rect 6604 19904 6610 19916
rect 6825 19907 6883 19913
rect 6825 19904 6837 19907
rect 6604 19876 6837 19904
rect 6604 19864 6610 19876
rect 6825 19873 6837 19876
rect 6871 19904 6883 19907
rect 8662 19904 8668 19916
rect 6871 19876 8668 19904
rect 6871 19873 6883 19876
rect 6825 19867 6883 19873
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 10152 19904 10180 19944
rect 12713 19941 12725 19944
rect 12759 19941 12771 19975
rect 12713 19935 12771 19941
rect 12820 19944 13308 19972
rect 12820 19904 12848 19944
rect 10152 19876 12848 19904
rect 13170 19864 13176 19916
rect 13228 19864 13234 19916
rect 13280 19913 13308 19944
rect 14090 19932 14096 19984
rect 14148 19972 14154 19984
rect 14274 19972 14280 19984
rect 14148 19944 14280 19972
rect 14148 19932 14154 19944
rect 14274 19932 14280 19944
rect 14332 19932 14338 19984
rect 16684 19972 16712 20012
rect 16850 20000 16856 20052
rect 16908 20040 16914 20052
rect 17586 20040 17592 20052
rect 16908 20012 17592 20040
rect 16908 20000 16914 20012
rect 17586 20000 17592 20012
rect 17644 20000 17650 20052
rect 17770 20000 17776 20052
rect 17828 20040 17834 20052
rect 19150 20040 19156 20052
rect 17828 20012 19156 20040
rect 17828 20000 17834 20012
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19242 20000 19248 20052
rect 19300 20040 19306 20052
rect 19705 20043 19763 20049
rect 19705 20040 19717 20043
rect 19300 20012 19717 20040
rect 19300 20000 19306 20012
rect 19705 20009 19717 20012
rect 19751 20009 19763 20043
rect 20622 20040 20628 20052
rect 19705 20003 19763 20009
rect 20364 20012 20628 20040
rect 17678 19972 17684 19984
rect 16684 19944 17264 19972
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19873 13323 19907
rect 13265 19867 13323 19873
rect 13446 19864 13452 19916
rect 13504 19904 13510 19916
rect 15286 19904 15292 19916
rect 13504 19876 15292 19904
rect 13504 19864 13510 19876
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 15654 19864 15660 19916
rect 15712 19904 15718 19916
rect 16758 19904 16764 19916
rect 15712 19876 16764 19904
rect 15712 19864 15718 19876
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 17236 19904 17264 19944
rect 17512 19944 17684 19972
rect 17512 19913 17540 19944
rect 17678 19932 17684 19944
rect 17736 19932 17742 19984
rect 20364 19972 20392 20012
rect 20622 20000 20628 20012
rect 20680 20000 20686 20052
rect 20714 20000 20720 20052
rect 20772 20040 20778 20052
rect 22002 20040 22008 20052
rect 20772 20012 22008 20040
rect 20772 20000 20778 20012
rect 22002 20000 22008 20012
rect 22060 20040 22066 20052
rect 23937 20043 23995 20049
rect 23937 20040 23949 20043
rect 22060 20012 23949 20040
rect 22060 20000 22066 20012
rect 23937 20009 23949 20012
rect 23983 20040 23995 20043
rect 24946 20040 24952 20052
rect 23983 20012 24952 20040
rect 23983 20009 23995 20012
rect 23937 20003 23995 20009
rect 24946 20000 24952 20012
rect 25004 20000 25010 20052
rect 27154 20040 27160 20052
rect 25056 20012 27160 20040
rect 17880 19944 20392 19972
rect 17880 19916 17908 19944
rect 22278 19932 22284 19984
rect 22336 19932 22342 19984
rect 22557 19975 22615 19981
rect 22557 19941 22569 19975
rect 22603 19972 22615 19975
rect 23106 19972 23112 19984
rect 22603 19944 23112 19972
rect 22603 19941 22615 19944
rect 22557 19935 22615 19941
rect 23106 19932 23112 19944
rect 23164 19932 23170 19984
rect 25056 19972 25084 20012
rect 27154 20000 27160 20012
rect 27212 20000 27218 20052
rect 27617 20043 27675 20049
rect 27617 20009 27629 20043
rect 27663 20040 27675 20043
rect 27706 20040 27712 20052
rect 27663 20012 27712 20040
rect 27663 20009 27675 20012
rect 27617 20003 27675 20009
rect 27706 20000 27712 20012
rect 27764 20000 27770 20052
rect 28442 20000 28448 20052
rect 28500 20040 28506 20052
rect 28997 20043 29055 20049
rect 28997 20040 29009 20043
rect 28500 20012 29009 20040
rect 28500 20000 28506 20012
rect 28997 20009 29009 20012
rect 29043 20009 29055 20043
rect 28997 20003 29055 20009
rect 29546 20000 29552 20052
rect 29604 20040 29610 20052
rect 31386 20040 31392 20052
rect 29604 20012 31392 20040
rect 29604 20000 29610 20012
rect 31386 20000 31392 20012
rect 31444 20000 31450 20052
rect 31938 20000 31944 20052
rect 31996 20040 32002 20052
rect 32582 20040 32588 20052
rect 31996 20012 32588 20040
rect 31996 20000 32002 20012
rect 32582 20000 32588 20012
rect 32640 20000 32646 20052
rect 35526 20000 35532 20052
rect 35584 20000 35590 20052
rect 38841 20043 38899 20049
rect 38841 20009 38853 20043
rect 38887 20040 38899 20043
rect 40034 20040 40040 20052
rect 38887 20012 40040 20040
rect 38887 20009 38899 20012
rect 38841 20003 38899 20009
rect 40034 20000 40040 20012
rect 40092 20000 40098 20052
rect 40144 20012 41092 20040
rect 31573 19975 31631 19981
rect 31573 19972 31585 19975
rect 23308 19944 25084 19972
rect 29196 19944 31585 19972
rect 17497 19907 17555 19913
rect 17497 19904 17509 19907
rect 16868 19876 17080 19904
rect 17236 19876 17509 19904
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 3694 19728 3700 19780
rect 3752 19768 3758 19780
rect 4154 19768 4160 19780
rect 3752 19740 4160 19768
rect 3752 19728 3758 19740
rect 4154 19728 4160 19740
rect 4212 19728 4218 19780
rect 4632 19768 4660 19799
rect 9214 19796 9220 19848
rect 9272 19836 9278 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 9272 19808 9413 19836
rect 9272 19796 9278 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 10045 19839 10103 19845
rect 10045 19836 10057 19839
rect 9640 19808 10057 19836
rect 9640 19796 9646 19808
rect 10045 19805 10057 19808
rect 10091 19805 10103 19839
rect 10045 19799 10103 19805
rect 11698 19796 11704 19848
rect 11756 19836 11762 19848
rect 11756 19808 13768 19836
rect 11756 19796 11762 19808
rect 4798 19768 4804 19780
rect 4632 19740 4804 19768
rect 4798 19728 4804 19740
rect 4856 19728 4862 19780
rect 4893 19771 4951 19777
rect 4893 19737 4905 19771
rect 4939 19737 4951 19771
rect 6822 19768 6828 19780
rect 6118 19740 6828 19768
rect 4893 19731 4951 19737
rect 3418 19660 3424 19712
rect 3476 19660 3482 19712
rect 4246 19660 4252 19712
rect 4304 19700 4310 19712
rect 4908 19700 4936 19731
rect 6822 19728 6828 19740
rect 6880 19728 6886 19780
rect 7098 19728 7104 19780
rect 7156 19728 7162 19780
rect 7484 19740 7590 19768
rect 4304 19672 4936 19700
rect 4304 19660 4310 19672
rect 5626 19660 5632 19712
rect 5684 19700 5690 19712
rect 6178 19700 6184 19712
rect 5684 19672 6184 19700
rect 5684 19660 5690 19672
rect 6178 19660 6184 19672
rect 6236 19660 6242 19712
rect 6365 19703 6423 19709
rect 6365 19669 6377 19703
rect 6411 19700 6423 19703
rect 6454 19700 6460 19712
rect 6411 19672 6460 19700
rect 6411 19669 6423 19672
rect 6365 19663 6423 19669
rect 6454 19660 6460 19672
rect 6512 19660 6518 19712
rect 6730 19660 6736 19712
rect 6788 19700 6794 19712
rect 7484 19700 7512 19740
rect 8662 19728 8668 19780
rect 8720 19768 8726 19780
rect 9600 19768 9628 19796
rect 8720 19740 9628 19768
rect 8720 19728 8726 19740
rect 10318 19728 10324 19780
rect 10376 19728 10382 19780
rect 10778 19768 10784 19780
rect 10704 19740 10784 19768
rect 6788 19672 7512 19700
rect 6788 19660 6794 19672
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 8573 19703 8631 19709
rect 8573 19700 8585 19703
rect 7800 19672 8585 19700
rect 7800 19660 7806 19672
rect 8573 19669 8585 19672
rect 8619 19669 8631 19703
rect 8573 19663 8631 19669
rect 9122 19660 9128 19712
rect 9180 19700 9186 19712
rect 9493 19703 9551 19709
rect 9493 19700 9505 19703
rect 9180 19672 9505 19700
rect 9180 19660 9186 19672
rect 9493 19669 9505 19672
rect 9539 19669 9551 19703
rect 10704 19700 10732 19740
rect 10778 19728 10784 19740
rect 10836 19728 10842 19780
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 12802 19768 12808 19780
rect 11940 19740 12808 19768
rect 11940 19728 11946 19740
rect 12802 19728 12808 19740
rect 12860 19728 12866 19780
rect 13081 19771 13139 19777
rect 13081 19737 13093 19771
rect 13127 19768 13139 19771
rect 13740 19768 13768 19808
rect 13814 19796 13820 19848
rect 13872 19796 13878 19848
rect 14366 19796 14372 19848
rect 14424 19796 14430 19848
rect 16669 19839 16727 19845
rect 16669 19805 16681 19839
rect 16715 19836 16727 19839
rect 16868 19836 16896 19876
rect 16715 19808 16896 19836
rect 16715 19805 16727 19808
rect 16669 19799 16727 19805
rect 16942 19796 16948 19848
rect 17000 19796 17006 19848
rect 14642 19768 14648 19780
rect 13127 19740 13584 19768
rect 13740 19740 14648 19768
rect 13127 19737 13139 19740
rect 13081 19731 13139 19737
rect 11330 19700 11336 19712
rect 10704 19672 11336 19700
rect 9493 19663 9551 19669
rect 11330 19660 11336 19672
rect 11388 19660 11394 19712
rect 11793 19703 11851 19709
rect 11793 19669 11805 19703
rect 11839 19700 11851 19703
rect 12066 19700 12072 19712
rect 11839 19672 12072 19700
rect 11839 19669 11851 19672
rect 11793 19663 11851 19669
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 12253 19703 12311 19709
rect 12253 19669 12265 19703
rect 12299 19700 12311 19703
rect 13446 19700 13452 19712
rect 12299 19672 13452 19700
rect 12299 19669 12311 19672
rect 12253 19663 12311 19669
rect 13446 19660 13452 19672
rect 13504 19660 13510 19712
rect 13556 19700 13584 19740
rect 14642 19728 14648 19740
rect 14700 19728 14706 19780
rect 15028 19740 15134 19768
rect 13722 19700 13728 19712
rect 13556 19672 13728 19700
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 14458 19660 14464 19712
rect 14516 19700 14522 19712
rect 15028 19700 15056 19740
rect 15470 19700 15476 19712
rect 14516 19672 15476 19700
rect 14516 19660 14522 19672
rect 15470 19660 15476 19672
rect 15528 19660 15534 19712
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 16960 19709 16988 19796
rect 17052 19768 17080 19876
rect 17497 19873 17509 19876
rect 17543 19873 17555 19907
rect 17497 19867 17555 19873
rect 17862 19864 17868 19916
rect 17920 19864 17926 19916
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19904 18843 19907
rect 19058 19904 19064 19916
rect 18831 19876 19064 19904
rect 18831 19873 18843 19876
rect 18785 19867 18843 19873
rect 19058 19864 19064 19876
rect 19116 19904 19122 19916
rect 19518 19904 19524 19916
rect 19116 19876 19524 19904
rect 19116 19864 19122 19876
rect 19518 19864 19524 19876
rect 19576 19864 19582 19916
rect 20070 19864 20076 19916
rect 20128 19904 20134 19916
rect 23308 19913 23336 19944
rect 23293 19907 23351 19913
rect 20128 19876 23244 19904
rect 20128 19864 20134 19876
rect 17310 19796 17316 19848
rect 17368 19796 17374 19848
rect 17402 19796 17408 19848
rect 17460 19796 17466 19848
rect 19610 19836 19616 19848
rect 17696 19808 19616 19836
rect 17696 19768 17724 19808
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 20254 19796 20260 19848
rect 20312 19796 20318 19848
rect 23216 19845 23244 19876
rect 23293 19873 23305 19907
rect 23339 19873 23351 19907
rect 23293 19867 23351 19873
rect 23477 19907 23535 19913
rect 23477 19873 23489 19907
rect 23523 19904 23535 19907
rect 23523 19876 25084 19904
rect 23523 19873 23535 19876
rect 23477 19867 23535 19873
rect 23201 19839 23259 19845
rect 22756 19808 23060 19836
rect 17052 19740 17724 19768
rect 17770 19728 17776 19780
rect 17828 19768 17834 19780
rect 19794 19768 19800 19780
rect 17828 19740 19800 19768
rect 17828 19728 17834 19740
rect 19794 19728 19800 19740
rect 19852 19728 19858 19780
rect 20530 19728 20536 19780
rect 20588 19728 20594 19780
rect 20990 19728 20996 19780
rect 21048 19728 21054 19780
rect 22756 19768 22784 19808
rect 22020 19740 22784 19768
rect 16117 19703 16175 19709
rect 16117 19700 16129 19703
rect 15712 19672 16129 19700
rect 15712 19660 15718 19672
rect 16117 19669 16129 19672
rect 16163 19669 16175 19703
rect 16117 19663 16175 19669
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 17402 19660 17408 19712
rect 17460 19700 17466 19712
rect 18141 19703 18199 19709
rect 18141 19700 18153 19703
rect 17460 19672 18153 19700
rect 17460 19660 17466 19672
rect 18141 19669 18153 19672
rect 18187 19669 18199 19703
rect 18141 19663 18199 19669
rect 18506 19660 18512 19712
rect 18564 19660 18570 19712
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 21174 19700 21180 19712
rect 18647 19672 21180 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 21174 19660 21180 19672
rect 21232 19660 21238 19712
rect 22020 19709 22048 19740
rect 22005 19703 22063 19709
rect 22005 19669 22017 19703
rect 22051 19669 22063 19703
rect 22005 19663 22063 19669
rect 22370 19660 22376 19712
rect 22428 19700 22434 19712
rect 22833 19703 22891 19709
rect 22833 19700 22845 19703
rect 22428 19672 22845 19700
rect 22428 19660 22434 19672
rect 22833 19669 22845 19672
rect 22879 19669 22891 19703
rect 23032 19700 23060 19808
rect 23201 19805 23213 19839
rect 23247 19805 23259 19839
rect 23201 19799 23259 19805
rect 25056 19768 25084 19876
rect 25222 19864 25228 19916
rect 25280 19864 25286 19916
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19904 26203 19907
rect 29196 19904 29224 19944
rect 31573 19941 31585 19944
rect 31619 19941 31631 19975
rect 31573 19935 31631 19941
rect 33134 19932 33140 19984
rect 33192 19972 33198 19984
rect 40144 19972 40172 20012
rect 33192 19944 40172 19972
rect 40313 19975 40371 19981
rect 33192 19932 33198 19944
rect 40313 19941 40325 19975
rect 40359 19972 40371 19975
rect 40954 19972 40960 19984
rect 40359 19944 40960 19972
rect 40359 19941 40371 19944
rect 40313 19935 40371 19941
rect 40954 19932 40960 19944
rect 41012 19932 41018 19984
rect 41064 19972 41092 20012
rect 41230 20000 41236 20052
rect 41288 20040 41294 20052
rect 41969 20043 42027 20049
rect 41969 20040 41981 20043
rect 41288 20012 41981 20040
rect 41288 20000 41294 20012
rect 41969 20009 41981 20012
rect 42015 20009 42027 20043
rect 41969 20003 42027 20009
rect 42150 20000 42156 20052
rect 42208 20040 42214 20052
rect 42337 20043 42395 20049
rect 42337 20040 42349 20043
rect 42208 20012 42349 20040
rect 42208 20000 42214 20012
rect 42337 20009 42349 20012
rect 42383 20009 42395 20043
rect 42337 20003 42395 20009
rect 46750 19972 46756 19984
rect 41064 19944 46756 19972
rect 46750 19932 46756 19944
rect 46808 19932 46814 19984
rect 26191 19876 29224 19904
rect 29365 19907 29423 19913
rect 26191 19873 26203 19876
rect 26145 19867 26203 19873
rect 29365 19873 29377 19907
rect 29411 19904 29423 19907
rect 29822 19904 29828 19916
rect 29411 19876 29828 19904
rect 29411 19873 29423 19876
rect 29365 19867 29423 19873
rect 29822 19864 29828 19876
rect 29880 19864 29886 19916
rect 30282 19864 30288 19916
rect 30340 19864 30346 19916
rect 31018 19864 31024 19916
rect 31076 19904 31082 19916
rect 31849 19907 31907 19913
rect 31849 19904 31861 19907
rect 31076 19876 31861 19904
rect 31076 19864 31082 19876
rect 31849 19873 31861 19876
rect 31895 19873 31907 19907
rect 34054 19904 34060 19916
rect 31849 19867 31907 19873
rect 32324 19876 34060 19904
rect 25133 19839 25191 19845
rect 25133 19805 25145 19839
rect 25179 19836 25191 19839
rect 25314 19836 25320 19848
rect 25179 19808 25320 19836
rect 25179 19805 25191 19808
rect 25133 19799 25191 19805
rect 25314 19796 25320 19808
rect 25372 19796 25378 19848
rect 25774 19796 25780 19848
rect 25832 19836 25838 19848
rect 25869 19839 25927 19845
rect 25869 19836 25881 19839
rect 25832 19808 25881 19836
rect 25832 19796 25838 19808
rect 25869 19805 25881 19808
rect 25915 19805 25927 19839
rect 25869 19799 25927 19805
rect 28077 19839 28135 19845
rect 28077 19805 28089 19839
rect 28123 19836 28135 19839
rect 30098 19836 30104 19848
rect 28123 19808 30104 19836
rect 28123 19805 28135 19808
rect 28077 19799 28135 19805
rect 30098 19796 30104 19808
rect 30156 19796 30162 19848
rect 30929 19839 30987 19845
rect 30929 19805 30941 19839
rect 30975 19836 30987 19839
rect 32214 19836 32220 19848
rect 30975 19808 32220 19836
rect 30975 19805 30987 19808
rect 30929 19799 30987 19805
rect 32214 19796 32220 19808
rect 32272 19796 32278 19848
rect 32324 19845 32352 19876
rect 34054 19864 34060 19876
rect 34112 19864 34118 19916
rect 46658 19904 46664 19916
rect 34164 19876 46664 19904
rect 32309 19839 32367 19845
rect 32309 19805 32321 19839
rect 32355 19805 32367 19839
rect 32309 19799 32367 19805
rect 32953 19839 33011 19845
rect 32953 19805 32965 19839
rect 32999 19836 33011 19839
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 32999 19808 33425 19836
rect 32999 19805 33011 19808
rect 32953 19799 33011 19805
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 25056 19740 26556 19768
rect 23842 19700 23848 19712
rect 23032 19672 23848 19700
rect 22833 19663 22891 19669
rect 23842 19660 23848 19672
rect 23900 19660 23906 19712
rect 24213 19703 24271 19709
rect 24213 19669 24225 19703
rect 24259 19700 24271 19703
rect 24302 19700 24308 19712
rect 24259 19672 24308 19700
rect 24259 19669 24271 19672
rect 24213 19663 24271 19669
rect 24302 19660 24308 19672
rect 24360 19660 24366 19712
rect 24670 19660 24676 19712
rect 24728 19660 24734 19712
rect 25038 19660 25044 19712
rect 25096 19660 25102 19712
rect 26528 19700 26556 19740
rect 26602 19728 26608 19780
rect 26660 19728 26666 19780
rect 27430 19728 27436 19780
rect 27488 19768 27494 19780
rect 28721 19771 28779 19777
rect 28721 19768 28733 19771
rect 27488 19740 28733 19768
rect 27488 19728 27494 19740
rect 28721 19737 28733 19740
rect 28767 19737 28779 19771
rect 30466 19768 30472 19780
rect 28721 19731 28779 19737
rect 29288 19740 30472 19768
rect 27154 19700 27160 19712
rect 26528 19672 27160 19700
rect 27154 19660 27160 19672
rect 27212 19700 27218 19712
rect 29288 19700 29316 19740
rect 30466 19728 30472 19740
rect 30524 19728 30530 19780
rect 30558 19728 30564 19780
rect 30616 19768 30622 19780
rect 33042 19768 33048 19780
rect 30616 19740 33048 19768
rect 30616 19728 30622 19740
rect 33042 19728 33048 19740
rect 33100 19728 33106 19780
rect 34164 19768 34192 19876
rect 46658 19864 46664 19876
rect 46716 19864 46722 19916
rect 34422 19796 34428 19848
rect 34480 19836 34486 19848
rect 34885 19839 34943 19845
rect 34885 19836 34897 19839
rect 34480 19808 34897 19836
rect 34480 19796 34486 19808
rect 34885 19805 34897 19808
rect 34931 19805 34943 19839
rect 35989 19839 36047 19845
rect 35989 19836 36001 19839
rect 34885 19799 34943 19805
rect 35176 19808 36001 19836
rect 33152 19740 34192 19768
rect 27212 19672 29316 19700
rect 27212 19660 27218 19672
rect 29362 19660 29368 19712
rect 29420 19700 29426 19712
rect 29733 19703 29791 19709
rect 29733 19700 29745 19703
rect 29420 19672 29745 19700
rect 29420 19660 29426 19672
rect 29733 19669 29745 19672
rect 29779 19669 29791 19703
rect 29733 19663 29791 19669
rect 29822 19660 29828 19712
rect 29880 19700 29886 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 29880 19672 30113 19700
rect 29880 19660 29886 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 30101 19663 30159 19669
rect 30190 19660 30196 19712
rect 30248 19660 30254 19712
rect 30926 19660 30932 19712
rect 30984 19700 30990 19712
rect 32122 19700 32128 19712
rect 30984 19672 32128 19700
rect 30984 19660 30990 19672
rect 32122 19660 32128 19672
rect 32180 19660 32186 19712
rect 32214 19660 32220 19712
rect 32272 19700 32278 19712
rect 33152 19700 33180 19740
rect 35176 19712 35204 19808
rect 35989 19805 36001 19808
rect 36035 19805 36047 19839
rect 35989 19799 36047 19805
rect 37090 19796 37096 19848
rect 37148 19796 37154 19848
rect 38197 19839 38255 19845
rect 38197 19836 38209 19839
rect 37200 19808 38209 19836
rect 36998 19728 37004 19780
rect 37056 19768 37062 19780
rect 37200 19768 37228 19808
rect 38197 19805 38209 19808
rect 38243 19805 38255 19839
rect 38197 19799 38255 19805
rect 39390 19796 39396 19848
rect 39448 19836 39454 19848
rect 39485 19839 39543 19845
rect 39485 19836 39497 19839
rect 39448 19808 39497 19836
rect 39448 19796 39454 19808
rect 39485 19805 39497 19808
rect 39531 19805 39543 19839
rect 39485 19799 39543 19805
rect 40862 19796 40868 19848
rect 40920 19796 40926 19848
rect 41690 19796 41696 19848
rect 41748 19836 41754 19848
rect 42153 19839 42211 19845
rect 42153 19836 42165 19839
rect 41748 19808 42165 19836
rect 41748 19796 41754 19808
rect 42153 19805 42165 19808
rect 42199 19805 42211 19839
rect 42153 19799 42211 19805
rect 37056 19740 37228 19768
rect 37056 19728 37062 19740
rect 37642 19728 37648 19780
rect 37700 19768 37706 19780
rect 38562 19768 38568 19780
rect 37700 19740 38568 19768
rect 37700 19728 37706 19740
rect 38562 19728 38568 19740
rect 38620 19728 38626 19780
rect 40129 19771 40187 19777
rect 40129 19737 40141 19771
rect 40175 19768 40187 19771
rect 40586 19768 40592 19780
rect 40175 19740 40592 19768
rect 40175 19737 40187 19740
rect 40129 19731 40187 19737
rect 40586 19728 40592 19740
rect 40644 19728 40650 19780
rect 32272 19672 33180 19700
rect 32272 19660 32278 19672
rect 34054 19660 34060 19712
rect 34112 19660 34118 19712
rect 34517 19703 34575 19709
rect 34517 19669 34529 19703
rect 34563 19700 34575 19703
rect 35158 19700 35164 19712
rect 34563 19672 35164 19700
rect 34563 19669 34575 19672
rect 34517 19663 34575 19669
rect 35158 19660 35164 19672
rect 35216 19660 35222 19712
rect 35986 19660 35992 19712
rect 36044 19700 36050 19712
rect 36633 19703 36691 19709
rect 36633 19700 36645 19703
rect 36044 19672 36645 19700
rect 36044 19660 36050 19672
rect 36633 19669 36645 19672
rect 36679 19669 36691 19703
rect 36633 19663 36691 19669
rect 37550 19660 37556 19712
rect 37608 19700 37614 19712
rect 37737 19703 37795 19709
rect 37737 19700 37749 19703
rect 37608 19672 37749 19700
rect 37608 19660 37614 19672
rect 37737 19669 37749 19672
rect 37783 19669 37795 19703
rect 37737 19663 37795 19669
rect 38654 19660 38660 19712
rect 38712 19700 38718 19712
rect 39301 19703 39359 19709
rect 39301 19700 39313 19703
rect 38712 19672 39313 19700
rect 38712 19660 38718 19672
rect 39301 19669 39313 19672
rect 39347 19669 39359 19703
rect 39301 19663 39359 19669
rect 40954 19660 40960 19712
rect 41012 19660 41018 19712
rect 41509 19703 41567 19709
rect 41509 19669 41521 19703
rect 41555 19700 41567 19703
rect 41598 19700 41604 19712
rect 41555 19672 41604 19700
rect 41555 19669 41567 19672
rect 41509 19663 41567 19669
rect 41598 19660 41604 19672
rect 41656 19660 41662 19712
rect 42518 19660 42524 19712
rect 42576 19660 42582 19712
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 5261 19499 5319 19505
rect 5261 19496 5273 19499
rect 2746 19468 5273 19496
rect 658 19388 664 19440
rect 716 19428 722 19440
rect 2746 19428 2774 19468
rect 5261 19465 5273 19468
rect 5307 19465 5319 19499
rect 5261 19459 5319 19465
rect 5718 19456 5724 19508
rect 5776 19456 5782 19508
rect 6178 19456 6184 19508
rect 6236 19496 6242 19508
rect 6730 19496 6736 19508
rect 6236 19468 6736 19496
rect 6236 19456 6242 19468
rect 6730 19456 6736 19468
rect 6788 19456 6794 19508
rect 7190 19456 7196 19508
rect 7248 19496 7254 19508
rect 7650 19496 7656 19508
rect 7248 19468 7656 19496
rect 7248 19456 7254 19468
rect 7650 19456 7656 19468
rect 7708 19496 7714 19508
rect 9122 19496 9128 19508
rect 7708 19468 9128 19496
rect 7708 19456 7714 19468
rect 9122 19456 9128 19468
rect 9180 19456 9186 19508
rect 9217 19499 9275 19505
rect 9217 19465 9229 19499
rect 9263 19465 9275 19499
rect 9217 19459 9275 19465
rect 716 19400 2774 19428
rect 716 19388 722 19400
rect 3694 19388 3700 19440
rect 3752 19428 3758 19440
rect 3970 19428 3976 19440
rect 3752 19400 3976 19428
rect 3752 19388 3758 19400
rect 3970 19388 3976 19400
rect 4028 19388 4034 19440
rect 4338 19388 4344 19440
rect 4396 19388 4402 19440
rect 5552 19400 5856 19428
rect 1765 19363 1823 19369
rect 1765 19329 1777 19363
rect 1811 19360 1823 19363
rect 2130 19360 2136 19372
rect 1811 19332 2136 19360
rect 1811 19329 1823 19332
rect 1765 19323 1823 19329
rect 2130 19320 2136 19332
rect 2188 19320 2194 19372
rect 3605 19363 3663 19369
rect 3605 19329 3617 19363
rect 3651 19360 3663 19363
rect 4614 19360 4620 19372
rect 3651 19332 4620 19360
rect 3651 19329 3663 19332
rect 3605 19323 3663 19329
rect 4614 19320 4620 19332
rect 4672 19320 4678 19372
rect 2038 19252 2044 19304
rect 2096 19252 2102 19304
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 5552 19292 5580 19400
rect 5629 19363 5687 19369
rect 5629 19329 5641 19363
rect 5675 19360 5687 19363
rect 5828 19360 5856 19400
rect 6362 19388 6368 19440
rect 6420 19428 6426 19440
rect 6825 19431 6883 19437
rect 6825 19428 6837 19431
rect 6420 19400 6837 19428
rect 6420 19388 6426 19400
rect 6825 19397 6837 19400
rect 6871 19397 6883 19431
rect 6825 19391 6883 19397
rect 7558 19388 7564 19440
rect 7616 19388 7622 19440
rect 9232 19428 9260 19459
rect 9490 19456 9496 19508
rect 9548 19496 9554 19508
rect 9585 19499 9643 19505
rect 9585 19496 9597 19499
rect 9548 19468 9597 19496
rect 9548 19456 9554 19468
rect 9585 19465 9597 19468
rect 9631 19465 9643 19499
rect 9585 19459 9643 19465
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19496 10471 19499
rect 10594 19496 10600 19508
rect 10459 19468 10600 19496
rect 10459 19465 10471 19468
rect 10413 19459 10471 19465
rect 10594 19456 10600 19468
rect 10652 19456 10658 19508
rect 10686 19456 10692 19508
rect 10744 19496 10750 19508
rect 10781 19499 10839 19505
rect 10781 19496 10793 19499
rect 10744 19468 10793 19496
rect 10744 19456 10750 19468
rect 10781 19465 10793 19468
rect 10827 19465 10839 19499
rect 17589 19499 17647 19505
rect 17589 19496 17601 19499
rect 10781 19459 10839 19465
rect 11716 19468 17601 19496
rect 9232 19400 11652 19428
rect 5675 19332 5764 19360
rect 5828 19332 5948 19360
rect 5675 19329 5687 19332
rect 5629 19323 5687 19329
rect 5736 19292 5764 19332
rect 2924 19264 5580 19292
rect 5644 19264 5764 19292
rect 5813 19295 5871 19301
rect 2924 19252 2930 19264
rect 2130 19116 2136 19168
rect 2188 19156 2194 19168
rect 5077 19159 5135 19165
rect 5077 19156 5089 19159
rect 2188 19128 5089 19156
rect 2188 19116 2194 19128
rect 5077 19125 5089 19128
rect 5123 19156 5135 19159
rect 5644 19156 5672 19264
rect 5813 19261 5825 19295
rect 5859 19261 5871 19295
rect 5920 19292 5948 19332
rect 6546 19320 6552 19372
rect 6604 19320 6610 19372
rect 8757 19363 8815 19369
rect 8757 19329 8769 19363
rect 8803 19360 8815 19363
rect 10318 19360 10324 19372
rect 8803 19332 10324 19360
rect 8803 19329 8815 19332
rect 8757 19323 8815 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 11514 19360 11520 19372
rect 10919 19332 11520 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 7834 19292 7840 19304
rect 5920 19264 7840 19292
rect 5813 19255 5871 19261
rect 5828 19224 5856 19255
rect 7834 19252 7840 19264
rect 7892 19252 7898 19304
rect 9122 19252 9128 19304
rect 9180 19292 9186 19304
rect 9677 19295 9735 19301
rect 9677 19292 9689 19295
rect 9180 19264 9689 19292
rect 9180 19252 9186 19264
rect 9677 19261 9689 19264
rect 9723 19261 9735 19295
rect 9677 19255 9735 19261
rect 9858 19252 9864 19304
rect 9916 19252 9922 19304
rect 10778 19252 10784 19304
rect 10836 19292 10842 19304
rect 10965 19295 11023 19301
rect 10965 19292 10977 19295
rect 10836 19264 10977 19292
rect 10836 19252 10842 19264
rect 10965 19261 10977 19264
rect 11011 19261 11023 19295
rect 11624 19292 11652 19400
rect 11716 19369 11744 19468
rect 17589 19465 17601 19468
rect 17635 19465 17647 19499
rect 17589 19459 17647 19465
rect 17696 19468 17816 19496
rect 11974 19388 11980 19440
rect 12032 19428 12038 19440
rect 12032 19400 12940 19428
rect 12032 19388 12038 19400
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11701 19323 11759 19329
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12345 19363 12403 19369
rect 12345 19360 12357 19363
rect 11940 19332 12357 19360
rect 11940 19320 11946 19332
rect 12345 19329 12357 19332
rect 12391 19329 12403 19363
rect 12345 19323 12403 19329
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12805 19363 12863 19369
rect 12805 19360 12817 19363
rect 12492 19332 12817 19360
rect 12492 19320 12498 19332
rect 12805 19329 12817 19332
rect 12851 19329 12863 19363
rect 12912 19360 12940 19400
rect 13538 19388 13544 19440
rect 13596 19388 13602 19440
rect 14737 19431 14795 19437
rect 14737 19397 14749 19431
rect 14783 19428 14795 19431
rect 16206 19428 16212 19440
rect 14783 19400 16212 19428
rect 14783 19397 14795 19400
rect 14737 19391 14795 19397
rect 16206 19388 16212 19400
rect 16264 19388 16270 19440
rect 16298 19388 16304 19440
rect 16356 19428 16362 19440
rect 17696 19428 17724 19468
rect 17788 19440 17816 19468
rect 18782 19456 18788 19508
rect 18840 19496 18846 19508
rect 19245 19499 19303 19505
rect 19245 19496 19257 19499
rect 18840 19468 19257 19496
rect 18840 19456 18846 19468
rect 19245 19465 19257 19468
rect 19291 19465 19303 19499
rect 19245 19459 19303 19465
rect 20346 19456 20352 19508
rect 20404 19456 20410 19508
rect 21450 19456 21456 19508
rect 21508 19456 21514 19508
rect 21910 19456 21916 19508
rect 21968 19496 21974 19508
rect 22005 19499 22063 19505
rect 22005 19496 22017 19499
rect 21968 19468 22017 19496
rect 21968 19456 21974 19468
rect 22005 19465 22017 19468
rect 22051 19465 22063 19499
rect 22005 19459 22063 19465
rect 22465 19499 22523 19505
rect 22465 19465 22477 19499
rect 22511 19496 22523 19499
rect 23290 19496 23296 19508
rect 22511 19468 23296 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 23290 19456 23296 19468
rect 23348 19456 23354 19508
rect 23474 19456 23480 19508
rect 23532 19496 23538 19508
rect 23753 19499 23811 19505
rect 23753 19496 23765 19499
rect 23532 19468 23765 19496
rect 23532 19456 23538 19468
rect 23753 19465 23765 19468
rect 23799 19465 23811 19499
rect 23753 19459 23811 19465
rect 24118 19456 24124 19508
rect 24176 19496 24182 19508
rect 24176 19468 24808 19496
rect 24176 19456 24182 19468
rect 16356 19400 17724 19428
rect 16356 19388 16362 19400
rect 17770 19388 17776 19440
rect 17828 19388 17834 19440
rect 19150 19388 19156 19440
rect 19208 19428 19214 19440
rect 20364 19428 20392 19456
rect 19208 19400 20392 19428
rect 19208 19388 19214 19400
rect 20990 19388 20996 19440
rect 21048 19388 21054 19440
rect 21266 19388 21272 19440
rect 21324 19428 21330 19440
rect 24670 19428 24676 19440
rect 21324 19400 24676 19428
rect 21324 19388 21330 19400
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 24780 19428 24808 19468
rect 24854 19456 24860 19508
rect 24912 19496 24918 19508
rect 27157 19499 27215 19505
rect 27157 19496 27169 19499
rect 24912 19468 27169 19496
rect 24912 19456 24918 19468
rect 27157 19465 27169 19468
rect 27203 19465 27215 19499
rect 27157 19459 27215 19465
rect 27525 19499 27583 19505
rect 27525 19465 27537 19499
rect 27571 19496 27583 19499
rect 29638 19496 29644 19508
rect 27571 19468 29644 19496
rect 27571 19465 27583 19468
rect 27525 19459 27583 19465
rect 29638 19456 29644 19468
rect 29696 19456 29702 19508
rect 30101 19499 30159 19505
rect 30101 19465 30113 19499
rect 30147 19465 30159 19499
rect 30101 19459 30159 19465
rect 31205 19499 31263 19505
rect 31205 19465 31217 19499
rect 31251 19496 31263 19499
rect 32306 19496 32312 19508
rect 31251 19468 32312 19496
rect 31251 19465 31263 19468
rect 31205 19459 31263 19465
rect 24780 19400 24900 19428
rect 14645 19363 14703 19369
rect 14645 19360 14657 19363
rect 12912 19332 14657 19360
rect 12805 19323 12863 19329
rect 14645 19329 14657 19332
rect 14691 19329 14703 19363
rect 14918 19360 14924 19372
rect 14645 19323 14703 19329
rect 14752 19332 14924 19360
rect 11974 19292 11980 19304
rect 11624 19264 11980 19292
rect 10965 19255 11023 19261
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12250 19252 12256 19304
rect 12308 19292 12314 19304
rect 14752 19292 14780 19332
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 15286 19320 15292 19372
rect 15344 19360 15350 19372
rect 15841 19363 15899 19369
rect 15841 19360 15853 19363
rect 15344 19332 15853 19360
rect 15344 19320 15350 19332
rect 15841 19329 15853 19332
rect 15887 19329 15899 19363
rect 15841 19323 15899 19329
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17586 19360 17592 19372
rect 16991 19332 17592 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17586 19320 17592 19332
rect 17644 19320 17650 19372
rect 17696 19332 18080 19360
rect 17696 19304 17724 19332
rect 12308 19264 14780 19292
rect 12308 19252 12314 19264
rect 14826 19252 14832 19304
rect 14884 19252 14890 19304
rect 15930 19252 15936 19304
rect 15988 19252 15994 19304
rect 16022 19252 16028 19304
rect 16080 19252 16086 19304
rect 16114 19252 16120 19304
rect 16172 19292 16178 19304
rect 17494 19292 17500 19304
rect 16172 19264 17500 19292
rect 16172 19252 16178 19264
rect 17494 19252 17500 19264
rect 17552 19252 17558 19304
rect 17678 19252 17684 19304
rect 17736 19252 17742 19304
rect 17954 19252 17960 19304
rect 18012 19252 18018 19304
rect 6086 19224 6092 19236
rect 5828 19196 6092 19224
rect 6086 19184 6092 19196
rect 6144 19184 6150 19236
rect 7852 19224 7880 19252
rect 11606 19224 11612 19236
rect 7852 19196 11612 19224
rect 11606 19184 11612 19196
rect 11664 19184 11670 19236
rect 13814 19224 13820 19236
rect 12268 19196 13820 19224
rect 5123 19128 5672 19156
rect 6104 19156 6132 19184
rect 8297 19159 8355 19165
rect 8297 19156 8309 19159
rect 6104 19128 8309 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 8297 19125 8309 19128
rect 8343 19125 8355 19159
rect 8297 19119 8355 19125
rect 8938 19116 8944 19168
rect 8996 19116 9002 19168
rect 9490 19116 9496 19168
rect 9548 19156 9554 19168
rect 12268 19156 12296 19196
rect 13814 19184 13820 19196
rect 13872 19184 13878 19236
rect 14274 19184 14280 19236
rect 14332 19184 14338 19236
rect 17972 19224 18000 19252
rect 14384 19196 18000 19224
rect 9548 19128 12296 19156
rect 9548 19116 9554 19128
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 14384 19156 14412 19196
rect 12584 19128 14412 19156
rect 15473 19159 15531 19165
rect 12584 19116 12590 19128
rect 15473 19125 15485 19159
rect 15519 19156 15531 19159
rect 16666 19156 16672 19168
rect 15519 19128 16672 19156
rect 15519 19125 15531 19128
rect 15473 19119 15531 19125
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 17862 19156 17868 19168
rect 16816 19128 17868 19156
rect 16816 19116 16822 19128
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 18052 19165 18080 19332
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 19610 19360 19616 19372
rect 18472 19332 19616 19360
rect 18472 19320 18478 19332
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 19702 19320 19708 19372
rect 19760 19320 19766 19372
rect 22370 19320 22376 19372
rect 22428 19320 22434 19372
rect 22572 19332 22876 19360
rect 18230 19252 18236 19304
rect 18288 19252 18294 19304
rect 18509 19295 18567 19301
rect 18509 19261 18521 19295
rect 18555 19261 18567 19295
rect 18509 19255 18567 19261
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19292 18659 19295
rect 18782 19292 18788 19304
rect 18647 19264 18788 19292
rect 18647 19261 18659 19264
rect 18601 19255 18659 19261
rect 18049 19159 18107 19165
rect 18049 19125 18061 19159
rect 18095 19125 18107 19159
rect 18248 19156 18276 19252
rect 18524 19224 18552 19255
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 18892 19264 19993 19292
rect 18690 19224 18696 19236
rect 18524 19196 18696 19224
rect 18690 19184 18696 19196
rect 18748 19184 18754 19236
rect 18892 19156 18920 19264
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 21358 19252 21364 19304
rect 21416 19292 21422 19304
rect 22572 19292 22600 19332
rect 21416 19264 22600 19292
rect 22649 19295 22707 19301
rect 21416 19252 21422 19264
rect 22649 19261 22661 19295
rect 22695 19292 22707 19295
rect 22738 19292 22744 19304
rect 22695 19264 22744 19292
rect 22695 19261 22707 19264
rect 22649 19255 22707 19261
rect 22738 19252 22744 19264
rect 22796 19252 22802 19304
rect 22848 19292 22876 19332
rect 22922 19320 22928 19372
rect 22980 19360 22986 19372
rect 24118 19360 24124 19372
rect 22980 19332 24124 19360
rect 22980 19320 22986 19332
rect 24118 19320 24124 19332
rect 24176 19320 24182 19372
rect 24213 19363 24271 19369
rect 24213 19329 24225 19363
rect 24259 19360 24271 19363
rect 24872 19360 24900 19400
rect 24946 19388 24952 19440
rect 25004 19388 25010 19440
rect 25498 19388 25504 19440
rect 25556 19428 25562 19440
rect 26421 19431 26479 19437
rect 25556 19400 26372 19428
rect 25556 19388 25562 19400
rect 25590 19360 25596 19372
rect 24259 19332 24808 19360
rect 24872 19332 25596 19360
rect 24259 19329 24271 19332
rect 24213 19323 24271 19329
rect 23293 19295 23351 19301
rect 23293 19292 23305 19295
rect 22848 19264 23305 19292
rect 23293 19261 23305 19264
rect 23339 19292 23351 19295
rect 24228 19292 24256 19323
rect 23339 19264 24256 19292
rect 23339 19261 23351 19264
rect 23293 19255 23351 19261
rect 24394 19252 24400 19304
rect 24452 19252 24458 19304
rect 24780 19292 24808 19332
rect 25590 19320 25596 19332
rect 25648 19320 25654 19372
rect 26344 19360 26372 19400
rect 26421 19397 26433 19431
rect 26467 19428 26479 19431
rect 26786 19428 26792 19440
rect 26467 19400 26792 19428
rect 26467 19397 26479 19400
rect 26421 19391 26479 19397
rect 26786 19388 26792 19400
rect 26844 19388 26850 19440
rect 27706 19388 27712 19440
rect 27764 19388 27770 19440
rect 28629 19431 28687 19437
rect 28629 19397 28641 19431
rect 28675 19428 28687 19431
rect 28902 19428 28908 19440
rect 28675 19400 28908 19428
rect 28675 19397 28687 19400
rect 28629 19391 28687 19397
rect 28902 19388 28908 19400
rect 28960 19388 28966 19440
rect 30116 19428 30144 19459
rect 32306 19456 32312 19468
rect 32364 19456 32370 19508
rect 36630 19456 36636 19508
rect 36688 19456 36694 19508
rect 40218 19496 40224 19508
rect 37752 19468 40224 19496
rect 31294 19428 31300 19440
rect 30116 19400 31300 19428
rect 31294 19388 31300 19400
rect 31352 19428 31358 19440
rect 37752 19428 37780 19468
rect 40218 19456 40224 19468
rect 40276 19456 40282 19508
rect 41230 19456 41236 19508
rect 41288 19496 41294 19508
rect 41325 19499 41383 19505
rect 41325 19496 41337 19499
rect 41288 19468 41337 19496
rect 41288 19456 41294 19468
rect 41325 19465 41337 19468
rect 41371 19496 41383 19499
rect 41506 19496 41512 19508
rect 41371 19468 41512 19496
rect 41371 19465 41383 19468
rect 41325 19459 41383 19465
rect 41506 19456 41512 19468
rect 41564 19456 41570 19508
rect 31352 19400 33456 19428
rect 31352 19388 31358 19400
rect 27724 19360 27752 19388
rect 25700 19332 25912 19360
rect 26344 19332 27752 19360
rect 25700 19292 25728 19332
rect 24780 19264 25728 19292
rect 25774 19252 25780 19304
rect 25832 19252 25838 19304
rect 25884 19292 25912 19332
rect 29730 19320 29736 19372
rect 29788 19320 29794 19372
rect 29840 19332 30420 19360
rect 25884 19264 26924 19292
rect 26786 19224 26792 19236
rect 21008 19196 26792 19224
rect 18248 19128 18920 19156
rect 19429 19159 19487 19165
rect 18049 19119 18107 19125
rect 19429 19125 19441 19159
rect 19475 19156 19487 19159
rect 19518 19156 19524 19168
rect 19475 19128 19524 19156
rect 19475 19125 19487 19128
rect 19429 19119 19487 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 19978 19116 19984 19168
rect 20036 19156 20042 19168
rect 21008 19156 21036 19196
rect 26786 19184 26792 19196
rect 26844 19184 26850 19236
rect 20036 19128 21036 19156
rect 20036 19116 20042 19128
rect 22646 19116 22652 19168
rect 22704 19156 22710 19168
rect 22830 19156 22836 19168
rect 22704 19128 22836 19156
rect 22704 19116 22710 19128
rect 22830 19116 22836 19128
rect 22888 19156 22894 19168
rect 23017 19159 23075 19165
rect 23017 19156 23029 19159
rect 22888 19128 23029 19156
rect 22888 19116 22894 19128
rect 23017 19125 23029 19128
rect 23063 19125 23075 19159
rect 23017 19119 23075 19125
rect 23477 19159 23535 19165
rect 23477 19125 23489 19159
rect 23523 19156 23535 19159
rect 23566 19156 23572 19168
rect 23523 19128 23572 19156
rect 23523 19125 23535 19128
rect 23477 19119 23535 19125
rect 23566 19116 23572 19128
rect 23624 19116 23630 19168
rect 24486 19116 24492 19168
rect 24544 19156 24550 19168
rect 26510 19156 26516 19168
rect 24544 19128 26516 19156
rect 24544 19116 24550 19128
rect 26510 19116 26516 19128
rect 26568 19116 26574 19168
rect 26896 19156 26924 19264
rect 27614 19252 27620 19304
rect 27672 19252 27678 19304
rect 27709 19295 27767 19301
rect 27709 19261 27721 19295
rect 27755 19261 27767 19295
rect 27709 19255 27767 19261
rect 27338 19184 27344 19236
rect 27396 19224 27402 19236
rect 27724 19224 27752 19255
rect 28350 19252 28356 19304
rect 28408 19252 28414 19304
rect 29270 19252 29276 19304
rect 29328 19292 29334 19304
rect 29840 19292 29868 19332
rect 29328 19264 29868 19292
rect 30392 19292 30420 19332
rect 30466 19320 30472 19372
rect 30524 19360 30530 19372
rect 30561 19363 30619 19369
rect 30561 19360 30573 19363
rect 30524 19332 30573 19360
rect 30524 19320 30530 19332
rect 30561 19329 30573 19332
rect 30607 19329 30619 19363
rect 30561 19323 30619 19329
rect 31573 19363 31631 19369
rect 31573 19329 31585 19363
rect 31619 19360 31631 19363
rect 31754 19360 31760 19372
rect 31619 19332 31760 19360
rect 31619 19329 31631 19332
rect 31573 19323 31631 19329
rect 31754 19320 31760 19332
rect 31812 19360 31818 19372
rect 32122 19360 32128 19372
rect 31812 19332 32128 19360
rect 31812 19320 31818 19332
rect 32122 19320 32128 19332
rect 32180 19320 32186 19372
rect 33428 19369 33456 19400
rect 34900 19400 37780 19428
rect 34900 19369 34928 19400
rect 38378 19388 38384 19440
rect 38436 19428 38442 19440
rect 38841 19431 38899 19437
rect 38841 19428 38853 19431
rect 38436 19400 38853 19428
rect 38436 19388 38442 19400
rect 38841 19397 38853 19400
rect 38887 19428 38899 19431
rect 40129 19431 40187 19437
rect 40129 19428 40141 19431
rect 38887 19400 40141 19428
rect 38887 19397 38899 19400
rect 38841 19391 38899 19397
rect 40129 19397 40141 19400
rect 40175 19397 40187 19431
rect 40129 19391 40187 19397
rect 40494 19388 40500 19440
rect 40552 19428 40558 19440
rect 40681 19431 40739 19437
rect 40681 19428 40693 19431
rect 40552 19400 40693 19428
rect 40552 19388 40558 19400
rect 40681 19397 40693 19400
rect 40727 19428 40739 19431
rect 41141 19431 41199 19437
rect 41141 19428 41153 19431
rect 40727 19400 41153 19428
rect 40727 19397 40739 19400
rect 40681 19391 40739 19397
rect 41141 19397 41153 19400
rect 41187 19397 41199 19431
rect 41141 19391 41199 19397
rect 32309 19363 32367 19369
rect 32309 19329 32321 19363
rect 32355 19360 32367 19363
rect 33413 19363 33471 19369
rect 32355 19332 33364 19360
rect 32355 19329 32367 19332
rect 32309 19323 32367 19329
rect 30392 19264 31524 19292
rect 29328 19252 29334 19264
rect 31496 19236 31524 19264
rect 31938 19252 31944 19304
rect 31996 19292 32002 19304
rect 33134 19292 33140 19304
rect 31996 19264 33140 19292
rect 31996 19252 32002 19264
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 33336 19292 33364 19332
rect 33413 19329 33425 19363
rect 33459 19329 33471 19363
rect 34057 19363 34115 19369
rect 34057 19360 34069 19363
rect 33413 19323 33471 19329
rect 33520 19332 34069 19360
rect 33520 19292 33548 19332
rect 34057 19329 34069 19332
rect 34103 19329 34115 19363
rect 34057 19323 34115 19329
rect 34885 19363 34943 19369
rect 34885 19329 34897 19363
rect 34931 19329 34943 19363
rect 34885 19323 34943 19329
rect 35526 19320 35532 19372
rect 35584 19320 35590 19372
rect 35986 19320 35992 19372
rect 36044 19320 36050 19372
rect 37737 19363 37795 19369
rect 37737 19329 37749 19363
rect 37783 19360 37795 19363
rect 38470 19360 38476 19372
rect 37783 19332 38476 19360
rect 37783 19329 37795 19332
rect 37737 19323 37795 19329
rect 38470 19320 38476 19332
rect 38528 19320 38534 19372
rect 38562 19320 38568 19372
rect 38620 19360 38626 19372
rect 39669 19363 39727 19369
rect 39669 19360 39681 19363
rect 38620 19332 39681 19360
rect 38620 19320 38626 19332
rect 39669 19329 39681 19332
rect 39715 19360 39727 19363
rect 40218 19360 40224 19372
rect 39715 19332 40224 19360
rect 39715 19329 39727 19332
rect 39669 19323 39727 19329
rect 40218 19320 40224 19332
rect 40276 19320 40282 19372
rect 33336 19264 33548 19292
rect 36630 19252 36636 19304
rect 36688 19292 36694 19304
rect 37461 19295 37519 19301
rect 37461 19292 37473 19295
rect 36688 19264 37473 19292
rect 36688 19252 36694 19264
rect 37461 19261 37473 19264
rect 37507 19261 37519 19295
rect 37461 19255 37519 19261
rect 39025 19295 39083 19301
rect 39025 19261 39037 19295
rect 39071 19292 39083 19295
rect 39114 19292 39120 19304
rect 39071 19264 39120 19292
rect 39071 19261 39083 19264
rect 39025 19255 39083 19261
rect 39114 19252 39120 19264
rect 39172 19252 39178 19304
rect 41601 19295 41659 19301
rect 39224 19264 41414 19292
rect 27396 19196 27752 19224
rect 27396 19184 27402 19196
rect 30926 19184 30932 19236
rect 30984 19224 30990 19236
rect 31294 19224 31300 19236
rect 30984 19196 31300 19224
rect 30984 19184 30990 19196
rect 31294 19184 31300 19196
rect 31352 19184 31358 19236
rect 31478 19184 31484 19236
rect 31536 19224 31542 19236
rect 31849 19227 31907 19233
rect 31849 19224 31861 19227
rect 31536 19196 31861 19224
rect 31536 19184 31542 19196
rect 31849 19193 31861 19196
rect 31895 19193 31907 19227
rect 31849 19187 31907 19193
rect 33042 19184 33048 19236
rect 33100 19224 33106 19236
rect 34517 19227 34575 19233
rect 34517 19224 34529 19227
rect 33100 19196 33548 19224
rect 33100 19184 33106 19196
rect 28810 19156 28816 19168
rect 26896 19128 28816 19156
rect 28810 19116 28816 19128
rect 28868 19116 28874 19168
rect 31754 19116 31760 19168
rect 31812 19116 31818 19168
rect 32306 19116 32312 19168
rect 32364 19156 32370 19168
rect 32953 19159 33011 19165
rect 32953 19156 32965 19159
rect 32364 19128 32965 19156
rect 32364 19116 32370 19128
rect 32953 19125 32965 19128
rect 32999 19125 33011 19159
rect 33520 19156 33548 19196
rect 33796 19196 34529 19224
rect 33796 19156 33824 19196
rect 34517 19193 34529 19196
rect 34563 19193 34575 19227
rect 34517 19187 34575 19193
rect 34606 19184 34612 19236
rect 34664 19224 34670 19236
rect 39224 19224 39252 19264
rect 34664 19196 39252 19224
rect 34664 19184 34670 19196
rect 39390 19184 39396 19236
rect 39448 19224 39454 19236
rect 40037 19227 40095 19233
rect 40037 19224 40049 19227
rect 39448 19196 40049 19224
rect 39448 19184 39454 19196
rect 40037 19193 40049 19196
rect 40083 19193 40095 19227
rect 41386 19224 41414 19264
rect 41601 19261 41613 19295
rect 41647 19292 41659 19295
rect 41782 19292 41788 19304
rect 41647 19264 41788 19292
rect 41647 19261 41659 19264
rect 41601 19255 41659 19261
rect 41782 19252 41788 19264
rect 41840 19252 41846 19304
rect 45462 19224 45468 19236
rect 41386 19196 45468 19224
rect 40037 19187 40095 19193
rect 45462 19184 45468 19196
rect 45520 19184 45526 19236
rect 33520 19128 33824 19156
rect 32953 19119 33011 19125
rect 34330 19116 34336 19168
rect 34388 19116 34394 19168
rect 36630 19116 36636 19168
rect 36688 19156 36694 19168
rect 37001 19159 37059 19165
rect 37001 19156 37013 19159
rect 36688 19128 37013 19156
rect 36688 19116 36694 19128
rect 37001 19125 37013 19128
rect 37047 19125 37059 19159
rect 37001 19119 37059 19125
rect 39482 19116 39488 19168
rect 39540 19116 39546 19168
rect 40770 19116 40776 19168
rect 40828 19116 40834 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 6730 18952 6736 18964
rect 2464 18924 6736 18952
rect 2464 18912 2470 18924
rect 6730 18912 6736 18924
rect 6788 18952 6794 18964
rect 6788 18924 7328 18952
rect 6788 18912 6794 18924
rect 474 18844 480 18896
rect 532 18884 538 18896
rect 6362 18884 6368 18896
rect 532 18856 6368 18884
rect 532 18844 538 18856
rect 6362 18844 6368 18856
rect 6420 18844 6426 18896
rect 1394 18776 1400 18828
rect 1452 18816 1458 18828
rect 2041 18819 2099 18825
rect 2041 18816 2053 18819
rect 1452 18788 2053 18816
rect 1452 18776 1458 18788
rect 2041 18785 2053 18788
rect 2087 18785 2099 18819
rect 2041 18779 2099 18785
rect 3418 18776 3424 18828
rect 3476 18776 3482 18828
rect 3602 18776 3608 18828
rect 3660 18816 3666 18828
rect 4433 18819 4491 18825
rect 4433 18816 4445 18819
rect 3660 18788 4445 18816
rect 3660 18776 3666 18788
rect 4433 18785 4445 18788
rect 4479 18785 4491 18819
rect 4433 18779 4491 18785
rect 6270 18776 6276 18828
rect 6328 18776 6334 18828
rect 7300 18816 7328 18924
rect 7374 18912 7380 18964
rect 7432 18952 7438 18964
rect 7834 18952 7840 18964
rect 7432 18924 7840 18952
rect 7432 18912 7438 18924
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8938 18912 8944 18964
rect 8996 18952 9002 18964
rect 10413 18955 10471 18961
rect 10413 18952 10425 18955
rect 8996 18924 10425 18952
rect 8996 18912 9002 18924
rect 10413 18921 10425 18924
rect 10459 18952 10471 18955
rect 12434 18952 12440 18964
rect 10459 18924 12440 18952
rect 10459 18921 10471 18924
rect 10413 18915 10471 18921
rect 12434 18912 12440 18924
rect 12492 18912 12498 18964
rect 12618 18912 12624 18964
rect 12676 18912 12682 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 13725 18955 13783 18961
rect 13725 18952 13737 18955
rect 13688 18924 13737 18952
rect 13688 18912 13694 18924
rect 13725 18921 13737 18924
rect 13771 18921 13783 18955
rect 13725 18915 13783 18921
rect 13906 18912 13912 18964
rect 13964 18952 13970 18964
rect 14826 18952 14832 18964
rect 13964 18924 14832 18952
rect 13964 18912 13970 18924
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 17218 18952 17224 18964
rect 16632 18924 17224 18952
rect 16632 18912 16638 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 17589 18955 17647 18961
rect 17589 18952 17601 18955
rect 17328 18924 17601 18952
rect 7926 18844 7932 18896
rect 7984 18884 7990 18896
rect 9950 18884 9956 18896
rect 7984 18856 9956 18884
rect 7984 18844 7990 18856
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 13998 18884 14004 18896
rect 12400 18856 14004 18884
rect 12400 18844 12406 18856
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 16206 18844 16212 18896
rect 16264 18884 16270 18896
rect 16264 18856 16988 18884
rect 16264 18844 16270 18856
rect 8205 18819 8263 18825
rect 8205 18816 8217 18819
rect 7300 18788 8217 18816
rect 8205 18785 8217 18788
rect 8251 18816 8263 18819
rect 8294 18816 8300 18828
rect 8251 18788 8300 18816
rect 8251 18785 8263 18788
rect 8205 18779 8263 18785
rect 8294 18776 8300 18788
rect 8352 18776 8358 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 9585 18819 9643 18825
rect 9585 18816 9597 18819
rect 8444 18788 9597 18816
rect 8444 18776 8450 18788
rect 9585 18785 9597 18788
rect 9631 18785 9643 18819
rect 9585 18779 9643 18785
rect 9677 18819 9735 18825
rect 9677 18785 9689 18819
rect 9723 18785 9735 18819
rect 9677 18779 9735 18785
rect 10873 18819 10931 18825
rect 10873 18785 10885 18819
rect 10919 18816 10931 18819
rect 11698 18816 11704 18828
rect 10919 18788 11704 18816
rect 10919 18785 10931 18788
rect 10873 18779 10931 18785
rect 1765 18751 1823 18757
rect 1765 18717 1777 18751
rect 1811 18748 1823 18751
rect 3510 18748 3516 18760
rect 1811 18720 3516 18748
rect 1811 18717 1823 18720
rect 1765 18711 1823 18717
rect 3510 18708 3516 18720
rect 3568 18708 3574 18760
rect 4157 18751 4215 18757
rect 4157 18717 4169 18751
rect 4203 18717 4215 18751
rect 4157 18711 4215 18717
rect 4172 18680 4200 18711
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 8312 18748 8340 18776
rect 9122 18748 9128 18760
rect 8312 18720 9128 18748
rect 9122 18708 9128 18720
rect 9180 18708 9186 18760
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9692 18748 9720 18779
rect 11698 18776 11704 18788
rect 11756 18816 11762 18828
rect 14366 18816 14372 18828
rect 11756 18788 14372 18816
rect 11756 18776 11762 18788
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 14458 18776 14464 18828
rect 14516 18776 14522 18828
rect 14737 18819 14795 18825
rect 14737 18785 14749 18819
rect 14783 18816 14795 18819
rect 15746 18816 15752 18828
rect 14783 18788 15752 18816
rect 14783 18785 14795 18788
rect 14737 18779 14795 18785
rect 15746 18776 15752 18788
rect 15804 18776 15810 18828
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16853 18819 16911 18825
rect 16853 18816 16865 18819
rect 16632 18788 16865 18816
rect 16632 18776 16638 18788
rect 16853 18785 16865 18788
rect 16899 18785 16911 18819
rect 16960 18816 16988 18856
rect 17328 18816 17356 18924
rect 17589 18921 17601 18924
rect 17635 18921 17647 18955
rect 17589 18915 17647 18921
rect 17678 18912 17684 18964
rect 17736 18952 17742 18964
rect 19886 18952 19892 18964
rect 17736 18924 19892 18952
rect 17736 18912 17742 18924
rect 19886 18912 19892 18924
rect 19944 18912 19950 18964
rect 22370 18912 22376 18964
rect 22428 18952 22434 18964
rect 23293 18955 23351 18961
rect 23293 18952 23305 18955
rect 22428 18924 23305 18952
rect 22428 18912 22434 18924
rect 23293 18921 23305 18924
rect 23339 18921 23351 18955
rect 23293 18915 23351 18921
rect 23382 18912 23388 18964
rect 23440 18952 23446 18964
rect 24762 18952 24768 18964
rect 23440 18924 24768 18952
rect 23440 18912 23446 18924
rect 24762 18912 24768 18924
rect 24820 18912 24826 18964
rect 25314 18952 25320 18964
rect 24872 18924 25320 18952
rect 17494 18844 17500 18896
rect 17552 18884 17558 18896
rect 17552 18856 21220 18884
rect 17552 18844 17558 18856
rect 16960 18788 17356 18816
rect 16853 18779 16911 18785
rect 9272 18720 9720 18748
rect 9272 18708 9278 18720
rect 12710 18708 12716 18760
rect 12768 18748 12774 18760
rect 13081 18751 13139 18757
rect 13081 18748 13093 18751
rect 12768 18720 13093 18748
rect 12768 18708 12774 18720
rect 13081 18717 13093 18720
rect 13127 18717 13139 18751
rect 16868 18748 16896 18779
rect 17770 18776 17776 18828
rect 17828 18816 17834 18828
rect 18049 18819 18107 18825
rect 18049 18816 18061 18819
rect 17828 18788 18061 18816
rect 17828 18776 17834 18788
rect 18049 18785 18061 18788
rect 18095 18785 18107 18819
rect 18049 18779 18107 18785
rect 18138 18776 18144 18828
rect 18196 18776 18202 18828
rect 18601 18819 18659 18825
rect 18601 18816 18613 18819
rect 18248 18788 18613 18816
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 16868 18720 16957 18748
rect 13081 18711 13139 18717
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17034 18708 17040 18760
rect 17092 18748 17098 18760
rect 18248 18748 18276 18788
rect 18601 18785 18613 18788
rect 18647 18816 18659 18819
rect 19978 18816 19984 18828
rect 18647 18788 19984 18816
rect 18647 18785 18659 18788
rect 18601 18779 18659 18785
rect 19978 18776 19984 18788
rect 20036 18776 20042 18828
rect 20254 18776 20260 18828
rect 20312 18816 20318 18828
rect 20349 18819 20407 18825
rect 20349 18816 20361 18819
rect 20312 18788 20361 18816
rect 20312 18776 20318 18788
rect 20349 18785 20361 18788
rect 20395 18785 20407 18819
rect 20349 18779 20407 18785
rect 20898 18776 20904 18828
rect 20956 18816 20962 18828
rect 21085 18819 21143 18825
rect 21085 18816 21097 18819
rect 20956 18788 21097 18816
rect 20956 18776 20962 18788
rect 21085 18785 21097 18788
rect 21131 18785 21143 18819
rect 21192 18816 21220 18856
rect 23566 18844 23572 18896
rect 23624 18884 23630 18896
rect 24872 18893 24900 18924
rect 25314 18912 25320 18924
rect 25372 18952 25378 18964
rect 25498 18952 25504 18964
rect 25372 18924 25504 18952
rect 25372 18912 25378 18924
rect 25498 18912 25504 18924
rect 25556 18912 25562 18964
rect 25764 18955 25822 18961
rect 25764 18921 25776 18955
rect 25810 18952 25822 18955
rect 27522 18952 27528 18964
rect 25810 18924 27528 18952
rect 25810 18921 25822 18924
rect 25764 18915 25822 18921
rect 27522 18912 27528 18924
rect 27580 18912 27586 18964
rect 27614 18912 27620 18964
rect 27672 18952 27678 18964
rect 28445 18955 28503 18961
rect 28445 18952 28457 18955
rect 27672 18924 28457 18952
rect 27672 18912 27678 18924
rect 28445 18921 28457 18924
rect 28491 18921 28503 18955
rect 28445 18915 28503 18921
rect 29822 18912 29828 18964
rect 29880 18952 29886 18964
rect 32033 18955 32091 18961
rect 32033 18952 32045 18955
rect 29880 18924 32045 18952
rect 29880 18912 29886 18924
rect 32033 18921 32045 18924
rect 32079 18952 32091 18955
rect 33318 18952 33324 18964
rect 32079 18924 33324 18952
rect 32079 18921 32091 18924
rect 32033 18915 32091 18921
rect 33318 18912 33324 18924
rect 33376 18912 33382 18964
rect 33413 18955 33471 18961
rect 33413 18921 33425 18955
rect 33459 18952 33471 18955
rect 33686 18952 33692 18964
rect 33459 18924 33692 18952
rect 33459 18921 33471 18924
rect 33413 18915 33471 18921
rect 33686 18912 33692 18924
rect 33744 18912 33750 18964
rect 34238 18912 34244 18964
rect 34296 18952 34302 18964
rect 35618 18952 35624 18964
rect 34296 18924 35624 18952
rect 34296 18912 34302 18924
rect 35618 18912 35624 18924
rect 35676 18912 35682 18964
rect 35710 18912 35716 18964
rect 35768 18952 35774 18964
rect 36817 18955 36875 18961
rect 35768 18924 36768 18952
rect 35768 18912 35774 18924
rect 24857 18887 24915 18893
rect 23624 18856 24808 18884
rect 23624 18844 23630 18856
rect 23109 18819 23167 18825
rect 23109 18816 23121 18819
rect 21192 18788 23121 18816
rect 21085 18779 21143 18785
rect 23109 18785 23121 18788
rect 23155 18816 23167 18819
rect 23155 18788 23704 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 17092 18720 18276 18748
rect 17092 18708 17098 18720
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 19426 18748 19432 18760
rect 19116 18720 19432 18748
rect 19116 18708 19122 18720
rect 19426 18708 19432 18720
rect 19484 18748 19490 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19484 18720 19625 18748
rect 19484 18708 19490 18720
rect 19613 18717 19625 18720
rect 19659 18748 19671 18751
rect 20714 18748 20720 18760
rect 19659 18720 20720 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 23566 18748 23572 18760
rect 22494 18720 23572 18748
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 23676 18757 23704 18788
rect 23842 18776 23848 18828
rect 23900 18816 23906 18828
rect 23937 18819 23995 18825
rect 23937 18816 23949 18819
rect 23900 18788 23949 18816
rect 23900 18776 23906 18788
rect 23937 18785 23949 18788
rect 23983 18816 23995 18819
rect 24670 18816 24676 18828
rect 23983 18788 24676 18816
rect 23983 18785 23995 18788
rect 23937 18779 23995 18785
rect 24670 18776 24676 18788
rect 24728 18776 24734 18828
rect 24780 18816 24808 18856
rect 24857 18853 24869 18887
rect 24903 18853 24915 18887
rect 24857 18847 24915 18853
rect 26786 18844 26792 18896
rect 26844 18884 26850 18896
rect 36740 18884 36768 18924
rect 36817 18921 36829 18955
rect 36863 18952 36875 18955
rect 37090 18952 37096 18964
rect 36863 18924 37096 18952
rect 36863 18921 36875 18924
rect 36817 18915 36875 18921
rect 37090 18912 37096 18924
rect 37148 18912 37154 18964
rect 39224 18924 39528 18952
rect 39224 18884 39252 18924
rect 26844 18856 36216 18884
rect 36740 18856 39252 18884
rect 39301 18887 39359 18893
rect 26844 18844 26850 18856
rect 25501 18819 25559 18825
rect 24780 18788 25452 18816
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18717 23719 18751
rect 23661 18711 23719 18717
rect 23768 18720 25360 18748
rect 7926 18680 7932 18692
rect 4172 18652 7932 18680
rect 7926 18640 7932 18652
rect 7984 18640 7990 18692
rect 8018 18640 8024 18692
rect 8076 18640 8082 18692
rect 9398 18640 9404 18692
rect 9456 18680 9462 18692
rect 9493 18683 9551 18689
rect 9493 18680 9505 18683
rect 9456 18652 9505 18680
rect 9456 18640 9462 18652
rect 9493 18649 9505 18652
rect 9539 18649 9551 18683
rect 9493 18643 9551 18649
rect 10594 18640 10600 18692
rect 10652 18640 10658 18692
rect 11146 18640 11152 18692
rect 11204 18640 11210 18692
rect 11348 18652 11638 18680
rect 11348 18624 11376 18652
rect 15010 18640 15016 18692
rect 15068 18640 15074 18692
rect 15470 18640 15476 18692
rect 15528 18640 15534 18692
rect 16298 18640 16304 18692
rect 16356 18680 16362 18692
rect 16356 18652 16620 18680
rect 16356 18640 16362 18652
rect 3602 18572 3608 18624
rect 3660 18572 3666 18624
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 7558 18612 7564 18624
rect 5776 18584 7564 18612
rect 5776 18572 5782 18584
rect 7558 18572 7564 18584
rect 7616 18572 7622 18624
rect 7650 18572 7656 18624
rect 7708 18572 7714 18624
rect 7834 18572 7840 18624
rect 7892 18612 7898 18624
rect 8113 18615 8171 18621
rect 8113 18612 8125 18615
rect 7892 18584 8125 18612
rect 7892 18572 7898 18584
rect 8113 18581 8125 18584
rect 8159 18581 8171 18615
rect 8113 18575 8171 18581
rect 8754 18572 8760 18624
rect 8812 18572 8818 18624
rect 8846 18572 8852 18624
rect 8904 18612 8910 18624
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 8904 18584 9137 18612
rect 8904 18572 8910 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 10229 18615 10287 18621
rect 10229 18581 10241 18615
rect 10275 18612 10287 18615
rect 10318 18612 10324 18624
rect 10275 18584 10324 18612
rect 10275 18581 10287 18584
rect 10229 18575 10287 18581
rect 10318 18572 10324 18584
rect 10376 18612 10382 18624
rect 11054 18612 11060 18624
rect 10376 18584 11060 18612
rect 10376 18572 10382 18584
rect 11054 18572 11060 18584
rect 11112 18572 11118 18624
rect 11330 18572 11336 18624
rect 11388 18612 11394 18624
rect 11974 18612 11980 18624
rect 11388 18584 11980 18612
rect 11388 18572 11394 18584
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 14277 18615 14335 18621
rect 14277 18581 14289 18615
rect 14323 18612 14335 18615
rect 15286 18612 15292 18624
rect 14323 18584 15292 18612
rect 14323 18581 14335 18584
rect 14277 18575 14335 18581
rect 15286 18572 15292 18584
rect 15344 18572 15350 18624
rect 15746 18572 15752 18624
rect 15804 18612 15810 18624
rect 16485 18615 16543 18621
rect 16485 18612 16497 18615
rect 15804 18584 16497 18612
rect 15804 18572 15810 18584
rect 16485 18581 16497 18584
rect 16531 18581 16543 18615
rect 16592 18612 16620 18652
rect 16758 18640 16764 18692
rect 16816 18680 16822 18692
rect 17862 18680 17868 18692
rect 16816 18652 17868 18680
rect 16816 18640 16822 18652
rect 17862 18640 17868 18652
rect 17920 18680 17926 18692
rect 17957 18683 18015 18689
rect 17957 18680 17969 18683
rect 17920 18652 17969 18680
rect 17920 18640 17926 18652
rect 17957 18649 17969 18652
rect 18003 18649 18015 18683
rect 21361 18683 21419 18689
rect 21361 18680 21373 18683
rect 17957 18643 18015 18649
rect 18052 18652 21373 18680
rect 18052 18612 18080 18652
rect 21361 18649 21373 18652
rect 21407 18649 21419 18683
rect 21361 18643 21419 18649
rect 22646 18640 22652 18692
rect 22704 18680 22710 18692
rect 23768 18680 23796 18720
rect 22704 18652 23796 18680
rect 22704 18640 22710 18652
rect 24302 18640 24308 18692
rect 24360 18680 24366 18692
rect 24673 18683 24731 18689
rect 24673 18680 24685 18683
rect 24360 18652 24685 18680
rect 24360 18640 24366 18652
rect 24673 18649 24685 18652
rect 24719 18680 24731 18683
rect 24946 18680 24952 18692
rect 24719 18652 24952 18680
rect 24719 18649 24731 18652
rect 24673 18643 24731 18649
rect 24946 18640 24952 18652
rect 25004 18640 25010 18692
rect 16592 18584 18080 18612
rect 16485 18575 16543 18581
rect 18230 18572 18236 18624
rect 18288 18612 18294 18624
rect 18414 18612 18420 18624
rect 18288 18584 18420 18612
rect 18288 18572 18294 18584
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 18782 18572 18788 18624
rect 18840 18572 18846 18624
rect 19061 18615 19119 18621
rect 19061 18581 19073 18615
rect 19107 18612 19119 18615
rect 19150 18612 19156 18624
rect 19107 18584 19156 18612
rect 19107 18581 19119 18584
rect 19061 18575 19119 18581
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19337 18615 19395 18621
rect 19337 18581 19349 18615
rect 19383 18612 19395 18615
rect 19426 18612 19432 18624
rect 19383 18584 19432 18612
rect 19383 18581 19395 18584
rect 19337 18575 19395 18581
rect 19426 18572 19432 18584
rect 19484 18612 19490 18624
rect 20622 18612 20628 18624
rect 19484 18584 20628 18612
rect 19484 18572 19490 18584
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 22738 18572 22744 18624
rect 22796 18612 22802 18624
rect 22833 18615 22891 18621
rect 22833 18612 22845 18615
rect 22796 18584 22845 18612
rect 22796 18572 22802 18584
rect 22833 18581 22845 18584
rect 22879 18581 22891 18615
rect 22833 18575 22891 18581
rect 23658 18572 23664 18624
rect 23716 18612 23722 18624
rect 23753 18615 23811 18621
rect 23753 18612 23765 18615
rect 23716 18584 23765 18612
rect 23716 18572 23722 18584
rect 23753 18581 23765 18584
rect 23799 18612 23811 18615
rect 23842 18612 23848 18624
rect 23799 18584 23848 18612
rect 23799 18581 23811 18584
rect 23753 18575 23811 18581
rect 23842 18572 23848 18584
rect 23900 18572 23906 18624
rect 25222 18572 25228 18624
rect 25280 18572 25286 18624
rect 25332 18612 25360 18720
rect 25424 18680 25452 18788
rect 25501 18785 25513 18819
rect 25547 18816 25559 18819
rect 25774 18816 25780 18828
rect 25547 18788 25780 18816
rect 25547 18785 25559 18788
rect 25501 18779 25559 18785
rect 25774 18776 25780 18788
rect 25832 18776 25838 18828
rect 25866 18776 25872 18828
rect 25924 18816 25930 18828
rect 26142 18816 26148 18828
rect 25924 18788 26148 18816
rect 25924 18776 25930 18788
rect 26142 18776 26148 18788
rect 26200 18776 26206 18828
rect 26234 18776 26240 18828
rect 26292 18816 26298 18828
rect 27709 18819 27767 18825
rect 27709 18816 27721 18819
rect 26292 18788 27721 18816
rect 26292 18776 26298 18788
rect 27709 18785 27721 18788
rect 27755 18785 27767 18819
rect 27709 18779 27767 18785
rect 28258 18776 28264 18828
rect 28316 18816 28322 18828
rect 28316 18788 29040 18816
rect 28316 18776 28322 18788
rect 28810 18708 28816 18760
rect 28868 18748 28874 18760
rect 28905 18751 28963 18757
rect 28905 18748 28917 18751
rect 28868 18720 28917 18748
rect 28868 18708 28874 18720
rect 28905 18717 28917 18720
rect 28951 18717 28963 18751
rect 29012 18748 29040 18788
rect 29086 18776 29092 18828
rect 29144 18776 29150 18828
rect 29454 18816 29460 18828
rect 29196 18788 29460 18816
rect 29196 18748 29224 18788
rect 29454 18776 29460 18788
rect 29512 18816 29518 18828
rect 29512 18788 30972 18816
rect 29512 18776 29518 18788
rect 29012 18720 29224 18748
rect 29733 18751 29791 18757
rect 28905 18711 28963 18717
rect 29733 18717 29745 18751
rect 29779 18717 29791 18751
rect 29733 18711 29791 18717
rect 26234 18680 26240 18692
rect 25424 18652 26240 18680
rect 26234 18640 26240 18652
rect 26292 18640 26298 18692
rect 29748 18680 29776 18711
rect 30834 18708 30840 18760
rect 30892 18708 30898 18760
rect 30944 18748 30972 18788
rect 31202 18776 31208 18828
rect 31260 18816 31266 18828
rect 31260 18788 35572 18816
rect 31260 18776 31266 18788
rect 32214 18748 32220 18760
rect 30944 18720 32220 18748
rect 32214 18708 32220 18720
rect 32272 18708 32278 18760
rect 32306 18708 32312 18760
rect 32364 18708 32370 18760
rect 32490 18708 32496 18760
rect 32548 18748 32554 18760
rect 33597 18751 33655 18757
rect 33597 18748 33609 18751
rect 32548 18720 33609 18748
rect 32548 18708 32554 18720
rect 33597 18717 33609 18720
rect 33643 18717 33655 18751
rect 33597 18711 33655 18717
rect 33778 18708 33784 18760
rect 33836 18748 33842 18760
rect 33836 18720 34468 18748
rect 33836 18708 33842 18720
rect 31481 18683 31539 18689
rect 31481 18680 31493 18683
rect 27080 18652 29776 18680
rect 31404 18652 31493 18680
rect 27080 18612 27108 18652
rect 25332 18584 27108 18612
rect 27154 18572 27160 18624
rect 27212 18612 27218 18624
rect 27249 18615 27307 18621
rect 27249 18612 27261 18615
rect 27212 18584 27261 18612
rect 27212 18572 27218 18584
rect 27249 18581 27261 18584
rect 27295 18581 27307 18615
rect 27249 18575 27307 18581
rect 27798 18572 27804 18624
rect 27856 18612 27862 18624
rect 28258 18612 28264 18624
rect 27856 18584 28264 18612
rect 27856 18572 27862 18584
rect 28258 18572 28264 18584
rect 28316 18612 28322 18624
rect 28813 18615 28871 18621
rect 28813 18612 28825 18615
rect 28316 18584 28825 18612
rect 28316 18572 28322 18584
rect 28813 18581 28825 18584
rect 28859 18581 28871 18615
rect 28813 18575 28871 18581
rect 29362 18572 29368 18624
rect 29420 18612 29426 18624
rect 30190 18612 30196 18624
rect 29420 18584 30196 18612
rect 29420 18572 29426 18584
rect 30190 18572 30196 18584
rect 30248 18572 30254 18624
rect 30374 18572 30380 18624
rect 30432 18572 30438 18624
rect 30558 18572 30564 18624
rect 30616 18612 30622 18624
rect 31404 18612 31432 18652
rect 31481 18649 31493 18652
rect 31527 18649 31539 18683
rect 31481 18643 31539 18649
rect 31754 18640 31760 18692
rect 31812 18640 31818 18692
rect 33686 18640 33692 18692
rect 33744 18680 33750 18692
rect 34149 18683 34207 18689
rect 34149 18680 34161 18683
rect 33744 18652 34161 18680
rect 33744 18640 33750 18652
rect 34149 18649 34161 18652
rect 34195 18680 34207 18683
rect 34330 18680 34336 18692
rect 34195 18652 34336 18680
rect 34195 18649 34207 18652
rect 34149 18643 34207 18649
rect 34330 18640 34336 18652
rect 34388 18640 34394 18692
rect 34440 18680 34468 18720
rect 34882 18708 34888 18760
rect 34940 18708 34946 18760
rect 35161 18751 35219 18757
rect 35161 18717 35173 18751
rect 35207 18717 35219 18751
rect 35161 18711 35219 18717
rect 35176 18680 35204 18711
rect 34440 18652 35204 18680
rect 35544 18680 35572 18788
rect 36188 18757 36216 18856
rect 39301 18853 39313 18887
rect 39347 18853 39359 18887
rect 39301 18847 39359 18853
rect 39500 18884 39528 18924
rect 39574 18912 39580 18964
rect 39632 18952 39638 18964
rect 43530 18952 43536 18964
rect 39632 18924 43536 18952
rect 39632 18912 39638 18924
rect 43530 18912 43536 18924
rect 43588 18912 43594 18964
rect 40037 18887 40095 18893
rect 40037 18884 40049 18887
rect 39500 18856 40049 18884
rect 39316 18816 39344 18847
rect 37200 18788 39344 18816
rect 36173 18751 36231 18757
rect 36173 18717 36185 18751
rect 36219 18748 36231 18751
rect 37093 18751 37151 18757
rect 37093 18748 37105 18751
rect 36219 18720 37105 18748
rect 36219 18717 36231 18720
rect 36173 18711 36231 18717
rect 37093 18717 37105 18720
rect 37139 18717 37151 18751
rect 37093 18711 37151 18717
rect 37200 18680 37228 18788
rect 37458 18708 37464 18760
rect 37516 18708 37522 18760
rect 39500 18757 39528 18856
rect 40037 18853 40049 18856
rect 40083 18853 40095 18887
rect 40037 18847 40095 18853
rect 40218 18844 40224 18896
rect 40276 18844 40282 18896
rect 39485 18751 39543 18757
rect 39485 18717 39497 18751
rect 39531 18717 39543 18751
rect 39485 18711 39543 18717
rect 38657 18683 38715 18689
rect 38657 18680 38669 18683
rect 35544 18652 37228 18680
rect 37292 18652 38669 18680
rect 30616 18584 31432 18612
rect 30616 18572 30622 18584
rect 32950 18572 32956 18624
rect 33008 18572 33014 18624
rect 33502 18572 33508 18624
rect 33560 18612 33566 18624
rect 34241 18615 34299 18621
rect 34241 18612 34253 18615
rect 33560 18584 34253 18612
rect 33560 18572 33566 18584
rect 34241 18581 34253 18584
rect 34287 18581 34299 18615
rect 34241 18575 34299 18581
rect 34793 18615 34851 18621
rect 34793 18581 34805 18615
rect 34839 18612 34851 18615
rect 34882 18612 34888 18624
rect 34839 18584 34888 18612
rect 34839 18581 34851 18584
rect 34793 18575 34851 18581
rect 34882 18572 34888 18584
rect 34940 18572 34946 18624
rect 35618 18572 35624 18624
rect 35676 18612 35682 18624
rect 37292 18612 37320 18652
rect 38657 18649 38669 18652
rect 38703 18680 38715 18683
rect 39853 18683 39911 18689
rect 39853 18680 39865 18683
rect 38703 18652 39865 18680
rect 38703 18649 38715 18652
rect 38657 18643 38715 18649
rect 39853 18649 39865 18652
rect 39899 18649 39911 18683
rect 39853 18643 39911 18649
rect 35676 18584 37320 18612
rect 35676 18572 35682 18584
rect 37826 18572 37832 18624
rect 37884 18612 37890 18624
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 37884 18584 38117 18612
rect 37884 18572 37890 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 38746 18572 38752 18624
rect 38804 18572 38810 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 10321 18411 10379 18417
rect 3476 18380 8892 18408
rect 3476 18368 3482 18380
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 5810 18340 5816 18352
rect 5675 18312 5816 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 5810 18300 5816 18312
rect 5868 18300 5874 18352
rect 7374 18340 7380 18352
rect 6656 18312 7380 18340
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 3326 18272 3332 18284
rect 1811 18244 3332 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 3326 18232 3332 18244
rect 3384 18232 3390 18284
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18272 3663 18275
rect 6656 18272 6684 18312
rect 7374 18300 7380 18312
rect 7432 18300 7438 18352
rect 7466 18300 7472 18352
rect 7524 18300 7530 18352
rect 7926 18300 7932 18352
rect 7984 18340 7990 18352
rect 7984 18312 8800 18340
rect 7984 18300 7990 18312
rect 3651 18244 6684 18272
rect 6733 18275 6791 18281
rect 3651 18241 3663 18244
rect 3605 18235 3663 18241
rect 6733 18241 6745 18275
rect 6779 18272 6791 18275
rect 6779 18244 8156 18272
rect 6779 18241 6791 18244
rect 6733 18235 6791 18241
rect 2038 18164 2044 18216
rect 2096 18164 2102 18216
rect 3878 18164 3884 18216
rect 3936 18164 3942 18216
rect 5718 18164 5724 18216
rect 5776 18164 5782 18216
rect 5902 18164 5908 18216
rect 5960 18164 5966 18216
rect 6086 18164 6092 18216
rect 6144 18204 6150 18216
rect 7282 18204 7288 18216
rect 6144 18176 7288 18204
rect 6144 18164 6150 18176
rect 7282 18164 7288 18176
rect 7340 18164 7346 18216
rect 5261 18139 5319 18145
rect 5261 18105 5273 18139
rect 5307 18136 5319 18139
rect 7926 18136 7932 18148
rect 5307 18108 7932 18136
rect 5307 18105 5319 18108
rect 5261 18099 5319 18105
rect 7926 18096 7932 18108
rect 7984 18096 7990 18148
rect 8128 18136 8156 18244
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 8260 18176 8401 18204
rect 8260 18164 8266 18176
rect 8389 18173 8401 18176
rect 8435 18173 8447 18207
rect 8772 18204 8800 18312
rect 8864 18272 8892 18380
rect 10321 18377 10333 18411
rect 10367 18408 10379 18411
rect 10870 18408 10876 18420
rect 10367 18380 10876 18408
rect 10367 18377 10379 18380
rect 10321 18371 10379 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 11514 18368 11520 18420
rect 11572 18408 11578 18420
rect 12253 18411 12311 18417
rect 12253 18408 12265 18411
rect 11572 18380 12265 18408
rect 11572 18368 11578 18380
rect 12253 18377 12265 18380
rect 12299 18377 12311 18411
rect 12253 18371 12311 18377
rect 12621 18411 12679 18417
rect 12621 18377 12633 18411
rect 12667 18408 12679 18411
rect 12894 18408 12900 18420
rect 12667 18380 12900 18408
rect 12667 18377 12679 18380
rect 12621 18371 12679 18377
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 14642 18408 14648 18420
rect 13832 18380 14648 18408
rect 9582 18300 9588 18352
rect 9640 18340 9646 18352
rect 9677 18343 9735 18349
rect 9677 18340 9689 18343
rect 9640 18312 9689 18340
rect 9640 18300 9646 18312
rect 9677 18309 9689 18312
rect 9723 18309 9735 18343
rect 9677 18303 9735 18309
rect 10612 18312 10824 18340
rect 8938 18272 8944 18284
rect 8864 18244 8944 18272
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9398 18232 9404 18284
rect 9456 18272 9462 18284
rect 10612 18272 10640 18312
rect 9456 18244 10640 18272
rect 9456 18232 9462 18244
rect 10686 18232 10692 18284
rect 10744 18232 10750 18284
rect 10796 18272 10824 18312
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 11701 18343 11759 18349
rect 11701 18340 11713 18343
rect 11664 18312 11713 18340
rect 11664 18300 11670 18312
rect 11701 18309 11713 18312
rect 11747 18309 11759 18343
rect 11701 18303 11759 18309
rect 11977 18343 12035 18349
rect 11977 18309 11989 18343
rect 12023 18340 12035 18343
rect 12434 18340 12440 18352
rect 12023 18312 12440 18340
rect 12023 18309 12035 18312
rect 11977 18303 12035 18309
rect 12434 18300 12440 18312
rect 12492 18340 12498 18352
rect 13449 18343 13507 18349
rect 13449 18340 13461 18343
rect 12492 18312 13461 18340
rect 12492 18300 12498 18312
rect 13449 18309 13461 18312
rect 13495 18309 13507 18343
rect 13449 18303 13507 18309
rect 12713 18275 12771 18281
rect 12713 18272 12725 18275
rect 10796 18244 12725 18272
rect 12713 18241 12725 18244
rect 12759 18272 12771 18275
rect 13832 18272 13860 18380
rect 14642 18368 14648 18380
rect 14700 18368 14706 18420
rect 14829 18411 14887 18417
rect 14829 18377 14841 18411
rect 14875 18408 14887 18411
rect 15102 18408 15108 18420
rect 14875 18380 15108 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 15102 18368 15108 18380
rect 15160 18368 15166 18420
rect 15289 18411 15347 18417
rect 15289 18377 15301 18411
rect 15335 18408 15347 18411
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 15335 18380 19165 18408
rect 15335 18377 15347 18380
rect 15289 18371 15347 18377
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 21453 18411 21511 18417
rect 21453 18408 21465 18411
rect 19153 18371 19211 18377
rect 19260 18380 21465 18408
rect 14277 18343 14335 18349
rect 14277 18309 14289 18343
rect 14323 18340 14335 18343
rect 14366 18340 14372 18352
rect 14323 18312 14372 18340
rect 14323 18309 14335 18312
rect 14277 18303 14335 18309
rect 14366 18300 14372 18312
rect 14424 18300 14430 18352
rect 17221 18343 17279 18349
rect 17221 18340 17233 18343
rect 14476 18312 17233 18340
rect 12759 18244 13860 18272
rect 12759 18241 12771 18244
rect 12713 18235 12771 18241
rect 13906 18232 13912 18284
rect 13964 18272 13970 18284
rect 14476 18272 14504 18312
rect 17221 18309 17233 18312
rect 17267 18309 17279 18343
rect 19260 18340 19288 18380
rect 21453 18377 21465 18380
rect 21499 18377 21511 18411
rect 24857 18411 24915 18417
rect 24857 18408 24869 18411
rect 21453 18371 21511 18377
rect 21560 18380 24869 18408
rect 17221 18303 17279 18309
rect 18064 18312 19288 18340
rect 13964 18244 14504 18272
rect 13964 18232 13970 18244
rect 15194 18232 15200 18284
rect 15252 18232 15258 18284
rect 15286 18232 15292 18284
rect 15344 18272 15350 18284
rect 15344 18244 16068 18272
rect 15344 18232 15350 18244
rect 10594 18204 10600 18216
rect 8772 18176 10600 18204
rect 8389 18167 8447 18173
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 10870 18204 10876 18216
rect 10827 18176 10876 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 10870 18164 10876 18176
rect 10928 18164 10934 18216
rect 10962 18164 10968 18216
rect 11020 18204 11026 18216
rect 12250 18204 12256 18216
rect 11020 18176 12256 18204
rect 11020 18164 11026 18176
rect 12250 18164 12256 18176
rect 12308 18164 12314 18216
rect 12897 18207 12955 18213
rect 12897 18173 12909 18207
rect 12943 18204 12955 18207
rect 13446 18204 13452 18216
rect 12943 18176 13452 18204
rect 12943 18173 12955 18176
rect 12897 18167 12955 18173
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 15746 18204 15752 18216
rect 15436 18176 15752 18204
rect 15436 18164 15442 18176
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 16040 18204 16068 18244
rect 16114 18232 16120 18284
rect 16172 18232 16178 18284
rect 16206 18232 16212 18284
rect 16264 18272 16270 18284
rect 17126 18272 17132 18284
rect 16264 18244 17132 18272
rect 16264 18232 16270 18244
rect 17126 18232 17132 18244
rect 17184 18232 17190 18284
rect 17313 18275 17371 18281
rect 17313 18241 17325 18275
rect 17359 18272 17371 18275
rect 17862 18272 17868 18284
rect 17359 18244 17868 18272
rect 17359 18241 17371 18244
rect 17313 18235 17371 18241
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 18064 18281 18092 18312
rect 19794 18300 19800 18352
rect 19852 18340 19858 18352
rect 21560 18340 21588 18380
rect 24857 18377 24869 18380
rect 24903 18377 24915 18411
rect 29362 18408 29368 18420
rect 24857 18371 24915 18377
rect 24964 18380 29368 18408
rect 19852 18312 21588 18340
rect 19852 18300 19858 18312
rect 22646 18300 22652 18352
rect 22704 18300 22710 18352
rect 23290 18300 23296 18352
rect 23348 18340 23354 18352
rect 23385 18343 23443 18349
rect 23385 18340 23397 18343
rect 23348 18312 23397 18340
rect 23348 18300 23354 18312
rect 23385 18309 23397 18312
rect 23431 18309 23443 18343
rect 23385 18303 23443 18309
rect 23842 18300 23848 18352
rect 23900 18300 23906 18352
rect 24670 18300 24676 18352
rect 24728 18340 24734 18352
rect 24964 18340 24992 18380
rect 29362 18368 29368 18380
rect 29420 18368 29426 18420
rect 29730 18408 29736 18420
rect 29472 18380 29736 18408
rect 24728 18312 24992 18340
rect 24728 18300 24734 18312
rect 25958 18300 25964 18352
rect 26016 18340 26022 18352
rect 26053 18343 26111 18349
rect 26053 18340 26065 18343
rect 26016 18312 26065 18340
rect 26016 18300 26022 18312
rect 26053 18309 26065 18312
rect 26099 18309 26111 18343
rect 26053 18303 26111 18309
rect 26142 18300 26148 18352
rect 26200 18340 26206 18352
rect 27614 18340 27620 18352
rect 26200 18312 27620 18340
rect 26200 18300 26206 18312
rect 27614 18300 27620 18312
rect 27672 18300 27678 18352
rect 28350 18340 28356 18352
rect 28092 18312 28356 18340
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18049 18235 18107 18241
rect 18138 18232 18144 18284
rect 18196 18272 18202 18284
rect 18966 18272 18972 18284
rect 18196 18244 18972 18272
rect 18196 18232 18202 18244
rect 18966 18232 18972 18244
rect 19024 18232 19030 18284
rect 19518 18232 19524 18284
rect 19576 18232 19582 18284
rect 20809 18275 20867 18281
rect 19628 18244 20760 18272
rect 16574 18204 16580 18216
rect 16040 18176 16580 18204
rect 16574 18164 16580 18176
rect 16632 18164 16638 18216
rect 17497 18207 17555 18213
rect 17497 18173 17509 18207
rect 17543 18204 17555 18207
rect 19150 18204 19156 18216
rect 17543 18176 19156 18204
rect 17543 18173 17555 18176
rect 17497 18167 17555 18173
rect 19150 18164 19156 18176
rect 19208 18164 19214 18216
rect 19242 18164 19248 18216
rect 19300 18204 19306 18216
rect 19628 18213 19656 18244
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 19300 18176 19625 18204
rect 19300 18164 19306 18176
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19613 18167 19671 18173
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18204 19763 18207
rect 19978 18204 19984 18216
rect 19751 18176 19984 18204
rect 19751 18173 19763 18176
rect 19705 18167 19763 18173
rect 19978 18164 19984 18176
rect 20036 18164 20042 18216
rect 16301 18139 16359 18145
rect 16301 18136 16313 18139
rect 8128 18108 16313 18136
rect 16301 18105 16313 18108
rect 16347 18105 16359 18139
rect 16301 18099 16359 18105
rect 16758 18096 16764 18148
rect 16816 18136 16822 18148
rect 16853 18139 16911 18145
rect 16853 18136 16865 18139
rect 16816 18108 16865 18136
rect 16816 18096 16822 18108
rect 16853 18105 16865 18108
rect 16899 18105 16911 18139
rect 16853 18099 16911 18105
rect 17126 18096 17132 18148
rect 17184 18136 17190 18148
rect 19518 18136 19524 18148
rect 17184 18108 19524 18136
rect 17184 18096 17190 18108
rect 19518 18096 19524 18108
rect 19576 18096 19582 18148
rect 20732 18136 20760 18244
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20824 18204 20852 18235
rect 22002 18232 22008 18284
rect 22060 18232 22066 18284
rect 23106 18232 23112 18284
rect 23164 18232 23170 18284
rect 25222 18232 25228 18284
rect 25280 18272 25286 18284
rect 25317 18275 25375 18281
rect 25317 18272 25329 18275
rect 25280 18244 25329 18272
rect 25280 18232 25286 18244
rect 25317 18241 25329 18244
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 27522 18232 27528 18284
rect 27580 18272 27586 18284
rect 27982 18272 27988 18284
rect 27580 18244 27988 18272
rect 27580 18232 27586 18244
rect 27982 18232 27988 18244
rect 28040 18272 28046 18284
rect 28092 18281 28120 18312
rect 28350 18300 28356 18312
rect 28408 18300 28414 18352
rect 29472 18284 29500 18380
rect 29730 18368 29736 18380
rect 29788 18368 29794 18420
rect 32122 18368 32128 18420
rect 32180 18368 32186 18420
rect 32769 18411 32827 18417
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 33594 18408 33600 18420
rect 32815 18380 33600 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 30098 18300 30104 18352
rect 30156 18340 30162 18352
rect 30929 18343 30987 18349
rect 30929 18340 30941 18343
rect 30156 18312 30941 18340
rect 30156 18300 30162 18312
rect 30929 18309 30941 18312
rect 30975 18309 30987 18343
rect 30929 18303 30987 18309
rect 31757 18343 31815 18349
rect 31757 18309 31769 18343
rect 31803 18340 31815 18343
rect 32030 18340 32036 18352
rect 31803 18312 32036 18340
rect 31803 18309 31815 18312
rect 31757 18303 31815 18309
rect 32030 18300 32036 18312
rect 32088 18300 32094 18352
rect 28077 18275 28135 18281
rect 28077 18272 28089 18275
rect 28040 18244 28089 18272
rect 28040 18232 28046 18244
rect 28077 18241 28089 18244
rect 28123 18241 28135 18275
rect 28077 18235 28135 18241
rect 29454 18232 29460 18284
rect 29512 18232 29518 18284
rect 30285 18275 30343 18281
rect 30285 18241 30297 18275
rect 30331 18272 30343 18275
rect 30558 18272 30564 18284
rect 30331 18244 30564 18272
rect 30331 18241 30343 18244
rect 30285 18235 30343 18241
rect 30558 18232 30564 18244
rect 30616 18232 30622 18284
rect 31573 18275 31631 18281
rect 31573 18241 31585 18275
rect 31619 18272 31631 18275
rect 32784 18272 32812 18371
rect 33594 18368 33600 18380
rect 33652 18368 33658 18420
rect 36906 18368 36912 18420
rect 36964 18408 36970 18420
rect 39393 18411 39451 18417
rect 39393 18408 39405 18411
rect 36964 18380 39405 18408
rect 36964 18368 36970 18380
rect 37734 18340 37740 18352
rect 33244 18312 37740 18340
rect 33244 18281 33272 18312
rect 37734 18300 37740 18312
rect 37792 18300 37798 18352
rect 31619 18244 32812 18272
rect 33229 18275 33287 18281
rect 31619 18241 31631 18244
rect 31573 18235 31631 18241
rect 33229 18241 33241 18275
rect 33275 18241 33287 18275
rect 33229 18235 33287 18241
rect 34238 18232 34244 18284
rect 34296 18272 34302 18284
rect 34793 18275 34851 18281
rect 34793 18272 34805 18275
rect 34296 18244 34805 18272
rect 34296 18232 34302 18244
rect 34793 18241 34805 18244
rect 34839 18241 34851 18275
rect 34793 18235 34851 18241
rect 35802 18232 35808 18284
rect 35860 18272 35866 18284
rect 36725 18275 36783 18281
rect 36725 18272 36737 18275
rect 35860 18244 36737 18272
rect 35860 18232 35866 18244
rect 36725 18241 36737 18244
rect 36771 18241 36783 18275
rect 36725 18235 36783 18241
rect 37182 18232 37188 18284
rect 37240 18272 37246 18284
rect 37553 18275 37611 18281
rect 37553 18272 37565 18275
rect 37240 18244 37565 18272
rect 37240 18232 37246 18244
rect 37553 18241 37565 18244
rect 37599 18241 37611 18275
rect 37553 18235 37611 18241
rect 38197 18275 38255 18281
rect 38197 18241 38209 18275
rect 38243 18272 38255 18275
rect 38654 18272 38660 18284
rect 38243 18244 38660 18272
rect 38243 18241 38255 18244
rect 38197 18235 38255 18241
rect 38654 18232 38660 18244
rect 38712 18232 38718 18284
rect 39132 18281 39160 18380
rect 39393 18377 39405 18380
rect 39439 18377 39451 18411
rect 39393 18371 39451 18377
rect 39117 18275 39175 18281
rect 39117 18241 39129 18275
rect 39163 18241 39175 18275
rect 39117 18235 39175 18241
rect 25130 18204 25136 18216
rect 20824 18176 25136 18204
rect 25130 18164 25136 18176
rect 25188 18204 25194 18216
rect 26142 18204 26148 18216
rect 25188 18176 26148 18204
rect 25188 18164 25194 18176
rect 26142 18164 26148 18176
rect 26200 18164 26206 18216
rect 27154 18164 27160 18216
rect 27212 18164 27218 18216
rect 28353 18207 28411 18213
rect 28353 18173 28365 18207
rect 28399 18204 28411 18207
rect 32950 18204 32956 18216
rect 28399 18176 32956 18204
rect 28399 18173 28411 18176
rect 28353 18167 28411 18173
rect 32950 18164 32956 18176
rect 33008 18164 33014 18216
rect 33410 18164 33416 18216
rect 33468 18204 33474 18216
rect 33505 18207 33563 18213
rect 33505 18204 33517 18207
rect 33468 18176 33517 18204
rect 33468 18164 33474 18176
rect 33505 18173 33517 18176
rect 33551 18173 33563 18207
rect 33505 18167 33563 18173
rect 34514 18164 34520 18216
rect 34572 18164 34578 18216
rect 34624 18176 36676 18204
rect 22462 18136 22468 18148
rect 20732 18108 22468 18136
rect 22462 18096 22468 18108
rect 22520 18096 22526 18148
rect 26510 18096 26516 18148
rect 26568 18136 26574 18148
rect 26568 18108 28212 18136
rect 26568 18096 26574 18108
rect 5994 18028 6000 18080
rect 6052 18068 6058 18080
rect 7098 18068 7104 18080
rect 6052 18040 7104 18068
rect 6052 18028 6058 18040
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 8110 18028 8116 18080
rect 8168 18068 8174 18080
rect 8205 18071 8263 18077
rect 8205 18068 8217 18071
rect 8168 18040 8217 18068
rect 8168 18028 8174 18040
rect 8205 18037 8217 18040
rect 8251 18068 8263 18071
rect 8570 18068 8576 18080
rect 8251 18040 8576 18068
rect 8251 18037 8263 18040
rect 8205 18031 8263 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 8662 18028 8668 18080
rect 8720 18028 8726 18080
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 8812 18040 11529 18068
rect 8812 18028 8818 18040
rect 11517 18037 11529 18040
rect 11563 18068 11575 18071
rect 12894 18068 12900 18080
rect 11563 18040 12900 18068
rect 11563 18037 11575 18040
rect 11517 18031 11575 18037
rect 12894 18028 12900 18040
rect 12952 18068 12958 18080
rect 14366 18068 14372 18080
rect 12952 18040 14372 18068
rect 12952 18028 12958 18040
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14918 18028 14924 18080
rect 14976 18068 14982 18080
rect 18414 18068 18420 18080
rect 14976 18040 18420 18068
rect 14976 18028 14982 18040
rect 18414 18028 18420 18040
rect 18472 18028 18478 18080
rect 18693 18071 18751 18077
rect 18693 18037 18705 18071
rect 18739 18068 18751 18071
rect 20070 18068 20076 18080
rect 18739 18040 20076 18068
rect 18739 18037 18751 18040
rect 18693 18031 18751 18037
rect 20070 18028 20076 18040
rect 20128 18028 20134 18080
rect 20162 18028 20168 18080
rect 20220 18028 20226 18080
rect 20346 18028 20352 18080
rect 20404 18068 20410 18080
rect 20441 18071 20499 18077
rect 20441 18068 20453 18071
rect 20404 18040 20453 18068
rect 20404 18028 20410 18040
rect 20441 18037 20453 18040
rect 20487 18037 20499 18071
rect 20441 18031 20499 18037
rect 23106 18028 23112 18080
rect 23164 18068 23170 18080
rect 23382 18068 23388 18080
rect 23164 18040 23388 18068
rect 23164 18028 23170 18040
rect 23382 18028 23388 18040
rect 23440 18028 23446 18080
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 25498 18068 25504 18080
rect 23532 18040 25504 18068
rect 23532 18028 23538 18040
rect 25498 18028 25504 18040
rect 25556 18028 25562 18080
rect 26605 18071 26663 18077
rect 26605 18037 26617 18071
rect 26651 18068 26663 18071
rect 26789 18071 26847 18077
rect 26789 18068 26801 18071
rect 26651 18040 26801 18068
rect 26651 18037 26663 18040
rect 26605 18031 26663 18037
rect 26789 18037 26801 18040
rect 26835 18068 26847 18071
rect 27062 18068 27068 18080
rect 26835 18040 27068 18068
rect 26835 18037 26847 18040
rect 26789 18031 26847 18037
rect 27062 18028 27068 18040
rect 27120 18028 27126 18080
rect 27709 18071 27767 18077
rect 27709 18037 27721 18071
rect 27755 18068 27767 18071
rect 27798 18068 27804 18080
rect 27755 18040 27804 18068
rect 27755 18037 27767 18040
rect 27709 18031 27767 18037
rect 27798 18028 27804 18040
rect 27856 18028 27862 18080
rect 28184 18068 28212 18108
rect 30558 18096 30564 18148
rect 30616 18136 30622 18148
rect 32401 18139 32459 18145
rect 32401 18136 32413 18139
rect 30616 18108 32413 18136
rect 30616 18096 30622 18108
rect 32401 18105 32413 18108
rect 32447 18136 32459 18139
rect 34624 18136 34652 18176
rect 32447 18108 34652 18136
rect 36648 18136 36676 18176
rect 36814 18164 36820 18216
rect 36872 18204 36878 18216
rect 39850 18204 39856 18216
rect 36872 18176 39856 18204
rect 36872 18164 36878 18176
rect 39850 18164 39856 18176
rect 39908 18164 39914 18216
rect 46842 18136 46848 18148
rect 36648 18108 46848 18136
rect 32447 18105 32459 18108
rect 32401 18099 32459 18105
rect 46842 18096 46848 18108
rect 46900 18096 46906 18148
rect 29825 18071 29883 18077
rect 29825 18068 29837 18071
rect 28184 18040 29837 18068
rect 29825 18037 29837 18040
rect 29871 18068 29883 18071
rect 30834 18068 30840 18080
rect 29871 18040 30840 18068
rect 29871 18037 29883 18040
rect 29825 18031 29883 18037
rect 30834 18028 30840 18040
rect 30892 18028 30898 18080
rect 31662 18028 31668 18080
rect 31720 18068 31726 18080
rect 32493 18071 32551 18077
rect 32493 18068 32505 18071
rect 31720 18040 32505 18068
rect 31720 18028 31726 18040
rect 32493 18037 32505 18040
rect 32539 18037 32551 18071
rect 32493 18031 32551 18037
rect 36446 18028 36452 18080
rect 36504 18028 36510 18080
rect 36722 18028 36728 18080
rect 36780 18068 36786 18080
rect 37001 18071 37059 18077
rect 37001 18068 37013 18071
rect 36780 18040 37013 18068
rect 36780 18028 36786 18040
rect 37001 18037 37013 18040
rect 37047 18068 37059 18071
rect 37182 18068 37188 18080
rect 37047 18040 37188 18068
rect 37047 18037 37059 18040
rect 37001 18031 37059 18037
rect 37182 18028 37188 18040
rect 37240 18028 37246 18080
rect 37642 18028 37648 18080
rect 37700 18028 37706 18080
rect 38378 18028 38384 18080
rect 38436 18028 38442 18080
rect 38930 18028 38936 18080
rect 38988 18028 38994 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 1302 17824 1308 17876
rect 1360 17864 1366 17876
rect 1578 17864 1584 17876
rect 1360 17836 1584 17864
rect 1360 17824 1366 17836
rect 1578 17824 1584 17836
rect 1636 17824 1642 17876
rect 2774 17824 2780 17876
rect 2832 17864 2838 17876
rect 7285 17867 7343 17873
rect 7285 17864 7297 17867
rect 2832 17836 7297 17864
rect 2832 17824 2838 17836
rect 7285 17833 7297 17836
rect 7331 17833 7343 17867
rect 7285 17827 7343 17833
rect 7466 17824 7472 17876
rect 7524 17864 7530 17876
rect 10962 17864 10968 17876
rect 7524 17836 10968 17864
rect 7524 17824 7530 17836
rect 10962 17824 10968 17836
rect 11020 17824 11026 17876
rect 11793 17867 11851 17873
rect 11793 17833 11805 17867
rect 11839 17864 11851 17867
rect 11839 17836 12756 17864
rect 11839 17833 11851 17836
rect 11793 17827 11851 17833
rect 4157 17799 4215 17805
rect 4157 17796 4169 17799
rect 2746 17768 4169 17796
rect 1210 17688 1216 17740
rect 1268 17728 1274 17740
rect 2041 17731 2099 17737
rect 2041 17728 2053 17731
rect 1268 17700 2053 17728
rect 1268 17688 1274 17700
rect 2041 17697 2053 17700
rect 2087 17697 2099 17731
rect 2041 17691 2099 17697
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 2746 17660 2774 17768
rect 4157 17765 4169 17768
rect 4203 17765 4215 17799
rect 4157 17759 4215 17765
rect 6546 17756 6552 17808
rect 6604 17796 6610 17808
rect 11882 17796 11888 17808
rect 6604 17768 11888 17796
rect 6604 17756 6610 17768
rect 11882 17756 11888 17768
rect 11940 17756 11946 17808
rect 12066 17756 12072 17808
rect 12124 17796 12130 17808
rect 12728 17796 12756 17836
rect 12802 17824 12808 17876
rect 12860 17864 12866 17876
rect 12897 17867 12955 17873
rect 12897 17864 12909 17867
rect 12860 17836 12909 17864
rect 12860 17824 12866 17836
rect 12897 17833 12909 17836
rect 12943 17833 12955 17867
rect 12897 17827 12955 17833
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 14550 17864 14556 17876
rect 14323 17836 14556 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 15286 17864 15292 17876
rect 14884 17836 15292 17864
rect 14884 17824 14890 17836
rect 15286 17824 15292 17836
rect 15344 17824 15350 17876
rect 15381 17867 15439 17873
rect 15381 17833 15393 17867
rect 15427 17864 15439 17867
rect 16298 17864 16304 17876
rect 15427 17836 16304 17864
rect 15427 17833 15439 17836
rect 15381 17827 15439 17833
rect 16298 17824 16304 17836
rect 16356 17824 16362 17876
rect 16574 17824 16580 17876
rect 16632 17864 16638 17876
rect 16632 17836 17172 17864
rect 16632 17824 16638 17836
rect 17144 17796 17172 17836
rect 17218 17824 17224 17876
rect 17276 17864 17282 17876
rect 18414 17864 18420 17876
rect 17276 17836 18420 17864
rect 17276 17824 17282 17836
rect 18414 17824 18420 17836
rect 18472 17824 18478 17876
rect 21174 17864 21180 17876
rect 18708 17836 21180 17864
rect 17678 17796 17684 17808
rect 12124 17768 12480 17796
rect 12728 17768 15976 17796
rect 17144 17768 17684 17796
rect 12124 17756 12130 17768
rect 3602 17688 3608 17740
rect 3660 17688 3666 17740
rect 4798 17688 4804 17740
rect 4856 17728 4862 17740
rect 4856 17700 6316 17728
rect 4856 17688 4862 17700
rect 1811 17632 2774 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 3878 17620 3884 17672
rect 3936 17620 3942 17672
rect 4338 17620 4344 17672
rect 4396 17620 4402 17672
rect 6178 17620 6184 17672
rect 6236 17620 6242 17672
rect 6288 17660 6316 17700
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 6972 17700 8401 17728
rect 6972 17688 6978 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9490 17728 9496 17740
rect 9180 17700 9496 17728
rect 9180 17688 9186 17700
rect 9490 17688 9496 17700
rect 9548 17688 9554 17740
rect 10594 17688 10600 17740
rect 10652 17728 10658 17740
rect 10965 17731 11023 17737
rect 10965 17728 10977 17731
rect 10652 17700 10977 17728
rect 10652 17688 10658 17700
rect 10965 17697 10977 17700
rect 11011 17697 11023 17731
rect 10965 17691 11023 17697
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17728 11207 17731
rect 11514 17728 11520 17740
rect 11195 17700 11520 17728
rect 11195 17697 11207 17700
rect 11149 17691 11207 17697
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11606 17688 11612 17740
rect 11664 17728 11670 17740
rect 11790 17728 11796 17740
rect 11664 17700 11796 17728
rect 11664 17688 11670 17700
rect 11790 17688 11796 17700
rect 11848 17688 11854 17740
rect 12342 17688 12348 17740
rect 12400 17688 12406 17740
rect 12452 17728 12480 17768
rect 13541 17731 13599 17737
rect 13541 17728 13553 17731
rect 12452 17700 13553 17728
rect 13541 17697 13553 17700
rect 13587 17728 13599 17731
rect 13722 17728 13728 17740
rect 13587 17700 13728 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 14461 17731 14519 17737
rect 14461 17697 14473 17731
rect 14507 17728 14519 17731
rect 14918 17728 14924 17740
rect 14507 17700 14924 17728
rect 14507 17697 14519 17700
rect 14461 17691 14519 17697
rect 14918 17688 14924 17700
rect 14976 17688 14982 17740
rect 15838 17688 15844 17740
rect 15896 17688 15902 17740
rect 15948 17728 15976 17768
rect 17678 17756 17684 17768
rect 17736 17796 17742 17808
rect 18138 17796 18144 17808
rect 17736 17768 18144 17796
rect 17736 17756 17742 17768
rect 18138 17756 18144 17768
rect 18196 17756 18202 17808
rect 18708 17796 18736 17836
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 22186 17824 22192 17876
rect 22244 17824 22250 17876
rect 22462 17824 22468 17876
rect 22520 17864 22526 17876
rect 24302 17864 24308 17876
rect 22520 17836 24308 17864
rect 22520 17824 22526 17836
rect 24302 17824 24308 17836
rect 24360 17824 24366 17876
rect 25120 17867 25178 17873
rect 25120 17833 25132 17867
rect 25166 17864 25178 17867
rect 30374 17864 30380 17876
rect 25166 17836 30380 17864
rect 25166 17833 25178 17836
rect 25120 17827 25178 17833
rect 30374 17824 30380 17836
rect 30432 17824 30438 17876
rect 35529 17867 35587 17873
rect 35529 17833 35541 17867
rect 35575 17864 35587 17867
rect 37458 17864 37464 17876
rect 35575 17836 37464 17864
rect 35575 17833 35587 17836
rect 35529 17827 35587 17833
rect 37458 17824 37464 17836
rect 37516 17824 37522 17876
rect 38654 17824 38660 17876
rect 38712 17864 38718 17876
rect 45370 17864 45376 17876
rect 38712 17836 45376 17864
rect 38712 17824 38718 17836
rect 45370 17824 45376 17836
rect 45428 17824 45434 17876
rect 20257 17799 20315 17805
rect 20257 17796 20269 17799
rect 18248 17768 18736 17796
rect 18800 17768 20269 17796
rect 17770 17728 17776 17740
rect 15948 17700 17776 17728
rect 17770 17688 17776 17700
rect 17828 17688 17834 17740
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 6288 17632 9873 17660
rect 9861 17629 9873 17632
rect 9907 17629 9919 17663
rect 9861 17623 9919 17629
rect 9950 17620 9956 17672
rect 10008 17660 10014 17672
rect 10008 17632 13492 17660
rect 10008 17620 10014 17632
rect 2498 17552 2504 17604
rect 2556 17592 2562 17604
rect 4246 17592 4252 17604
rect 2556 17564 4252 17592
rect 2556 17552 2562 17564
rect 4246 17552 4252 17564
rect 4304 17552 4310 17604
rect 5077 17595 5135 17601
rect 5077 17561 5089 17595
rect 5123 17592 5135 17595
rect 5166 17592 5172 17604
rect 5123 17564 5172 17592
rect 5123 17561 5135 17564
rect 5077 17555 5135 17561
rect 5166 17552 5172 17564
rect 5224 17552 5230 17604
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17561 7251 17595
rect 7193 17555 7251 17561
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8846 17592 8852 17604
rect 8251 17564 8852 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 1394 17484 1400 17536
rect 1452 17524 1458 17536
rect 3329 17527 3387 17533
rect 3329 17524 3341 17527
rect 1452 17496 3341 17524
rect 1452 17484 1458 17496
rect 3329 17493 3341 17496
rect 3375 17524 3387 17527
rect 6549 17527 6607 17533
rect 6549 17524 6561 17527
rect 3375 17496 6561 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 6549 17493 6561 17496
rect 6595 17524 6607 17527
rect 6822 17524 6828 17536
rect 6595 17496 6828 17524
rect 6595 17493 6607 17496
rect 6549 17487 6607 17493
rect 6822 17484 6828 17496
rect 6880 17484 6886 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7210 17524 7238 17555
rect 8846 17552 8852 17564
rect 8904 17552 8910 17604
rect 8938 17552 8944 17604
rect 8996 17592 9002 17604
rect 9122 17592 9128 17604
rect 8996 17564 9128 17592
rect 8996 17552 9002 17564
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 9214 17552 9220 17604
rect 9272 17592 9278 17604
rect 11514 17592 11520 17604
rect 9272 17564 11520 17592
rect 9272 17552 9278 17564
rect 11514 17552 11520 17564
rect 11572 17552 11578 17604
rect 11609 17595 11667 17601
rect 11609 17561 11621 17595
rect 11655 17592 11667 17595
rect 12069 17595 12127 17601
rect 12069 17592 12081 17595
rect 11655 17564 12081 17592
rect 11655 17561 11667 17564
rect 11609 17555 11667 17561
rect 12069 17561 12081 17564
rect 12115 17592 12127 17595
rect 12115 17564 12480 17592
rect 12115 17561 12127 17564
rect 12069 17555 12127 17561
rect 6972 17496 7238 17524
rect 6972 17484 6978 17496
rect 7834 17484 7840 17536
rect 7892 17484 7898 17536
rect 8297 17527 8355 17533
rect 8297 17493 8309 17527
rect 8343 17524 8355 17527
rect 10505 17527 10563 17533
rect 10505 17524 10517 17527
rect 8343 17496 10517 17524
rect 8343 17493 8355 17496
rect 8297 17487 8355 17493
rect 10505 17493 10517 17496
rect 10551 17493 10563 17527
rect 10505 17487 10563 17493
rect 10594 17484 10600 17536
rect 10652 17524 10658 17536
rect 10873 17527 10931 17533
rect 10873 17524 10885 17527
rect 10652 17496 10885 17524
rect 10652 17484 10658 17496
rect 10873 17493 10885 17496
rect 10919 17493 10931 17527
rect 10873 17487 10931 17493
rect 12250 17484 12256 17536
rect 12308 17484 12314 17536
rect 12452 17524 12480 17564
rect 12526 17552 12532 17604
rect 12584 17592 12590 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 12584 17564 13369 17592
rect 12584 17552 12590 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13464 17592 13492 17632
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 14737 17663 14795 17669
rect 14737 17660 14749 17663
rect 14608 17632 14749 17660
rect 14608 17620 14614 17632
rect 14737 17629 14749 17632
rect 14783 17629 14795 17663
rect 14737 17623 14795 17629
rect 17402 17620 17408 17672
rect 17460 17660 17466 17672
rect 18138 17660 18144 17672
rect 17460 17632 18144 17660
rect 17460 17620 17466 17632
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 18248 17669 18276 17768
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 15838 17592 15844 17604
rect 13464 17564 15844 17592
rect 13357 17555 13415 17561
rect 15838 17552 15844 17564
rect 15896 17552 15902 17604
rect 16114 17552 16120 17604
rect 16172 17552 16178 17604
rect 17494 17592 17500 17604
rect 17342 17564 17500 17592
rect 17494 17552 17500 17564
rect 17552 17552 17558 17604
rect 17862 17552 17868 17604
rect 17920 17592 17926 17604
rect 18800 17592 18828 17768
rect 20257 17765 20269 17768
rect 20303 17765 20315 17799
rect 22002 17796 22008 17808
rect 20257 17759 20315 17765
rect 20456 17768 22008 17796
rect 18877 17731 18935 17737
rect 18877 17697 18889 17731
rect 18923 17728 18935 17731
rect 20456 17728 20484 17768
rect 22002 17756 22008 17768
rect 22060 17756 22066 17808
rect 18923 17700 20484 17728
rect 18923 17697 18935 17700
rect 18877 17691 18935 17697
rect 20622 17688 20628 17740
rect 20680 17728 20686 17740
rect 20901 17731 20959 17737
rect 20901 17728 20913 17731
rect 20680 17700 20913 17728
rect 20680 17688 20686 17700
rect 20901 17697 20913 17700
rect 20947 17728 20959 17731
rect 22204 17728 22232 17824
rect 26142 17756 26148 17808
rect 26200 17796 26206 17808
rect 26605 17799 26663 17805
rect 26605 17796 26617 17799
rect 26200 17768 26617 17796
rect 26200 17756 26206 17768
rect 26605 17765 26617 17768
rect 26651 17765 26663 17799
rect 26605 17759 26663 17765
rect 28442 17756 28448 17808
rect 28500 17796 28506 17808
rect 28813 17799 28871 17805
rect 28500 17768 28764 17796
rect 28500 17756 28506 17768
rect 22373 17731 22431 17737
rect 22373 17728 22385 17731
rect 20947 17700 21864 17728
rect 22204 17700 22385 17728
rect 20947 17697 20959 17700
rect 20901 17691 20959 17697
rect 18966 17620 18972 17672
rect 19024 17660 19030 17672
rect 21634 17660 21640 17672
rect 19024 17632 21640 17660
rect 19024 17620 19030 17632
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 17920 17564 18828 17592
rect 17920 17552 17926 17564
rect 18874 17552 18880 17604
rect 18932 17592 18938 17604
rect 19242 17592 19248 17604
rect 18932 17564 19248 17592
rect 18932 17552 18938 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19521 17595 19579 17601
rect 19521 17561 19533 17595
rect 19567 17592 19579 17595
rect 21266 17592 21272 17604
rect 19567 17564 21272 17592
rect 19567 17561 19579 17564
rect 19521 17555 19579 17561
rect 21266 17552 21272 17564
rect 21324 17552 21330 17604
rect 21836 17592 21864 17700
rect 22373 17697 22385 17700
rect 22419 17697 22431 17731
rect 24670 17728 24676 17740
rect 22373 17691 22431 17697
rect 23400 17700 24676 17728
rect 23400 17672 23428 17700
rect 24670 17688 24676 17700
rect 24728 17728 24734 17740
rect 24857 17731 24915 17737
rect 24857 17728 24869 17731
rect 24728 17700 24869 17728
rect 24728 17688 24734 17700
rect 24857 17697 24869 17700
rect 24903 17728 24915 17731
rect 25774 17728 25780 17740
rect 24903 17700 25780 17728
rect 24903 17697 24915 17700
rect 24857 17691 24915 17697
rect 25774 17688 25780 17700
rect 25832 17728 25838 17740
rect 27065 17731 27123 17737
rect 27065 17728 27077 17731
rect 25832 17700 27077 17728
rect 25832 17688 25838 17700
rect 27065 17697 27077 17700
rect 27111 17728 27123 17731
rect 27982 17728 27988 17740
rect 27111 17700 27988 17728
rect 27111 17697 27123 17700
rect 27065 17691 27123 17697
rect 27982 17688 27988 17700
rect 28040 17688 28046 17740
rect 28736 17728 28764 17768
rect 28813 17765 28825 17799
rect 28859 17796 28871 17799
rect 30190 17796 30196 17808
rect 28859 17768 30196 17796
rect 28859 17765 28871 17768
rect 28813 17759 28871 17765
rect 30190 17756 30196 17768
rect 30248 17756 30254 17808
rect 31570 17756 31576 17808
rect 31628 17796 31634 17808
rect 31628 17768 32812 17796
rect 31628 17756 31634 17768
rect 29181 17731 29239 17737
rect 29181 17728 29193 17731
rect 28736 17700 29193 17728
rect 29181 17697 29193 17700
rect 29227 17728 29239 17731
rect 29454 17728 29460 17740
rect 29227 17700 29460 17728
rect 29227 17697 29239 17700
rect 29181 17691 29239 17697
rect 29454 17688 29460 17700
rect 29512 17688 29518 17740
rect 30285 17731 30343 17737
rect 30285 17697 30297 17731
rect 30331 17728 30343 17731
rect 31018 17728 31024 17740
rect 30331 17700 31024 17728
rect 30331 17697 30343 17700
rect 30285 17691 30343 17697
rect 31018 17688 31024 17700
rect 31076 17688 31082 17740
rect 22002 17620 22008 17672
rect 22060 17660 22066 17672
rect 22097 17663 22155 17669
rect 22097 17660 22109 17663
rect 22060 17632 22109 17660
rect 22060 17620 22066 17632
rect 22097 17629 22109 17632
rect 22143 17629 22155 17663
rect 22097 17623 22155 17629
rect 23382 17620 23388 17672
rect 23440 17620 23446 17672
rect 23658 17660 23664 17672
rect 23506 17632 23664 17660
rect 23658 17620 23664 17632
rect 23716 17620 23722 17672
rect 23750 17620 23756 17672
rect 23808 17660 23814 17672
rect 24397 17663 24455 17669
rect 24397 17660 24409 17663
rect 23808 17632 24409 17660
rect 23808 17620 23814 17632
rect 24397 17629 24409 17632
rect 24443 17629 24455 17663
rect 24397 17623 24455 17629
rect 26786 17620 26792 17672
rect 26844 17660 26850 17672
rect 26970 17660 26976 17672
rect 26844 17632 26976 17660
rect 26844 17620 26850 17632
rect 26970 17620 26976 17632
rect 27028 17620 27034 17672
rect 28442 17620 28448 17672
rect 28500 17620 28506 17672
rect 30834 17620 30840 17672
rect 30892 17660 30898 17672
rect 30929 17663 30987 17669
rect 30929 17660 30941 17663
rect 30892 17632 30941 17660
rect 30892 17620 30898 17632
rect 30929 17629 30941 17632
rect 30975 17629 30987 17663
rect 30929 17623 30987 17629
rect 32030 17620 32036 17672
rect 32088 17620 32094 17672
rect 27062 17592 27068 17604
rect 21836 17564 22600 17592
rect 12618 17524 12624 17536
rect 12452 17496 12624 17524
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 14366 17524 14372 17536
rect 13320 17496 14372 17524
rect 13320 17484 13326 17496
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 16850 17524 16856 17536
rect 14516 17496 16856 17524
rect 14516 17484 14522 17496
rect 16850 17484 16856 17496
rect 16908 17484 16914 17536
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 19426 17524 19432 17536
rect 17644 17496 19432 17524
rect 17644 17484 17650 17496
rect 19426 17484 19432 17496
rect 19484 17484 19490 17536
rect 19610 17484 19616 17536
rect 19668 17484 19674 17536
rect 20254 17484 20260 17536
rect 20312 17524 20318 17536
rect 20622 17524 20628 17536
rect 20312 17496 20628 17524
rect 20312 17484 20318 17496
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 20717 17527 20775 17533
rect 20717 17493 20729 17527
rect 20763 17524 20775 17527
rect 20898 17524 20904 17536
rect 20763 17496 20904 17524
rect 20763 17493 20775 17496
rect 20717 17487 20775 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 21453 17527 21511 17533
rect 21453 17493 21465 17527
rect 21499 17524 21511 17527
rect 22462 17524 22468 17536
rect 21499 17496 22468 17524
rect 21499 17493 21511 17496
rect 21453 17487 21511 17493
rect 22462 17484 22468 17496
rect 22520 17484 22526 17536
rect 22572 17524 22600 17564
rect 23676 17564 24440 17592
rect 26358 17564 27068 17592
rect 23676 17524 23704 17564
rect 22572 17496 23704 17524
rect 23842 17484 23848 17536
rect 23900 17484 23906 17536
rect 24213 17527 24271 17533
rect 24213 17493 24225 17527
rect 24259 17524 24271 17527
rect 24302 17524 24308 17536
rect 24259 17496 24308 17524
rect 24259 17493 24271 17496
rect 24213 17487 24271 17493
rect 24302 17484 24308 17496
rect 24360 17484 24366 17536
rect 24412 17524 24440 17564
rect 27062 17552 27068 17564
rect 27120 17552 27126 17604
rect 27341 17595 27399 17601
rect 27341 17561 27353 17595
rect 27387 17592 27399 17595
rect 27430 17592 27436 17604
rect 27387 17564 27436 17592
rect 27387 17561 27399 17564
rect 27341 17555 27399 17561
rect 27430 17552 27436 17564
rect 27488 17552 27494 17604
rect 29270 17552 29276 17604
rect 29328 17552 29334 17604
rect 32784 17592 32812 17768
rect 32858 17756 32864 17808
rect 32916 17796 32922 17808
rect 36630 17796 36636 17808
rect 32916 17768 36636 17796
rect 32916 17756 32922 17768
rect 36630 17756 36636 17768
rect 36688 17756 36694 17808
rect 36906 17756 36912 17808
rect 36964 17756 36970 17808
rect 33781 17731 33839 17737
rect 33781 17697 33793 17731
rect 33827 17728 33839 17731
rect 36262 17728 36268 17740
rect 33827 17700 36268 17728
rect 33827 17697 33839 17700
rect 33781 17691 33839 17697
rect 36262 17688 36268 17700
rect 36320 17688 36326 17740
rect 33137 17663 33195 17669
rect 33137 17629 33149 17663
rect 33183 17660 33195 17663
rect 33318 17660 33324 17672
rect 33183 17632 33324 17660
rect 33183 17629 33195 17632
rect 33137 17623 33195 17629
rect 33318 17620 33324 17632
rect 33376 17660 33382 17672
rect 34241 17663 34299 17669
rect 34241 17660 34253 17663
rect 33376 17632 34253 17660
rect 33376 17620 33382 17632
rect 34241 17629 34253 17632
rect 34287 17629 34299 17663
rect 34241 17623 34299 17629
rect 34606 17620 34612 17672
rect 34664 17660 34670 17672
rect 34885 17663 34943 17669
rect 34885 17660 34897 17663
rect 34664 17632 34897 17660
rect 34664 17620 34670 17632
rect 34885 17629 34897 17632
rect 34931 17629 34943 17663
rect 34885 17623 34943 17629
rect 35894 17620 35900 17672
rect 35952 17660 35958 17672
rect 36173 17663 36231 17669
rect 36173 17660 36185 17663
rect 35952 17632 36185 17660
rect 35952 17620 35958 17632
rect 36173 17629 36185 17632
rect 36219 17629 36231 17663
rect 36998 17660 37004 17672
rect 36173 17623 36231 17629
rect 36648 17632 37004 17660
rect 36648 17592 36676 17632
rect 36998 17620 37004 17632
rect 37056 17620 37062 17672
rect 37458 17620 37464 17672
rect 37516 17660 37522 17672
rect 37553 17663 37611 17669
rect 37553 17660 37565 17663
rect 37516 17632 37565 17660
rect 37516 17620 37522 17632
rect 37553 17629 37565 17632
rect 37599 17660 37611 17663
rect 37829 17663 37887 17669
rect 37829 17660 37841 17663
rect 37599 17632 37841 17660
rect 37599 17629 37611 17632
rect 37553 17623 37611 17629
rect 37829 17629 37841 17632
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 32784 17564 36676 17592
rect 36725 17595 36783 17601
rect 36725 17561 36737 17595
rect 36771 17592 36783 17595
rect 39298 17592 39304 17604
rect 36771 17564 39304 17592
rect 36771 17561 36783 17564
rect 36725 17555 36783 17561
rect 39298 17552 39304 17564
rect 39356 17552 39362 17604
rect 28258 17524 28264 17536
rect 24412 17496 28264 17524
rect 28258 17484 28264 17496
rect 28316 17484 28322 17536
rect 29638 17484 29644 17536
rect 29696 17524 29702 17536
rect 29733 17527 29791 17533
rect 29733 17524 29745 17527
rect 29696 17496 29745 17524
rect 29696 17484 29702 17496
rect 29733 17493 29745 17496
rect 29779 17493 29791 17527
rect 29733 17487 29791 17493
rect 30098 17484 30104 17536
rect 30156 17484 30162 17536
rect 30190 17484 30196 17536
rect 30248 17524 30254 17536
rect 30558 17524 30564 17536
rect 30248 17496 30564 17524
rect 30248 17484 30254 17496
rect 30558 17484 30564 17496
rect 30616 17484 30622 17536
rect 31202 17484 31208 17536
rect 31260 17524 31266 17536
rect 31573 17527 31631 17533
rect 31573 17524 31585 17527
rect 31260 17496 31585 17524
rect 31260 17484 31266 17496
rect 31573 17493 31585 17496
rect 31619 17493 31631 17527
rect 31573 17487 31631 17493
rect 32674 17484 32680 17536
rect 32732 17484 32738 17536
rect 34054 17484 34060 17536
rect 34112 17484 34118 17536
rect 34517 17527 34575 17533
rect 34517 17493 34529 17527
rect 34563 17524 34575 17527
rect 34606 17524 34612 17536
rect 34563 17496 34612 17524
rect 34563 17493 34575 17496
rect 34517 17487 34575 17493
rect 34606 17484 34612 17496
rect 34664 17484 34670 17536
rect 35989 17527 36047 17533
rect 35989 17493 36001 17527
rect 36035 17524 36047 17527
rect 36078 17524 36084 17536
rect 36035 17496 36084 17524
rect 36035 17493 36047 17496
rect 35989 17487 36047 17493
rect 36078 17484 36084 17496
rect 36136 17484 36142 17536
rect 37366 17484 37372 17536
rect 37424 17484 37430 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 5261 17323 5319 17329
rect 5261 17289 5273 17323
rect 5307 17289 5319 17323
rect 5261 17283 5319 17289
rect 5721 17323 5779 17329
rect 5721 17289 5733 17323
rect 5767 17320 5779 17323
rect 7650 17320 7656 17332
rect 5767 17292 7656 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 5276 17252 5304 17283
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 8018 17280 8024 17332
rect 8076 17280 8082 17332
rect 8570 17280 8576 17332
rect 8628 17320 8634 17332
rect 9858 17320 9864 17332
rect 8628 17292 9864 17320
rect 8628 17280 8634 17292
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 9953 17323 10011 17329
rect 9953 17289 9965 17323
rect 9999 17320 10011 17323
rect 10226 17320 10232 17332
rect 9999 17292 10232 17320
rect 9999 17289 10011 17292
rect 9953 17283 10011 17289
rect 10226 17280 10232 17292
rect 10284 17320 10290 17332
rect 10781 17323 10839 17329
rect 10781 17320 10793 17323
rect 10284 17292 10793 17320
rect 10284 17280 10290 17292
rect 10781 17289 10793 17292
rect 10827 17289 10839 17323
rect 10781 17283 10839 17289
rect 10962 17280 10968 17332
rect 11020 17320 11026 17332
rect 14090 17320 14096 17332
rect 11020 17292 14096 17320
rect 11020 17280 11026 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14182 17280 14188 17332
rect 14240 17320 14246 17332
rect 14737 17323 14795 17329
rect 14737 17320 14749 17323
rect 14240 17292 14749 17320
rect 14240 17280 14246 17292
rect 14737 17289 14749 17292
rect 14783 17289 14795 17323
rect 14737 17283 14795 17289
rect 14826 17280 14832 17332
rect 14884 17320 14890 17332
rect 17037 17323 17095 17329
rect 17037 17320 17049 17323
rect 14884 17292 17049 17320
rect 14884 17280 14890 17292
rect 17037 17289 17049 17292
rect 17083 17289 17095 17323
rect 17037 17283 17095 17289
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 17552 17292 18276 17320
rect 17552 17280 17558 17292
rect 10594 17252 10600 17264
rect 5276 17224 10600 17252
rect 10594 17212 10600 17224
rect 10652 17212 10658 17264
rect 10980 17252 11008 17280
rect 10704 17224 11008 17252
rect 1762 17144 1768 17196
rect 1820 17144 1826 17196
rect 3605 17187 3663 17193
rect 3605 17153 3617 17187
rect 3651 17184 3663 17187
rect 4246 17184 4252 17196
rect 3651 17156 4252 17184
rect 3651 17153 3663 17156
rect 3605 17147 3663 17153
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 5629 17187 5687 17193
rect 5629 17153 5641 17187
rect 5675 17184 5687 17187
rect 6362 17184 6368 17196
rect 5675 17156 6368 17184
rect 5675 17153 5687 17156
rect 5629 17147 5687 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 6546 17144 6552 17196
rect 6604 17144 6610 17196
rect 7190 17144 7196 17196
rect 7248 17144 7254 17196
rect 8570 17184 8576 17196
rect 7392 17156 8576 17184
rect 1302 17076 1308 17128
rect 1360 17116 1366 17128
rect 2041 17119 2099 17125
rect 2041 17116 2053 17119
rect 1360 17088 2053 17116
rect 1360 17076 1366 17088
rect 2041 17085 2053 17088
rect 2087 17085 2099 17119
rect 2041 17079 2099 17085
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 5902 17076 5908 17128
rect 5960 17116 5966 17128
rect 6822 17116 6828 17128
rect 5960 17088 6828 17116
rect 5960 17076 5966 17088
rect 6822 17076 6828 17088
rect 6880 17076 6886 17128
rect 6914 17076 6920 17128
rect 6972 17116 6978 17128
rect 7392 17116 7420 17156
rect 8570 17144 8576 17156
rect 8628 17144 8634 17196
rect 9217 17187 9275 17193
rect 9217 17153 9229 17187
rect 9263 17184 9275 17187
rect 10704 17184 10732 17224
rect 11974 17212 11980 17264
rect 12032 17252 12038 17264
rect 14108 17252 14136 17280
rect 15102 17252 15108 17264
rect 12032 17224 12466 17252
rect 14108 17224 15108 17252
rect 12032 17212 12038 17224
rect 15102 17212 15108 17224
rect 15160 17212 15166 17264
rect 15473 17255 15531 17261
rect 15473 17221 15485 17255
rect 15519 17252 15531 17255
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 15519 17224 15945 17252
rect 15519 17221 15531 17224
rect 15473 17215 15531 17221
rect 15933 17221 15945 17224
rect 15979 17252 15991 17255
rect 17126 17252 17132 17264
rect 15979 17224 17132 17252
rect 15979 17221 15991 17224
rect 15933 17215 15991 17221
rect 17126 17212 17132 17224
rect 17184 17212 17190 17264
rect 17218 17212 17224 17264
rect 17276 17252 17282 17264
rect 17276 17224 17724 17252
rect 17276 17212 17282 17224
rect 9263 17156 10732 17184
rect 10873 17187 10931 17193
rect 9263 17153 9275 17156
rect 9217 17147 9275 17153
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 11054 17184 11060 17196
rect 10919 17156 11060 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11698 17144 11704 17196
rect 11756 17144 11762 17196
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 15654 17184 15660 17196
rect 14332 17156 15660 17184
rect 14332 17144 14338 17156
rect 15654 17144 15660 17156
rect 15712 17144 15718 17196
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17405 17187 17463 17193
rect 17405 17184 17417 17187
rect 17000 17156 17417 17184
rect 17000 17144 17006 17156
rect 17405 17153 17417 17156
rect 17451 17153 17463 17187
rect 17405 17147 17463 17153
rect 6972 17088 7420 17116
rect 6972 17076 6978 17088
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 8113 17119 8171 17125
rect 8113 17116 8125 17119
rect 7524 17088 8125 17116
rect 7524 17076 7530 17088
rect 8113 17085 8125 17088
rect 8159 17085 8171 17119
rect 8113 17079 8171 17085
rect 8202 17076 8208 17128
rect 8260 17076 8266 17128
rect 9306 17076 9312 17128
rect 9364 17076 9370 17128
rect 9490 17076 9496 17128
rect 9548 17076 9554 17128
rect 10318 17076 10324 17128
rect 10376 17116 10382 17128
rect 10594 17116 10600 17128
rect 10376 17088 10600 17116
rect 10376 17076 10382 17088
rect 10594 17076 10600 17088
rect 10652 17116 10658 17128
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10652 17088 10977 17116
rect 10652 17076 10658 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 10965 17079 11023 17085
rect 11072 17088 11989 17116
rect 5718 17008 5724 17060
rect 5776 17048 5782 17060
rect 8849 17051 8907 17057
rect 8849 17048 8861 17051
rect 5776 17020 8861 17048
rect 5776 17008 5782 17020
rect 8849 17017 8861 17020
rect 8895 17017 8907 17051
rect 8849 17011 8907 17017
rect 10778 17008 10784 17060
rect 10836 17048 10842 17060
rect 11072 17048 11100 17088
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 11977 17079 12035 17085
rect 12618 17076 12624 17128
rect 12676 17116 12682 17128
rect 14642 17116 14648 17128
rect 12676 17088 14648 17116
rect 12676 17076 12682 17088
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 14826 17076 14832 17128
rect 14884 17076 14890 17128
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 15746 17116 15752 17128
rect 15059 17088 15752 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 16022 17076 16028 17128
rect 16080 17076 16086 17128
rect 16206 17076 16212 17128
rect 16264 17076 16270 17128
rect 17696 17116 17724 17224
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 18141 17255 18199 17261
rect 18141 17252 18153 17255
rect 17920 17224 18153 17252
rect 17920 17212 17926 17224
rect 18141 17221 18153 17224
rect 18187 17221 18199 17255
rect 18248 17252 18276 17292
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 18380 17292 20576 17320
rect 18380 17280 18386 17292
rect 18248 17224 18630 17252
rect 18141 17215 18199 17221
rect 19794 17212 19800 17264
rect 19852 17252 19858 17264
rect 20346 17252 20352 17264
rect 19852 17224 20352 17252
rect 19852 17212 19858 17224
rect 20346 17212 20352 17224
rect 20404 17212 20410 17264
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20441 17187 20499 17193
rect 20441 17184 20453 17187
rect 19668 17156 20453 17184
rect 19668 17144 19674 17156
rect 20441 17153 20453 17156
rect 20487 17153 20499 17187
rect 20548 17184 20576 17292
rect 20714 17280 20720 17332
rect 20772 17320 20778 17332
rect 21269 17323 21327 17329
rect 21269 17320 21281 17323
rect 20772 17292 21281 17320
rect 20772 17280 20778 17292
rect 21269 17289 21281 17292
rect 21315 17289 21327 17323
rect 22186 17320 22192 17332
rect 21269 17283 21327 17289
rect 21468 17292 22192 17320
rect 21174 17212 21180 17264
rect 21232 17252 21238 17264
rect 21468 17252 21496 17292
rect 22186 17280 22192 17292
rect 22244 17280 22250 17332
rect 22462 17280 22468 17332
rect 22520 17280 22526 17332
rect 22557 17323 22615 17329
rect 22557 17289 22569 17323
rect 22603 17320 22615 17323
rect 23198 17320 23204 17332
rect 22603 17292 23204 17320
rect 22603 17289 22615 17292
rect 22557 17283 22615 17289
rect 23198 17280 23204 17292
rect 23256 17280 23262 17332
rect 23750 17280 23756 17332
rect 23808 17320 23814 17332
rect 23845 17323 23903 17329
rect 23845 17320 23857 17323
rect 23808 17292 23857 17320
rect 23808 17280 23814 17292
rect 23845 17289 23857 17292
rect 23891 17289 23903 17323
rect 27338 17320 27344 17332
rect 23845 17283 23903 17289
rect 24596 17292 27344 17320
rect 23937 17255 23995 17261
rect 21232 17224 21496 17252
rect 21560 17224 23888 17252
rect 21232 17212 21238 17224
rect 21453 17187 21511 17193
rect 21453 17184 21465 17187
rect 20548 17156 21465 17184
rect 20441 17147 20499 17153
rect 21453 17153 21465 17156
rect 21499 17153 21511 17187
rect 21453 17147 21511 17153
rect 17865 17119 17923 17125
rect 17865 17116 17877 17119
rect 17696 17088 17877 17116
rect 17865 17085 17877 17088
rect 17911 17085 17923 17119
rect 20162 17116 20168 17128
rect 17865 17079 17923 17085
rect 19720 17088 20168 17116
rect 10836 17020 11100 17048
rect 13909 17051 13967 17057
rect 10836 17008 10842 17020
rect 13909 17017 13921 17051
rect 13955 17048 13967 17051
rect 14369 17051 14427 17057
rect 13955 17020 14228 17048
rect 13955 17017 13967 17020
rect 13909 17011 13967 17017
rect 7653 16983 7711 16989
rect 7653 16949 7665 16983
rect 7699 16980 7711 16983
rect 9950 16980 9956 16992
rect 7699 16952 9956 16980
rect 7699 16949 7711 16952
rect 7653 16943 7711 16949
rect 9950 16940 9956 16952
rect 10008 16940 10014 16992
rect 10045 16983 10103 16989
rect 10045 16949 10057 16983
rect 10091 16980 10103 16983
rect 10318 16980 10324 16992
rect 10091 16952 10324 16980
rect 10091 16949 10103 16952
rect 10045 16943 10103 16949
rect 10318 16940 10324 16952
rect 10376 16940 10382 16992
rect 10410 16940 10416 16992
rect 10468 16940 10474 16992
rect 11974 16940 11980 16992
rect 12032 16980 12038 16992
rect 12618 16980 12624 16992
rect 12032 16952 12624 16980
rect 12032 16940 12038 16952
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 13446 16940 13452 16992
rect 13504 16940 13510 16992
rect 13630 16940 13636 16992
rect 13688 16980 13694 16992
rect 13924 16980 13952 17011
rect 13688 16952 13952 16980
rect 13688 16940 13694 16952
rect 14090 16940 14096 16992
rect 14148 16940 14154 16992
rect 14200 16980 14228 17020
rect 14369 17017 14381 17051
rect 14415 17048 14427 17051
rect 15378 17048 15384 17060
rect 14415 17020 15384 17048
rect 14415 17017 14427 17020
rect 14369 17011 14427 17017
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 17586 17048 17592 17060
rect 15488 17020 17592 17048
rect 15488 16980 15516 17020
rect 17586 17008 17592 17020
rect 17644 17008 17650 17060
rect 19150 17008 19156 17060
rect 19208 17048 19214 17060
rect 19613 17051 19671 17057
rect 19613 17048 19625 17051
rect 19208 17020 19625 17048
rect 19208 17008 19214 17020
rect 19613 17017 19625 17020
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 14200 16952 15516 16980
rect 15565 16983 15623 16989
rect 15565 16949 15577 16983
rect 15611 16980 15623 16983
rect 16758 16980 16764 16992
rect 15611 16952 16764 16980
rect 15611 16949 15623 16952
rect 15565 16943 15623 16949
rect 16758 16940 16764 16952
rect 16816 16940 16822 16992
rect 16850 16940 16856 16992
rect 16908 16980 16914 16992
rect 19720 16980 19748 17088
rect 20162 17076 20168 17088
rect 20220 17116 20226 17128
rect 20533 17119 20591 17125
rect 20533 17116 20545 17119
rect 20220 17088 20545 17116
rect 20220 17076 20226 17088
rect 20533 17085 20545 17088
rect 20579 17085 20591 17119
rect 20533 17079 20591 17085
rect 20625 17119 20683 17125
rect 20625 17085 20637 17119
rect 20671 17116 20683 17119
rect 21560 17116 21588 17224
rect 21634 17144 21640 17196
rect 21692 17184 21698 17196
rect 23750 17184 23756 17196
rect 21692 17156 23756 17184
rect 21692 17144 21698 17156
rect 23750 17144 23756 17156
rect 23808 17144 23814 17196
rect 23860 17184 23888 17224
rect 23937 17221 23949 17255
rect 23983 17252 23995 17255
rect 24302 17252 24308 17264
rect 23983 17224 24308 17252
rect 23983 17221 23995 17224
rect 23937 17215 23995 17221
rect 24302 17212 24308 17224
rect 24360 17212 24366 17264
rect 24596 17184 24624 17292
rect 27338 17280 27344 17292
rect 27396 17320 27402 17332
rect 29641 17323 29699 17329
rect 29641 17320 29653 17323
rect 27396 17292 29653 17320
rect 27396 17280 27402 17292
rect 29641 17289 29653 17292
rect 29687 17289 29699 17323
rect 29641 17283 29699 17289
rect 30745 17323 30803 17329
rect 30745 17289 30757 17323
rect 30791 17320 30803 17323
rect 32030 17320 32036 17332
rect 30791 17292 32036 17320
rect 30791 17289 30803 17292
rect 30745 17283 30803 17289
rect 27062 17252 27068 17264
rect 26174 17224 27068 17252
rect 27062 17212 27068 17224
rect 27120 17252 27126 17264
rect 28442 17252 28448 17264
rect 27120 17224 28448 17252
rect 27120 17212 27126 17224
rect 28442 17212 28448 17224
rect 28500 17212 28506 17264
rect 29454 17252 29460 17264
rect 29394 17224 29460 17252
rect 29454 17212 29460 17224
rect 29512 17212 29518 17264
rect 29656 17252 29684 17283
rect 32030 17280 32036 17292
rect 32088 17280 32094 17332
rect 34057 17323 34115 17329
rect 34057 17289 34069 17323
rect 34103 17320 34115 17323
rect 34514 17320 34520 17332
rect 34103 17292 34520 17320
rect 34103 17289 34115 17292
rect 34057 17283 34115 17289
rect 34514 17280 34520 17292
rect 34572 17280 34578 17332
rect 35894 17280 35900 17332
rect 35952 17280 35958 17332
rect 41598 17320 41604 17332
rect 36004 17292 41604 17320
rect 30834 17252 30840 17264
rect 29656 17224 30840 17252
rect 30834 17212 30840 17224
rect 30892 17212 30898 17264
rect 31573 17255 31631 17261
rect 31573 17221 31585 17255
rect 31619 17252 31631 17255
rect 31662 17252 31668 17264
rect 31619 17224 31668 17252
rect 31619 17221 31631 17224
rect 31573 17215 31631 17221
rect 31662 17212 31668 17224
rect 31720 17212 31726 17264
rect 32232 17224 32720 17252
rect 23860 17156 24624 17184
rect 24670 17144 24676 17196
rect 24728 17144 24734 17196
rect 26786 17144 26792 17196
rect 26844 17144 26850 17196
rect 27522 17144 27528 17196
rect 27580 17184 27586 17196
rect 27893 17187 27951 17193
rect 27893 17184 27905 17187
rect 27580 17156 27905 17184
rect 27580 17144 27586 17156
rect 27893 17153 27905 17156
rect 27939 17153 27951 17187
rect 27893 17147 27951 17153
rect 30101 17187 30159 17193
rect 30101 17153 30113 17187
rect 30147 17184 30159 17187
rect 30282 17184 30288 17196
rect 30147 17156 30288 17184
rect 30147 17153 30159 17156
rect 30101 17147 30159 17153
rect 30282 17144 30288 17156
rect 30340 17144 30346 17196
rect 31110 17144 31116 17196
rect 31168 17184 31174 17196
rect 32232 17184 32260 17224
rect 31168 17156 32260 17184
rect 32309 17187 32367 17193
rect 31168 17144 31174 17156
rect 32309 17153 32321 17187
rect 32355 17153 32367 17187
rect 32309 17147 32367 17153
rect 22462 17116 22468 17128
rect 20671 17088 21588 17116
rect 21652 17088 22468 17116
rect 20671 17085 20683 17088
rect 20625 17079 20683 17085
rect 20073 17051 20131 17057
rect 20073 17017 20085 17051
rect 20119 17048 20131 17051
rect 20119 17020 21404 17048
rect 20119 17017 20131 17020
rect 20073 17011 20131 17017
rect 16908 16952 19748 16980
rect 16908 16940 16914 16952
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 20898 16980 20904 16992
rect 20312 16952 20904 16980
rect 20312 16940 20318 16952
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 21376 16980 21404 17020
rect 21450 17008 21456 17060
rect 21508 17048 21514 17060
rect 21652 17048 21680 17088
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 22741 17119 22799 17125
rect 22741 17085 22753 17119
rect 22787 17116 22799 17119
rect 22787 17088 24072 17116
rect 22787 17085 22799 17088
rect 22741 17079 22799 17085
rect 21508 17020 21680 17048
rect 21508 17008 21514 17020
rect 22094 17008 22100 17060
rect 22152 17008 22158 17060
rect 23201 17051 23259 17057
rect 23201 17017 23213 17051
rect 23247 17048 23259 17051
rect 23658 17048 23664 17060
rect 23247 17020 23664 17048
rect 23247 17017 23259 17020
rect 23201 17011 23259 17017
rect 23658 17008 23664 17020
rect 23716 17008 23722 17060
rect 22738 16980 22744 16992
rect 21376 16952 22744 16980
rect 22738 16940 22744 16952
rect 22796 16940 22802 16992
rect 23474 16940 23480 16992
rect 23532 16940 23538 16992
rect 24044 16980 24072 17088
rect 24118 17076 24124 17128
rect 24176 17116 24182 17128
rect 24394 17116 24400 17128
rect 24176 17088 24400 17116
rect 24176 17076 24182 17088
rect 24394 17076 24400 17088
rect 24452 17076 24458 17128
rect 24949 17119 25007 17125
rect 24949 17085 24961 17119
rect 24995 17116 25007 17119
rect 26142 17116 26148 17128
rect 24995 17088 26148 17116
rect 24995 17085 25007 17088
rect 24949 17079 25007 17085
rect 26142 17076 26148 17088
rect 26200 17076 26206 17128
rect 27246 17076 27252 17128
rect 27304 17076 27310 17128
rect 28169 17119 28227 17125
rect 28169 17085 28181 17119
rect 28215 17116 28227 17119
rect 28902 17116 28908 17128
rect 28215 17088 28908 17116
rect 28215 17085 28227 17088
rect 28169 17079 28227 17085
rect 28902 17076 28908 17088
rect 28960 17076 28966 17128
rect 29178 17076 29184 17128
rect 29236 17116 29242 17128
rect 31294 17116 31300 17128
rect 29236 17088 31300 17116
rect 29236 17076 29242 17088
rect 31294 17076 31300 17088
rect 31352 17076 31358 17128
rect 32324 17116 32352 17147
rect 31404 17088 32352 17116
rect 26421 17051 26479 17057
rect 26421 17017 26433 17051
rect 26467 17017 26479 17051
rect 31404 17048 31432 17088
rect 26421 17011 26479 17017
rect 30484 17020 31432 17048
rect 31757 17051 31815 17057
rect 26436 16980 26464 17011
rect 30484 16980 30512 17020
rect 31757 17017 31769 17051
rect 31803 17048 31815 17051
rect 31938 17048 31944 17060
rect 31803 17020 31944 17048
rect 31803 17017 31815 17020
rect 31757 17011 31815 17017
rect 31938 17008 31944 17020
rect 31996 17008 32002 17060
rect 32692 17048 32720 17224
rect 33413 17187 33471 17193
rect 33413 17153 33425 17187
rect 33459 17184 33471 17187
rect 34054 17184 34060 17196
rect 33459 17156 34060 17184
rect 33459 17153 33471 17156
rect 33413 17147 33471 17153
rect 34054 17144 34060 17156
rect 34112 17144 34118 17196
rect 34514 17144 34520 17196
rect 34572 17184 34578 17196
rect 34609 17187 34667 17193
rect 34609 17184 34621 17187
rect 34572 17156 34621 17184
rect 34572 17144 34578 17156
rect 34609 17153 34621 17156
rect 34655 17153 34667 17187
rect 36004 17184 36032 17292
rect 41598 17280 41604 17292
rect 41656 17280 41662 17332
rect 47394 17252 47400 17264
rect 41386 17224 47400 17252
rect 34609 17147 34667 17153
rect 34716 17156 36032 17184
rect 32766 17076 32772 17128
rect 32824 17116 32830 17128
rect 34716 17116 34744 17156
rect 37274 17144 37280 17196
rect 37332 17184 37338 17196
rect 41386 17184 41414 17224
rect 47394 17212 47400 17224
rect 47452 17212 47458 17264
rect 37332 17156 41414 17184
rect 37332 17144 37338 17156
rect 32824 17088 34744 17116
rect 32824 17076 32830 17088
rect 34790 17076 34796 17128
rect 34848 17116 34854 17128
rect 35253 17119 35311 17125
rect 35253 17116 35265 17119
rect 34848 17088 35265 17116
rect 34848 17076 34854 17088
rect 35253 17085 35265 17088
rect 35299 17085 35311 17119
rect 35253 17079 35311 17085
rect 35986 17076 35992 17128
rect 36044 17116 36050 17128
rect 39206 17116 39212 17128
rect 36044 17088 39212 17116
rect 36044 17076 36050 17088
rect 39206 17076 39212 17088
rect 39264 17076 39270 17128
rect 38930 17048 38936 17060
rect 32692 17020 38936 17048
rect 38930 17008 38936 17020
rect 38988 17008 38994 17060
rect 24044 16952 30512 16980
rect 30558 16940 30564 16992
rect 30616 16980 30622 16992
rect 31021 16983 31079 16989
rect 31021 16980 31033 16983
rect 30616 16952 31033 16980
rect 30616 16940 30622 16952
rect 31021 16949 31033 16952
rect 31067 16949 31079 16983
rect 31021 16943 31079 16949
rect 32398 16940 32404 16992
rect 32456 16980 32462 16992
rect 32953 16983 33011 16989
rect 32953 16980 32965 16983
rect 32456 16952 32965 16980
rect 32456 16940 32462 16952
rect 32953 16949 32965 16952
rect 32999 16949 33011 16983
rect 32953 16943 33011 16949
rect 34698 16940 34704 16992
rect 34756 16940 34762 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 6089 16779 6147 16785
rect 6089 16776 6101 16779
rect 1780 16748 6101 16776
rect 1780 16581 1808 16748
rect 6089 16745 6101 16748
rect 6135 16745 6147 16779
rect 9217 16779 9275 16785
rect 6089 16739 6147 16745
rect 8036 16748 8708 16776
rect 3418 16668 3424 16720
rect 3476 16668 3482 16720
rect 3602 16668 3608 16720
rect 3660 16708 3666 16720
rect 8036 16708 8064 16748
rect 3660 16680 8064 16708
rect 3660 16668 3666 16680
rect 8110 16668 8116 16720
rect 8168 16708 8174 16720
rect 8570 16708 8576 16720
rect 8168 16680 8576 16708
rect 8168 16668 8174 16680
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 2406 16600 2412 16652
rect 2464 16640 2470 16652
rect 3513 16643 3571 16649
rect 3513 16640 3525 16643
rect 2464 16612 3525 16640
rect 2464 16600 2470 16612
rect 3513 16609 3525 16612
rect 3559 16609 3571 16643
rect 3513 16603 3571 16609
rect 3786 16600 3792 16652
rect 3844 16640 3850 16652
rect 3844 16612 7144 16640
rect 3844 16600 3850 16612
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16541 1823 16575
rect 1765 16535 1823 16541
rect 4157 16575 4215 16581
rect 4157 16541 4169 16575
rect 4203 16541 4215 16575
rect 4157 16535 4215 16541
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 2501 16507 2559 16513
rect 2501 16504 2513 16507
rect 1360 16476 2513 16504
rect 1360 16464 1366 16476
rect 2501 16473 2513 16476
rect 2547 16473 2559 16507
rect 4172 16504 4200 16535
rect 4982 16532 4988 16584
rect 5040 16532 5046 16584
rect 7116 16581 7144 16612
rect 7190 16600 7196 16652
rect 7248 16600 7254 16652
rect 8481 16643 8539 16649
rect 7300 16612 8156 16640
rect 7101 16575 7159 16581
rect 7101 16541 7113 16575
rect 7147 16572 7159 16575
rect 7300 16572 7328 16612
rect 7147 16544 7328 16572
rect 8128 16572 8156 16612
rect 8481 16609 8493 16643
rect 8527 16640 8539 16643
rect 8680 16640 8708 16748
rect 9217 16745 9229 16779
rect 9263 16776 9275 16779
rect 9398 16776 9404 16788
rect 9263 16748 9404 16776
rect 9263 16745 9275 16748
rect 9217 16739 9275 16745
rect 9398 16736 9404 16748
rect 9456 16736 9462 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 13354 16776 13360 16788
rect 11112 16748 13360 16776
rect 11112 16736 11118 16748
rect 13354 16736 13360 16748
rect 13412 16736 13418 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 14792 16748 15393 16776
rect 14792 16736 14798 16748
rect 15381 16745 15393 16748
rect 15427 16776 15439 16779
rect 15562 16776 15568 16788
rect 15427 16748 15568 16776
rect 15427 16745 15439 16748
rect 15381 16739 15439 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15749 16779 15807 16785
rect 15749 16745 15761 16779
rect 15795 16776 15807 16779
rect 15838 16776 15844 16788
rect 15795 16748 15844 16776
rect 15795 16745 15807 16748
rect 15749 16739 15807 16745
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 16669 16779 16727 16785
rect 16669 16745 16681 16779
rect 16715 16776 16727 16779
rect 19686 16779 19744 16785
rect 19686 16776 19698 16779
rect 16715 16748 19698 16776
rect 16715 16745 16727 16748
rect 16669 16739 16727 16745
rect 19686 16745 19698 16748
rect 19732 16745 19744 16779
rect 19686 16739 19744 16745
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20128 16748 22232 16776
rect 20128 16736 20134 16748
rect 9306 16668 9312 16720
rect 9364 16708 9370 16720
rect 16850 16708 16856 16720
rect 9364 16680 11744 16708
rect 9364 16668 9370 16680
rect 8527 16612 8708 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 8496 16572 8524 16603
rect 8754 16600 8760 16652
rect 8812 16640 8818 16652
rect 9677 16643 9735 16649
rect 9677 16640 9689 16643
rect 8812 16612 9689 16640
rect 8812 16600 8818 16612
rect 9677 16609 9689 16612
rect 9723 16609 9735 16643
rect 9677 16603 9735 16609
rect 9861 16643 9919 16649
rect 9861 16609 9873 16643
rect 9907 16640 9919 16643
rect 9950 16640 9956 16652
rect 9907 16612 9956 16640
rect 9907 16609 9919 16612
rect 9861 16603 9919 16609
rect 9950 16600 9956 16612
rect 10008 16600 10014 16652
rect 10318 16600 10324 16652
rect 10376 16640 10382 16652
rect 10870 16640 10876 16652
rect 10376 16612 10876 16640
rect 10376 16600 10382 16612
rect 10870 16600 10876 16612
rect 10928 16600 10934 16652
rect 11054 16600 11060 16652
rect 11112 16600 11118 16652
rect 11716 16640 11744 16680
rect 11900 16680 16856 16708
rect 11900 16640 11928 16680
rect 16850 16668 16856 16680
rect 16908 16668 16914 16720
rect 17126 16668 17132 16720
rect 17184 16668 17190 16720
rect 19242 16708 19248 16720
rect 17604 16680 19248 16708
rect 11716 16612 11928 16640
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12986 16640 12992 16652
rect 12483 16612 12992 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 12986 16600 12992 16612
rect 13044 16640 13050 16652
rect 13044 16612 13584 16640
rect 13044 16600 13050 16612
rect 9490 16572 9496 16584
rect 8128 16544 8340 16572
rect 8496 16544 9496 16572
rect 7147 16541 7159 16544
rect 7101 16535 7159 16541
rect 5810 16504 5816 16516
rect 4172 16476 5816 16504
rect 2501 16467 2559 16473
rect 5810 16464 5816 16476
rect 5868 16464 5874 16516
rect 5997 16507 6055 16513
rect 5997 16473 6009 16507
rect 6043 16504 6055 16507
rect 6454 16504 6460 16516
rect 6043 16476 6460 16504
rect 6043 16473 6055 16476
rect 5997 16467 6055 16473
rect 6454 16464 6460 16476
rect 6512 16464 6518 16516
rect 7009 16507 7067 16513
rect 7009 16504 7021 16507
rect 6564 16476 7021 16504
rect 4614 16396 4620 16448
rect 4672 16436 4678 16448
rect 5258 16436 5264 16448
rect 4672 16408 5264 16436
rect 4672 16396 4678 16408
rect 5258 16396 5264 16408
rect 5316 16396 5322 16448
rect 6086 16396 6092 16448
rect 6144 16436 6150 16448
rect 6564 16436 6592 16476
rect 7009 16473 7021 16476
rect 7055 16473 7067 16507
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7009 16467 7067 16473
rect 7576 16476 8217 16504
rect 6144 16408 6592 16436
rect 6641 16439 6699 16445
rect 6144 16396 6150 16408
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 6914 16436 6920 16448
rect 6687 16408 6920 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 6914 16396 6920 16408
rect 6972 16396 6978 16448
rect 7282 16396 7288 16448
rect 7340 16436 7346 16448
rect 7576 16436 7604 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 8312 16504 8340 16544
rect 9490 16532 9496 16544
rect 9548 16532 9554 16584
rect 9582 16532 9588 16584
rect 9640 16572 9646 16584
rect 11517 16575 11575 16581
rect 11517 16572 11529 16575
rect 9640 16544 11529 16572
rect 9640 16532 9646 16544
rect 11517 16541 11529 16544
rect 11563 16572 11575 16575
rect 12253 16575 12311 16581
rect 12253 16572 12265 16575
rect 11563 16544 12265 16572
rect 11563 16541 11575 16544
rect 11517 16535 11575 16541
rect 12253 16541 12265 16544
rect 12299 16572 12311 16575
rect 13262 16572 13268 16584
rect 12299 16544 13268 16572
rect 12299 16541 12311 16544
rect 12253 16535 12311 16541
rect 13262 16532 13268 16544
rect 13320 16532 13326 16584
rect 13354 16532 13360 16584
rect 13412 16532 13418 16584
rect 13556 16572 13584 16612
rect 13630 16600 13636 16652
rect 13688 16600 13694 16652
rect 13814 16600 13820 16652
rect 13872 16640 13878 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 13872 16612 14841 16640
rect 13872 16600 13878 16612
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 15010 16600 15016 16652
rect 15068 16640 15074 16652
rect 16390 16640 16396 16652
rect 15068 16612 16396 16640
rect 15068 16600 15074 16612
rect 16390 16600 16396 16612
rect 16448 16600 16454 16652
rect 17604 16649 17632 16680
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 20714 16668 20720 16720
rect 20772 16708 20778 16720
rect 21450 16708 21456 16720
rect 20772 16680 21456 16708
rect 20772 16668 20778 16680
rect 21450 16668 21456 16680
rect 21508 16708 21514 16720
rect 21821 16711 21879 16717
rect 21821 16708 21833 16711
rect 21508 16680 21833 16708
rect 21508 16668 21514 16680
rect 21821 16677 21833 16680
rect 21867 16677 21879 16711
rect 21821 16671 21879 16677
rect 17589 16643 17647 16649
rect 17589 16609 17601 16643
rect 17635 16609 17647 16643
rect 17589 16603 17647 16609
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16640 17831 16643
rect 18874 16640 18880 16652
rect 17819 16612 18880 16640
rect 17819 16609 17831 16612
rect 17773 16603 17831 16609
rect 18874 16600 18880 16612
rect 18932 16600 18938 16652
rect 18966 16600 18972 16652
rect 19024 16600 19030 16652
rect 19429 16643 19487 16649
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19702 16640 19708 16652
rect 19475 16612 19708 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20990 16640 20996 16652
rect 20824 16612 20996 16640
rect 14274 16572 14280 16584
rect 13556 16544 14280 16572
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 15565 16575 15623 16581
rect 15565 16541 15577 16575
rect 15611 16572 15623 16575
rect 15930 16572 15936 16584
rect 15611 16544 15936 16572
rect 15611 16541 15623 16544
rect 15565 16535 15623 16541
rect 15930 16532 15936 16544
rect 15988 16532 15994 16584
rect 16025 16575 16083 16581
rect 16025 16541 16037 16575
rect 16071 16572 16083 16575
rect 16114 16572 16120 16584
rect 16071 16544 16120 16572
rect 16071 16541 16083 16544
rect 16025 16535 16083 16541
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 16298 16532 16304 16584
rect 16356 16572 16362 16584
rect 17862 16572 17868 16584
rect 16356 16544 17868 16572
rect 16356 16532 16362 16544
rect 17862 16532 17868 16544
rect 17920 16532 17926 16584
rect 18417 16575 18475 16581
rect 18417 16541 18429 16575
rect 18463 16572 18475 16575
rect 18984 16572 19012 16600
rect 18463 16544 19012 16572
rect 18463 16541 18475 16544
rect 18417 16535 18475 16541
rect 9030 16504 9036 16516
rect 8312 16476 9036 16504
rect 8205 16467 8263 16473
rect 9030 16464 9036 16476
rect 9088 16504 9094 16516
rect 10870 16504 10876 16516
rect 9088 16476 10876 16504
rect 9088 16464 9094 16476
rect 10870 16464 10876 16476
rect 10928 16464 10934 16516
rect 13906 16504 13912 16516
rect 13004 16476 13912 16504
rect 7340 16408 7604 16436
rect 7340 16396 7346 16408
rect 7834 16396 7840 16448
rect 7892 16396 7898 16448
rect 8294 16396 8300 16448
rect 8352 16396 8358 16448
rect 8754 16396 8760 16448
rect 8812 16436 8818 16448
rect 9585 16439 9643 16445
rect 9585 16436 9597 16439
rect 8812 16408 9597 16436
rect 8812 16396 8818 16408
rect 9585 16405 9597 16408
rect 9631 16405 9643 16439
rect 9585 16399 9643 16405
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 10413 16439 10471 16445
rect 10413 16436 10425 16439
rect 9732 16408 10425 16436
rect 9732 16396 9738 16408
rect 10413 16405 10425 16408
rect 10459 16405 10471 16439
rect 10413 16399 10471 16405
rect 10502 16396 10508 16448
rect 10560 16436 10566 16448
rect 10781 16439 10839 16445
rect 10781 16436 10793 16439
rect 10560 16408 10793 16436
rect 10560 16396 10566 16408
rect 10781 16405 10793 16408
rect 10827 16405 10839 16439
rect 10781 16399 10839 16405
rect 11790 16396 11796 16448
rect 11848 16396 11854 16448
rect 11974 16396 11980 16448
rect 12032 16436 12038 16448
rect 13004 16445 13032 16476
rect 13906 16464 13912 16476
rect 13964 16464 13970 16516
rect 14645 16507 14703 16513
rect 14645 16504 14657 16507
rect 14108 16476 14657 16504
rect 14108 16448 14136 16476
rect 14645 16473 14657 16476
rect 14691 16473 14703 16507
rect 14645 16467 14703 16473
rect 14734 16464 14740 16516
rect 14792 16464 14798 16516
rect 14918 16464 14924 16516
rect 14976 16504 14982 16516
rect 17497 16507 17555 16513
rect 17497 16504 17509 16507
rect 14976 16476 17509 16504
rect 14976 16464 14982 16476
rect 17497 16473 17509 16476
rect 17543 16473 17555 16507
rect 17497 16467 17555 16473
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 17736 16476 20116 16504
rect 17736 16464 17742 16476
rect 12161 16439 12219 16445
rect 12161 16436 12173 16439
rect 12032 16408 12173 16436
rect 12032 16396 12038 16408
rect 12161 16405 12173 16408
rect 12207 16405 12219 16439
rect 12161 16399 12219 16405
rect 12989 16439 13047 16445
rect 12989 16405 13001 16439
rect 13035 16405 13047 16439
rect 12989 16399 13047 16405
rect 13449 16439 13507 16445
rect 13449 16405 13461 16439
rect 13495 16436 13507 16439
rect 13998 16436 14004 16448
rect 13495 16408 14004 16436
rect 13495 16405 13507 16408
rect 13449 16399 13507 16405
rect 13998 16396 14004 16408
rect 14056 16396 14062 16448
rect 14090 16396 14096 16448
rect 14148 16396 14154 16448
rect 14274 16396 14280 16448
rect 14332 16396 14338 16448
rect 15286 16396 15292 16448
rect 15344 16436 15350 16448
rect 18322 16436 18328 16448
rect 15344 16408 18328 16436
rect 15344 16396 15350 16408
rect 18322 16396 18328 16408
rect 18380 16396 18386 16448
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 18966 16396 18972 16448
rect 19024 16436 19030 16448
rect 19978 16436 19984 16448
rect 19024 16408 19984 16436
rect 19024 16396 19030 16408
rect 19978 16396 19984 16408
rect 20036 16396 20042 16448
rect 20088 16436 20116 16476
rect 20824 16436 20852 16612
rect 20990 16600 20996 16612
rect 21048 16640 21054 16652
rect 21048 16612 21680 16640
rect 21048 16600 21054 16612
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16572 21511 16575
rect 21542 16572 21548 16584
rect 21499 16544 21548 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 21542 16532 21548 16544
rect 21600 16532 21606 16584
rect 21652 16572 21680 16612
rect 21726 16600 21732 16652
rect 21784 16640 21790 16652
rect 22094 16640 22100 16652
rect 21784 16612 22100 16640
rect 21784 16600 21790 16612
rect 22094 16600 22100 16612
rect 22152 16600 22158 16652
rect 22204 16581 22232 16748
rect 22554 16736 22560 16788
rect 22612 16776 22618 16788
rect 23566 16776 23572 16788
rect 22612 16748 23572 16776
rect 22612 16736 22618 16748
rect 23566 16736 23572 16748
rect 23624 16736 23630 16788
rect 23658 16736 23664 16788
rect 23716 16776 23722 16788
rect 24118 16776 24124 16788
rect 23716 16748 24124 16776
rect 23716 16736 23722 16748
rect 24118 16736 24124 16748
rect 24176 16736 24182 16788
rect 25038 16736 25044 16788
rect 25096 16776 25102 16788
rect 27433 16779 27491 16785
rect 27433 16776 27445 16779
rect 25096 16748 27445 16776
rect 25096 16736 25102 16748
rect 27433 16745 27445 16748
rect 27479 16745 27491 16779
rect 27433 16739 27491 16745
rect 27614 16736 27620 16788
rect 27672 16776 27678 16788
rect 28902 16776 28908 16788
rect 27672 16748 28908 16776
rect 27672 16736 27678 16748
rect 28902 16736 28908 16748
rect 28960 16736 28966 16788
rect 29365 16779 29423 16785
rect 29365 16745 29377 16779
rect 29411 16776 29423 16779
rect 29454 16776 29460 16788
rect 29411 16748 29460 16776
rect 29411 16745 29423 16748
rect 29365 16739 29423 16745
rect 29454 16736 29460 16748
rect 29512 16736 29518 16788
rect 29638 16736 29644 16788
rect 29696 16736 29702 16788
rect 31294 16736 31300 16788
rect 31352 16776 31358 16788
rect 35158 16776 35164 16788
rect 31352 16748 35164 16776
rect 31352 16736 31358 16748
rect 35158 16736 35164 16748
rect 35216 16736 35222 16788
rect 24854 16708 24860 16720
rect 23768 16680 24860 16708
rect 22462 16600 22468 16652
rect 22520 16640 22526 16652
rect 23768 16649 23796 16680
rect 24854 16668 24860 16680
rect 24912 16668 24918 16720
rect 26602 16668 26608 16720
rect 26660 16708 26666 16720
rect 30466 16708 30472 16720
rect 26660 16680 30472 16708
rect 26660 16668 26666 16680
rect 30466 16668 30472 16680
rect 30524 16668 30530 16720
rect 37826 16708 37832 16720
rect 33244 16680 37832 16708
rect 23753 16643 23811 16649
rect 22520 16612 23428 16640
rect 22520 16600 22526 16612
rect 22189 16575 22247 16581
rect 21652 16544 21956 16572
rect 21560 16504 21588 16532
rect 21928 16516 21956 16544
rect 22189 16541 22201 16575
rect 22235 16541 22247 16575
rect 22189 16535 22247 16541
rect 22833 16575 22891 16581
rect 22833 16541 22845 16575
rect 22879 16572 22891 16575
rect 23290 16572 23296 16584
rect 22879 16544 23296 16572
rect 22879 16541 22891 16544
rect 22833 16535 22891 16541
rect 23290 16532 23296 16544
rect 23348 16532 23354 16584
rect 23400 16572 23428 16612
rect 23753 16609 23765 16643
rect 23799 16609 23811 16643
rect 23753 16603 23811 16609
rect 23934 16600 23940 16652
rect 23992 16600 23998 16652
rect 24489 16643 24547 16649
rect 24489 16640 24501 16643
rect 24044 16612 24501 16640
rect 23400 16544 23796 16572
rect 21560 16476 21864 16504
rect 20088 16408 20852 16436
rect 21836 16436 21864 16476
rect 21910 16464 21916 16516
rect 21968 16504 21974 16516
rect 22278 16504 22284 16516
rect 21968 16476 22284 16504
rect 21968 16464 21974 16476
rect 22278 16464 22284 16476
rect 22336 16464 22342 16516
rect 22738 16464 22744 16516
rect 22796 16504 22802 16516
rect 23661 16507 23719 16513
rect 23661 16504 23673 16507
rect 22796 16476 23673 16504
rect 22796 16464 22802 16476
rect 23661 16473 23673 16476
rect 23707 16473 23719 16507
rect 23768 16504 23796 16544
rect 23842 16532 23848 16584
rect 23900 16572 23906 16584
rect 24044 16572 24072 16612
rect 24489 16609 24501 16612
rect 24535 16640 24547 16643
rect 24535 16612 25176 16640
rect 24535 16609 24547 16612
rect 24489 16603 24547 16609
rect 25148 16584 25176 16612
rect 25314 16600 25320 16652
rect 25372 16600 25378 16652
rect 26510 16600 26516 16652
rect 26568 16600 26574 16652
rect 26786 16600 26792 16652
rect 26844 16640 26850 16652
rect 27430 16640 27436 16652
rect 26844 16612 27436 16640
rect 26844 16600 26850 16612
rect 27430 16600 27436 16612
rect 27488 16640 27494 16652
rect 27893 16643 27951 16649
rect 27893 16640 27905 16643
rect 27488 16612 27905 16640
rect 27488 16600 27494 16612
rect 27893 16609 27905 16612
rect 27939 16609 27951 16643
rect 27893 16603 27951 16609
rect 27982 16600 27988 16652
rect 28040 16640 28046 16652
rect 28077 16643 28135 16649
rect 28077 16640 28089 16643
rect 28040 16612 28089 16640
rect 28040 16600 28046 16612
rect 28077 16609 28089 16612
rect 28123 16640 28135 16643
rect 29178 16640 29184 16652
rect 28123 16612 29184 16640
rect 28123 16609 28135 16612
rect 28077 16603 28135 16609
rect 29178 16600 29184 16612
rect 29236 16600 29242 16652
rect 29638 16600 29644 16652
rect 29696 16640 29702 16652
rect 29696 16612 30236 16640
rect 29696 16600 29702 16612
rect 23900 16544 24072 16572
rect 23900 16532 23906 16544
rect 25130 16532 25136 16584
rect 25188 16532 25194 16584
rect 26329 16575 26387 16581
rect 26329 16541 26341 16575
rect 26375 16572 26387 16575
rect 27154 16572 27160 16584
rect 26375 16544 27160 16572
rect 26375 16541 26387 16544
rect 26329 16535 26387 16541
rect 27154 16532 27160 16544
rect 27212 16532 27218 16584
rect 27246 16532 27252 16584
rect 27304 16572 27310 16584
rect 27801 16575 27859 16581
rect 27801 16572 27813 16575
rect 27304 16544 27813 16572
rect 27304 16532 27310 16544
rect 27801 16541 27813 16544
rect 27847 16541 27859 16575
rect 27801 16535 27859 16541
rect 28350 16532 28356 16584
rect 28408 16572 28414 16584
rect 28813 16575 28871 16581
rect 28813 16572 28825 16575
rect 28408 16544 28825 16572
rect 28408 16532 28414 16544
rect 28813 16541 28825 16544
rect 28859 16541 28871 16575
rect 28813 16535 28871 16541
rect 28902 16532 28908 16584
rect 28960 16572 28966 16584
rect 29730 16572 29736 16584
rect 28960 16544 29736 16572
rect 28960 16532 28966 16544
rect 29730 16532 29736 16544
rect 29788 16532 29794 16584
rect 30208 16581 30236 16612
rect 30650 16600 30656 16652
rect 30708 16600 30714 16652
rect 30929 16643 30987 16649
rect 30929 16609 30941 16643
rect 30975 16640 30987 16643
rect 31386 16640 31392 16652
rect 30975 16612 31392 16640
rect 30975 16609 30987 16612
rect 30929 16603 30987 16609
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 32217 16643 32275 16649
rect 32217 16609 32229 16643
rect 32263 16640 32275 16643
rect 32306 16640 32312 16652
rect 32263 16612 32312 16640
rect 32263 16609 32275 16612
rect 32217 16603 32275 16609
rect 32306 16600 32312 16612
rect 32364 16600 32370 16652
rect 33244 16649 33272 16680
rect 37826 16668 37832 16680
rect 37884 16668 37890 16720
rect 33229 16643 33287 16649
rect 33229 16609 33241 16643
rect 33275 16609 33287 16643
rect 33229 16603 33287 16609
rect 33505 16643 33563 16649
rect 33505 16609 33517 16643
rect 33551 16640 33563 16643
rect 33870 16640 33876 16652
rect 33551 16612 33876 16640
rect 33551 16609 33563 16612
rect 33505 16603 33563 16609
rect 33870 16600 33876 16612
rect 33928 16600 33934 16652
rect 30193 16575 30251 16581
rect 30193 16541 30205 16575
rect 30239 16541 30251 16575
rect 30193 16535 30251 16541
rect 31941 16575 31999 16581
rect 31941 16541 31953 16575
rect 31987 16572 31999 16575
rect 32582 16572 32588 16584
rect 31987 16544 32588 16572
rect 31987 16541 31999 16544
rect 31941 16535 31999 16541
rect 32582 16532 32588 16544
rect 32640 16532 32646 16584
rect 33318 16532 33324 16584
rect 33376 16572 33382 16584
rect 34606 16572 34612 16584
rect 33376 16544 34612 16572
rect 33376 16532 33382 16544
rect 34606 16532 34612 16544
rect 34664 16532 34670 16584
rect 23768 16476 27752 16504
rect 23661 16467 23719 16473
rect 22462 16436 22468 16448
rect 21836 16408 22468 16436
rect 22462 16396 22468 16408
rect 22520 16396 22526 16448
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22888 16408 23305 16436
rect 22888 16396 22894 16408
rect 23293 16405 23305 16408
rect 23339 16405 23351 16439
rect 23293 16399 23351 16405
rect 24762 16396 24768 16448
rect 24820 16396 24826 16448
rect 25130 16396 25136 16448
rect 25188 16396 25194 16448
rect 25225 16439 25283 16445
rect 25225 16405 25237 16439
rect 25271 16436 25283 16439
rect 25406 16436 25412 16448
rect 25271 16408 25412 16436
rect 25271 16405 25283 16408
rect 25225 16399 25283 16405
rect 25406 16396 25412 16408
rect 25464 16396 25470 16448
rect 25498 16396 25504 16448
rect 25556 16436 25562 16448
rect 25682 16436 25688 16448
rect 25556 16408 25688 16436
rect 25556 16396 25562 16408
rect 25682 16396 25688 16408
rect 25740 16396 25746 16448
rect 25774 16396 25780 16448
rect 25832 16436 25838 16448
rect 25961 16439 26019 16445
rect 25961 16436 25973 16439
rect 25832 16408 25973 16436
rect 25832 16396 25838 16408
rect 25961 16405 25973 16408
rect 26007 16405 26019 16439
rect 25961 16399 26019 16405
rect 26421 16439 26479 16445
rect 26421 16405 26433 16439
rect 26467 16436 26479 16439
rect 26602 16436 26608 16448
rect 26467 16408 26608 16436
rect 26467 16405 26479 16408
rect 26421 16399 26479 16405
rect 26602 16396 26608 16408
rect 26660 16396 26666 16448
rect 27062 16396 27068 16448
rect 27120 16396 27126 16448
rect 27724 16436 27752 16476
rect 28718 16464 28724 16516
rect 28776 16504 28782 16516
rect 28776 16476 30052 16504
rect 28776 16464 28782 16476
rect 28442 16436 28448 16448
rect 27724 16408 28448 16436
rect 28442 16396 28448 16408
rect 28500 16396 28506 16448
rect 28629 16439 28687 16445
rect 28629 16405 28641 16439
rect 28675 16436 28687 16439
rect 28810 16436 28816 16448
rect 28675 16408 28816 16436
rect 28675 16405 28687 16408
rect 28629 16399 28687 16405
rect 28810 16396 28816 16408
rect 28868 16396 28874 16448
rect 29086 16396 29092 16448
rect 29144 16396 29150 16448
rect 30024 16445 30052 16476
rect 34974 16464 34980 16516
rect 35032 16504 35038 16516
rect 35437 16507 35495 16513
rect 35437 16504 35449 16507
rect 35032 16476 35449 16504
rect 35032 16464 35038 16476
rect 35437 16473 35449 16476
rect 35483 16473 35495 16507
rect 35437 16467 35495 16473
rect 30009 16439 30067 16445
rect 30009 16405 30021 16439
rect 30055 16405 30067 16439
rect 30009 16399 30067 16405
rect 30098 16396 30104 16448
rect 30156 16436 30162 16448
rect 33226 16436 33232 16448
rect 30156 16408 33232 16436
rect 30156 16396 30162 16408
rect 33226 16396 33232 16408
rect 33284 16396 33290 16448
rect 35066 16396 35072 16448
rect 35124 16396 35130 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 8662 16232 8668 16244
rect 5675 16204 8668 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 8662 16192 8668 16204
rect 8720 16192 8726 16244
rect 9030 16192 9036 16244
rect 9088 16232 9094 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 9088 16204 9137 16232
rect 9088 16192 9094 16204
rect 9125 16201 9137 16204
rect 9171 16201 9183 16235
rect 9125 16195 9183 16201
rect 9214 16192 9220 16244
rect 9272 16192 9278 16244
rect 9490 16232 9496 16244
rect 9416 16204 9496 16232
rect 4617 16167 4675 16173
rect 4617 16133 4629 16167
rect 4663 16164 4675 16167
rect 4706 16164 4712 16176
rect 4663 16136 4712 16164
rect 4663 16133 4675 16136
rect 4617 16127 4675 16133
rect 4706 16124 4712 16136
rect 4764 16124 4770 16176
rect 5721 16167 5779 16173
rect 5721 16133 5733 16167
rect 5767 16164 5779 16167
rect 9416 16164 9444 16204
rect 9490 16192 9496 16204
rect 9548 16232 9554 16244
rect 10413 16235 10471 16241
rect 9548 16204 9628 16232
rect 9548 16192 9554 16204
rect 5767 16136 9076 16164
rect 5767 16133 5779 16136
rect 5721 16127 5779 16133
rect 1762 16056 1768 16108
rect 1820 16056 1826 16108
rect 3605 16099 3663 16105
rect 3605 16065 3617 16099
rect 3651 16096 3663 16099
rect 6546 16096 6552 16108
rect 3651 16068 6552 16096
rect 3651 16065 3663 16068
rect 3605 16059 3663 16065
rect 6546 16056 6552 16068
rect 6604 16056 6610 16108
rect 6638 16056 6644 16108
rect 6696 16096 6702 16108
rect 6917 16099 6975 16105
rect 6917 16096 6929 16099
rect 6696 16068 6929 16096
rect 6696 16056 6702 16068
rect 6917 16065 6929 16068
rect 6963 16065 6975 16099
rect 6917 16059 6975 16065
rect 7926 16056 7932 16108
rect 7984 16056 7990 16108
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 4706 15988 4712 16040
rect 4764 16028 4770 16040
rect 5813 16031 5871 16037
rect 5813 16028 5825 16031
rect 4764 16000 5825 16028
rect 4764 15988 4770 16000
rect 5813 15997 5825 16000
rect 5859 15997 5871 16031
rect 5813 15991 5871 15997
rect 7650 15988 7656 16040
rect 7708 16028 7714 16040
rect 8021 16031 8079 16037
rect 8021 16028 8033 16031
rect 7708 16000 8033 16028
rect 7708 15988 7714 16000
rect 8021 15997 8033 16000
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 1854 15920 1860 15972
rect 1912 15960 1918 15972
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 1912 15932 7113 15960
rect 1912 15920 1918 15932
rect 7101 15929 7113 15932
rect 7147 15929 7159 15963
rect 7101 15923 7159 15929
rect 7558 15920 7564 15972
rect 7616 15920 7622 15972
rect 7742 15920 7748 15972
rect 7800 15960 7806 15972
rect 8128 15960 8156 15991
rect 9048 15960 9076 16136
rect 9324 16136 9444 16164
rect 9600 16164 9628 16204
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10962 16232 10968 16244
rect 10459 16204 10968 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10962 16192 10968 16204
rect 11020 16192 11026 16244
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16232 11391 16235
rect 11422 16232 11428 16244
rect 11379 16204 11428 16232
rect 11379 16201 11391 16204
rect 11333 16195 11391 16201
rect 11422 16192 11428 16204
rect 11480 16192 11486 16244
rect 11701 16235 11759 16241
rect 11701 16201 11713 16235
rect 11747 16232 11759 16235
rect 12986 16232 12992 16244
rect 11747 16204 12992 16232
rect 11747 16201 11759 16204
rect 11701 16195 11759 16201
rect 12986 16192 12992 16204
rect 13044 16192 13050 16244
rect 14366 16192 14372 16244
rect 14424 16232 14430 16244
rect 14642 16232 14648 16244
rect 14424 16204 14648 16232
rect 14424 16192 14430 16204
rect 14642 16192 14648 16204
rect 14700 16192 14706 16244
rect 18966 16232 18972 16244
rect 15672 16204 18972 16232
rect 10594 16164 10600 16176
rect 9600 16136 10600 16164
rect 9324 16037 9352 16136
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11974 16164 11980 16176
rect 11112 16136 11980 16164
rect 11112 16124 11118 16136
rect 11974 16124 11980 16136
rect 12032 16124 12038 16176
rect 12437 16167 12495 16173
rect 12437 16164 12449 16167
rect 12084 16136 12449 16164
rect 12084 16108 12112 16136
rect 12437 16133 12449 16136
rect 12483 16133 12495 16167
rect 12437 16127 12495 16133
rect 12894 16124 12900 16176
rect 12952 16164 12958 16176
rect 14274 16164 14280 16176
rect 12952 16136 14280 16164
rect 12952 16124 12958 16136
rect 14274 16124 14280 16136
rect 14332 16124 14338 16176
rect 12066 16056 12072 16108
rect 12124 16056 12130 16108
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16065 12403 16099
rect 12345 16059 12403 16065
rect 9309 16031 9367 16037
rect 9309 15997 9321 16031
rect 9355 15997 9367 16031
rect 9309 15991 9367 15997
rect 9582 15988 9588 16040
rect 9640 16028 9646 16040
rect 10505 16031 10563 16037
rect 10505 16028 10517 16031
rect 9640 16000 10517 16028
rect 9640 15988 9646 16000
rect 10505 15997 10517 16000
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 10594 15988 10600 16040
rect 10652 15988 10658 16040
rect 11422 15988 11428 16040
rect 11480 16028 11486 16040
rect 11793 16031 11851 16037
rect 11793 16028 11805 16031
rect 11480 16000 11805 16028
rect 11480 15988 11486 16000
rect 11793 15997 11805 16000
rect 11839 16028 11851 16031
rect 12360 16028 12388 16059
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14292 16068 14841 16096
rect 11839 16000 12388 16028
rect 12621 16031 12679 16037
rect 11839 15997 11851 16000
rect 11793 15991 11851 15997
rect 12621 15997 12633 16031
rect 12667 16028 12679 16031
rect 13906 16028 13912 16040
rect 12667 16000 13912 16028
rect 12667 15997 12679 16000
rect 12621 15991 12679 15997
rect 13906 15988 13912 16000
rect 13964 15988 13970 16040
rect 9674 15960 9680 15972
rect 7800 15932 8156 15960
rect 8266 15932 8892 15960
rect 9048 15932 9680 15960
rect 7800 15920 7806 15932
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5261 15895 5319 15901
rect 5261 15892 5273 15895
rect 5040 15864 5273 15892
rect 5040 15852 5046 15864
rect 5261 15861 5273 15864
rect 5307 15861 5319 15895
rect 5261 15855 5319 15861
rect 6549 15895 6607 15901
rect 6549 15861 6561 15895
rect 6595 15892 6607 15895
rect 8266 15892 8294 15932
rect 6595 15864 8294 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 8754 15852 8760 15904
rect 8812 15852 8818 15904
rect 8864 15892 8892 15932
rect 9674 15920 9680 15932
rect 9732 15920 9738 15972
rect 11977 15963 12035 15969
rect 11977 15960 11989 15963
rect 11808 15932 11989 15960
rect 11808 15904 11836 15932
rect 11977 15929 11989 15932
rect 12023 15929 12035 15963
rect 11977 15923 12035 15929
rect 14292 15904 14320 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 14921 16099 14979 16105
rect 14921 16065 14933 16099
rect 14967 16096 14979 16099
rect 15194 16096 15200 16108
rect 14967 16068 15200 16096
rect 14967 16065 14979 16068
rect 14921 16059 14979 16065
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 15672 16105 15700 16204
rect 18966 16192 18972 16204
rect 19024 16192 19030 16244
rect 19337 16235 19395 16241
rect 19337 16201 19349 16235
rect 19383 16232 19395 16235
rect 19426 16232 19432 16244
rect 19383 16204 19432 16232
rect 19383 16201 19395 16204
rect 19337 16195 19395 16201
rect 19426 16192 19432 16204
rect 19484 16192 19490 16244
rect 19797 16235 19855 16241
rect 19797 16201 19809 16235
rect 19843 16232 19855 16235
rect 22005 16235 22063 16241
rect 22005 16232 22017 16235
rect 19843 16204 22017 16232
rect 19843 16201 19855 16204
rect 19797 16195 19855 16201
rect 22005 16201 22017 16204
rect 22051 16201 22063 16235
rect 22005 16195 22063 16201
rect 22373 16235 22431 16241
rect 22373 16201 22385 16235
rect 22419 16232 22431 16235
rect 23474 16232 23480 16244
rect 22419 16204 23480 16232
rect 22419 16201 22431 16204
rect 22373 16195 22431 16201
rect 23474 16192 23480 16204
rect 23532 16192 23538 16244
rect 23934 16232 23940 16244
rect 23768 16204 23940 16232
rect 17218 16164 17224 16176
rect 16868 16136 17224 16164
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16065 15715 16099
rect 15657 16059 15715 16065
rect 16868 16040 16896 16136
rect 17218 16124 17224 16136
rect 17276 16124 17282 16176
rect 17678 16124 17684 16176
rect 17736 16124 17742 16176
rect 20993 16167 21051 16173
rect 20993 16164 21005 16167
rect 19306 16136 21005 16164
rect 19306 16096 19334 16136
rect 20993 16133 21005 16136
rect 21039 16164 21051 16167
rect 22278 16164 22284 16176
rect 21039 16136 22284 16164
rect 21039 16133 21051 16136
rect 20993 16127 21051 16133
rect 22278 16124 22284 16136
rect 22336 16124 22342 16176
rect 22465 16167 22523 16173
rect 22465 16133 22477 16167
rect 22511 16164 22523 16167
rect 23382 16164 23388 16176
rect 22511 16136 23388 16164
rect 22511 16133 22523 16136
rect 22465 16127 22523 16133
rect 23382 16124 23388 16136
rect 23440 16124 23446 16176
rect 18340 16068 19334 16096
rect 15105 16031 15163 16037
rect 15105 15997 15117 16031
rect 15151 16028 15163 16031
rect 15930 16028 15936 16040
rect 15151 16000 15936 16028
rect 15151 15997 15163 16000
rect 15105 15991 15163 15997
rect 15930 15988 15936 16000
rect 15988 15988 15994 16040
rect 16850 15988 16856 16040
rect 16908 15988 16914 16040
rect 17126 15988 17132 16040
rect 17184 15988 17190 16040
rect 17494 15988 17500 16040
rect 17552 16028 17558 16040
rect 18340 16028 18368 16068
rect 19426 16056 19432 16108
rect 19484 16096 19490 16108
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 19484 16068 19717 16096
rect 19484 16056 19490 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 19705 16059 19763 16065
rect 20901 16099 20959 16105
rect 20901 16065 20913 16099
rect 20947 16096 20959 16099
rect 21450 16096 21456 16108
rect 20947 16068 21456 16096
rect 20947 16065 20959 16068
rect 20901 16059 20959 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 23106 16096 23112 16108
rect 22152 16068 23112 16096
rect 22152 16056 22158 16068
rect 23106 16056 23112 16068
rect 23164 16056 23170 16108
rect 23198 16056 23204 16108
rect 23256 16056 23262 16108
rect 23477 16099 23535 16105
rect 23477 16065 23489 16099
rect 23523 16096 23535 16099
rect 23566 16096 23572 16108
rect 23523 16068 23572 16096
rect 23523 16065 23535 16068
rect 23477 16059 23535 16065
rect 23566 16056 23572 16068
rect 23624 16056 23630 16108
rect 23768 16105 23796 16204
rect 23934 16192 23940 16204
rect 23992 16232 23998 16244
rect 26605 16235 26663 16241
rect 26605 16232 26617 16235
rect 23992 16204 26617 16232
rect 23992 16192 23998 16204
rect 26605 16201 26617 16204
rect 26651 16201 26663 16235
rect 26605 16195 26663 16201
rect 27154 16192 27160 16244
rect 27212 16232 27218 16244
rect 31202 16232 31208 16244
rect 27212 16204 31208 16232
rect 27212 16192 27218 16204
rect 31202 16192 31208 16204
rect 31260 16192 31266 16244
rect 31846 16192 31852 16244
rect 31904 16232 31910 16244
rect 32674 16232 32680 16244
rect 31904 16204 32680 16232
rect 31904 16192 31910 16204
rect 32674 16192 32680 16204
rect 32732 16192 32738 16244
rect 26694 16124 26700 16176
rect 26752 16164 26758 16176
rect 26752 16136 27384 16164
rect 26752 16124 26758 16136
rect 23753 16099 23811 16105
rect 23753 16065 23765 16099
rect 23799 16065 23811 16099
rect 23753 16059 23811 16065
rect 24670 16056 24676 16108
rect 24728 16096 24734 16108
rect 24857 16099 24915 16105
rect 24857 16096 24869 16099
rect 24728 16068 24869 16096
rect 24728 16056 24734 16068
rect 24857 16065 24869 16068
rect 24903 16065 24915 16099
rect 27062 16096 27068 16108
rect 26266 16068 27068 16096
rect 24857 16059 24915 16065
rect 27062 16056 27068 16068
rect 27120 16056 27126 16108
rect 27154 16056 27160 16108
rect 27212 16056 27218 16108
rect 27356 16096 27384 16136
rect 27522 16124 27528 16176
rect 27580 16164 27586 16176
rect 31113 16167 31171 16173
rect 31113 16164 31125 16167
rect 27580 16136 31125 16164
rect 27580 16124 27586 16136
rect 31113 16133 31125 16136
rect 31159 16133 31171 16167
rect 31113 16127 31171 16133
rect 31220 16136 33824 16164
rect 27356 16068 27936 16096
rect 17552 16000 18368 16028
rect 17552 15988 17558 16000
rect 18966 15988 18972 16040
rect 19024 16028 19030 16040
rect 19889 16031 19947 16037
rect 19889 16028 19901 16031
rect 19024 16000 19901 16028
rect 19024 15988 19030 16000
rect 19889 15997 19901 16000
rect 19935 16028 19947 16031
rect 20622 16028 20628 16040
rect 19935 16000 20628 16028
rect 19935 15997 19947 16000
rect 19889 15991 19947 15997
rect 20622 15988 20628 16000
rect 20680 15988 20686 16040
rect 21174 15988 21180 16040
rect 21232 15988 21238 16040
rect 22557 16031 22615 16037
rect 22557 16028 22569 16031
rect 21652 16000 22569 16028
rect 21652 15972 21680 16000
rect 22557 15997 22569 16000
rect 22603 15997 22615 16031
rect 22557 15991 22615 15997
rect 22738 15988 22744 16040
rect 22796 16028 22802 16040
rect 24762 16028 24768 16040
rect 22796 16000 24768 16028
rect 22796 15988 22802 16000
rect 24762 15988 24768 16000
rect 24820 15988 24826 16040
rect 25133 16031 25191 16037
rect 25133 15997 25145 16031
rect 25179 16028 25191 16031
rect 27801 16031 27859 16037
rect 27801 16028 27813 16031
rect 25179 16000 27813 16028
rect 25179 15997 25191 16000
rect 25133 15991 25191 15997
rect 27801 15997 27813 16000
rect 27847 15997 27859 16031
rect 27908 16028 27936 16068
rect 28258 16056 28264 16108
rect 28316 16056 28322 16108
rect 30098 16096 30104 16108
rect 28368 16068 30104 16096
rect 28368 16028 28396 16068
rect 30098 16056 30104 16068
rect 30156 16056 30162 16108
rect 30469 16099 30527 16105
rect 30469 16065 30481 16099
rect 30515 16096 30527 16099
rect 30558 16096 30564 16108
rect 30515 16068 30564 16096
rect 30515 16065 30527 16068
rect 30469 16059 30527 16065
rect 30558 16056 30564 16068
rect 30616 16056 30622 16108
rect 30926 16056 30932 16108
rect 30984 16096 30990 16108
rect 31220 16096 31248 16136
rect 30984 16068 31248 16096
rect 30984 16056 30990 16068
rect 31662 16056 31668 16108
rect 31720 16096 31726 16108
rect 31754 16096 31760 16108
rect 31720 16068 31760 16096
rect 31720 16056 31726 16068
rect 31754 16056 31760 16068
rect 31812 16056 31818 16108
rect 33796 16105 33824 16136
rect 32585 16099 32643 16105
rect 32585 16096 32597 16099
rect 31864 16068 32597 16096
rect 27908 16000 28396 16028
rect 29457 16031 29515 16037
rect 27801 15991 27859 15997
rect 29457 15997 29469 16031
rect 29503 15997 29515 16031
rect 29457 15991 29515 15997
rect 14458 15920 14464 15972
rect 14516 15920 14522 15972
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 15068 15932 16436 15960
rect 15068 15920 15074 15932
rect 9214 15892 9220 15904
rect 8864 15864 9220 15892
rect 9214 15852 9220 15864
rect 9272 15852 9278 15904
rect 10042 15852 10048 15904
rect 10100 15852 10106 15904
rect 11790 15852 11796 15904
rect 11848 15852 11854 15904
rect 12434 15852 12440 15904
rect 12492 15892 12498 15904
rect 13081 15895 13139 15901
rect 13081 15892 13093 15895
rect 12492 15864 13093 15892
rect 12492 15852 12498 15864
rect 13081 15861 13093 15864
rect 13127 15892 13139 15895
rect 13814 15892 13820 15904
rect 13127 15864 13820 15892
rect 13127 15861 13139 15864
rect 13081 15855 13139 15861
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14182 15892 14188 15904
rect 14047 15864 14188 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14182 15852 14188 15864
rect 14240 15852 14246 15904
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 16298 15852 16304 15904
rect 16356 15852 16362 15904
rect 16408 15892 16436 15932
rect 19058 15920 19064 15972
rect 19116 15920 19122 15972
rect 19242 15920 19248 15972
rect 19300 15960 19306 15972
rect 20533 15963 20591 15969
rect 20533 15960 20545 15963
rect 19300 15932 20545 15960
rect 19300 15920 19306 15932
rect 20533 15929 20545 15932
rect 20579 15929 20591 15963
rect 20533 15923 20591 15929
rect 21634 15920 21640 15972
rect 21692 15920 21698 15972
rect 22278 15920 22284 15972
rect 22336 15960 22342 15972
rect 22336 15932 22876 15960
rect 22336 15920 22342 15932
rect 18601 15895 18659 15901
rect 18601 15892 18613 15895
rect 16408 15864 18613 15892
rect 18601 15861 18613 15864
rect 18647 15892 18659 15895
rect 19978 15892 19984 15904
rect 18647 15864 19984 15892
rect 18647 15861 18659 15864
rect 18601 15855 18659 15861
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 20070 15852 20076 15904
rect 20128 15892 20134 15904
rect 22554 15892 22560 15904
rect 20128 15864 22560 15892
rect 20128 15852 20134 15864
rect 22554 15852 22560 15864
rect 22612 15852 22618 15904
rect 22848 15892 22876 15932
rect 24320 15932 24992 15960
rect 23014 15892 23020 15904
rect 22848 15864 23020 15892
rect 23014 15852 23020 15864
rect 23072 15852 23078 15904
rect 23106 15852 23112 15904
rect 23164 15892 23170 15904
rect 24320 15892 24348 15932
rect 23164 15864 24348 15892
rect 23164 15852 23170 15864
rect 24394 15852 24400 15904
rect 24452 15852 24458 15904
rect 24486 15852 24492 15904
rect 24544 15892 24550 15904
rect 24762 15892 24768 15904
rect 24544 15864 24768 15892
rect 24544 15852 24550 15864
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 24964 15892 24992 15932
rect 26142 15920 26148 15972
rect 26200 15960 26206 15972
rect 28905 15963 28963 15969
rect 28905 15960 28917 15963
rect 26200 15932 28917 15960
rect 26200 15920 26206 15932
rect 28905 15929 28917 15932
rect 28951 15929 28963 15963
rect 29472 15960 29500 15991
rect 31478 15988 31484 16040
rect 31536 16028 31542 16040
rect 31864 16028 31892 16068
rect 32585 16065 32597 16068
rect 32631 16065 32643 16099
rect 32585 16059 32643 16065
rect 33781 16099 33839 16105
rect 33781 16065 33793 16099
rect 33827 16096 33839 16099
rect 34057 16099 34115 16105
rect 34057 16096 34069 16099
rect 33827 16068 34069 16096
rect 33827 16065 33839 16068
rect 33781 16059 33839 16065
rect 34057 16065 34069 16068
rect 34103 16065 34115 16099
rect 34057 16059 34115 16065
rect 31536 16000 31892 16028
rect 32309 16031 32367 16037
rect 31536 15988 31542 16000
rect 32309 15997 32321 16031
rect 32355 16028 32367 16031
rect 36446 16028 36452 16040
rect 32355 16000 36452 16028
rect 32355 15997 32367 16000
rect 32309 15991 32367 15997
rect 36446 15988 36452 16000
rect 36504 15988 36510 16040
rect 32398 15960 32404 15972
rect 29472 15932 32404 15960
rect 28905 15923 28963 15929
rect 32398 15920 32404 15932
rect 32456 15920 32462 15972
rect 28994 15892 29000 15904
rect 24964 15864 29000 15892
rect 28994 15852 29000 15864
rect 29052 15852 29058 15904
rect 29546 15852 29552 15904
rect 29604 15892 29610 15904
rect 30009 15895 30067 15901
rect 30009 15892 30021 15895
rect 29604 15864 30021 15892
rect 29604 15852 29610 15864
rect 30009 15861 30021 15864
rect 30055 15861 30067 15895
rect 30009 15855 30067 15861
rect 31570 15852 31576 15904
rect 31628 15852 31634 15904
rect 31662 15852 31668 15904
rect 31720 15892 31726 15904
rect 33597 15895 33655 15901
rect 33597 15892 33609 15895
rect 31720 15864 33609 15892
rect 31720 15852 31726 15864
rect 33597 15861 33609 15864
rect 33643 15861 33655 15895
rect 33597 15855 33655 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 2866 15688 2872 15700
rect 1176 15660 2872 15688
rect 1176 15648 1182 15660
rect 2866 15648 2872 15660
rect 2924 15648 2930 15700
rect 6362 15648 6368 15700
rect 6420 15688 6426 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 6420 15660 7573 15688
rect 6420 15648 6426 15660
rect 7561 15657 7573 15660
rect 7607 15657 7619 15691
rect 14274 15688 14280 15700
rect 7561 15651 7619 15657
rect 7668 15660 14280 15688
rect 3602 15580 3608 15632
rect 3660 15580 3666 15632
rect 3988 15592 5120 15620
rect 1302 15512 1308 15564
rect 1360 15552 1366 15564
rect 2041 15555 2099 15561
rect 2041 15552 2053 15555
rect 1360 15524 2053 15552
rect 1360 15512 1366 15524
rect 2041 15521 2053 15524
rect 2087 15521 2099 15555
rect 2041 15515 2099 15521
rect 2314 15512 2320 15564
rect 2372 15552 2378 15564
rect 3988 15552 4016 15592
rect 2372 15524 4016 15552
rect 2372 15512 2378 15524
rect 4798 15512 4804 15564
rect 4856 15552 4862 15564
rect 4985 15555 5043 15561
rect 4985 15552 4997 15555
rect 4856 15524 4997 15552
rect 4856 15512 4862 15524
rect 4985 15521 4997 15524
rect 5031 15521 5043 15555
rect 5092 15552 5120 15592
rect 6270 15580 6276 15632
rect 6328 15620 6334 15632
rect 7668 15620 7696 15660
rect 14274 15648 14280 15660
rect 14332 15648 14338 15700
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 15010 15688 15016 15700
rect 14507 15660 15016 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 15010 15648 15016 15660
rect 15068 15648 15074 15700
rect 15746 15648 15752 15700
rect 15804 15688 15810 15700
rect 16485 15691 16543 15697
rect 16485 15688 16497 15691
rect 15804 15660 16497 15688
rect 15804 15648 15810 15660
rect 16485 15657 16497 15660
rect 16531 15657 16543 15691
rect 16485 15651 16543 15657
rect 16666 15648 16672 15700
rect 16724 15688 16730 15700
rect 18966 15688 18972 15700
rect 16724 15660 18972 15688
rect 16724 15648 16730 15660
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19334 15648 19340 15700
rect 19392 15688 19398 15700
rect 19521 15691 19579 15697
rect 19521 15688 19533 15691
rect 19392 15660 19533 15688
rect 19392 15648 19398 15660
rect 19521 15657 19533 15660
rect 19567 15657 19579 15691
rect 19521 15651 19579 15657
rect 19886 15648 19892 15700
rect 19944 15688 19950 15700
rect 19944 15660 24624 15688
rect 19944 15648 19950 15660
rect 9490 15620 9496 15632
rect 6328 15592 7696 15620
rect 8680 15592 9496 15620
rect 6328 15580 6334 15592
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5092 15524 5273 15552
rect 4985 15515 5043 15521
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 7650 15512 7656 15564
rect 7708 15552 7714 15564
rect 8021 15555 8079 15561
rect 8021 15552 8033 15555
rect 7708 15524 8033 15552
rect 7708 15512 7714 15524
rect 8021 15521 8033 15524
rect 8067 15521 8079 15555
rect 8021 15515 8079 15521
rect 8113 15555 8171 15561
rect 8113 15521 8125 15555
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15484 1823 15487
rect 1854 15484 1860 15496
rect 1811 15456 1860 15484
rect 1811 15453 1823 15456
rect 1765 15447 1823 15453
rect 1854 15444 1860 15456
rect 1912 15444 1918 15496
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 2746 15456 4353 15484
rect 934 15376 940 15428
rect 992 15416 998 15428
rect 2746 15416 2774 15456
rect 4341 15453 4353 15456
rect 4387 15484 4399 15487
rect 4890 15484 4896 15496
rect 4387 15456 4896 15484
rect 4387 15453 4399 15456
rect 4341 15447 4399 15453
rect 4890 15444 4896 15456
rect 4948 15444 4954 15496
rect 6730 15444 6736 15496
rect 6788 15484 6794 15496
rect 8128 15484 8156 15515
rect 8680 15493 8708 15592
rect 9490 15580 9496 15592
rect 9548 15620 9554 15632
rect 9548 15592 9812 15620
rect 9548 15580 9554 15592
rect 9398 15512 9404 15564
rect 9456 15552 9462 15564
rect 9677 15555 9735 15561
rect 9677 15552 9689 15555
rect 9456 15524 9689 15552
rect 9456 15512 9462 15524
rect 9677 15521 9689 15524
rect 9723 15521 9735 15555
rect 9784 15552 9812 15592
rect 9858 15580 9864 15632
rect 9916 15620 9922 15632
rect 9916 15592 11100 15620
rect 9916 15580 9922 15592
rect 10965 15555 11023 15561
rect 10965 15552 10977 15555
rect 9784 15524 10977 15552
rect 9677 15515 9735 15521
rect 10965 15521 10977 15524
rect 11011 15521 11023 15555
rect 11072 15552 11100 15592
rect 16390 15580 16396 15632
rect 16448 15620 16454 15632
rect 16448 15592 17080 15620
rect 16448 15580 16454 15592
rect 13998 15552 14004 15564
rect 11072 15524 14004 15552
rect 10965 15515 11023 15521
rect 13998 15512 14004 15524
rect 14056 15512 14062 15564
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 17052 15552 17080 15592
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 18380 15592 20300 15620
rect 18380 15580 18386 15592
rect 14783 15524 16988 15552
rect 17052 15524 18736 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 16960 15496 16988 15524
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 6788 15456 8677 15484
rect 6788 15444 6794 15456
rect 8665 15453 8677 15456
rect 8711 15453 8723 15487
rect 9306 15484 9312 15496
rect 8665 15447 8723 15453
rect 8864 15456 9312 15484
rect 992 15388 2774 15416
rect 992 15376 998 15388
rect 3418 15376 3424 15428
rect 3476 15376 3482 15428
rect 3602 15376 3608 15428
rect 3660 15416 3666 15428
rect 6546 15416 6552 15428
rect 3660 15388 4200 15416
rect 6486 15388 6552 15416
rect 3660 15376 3666 15388
rect 2406 15308 2412 15360
rect 2464 15348 2470 15360
rect 3436 15348 3464 15376
rect 2464 15320 3464 15348
rect 3973 15351 4031 15357
rect 2464 15308 2470 15320
rect 3973 15317 3985 15351
rect 4019 15348 4031 15351
rect 4062 15348 4068 15360
rect 4019 15320 4068 15348
rect 4019 15317 4031 15320
rect 3973 15311 4031 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4172 15348 4200 15388
rect 6546 15376 6552 15388
rect 6604 15376 6610 15428
rect 6822 15376 6828 15428
rect 6880 15416 6886 15428
rect 7006 15416 7012 15428
rect 6880 15388 7012 15416
rect 6880 15376 6886 15388
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7926 15376 7932 15428
rect 7984 15376 7990 15428
rect 4433 15351 4491 15357
rect 4433 15348 4445 15351
rect 4172 15320 4445 15348
rect 4433 15317 4445 15320
rect 4479 15317 4491 15351
rect 4433 15311 4491 15317
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 6564 15348 6592 15376
rect 6236 15320 6592 15348
rect 6236 15308 6242 15320
rect 7190 15308 7196 15360
rect 7248 15348 7254 15360
rect 8864 15348 8892 15456
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15484 9551 15487
rect 11330 15484 11336 15496
rect 9539 15456 11336 15484
rect 9539 15453 9551 15456
rect 9493 15447 9551 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11609 15487 11667 15493
rect 11609 15453 11621 15487
rect 11655 15453 11667 15487
rect 11609 15447 11667 15453
rect 9030 15376 9036 15428
rect 9088 15416 9094 15428
rect 10873 15419 10931 15425
rect 10873 15416 10885 15419
rect 9088 15388 10885 15416
rect 9088 15376 9094 15388
rect 10873 15385 10885 15388
rect 10919 15385 10931 15419
rect 11624 15416 11652 15447
rect 13262 15444 13268 15496
rect 13320 15484 13326 15496
rect 13909 15487 13967 15493
rect 13909 15484 13921 15487
rect 13320 15456 13921 15484
rect 13320 15444 13326 15456
rect 13909 15453 13921 15456
rect 13955 15484 13967 15487
rect 14642 15484 14648 15496
rect 13955 15456 14648 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 16942 15444 16948 15496
rect 17000 15444 17006 15496
rect 18708 15484 18736 15524
rect 18782 15512 18788 15564
rect 18840 15552 18846 15564
rect 19061 15555 19119 15561
rect 19061 15552 19073 15555
rect 18840 15524 19073 15552
rect 18840 15512 18846 15524
rect 19061 15521 19073 15524
rect 19107 15552 19119 15555
rect 20070 15552 20076 15564
rect 19107 15524 20076 15552
rect 19107 15521 19119 15524
rect 19061 15515 19119 15521
rect 20070 15512 20076 15524
rect 20128 15512 20134 15564
rect 20162 15512 20168 15564
rect 20220 15512 20226 15564
rect 20272 15552 20300 15592
rect 20530 15580 20536 15632
rect 20588 15580 20594 15632
rect 20898 15552 20904 15564
rect 20272 15524 20904 15552
rect 20898 15512 20904 15524
rect 20956 15512 20962 15564
rect 22002 15552 22008 15564
rect 21008 15524 22008 15552
rect 19242 15484 19248 15496
rect 18708 15456 19248 15484
rect 19242 15444 19248 15456
rect 19300 15444 19306 15496
rect 19702 15444 19708 15496
rect 19760 15484 19766 15496
rect 21008 15493 21036 15524
rect 22002 15512 22008 15524
rect 22060 15552 22066 15564
rect 22278 15552 22284 15564
rect 22060 15524 22284 15552
rect 22060 15512 22066 15524
rect 22278 15512 22284 15524
rect 22336 15512 22342 15564
rect 23934 15512 23940 15564
rect 23992 15512 23998 15564
rect 24596 15561 24624 15660
rect 25130 15648 25136 15700
rect 25188 15688 25194 15700
rect 25188 15660 27108 15688
rect 25188 15648 25194 15660
rect 24581 15555 24639 15561
rect 24581 15521 24593 15555
rect 24627 15521 24639 15555
rect 24581 15515 24639 15521
rect 24854 15512 24860 15564
rect 24912 15512 24918 15564
rect 25682 15512 25688 15564
rect 25740 15552 25746 15564
rect 25961 15555 26019 15561
rect 25961 15552 25973 15555
rect 25740 15524 25973 15552
rect 25740 15512 25746 15524
rect 25961 15521 25973 15524
rect 26007 15521 26019 15555
rect 25961 15515 26019 15521
rect 26602 15512 26608 15564
rect 26660 15552 26666 15564
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 26660 15524 26985 15552
rect 26660 15512 26666 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 27080 15552 27108 15660
rect 27798 15648 27804 15700
rect 27856 15648 27862 15700
rect 27982 15648 27988 15700
rect 28040 15648 28046 15700
rect 31662 15688 31668 15700
rect 28184 15660 31668 15688
rect 27338 15580 27344 15632
rect 27396 15620 27402 15632
rect 28184 15620 28212 15660
rect 31662 15648 31668 15660
rect 31720 15648 31726 15700
rect 31754 15648 31760 15700
rect 31812 15688 31818 15700
rect 32401 15691 32459 15697
rect 32401 15688 32413 15691
rect 31812 15660 32413 15688
rect 31812 15648 31818 15660
rect 32401 15657 32413 15660
rect 32447 15657 32459 15691
rect 32401 15651 32459 15657
rect 27396 15592 28212 15620
rect 27396 15580 27402 15592
rect 28258 15580 28264 15632
rect 28316 15620 28322 15632
rect 31846 15620 31852 15632
rect 28316 15592 31852 15620
rect 28316 15580 28322 15592
rect 31846 15580 31852 15592
rect 31904 15580 31910 15632
rect 31941 15623 31999 15629
rect 31941 15589 31953 15623
rect 31987 15620 31999 15623
rect 32214 15620 32220 15632
rect 31987 15592 32220 15620
rect 31987 15589 31999 15592
rect 31941 15583 31999 15589
rect 32214 15580 32220 15592
rect 32272 15580 32278 15632
rect 27525 15555 27583 15561
rect 27525 15552 27537 15555
rect 27080 15524 27537 15552
rect 26973 15515 27031 15521
rect 27525 15521 27537 15524
rect 27571 15552 27583 15555
rect 37274 15552 37280 15564
rect 27571 15524 37280 15552
rect 27571 15521 27583 15524
rect 27525 15515 27583 15521
rect 20993 15487 21051 15493
rect 20993 15484 21005 15487
rect 19760 15456 21005 15484
rect 19760 15444 19766 15456
rect 20993 15453 21005 15456
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 23198 15444 23204 15496
rect 23256 15484 23262 15496
rect 23256 15456 24532 15484
rect 23256 15444 23262 15456
rect 11624 15388 11744 15416
rect 10873 15379 10931 15385
rect 7248 15320 8892 15348
rect 7248 15308 7254 15320
rect 8938 15308 8944 15360
rect 8996 15348 9002 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8996 15320 9137 15348
rect 8996 15308 9002 15320
rect 9125 15317 9137 15320
rect 9171 15317 9183 15351
rect 9125 15311 9183 15317
rect 9582 15308 9588 15360
rect 9640 15308 9646 15360
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 10413 15351 10471 15357
rect 10413 15348 10425 15351
rect 9732 15320 10425 15348
rect 9732 15308 9738 15320
rect 10413 15317 10425 15320
rect 10459 15317 10471 15351
rect 10413 15311 10471 15317
rect 10686 15308 10692 15360
rect 10744 15348 10750 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10744 15320 10793 15348
rect 10744 15308 10750 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10888 15348 10916 15379
rect 11716 15360 11744 15388
rect 11882 15376 11888 15428
rect 11940 15376 11946 15428
rect 12618 15376 12624 15428
rect 12676 15376 12682 15428
rect 13170 15376 13176 15428
rect 13228 15416 13234 15428
rect 13725 15419 13783 15425
rect 13725 15416 13737 15419
rect 13228 15388 13737 15416
rect 13228 15376 13234 15388
rect 13725 15385 13737 15388
rect 13771 15416 13783 15419
rect 14550 15416 14556 15428
rect 13771 15388 14556 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 14550 15376 14556 15388
rect 14608 15376 14614 15428
rect 15013 15419 15071 15425
rect 15013 15385 15025 15419
rect 15059 15416 15071 15419
rect 15102 15416 15108 15428
rect 15059 15388 15108 15416
rect 15059 15385 15071 15388
rect 15013 15379 15071 15385
rect 15102 15376 15108 15388
rect 15160 15376 15166 15428
rect 15654 15376 15660 15428
rect 15712 15376 15718 15428
rect 16850 15376 16856 15428
rect 16908 15416 16914 15428
rect 17208 15419 17266 15425
rect 17208 15416 17220 15419
rect 16908 15388 17220 15416
rect 16908 15376 16914 15388
rect 17208 15385 17220 15388
rect 17254 15385 17266 15419
rect 17208 15379 17266 15385
rect 17678 15376 17684 15428
rect 17736 15376 17742 15428
rect 19981 15419 20039 15425
rect 19981 15385 19993 15419
rect 20027 15416 20039 15419
rect 20806 15416 20812 15428
rect 20027 15388 20812 15416
rect 20027 15385 20039 15388
rect 19981 15379 20039 15385
rect 20806 15376 20812 15388
rect 20864 15376 20870 15428
rect 21269 15419 21327 15425
rect 21269 15416 21281 15419
rect 21100 15388 21281 15416
rect 21100 15360 21128 15388
rect 21269 15385 21281 15388
rect 21315 15385 21327 15419
rect 21269 15379 21327 15385
rect 21910 15376 21916 15428
rect 21968 15376 21974 15428
rect 22554 15376 22560 15428
rect 22612 15416 22618 15428
rect 23661 15419 23719 15425
rect 23661 15416 23673 15419
rect 22612 15388 23673 15416
rect 22612 15376 22618 15388
rect 23661 15385 23673 15388
rect 23707 15416 23719 15419
rect 24210 15416 24216 15428
rect 23707 15388 24216 15416
rect 23707 15385 23719 15388
rect 23661 15379 23719 15385
rect 24210 15376 24216 15388
rect 24268 15376 24274 15428
rect 24504 15416 24532 15456
rect 25406 15444 25412 15496
rect 25464 15484 25470 15496
rect 25869 15487 25927 15493
rect 25869 15484 25881 15487
rect 25464 15456 25881 15484
rect 25464 15444 25470 15456
rect 25869 15453 25881 15456
rect 25915 15484 25927 15487
rect 26881 15487 26939 15493
rect 26881 15484 26893 15487
rect 25915 15456 26893 15484
rect 25915 15453 25927 15456
rect 25869 15447 25927 15453
rect 26881 15453 26893 15456
rect 26927 15484 26939 15487
rect 27706 15484 27712 15496
rect 26927 15456 27712 15484
rect 26927 15453 26939 15456
rect 26881 15447 26939 15453
rect 27706 15444 27712 15456
rect 27764 15444 27770 15496
rect 25424 15416 25452 15444
rect 27246 15416 27252 15428
rect 24504 15388 25452 15416
rect 25516 15388 27252 15416
rect 11146 15348 11152 15360
rect 10888 15320 11152 15348
rect 10781 15311 10839 15317
rect 11146 15308 11152 15320
rect 11204 15308 11210 15360
rect 11698 15308 11704 15360
rect 11756 15308 11762 15360
rect 12526 15308 12532 15360
rect 12584 15348 12590 15360
rect 13357 15351 13415 15357
rect 13357 15348 13369 15351
rect 12584 15320 13369 15348
rect 12584 15308 12590 15320
rect 13357 15317 13369 15320
rect 13403 15317 13415 15351
rect 13357 15311 13415 15317
rect 14090 15308 14096 15360
rect 14148 15308 14154 15360
rect 16758 15308 16764 15360
rect 16816 15348 16822 15360
rect 18506 15348 18512 15360
rect 16816 15320 18512 15348
rect 16816 15308 16822 15320
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 18690 15308 18696 15360
rect 18748 15308 18754 15360
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20438 15348 20444 15360
rect 19935 15320 20444 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20438 15308 20444 15320
rect 20496 15308 20502 15360
rect 21082 15308 21088 15360
rect 21140 15308 21146 15360
rect 21634 15308 21640 15360
rect 21692 15348 21698 15360
rect 22741 15351 22799 15357
rect 22741 15348 22753 15351
rect 21692 15320 22753 15348
rect 21692 15308 21698 15320
rect 22741 15317 22753 15320
rect 22787 15317 22799 15351
rect 22741 15311 22799 15317
rect 23293 15351 23351 15357
rect 23293 15317 23305 15351
rect 23339 15348 23351 15351
rect 23382 15348 23388 15360
rect 23339 15320 23388 15348
rect 23339 15317 23351 15320
rect 23293 15311 23351 15317
rect 23382 15308 23388 15320
rect 23440 15308 23446 15360
rect 23750 15308 23756 15360
rect 23808 15348 23814 15360
rect 24762 15348 24768 15360
rect 23808 15320 24768 15348
rect 23808 15308 23814 15320
rect 24762 15308 24768 15320
rect 24820 15348 24826 15360
rect 25516 15348 25544 15388
rect 27246 15376 27252 15388
rect 27304 15376 27310 15428
rect 24820 15320 25544 15348
rect 24820 15308 24826 15320
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 26421 15351 26479 15357
rect 26421 15348 26433 15351
rect 26384 15320 26433 15348
rect 26384 15308 26390 15320
rect 26421 15317 26433 15320
rect 26467 15317 26479 15351
rect 26421 15311 26479 15317
rect 26789 15351 26847 15357
rect 26789 15317 26801 15351
rect 26835 15348 26847 15351
rect 27816 15348 27844 15524
rect 37274 15512 37280 15524
rect 37332 15512 37338 15564
rect 27982 15444 27988 15496
rect 28040 15484 28046 15496
rect 28353 15487 28411 15493
rect 28353 15484 28365 15487
rect 28040 15456 28365 15484
rect 28040 15444 28046 15456
rect 28353 15453 28365 15456
rect 28399 15453 28411 15487
rect 28353 15447 28411 15453
rect 28626 15444 28632 15496
rect 28684 15444 28690 15496
rect 29638 15444 29644 15496
rect 29696 15484 29702 15496
rect 29733 15487 29791 15493
rect 29733 15484 29745 15487
rect 29696 15456 29745 15484
rect 29696 15444 29702 15456
rect 29733 15453 29745 15456
rect 29779 15453 29791 15487
rect 29733 15447 29791 15453
rect 29748 15416 29776 15447
rect 30006 15444 30012 15496
rect 30064 15444 30070 15496
rect 30098 15444 30104 15496
rect 30156 15484 30162 15496
rect 31481 15487 31539 15493
rect 30156 15456 31248 15484
rect 30156 15444 30162 15456
rect 30837 15419 30895 15425
rect 30837 15416 30849 15419
rect 29748 15388 30849 15416
rect 30837 15385 30849 15388
rect 30883 15385 30895 15419
rect 31110 15416 31116 15428
rect 30837 15379 30895 15385
rect 30944 15388 31116 15416
rect 26835 15320 27844 15348
rect 26835 15317 26847 15320
rect 26789 15311 26847 15317
rect 28718 15308 28724 15360
rect 28776 15348 28782 15360
rect 30944 15348 30972 15388
rect 31110 15376 31116 15388
rect 31168 15376 31174 15428
rect 31220 15416 31248 15456
rect 31481 15453 31493 15487
rect 31527 15484 31539 15487
rect 31662 15484 31668 15496
rect 31527 15456 31668 15484
rect 31527 15453 31539 15456
rect 31481 15447 31539 15453
rect 31662 15444 31668 15456
rect 31720 15444 31726 15496
rect 32030 15444 32036 15496
rect 32088 15484 32094 15496
rect 32125 15487 32183 15493
rect 32125 15484 32137 15487
rect 32088 15456 32137 15484
rect 32088 15444 32094 15456
rect 32125 15453 32137 15456
rect 32171 15484 32183 15487
rect 32769 15487 32827 15493
rect 32769 15484 32781 15487
rect 32171 15456 32781 15484
rect 32171 15453 32183 15456
rect 32125 15447 32183 15453
rect 32769 15453 32781 15456
rect 32815 15453 32827 15487
rect 32769 15447 32827 15453
rect 33870 15444 33876 15496
rect 33928 15484 33934 15496
rect 38746 15484 38752 15496
rect 33928 15456 38752 15484
rect 33928 15444 33934 15456
rect 38746 15444 38752 15456
rect 38804 15444 38810 15496
rect 41230 15416 41236 15428
rect 31220 15388 41236 15416
rect 41230 15376 41236 15388
rect 41288 15376 41294 15428
rect 28776 15320 30972 15348
rect 28776 15308 28782 15320
rect 31018 15308 31024 15360
rect 31076 15348 31082 15360
rect 31297 15351 31355 15357
rect 31297 15348 31309 15351
rect 31076 15320 31309 15348
rect 31076 15308 31082 15320
rect 31297 15317 31309 15320
rect 31343 15317 31355 15351
rect 31297 15311 31355 15317
rect 32214 15308 32220 15360
rect 32272 15348 32278 15360
rect 32490 15348 32496 15360
rect 32272 15320 32496 15348
rect 32272 15308 32278 15320
rect 32490 15308 32496 15320
rect 32548 15308 32554 15360
rect 32582 15308 32588 15360
rect 32640 15308 32646 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 4525 15147 4583 15153
rect 4525 15144 4537 15147
rect 4488 15116 4537 15144
rect 4488 15104 4494 15116
rect 4525 15113 4537 15116
rect 4571 15113 4583 15147
rect 4525 15107 4583 15113
rect 5718 15104 5724 15156
rect 5776 15104 5782 15156
rect 7650 15104 7656 15156
rect 7708 15144 7714 15156
rect 7926 15144 7932 15156
rect 7708 15116 7932 15144
rect 7708 15104 7714 15116
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8018 15104 8024 15156
rect 8076 15104 8082 15156
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9677 15147 9735 15153
rect 9677 15144 9689 15147
rect 8812 15116 9689 15144
rect 8812 15104 8818 15116
rect 9677 15113 9689 15116
rect 9723 15113 9735 15147
rect 9677 15107 9735 15113
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 11609 15147 11667 15153
rect 11609 15144 11621 15147
rect 10652 15116 11621 15144
rect 10652 15104 10658 15116
rect 11609 15113 11621 15116
rect 11655 15144 11667 15147
rect 11698 15144 11704 15156
rect 11655 15116 11704 15144
rect 11655 15113 11667 15116
rect 11609 15107 11667 15113
rect 11698 15104 11704 15116
rect 11756 15104 11762 15156
rect 12250 15104 12256 15156
rect 12308 15104 12314 15156
rect 12713 15147 12771 15153
rect 12713 15113 12725 15147
rect 12759 15144 12771 15147
rect 14090 15144 14096 15156
rect 12759 15116 14096 15144
rect 12759 15113 12771 15116
rect 12713 15107 12771 15113
rect 14090 15104 14096 15116
rect 14148 15104 14154 15156
rect 14182 15104 14188 15156
rect 14240 15104 14246 15156
rect 14369 15147 14427 15153
rect 14369 15113 14381 15147
rect 14415 15144 14427 15147
rect 14826 15144 14832 15156
rect 14415 15116 14832 15144
rect 14415 15113 14427 15116
rect 14369 15107 14427 15113
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15565 15147 15623 15153
rect 15565 15113 15577 15147
rect 15611 15144 15623 15147
rect 16022 15144 16028 15156
rect 15611 15116 16028 15144
rect 15611 15113 15623 15116
rect 15565 15107 15623 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 16758 15144 16764 15156
rect 16540 15116 16764 15144
rect 16540 15104 16546 15116
rect 16758 15104 16764 15116
rect 16816 15104 16822 15156
rect 17310 15104 17316 15156
rect 17368 15144 17374 15156
rect 18230 15144 18236 15156
rect 17368 15116 18236 15144
rect 17368 15104 17374 15116
rect 18230 15104 18236 15116
rect 18288 15104 18294 15156
rect 18432 15116 20024 15144
rect 658 15036 664 15088
rect 716 15076 722 15088
rect 5534 15076 5540 15088
rect 716 15048 5540 15076
rect 716 15036 722 15048
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 5629 15079 5687 15085
rect 5629 15045 5641 15079
rect 5675 15076 5687 15079
rect 8938 15076 8944 15088
rect 5675 15048 8944 15076
rect 5675 15045 5687 15048
rect 5629 15039 5687 15045
rect 8938 15036 8944 15048
rect 8996 15036 9002 15088
rect 9585 15079 9643 15085
rect 9585 15045 9597 15079
rect 9631 15076 9643 15079
rect 10410 15076 10416 15088
rect 9631 15048 10416 15076
rect 9631 15045 9643 15048
rect 9585 15039 9643 15045
rect 10410 15036 10416 15048
rect 10468 15036 10474 15088
rect 12621 15079 12679 15085
rect 12621 15076 12633 15079
rect 10704 15048 11192 15076
rect 1765 15011 1823 15017
rect 1765 14977 1777 15011
rect 1811 15008 1823 15011
rect 2682 15008 2688 15020
rect 1811 14980 2688 15008
rect 1811 14977 1823 14980
rect 1765 14971 1823 14977
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 1302 14900 1308 14952
rect 1360 14940 1366 14952
rect 2041 14943 2099 14949
rect 2041 14940 2053 14943
rect 1360 14912 2053 14940
rect 1360 14900 1366 14912
rect 2041 14909 2053 14912
rect 2087 14909 2099 14943
rect 3620 14940 3648 14971
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 4433 15011 4491 15017
rect 4433 15008 4445 15011
rect 3752 14980 4445 15008
rect 3752 14968 3758 14980
rect 4433 14977 4445 14980
rect 4479 14977 4491 15011
rect 6641 15011 6699 15017
rect 4433 14971 4491 14977
rect 4632 14980 6040 15008
rect 3970 14940 3976 14952
rect 3620 14912 3976 14940
rect 2041 14903 2099 14909
rect 3970 14900 3976 14912
rect 4028 14900 4034 14952
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4632 14940 4660 14980
rect 4120 14912 4660 14940
rect 4120 14900 4126 14912
rect 4706 14900 4712 14952
rect 4764 14900 4770 14952
rect 5350 14900 5356 14952
rect 5408 14940 5414 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 5408 14912 5825 14940
rect 5408 14900 5414 14912
rect 5813 14909 5825 14912
rect 5859 14909 5871 14943
rect 6012 14940 6040 14980
rect 6641 14977 6653 15011
rect 6687 15008 6699 15011
rect 6822 15008 6828 15020
rect 6687 14980 6828 15008
rect 6687 14977 6699 14980
rect 6641 14971 6699 14977
rect 6822 14968 6828 14980
rect 6880 14968 6886 15020
rect 7650 14968 7656 15020
rect 7708 15008 7714 15020
rect 7929 15011 7987 15017
rect 7929 15008 7941 15011
rect 7708 14980 7941 15008
rect 7708 14968 7714 14980
rect 7929 14977 7941 14980
rect 7975 14977 7987 15011
rect 7929 14971 7987 14977
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9272 14980 9812 15008
rect 9272 14968 9278 14980
rect 7098 14940 7104 14952
rect 6012 14912 7104 14940
rect 5813 14903 5871 14909
rect 7098 14900 7104 14912
rect 7156 14940 7162 14952
rect 8113 14943 8171 14949
rect 8113 14940 8125 14943
rect 7156 14912 8125 14940
rect 7156 14900 7162 14912
rect 8113 14909 8125 14912
rect 8159 14940 8171 14943
rect 8570 14940 8576 14952
rect 8159 14912 8576 14940
rect 8159 14909 8171 14912
rect 8113 14903 8171 14909
rect 8570 14900 8576 14912
rect 8628 14900 8634 14952
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14940 8999 14943
rect 9582 14940 9588 14952
rect 8987 14912 9588 14940
rect 8987 14909 8999 14912
rect 8941 14903 8999 14909
rect 9582 14900 9588 14912
rect 9640 14900 9646 14952
rect 9784 14949 9812 14980
rect 9858 14968 9864 15020
rect 9916 15008 9922 15020
rect 10704 15008 10732 15048
rect 9916 14980 10732 15008
rect 10781 15011 10839 15017
rect 9916 14968 9922 14980
rect 10428 14952 10456 14980
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10962 15008 10968 15020
rect 10827 14980 10968 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 9769 14943 9827 14949
rect 9769 14909 9781 14943
rect 9815 14909 9827 14943
rect 9769 14903 9827 14909
rect 10410 14900 10416 14952
rect 10468 14900 10474 14952
rect 10594 14900 10600 14952
rect 10652 14940 10658 14952
rect 10873 14943 10931 14949
rect 10873 14940 10885 14943
rect 10652 14912 10885 14940
rect 10652 14900 10658 14912
rect 10873 14909 10885 14912
rect 10919 14909 10931 14943
rect 10873 14903 10931 14909
rect 11057 14943 11115 14949
rect 11057 14909 11069 14943
rect 11103 14940 11115 14943
rect 11164 14940 11192 15048
rect 11103 14912 11192 14940
rect 11256 15048 12633 15076
rect 11103 14909 11115 14912
rect 11057 14903 11115 14909
rect 1762 14832 1768 14884
rect 1820 14872 1826 14884
rect 6825 14875 6883 14881
rect 6825 14872 6837 14875
rect 1820 14844 6837 14872
rect 1820 14832 1826 14844
rect 6825 14841 6837 14844
rect 6871 14841 6883 14875
rect 6825 14835 6883 14841
rect 8018 14832 8024 14884
rect 8076 14872 8082 14884
rect 11256 14872 11284 15048
rect 12621 15045 12633 15048
rect 12667 15076 12679 15079
rect 13170 15076 13176 15088
rect 12667 15048 13176 15076
rect 12667 15045 12679 15048
rect 12621 15039 12679 15045
rect 13170 15036 13176 15048
rect 13228 15036 13234 15088
rect 13630 15036 13636 15088
rect 13688 15076 13694 15088
rect 13725 15079 13783 15085
rect 13725 15076 13737 15079
rect 13688 15048 13737 15076
rect 13688 15036 13694 15048
rect 13725 15045 13737 15048
rect 13771 15045 13783 15079
rect 14200 15076 14228 15104
rect 18432 15076 18460 15116
rect 19996 15085 20024 15116
rect 20622 15104 20628 15156
rect 20680 15144 20686 15156
rect 21453 15147 21511 15153
rect 21453 15144 21465 15147
rect 20680 15116 21465 15144
rect 20680 15104 20686 15116
rect 21453 15113 21465 15116
rect 21499 15113 21511 15147
rect 21453 15107 21511 15113
rect 21542 15104 21548 15156
rect 21600 15144 21606 15156
rect 28626 15144 28632 15156
rect 21600 15116 28632 15144
rect 21600 15104 21606 15116
rect 28626 15104 28632 15116
rect 28684 15104 28690 15156
rect 29178 15104 29184 15156
rect 29236 15144 29242 15156
rect 33502 15144 33508 15156
rect 29236 15116 33508 15144
rect 29236 15104 29242 15116
rect 33502 15104 33508 15116
rect 33560 15104 33566 15156
rect 14200 15048 18460 15076
rect 19981 15079 20039 15085
rect 13725 15039 13783 15045
rect 19981 15045 19993 15079
rect 20027 15045 20039 15079
rect 19981 15039 20039 15045
rect 20990 15036 20996 15088
rect 21048 15036 21054 15088
rect 23842 15076 23848 15088
rect 23782 15048 23848 15076
rect 23842 15036 23848 15048
rect 23900 15076 23906 15088
rect 24302 15076 24308 15088
rect 23900 15048 24308 15076
rect 23900 15036 23906 15048
rect 24302 15036 24308 15048
rect 24360 15076 24366 15088
rect 24581 15079 24639 15085
rect 24360 15048 24532 15076
rect 24360 15036 24366 15048
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 12492 14980 13553 15008
rect 12492 14968 12498 14980
rect 13541 14977 13553 14980
rect 13587 15008 13599 15011
rect 13906 15008 13912 15020
rect 13587 14980 13912 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14182 14968 14188 15020
rect 14240 15008 14246 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 14240 14980 14749 15008
rect 14240 14968 14246 14980
rect 14737 14977 14749 14980
rect 14783 14977 14795 15011
rect 14737 14971 14795 14977
rect 15933 15011 15991 15017
rect 15933 14977 15945 15011
rect 15979 14977 15991 15011
rect 15933 14971 15991 14977
rect 16025 15011 16083 15017
rect 16025 14977 16037 15011
rect 16071 15008 16083 15011
rect 16574 15008 16580 15020
rect 16071 14980 16580 15008
rect 16071 14977 16083 14980
rect 16025 14971 16083 14977
rect 12526 14900 12532 14952
rect 12584 14940 12590 14952
rect 12805 14943 12863 14949
rect 12805 14940 12817 14943
rect 12584 14912 12817 14940
rect 12584 14900 12590 14912
rect 12805 14909 12817 14912
rect 12851 14909 12863 14943
rect 12805 14903 12863 14909
rect 14093 14943 14151 14949
rect 14093 14909 14105 14943
rect 14139 14940 14151 14943
rect 14458 14940 14464 14952
rect 14139 14912 14464 14940
rect 14139 14909 14151 14912
rect 14093 14903 14151 14909
rect 14458 14900 14464 14912
rect 14516 14940 14522 14952
rect 14829 14943 14887 14949
rect 14829 14940 14841 14943
rect 14516 14912 14841 14940
rect 14516 14900 14522 14912
rect 14829 14909 14841 14912
rect 14875 14909 14887 14943
rect 14829 14903 14887 14909
rect 15010 14900 15016 14952
rect 15068 14900 15074 14952
rect 15948 14872 15976 14971
rect 16574 14968 16580 14980
rect 16632 15008 16638 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 17221 15011 17279 15017
rect 17221 14977 17233 15011
rect 17267 15008 17279 15011
rect 17267 14980 19380 15008
rect 17267 14977 17279 14980
rect 17221 14971 17279 14977
rect 16209 14943 16267 14949
rect 16209 14909 16221 14943
rect 16255 14940 16267 14943
rect 18782 14940 18788 14952
rect 16255 14912 18788 14940
rect 16255 14909 16267 14912
rect 16209 14903 16267 14909
rect 18782 14900 18788 14912
rect 18840 14900 18846 14952
rect 18969 14943 19027 14949
rect 18969 14909 18981 14943
rect 19015 14940 19027 14943
rect 19058 14940 19064 14952
rect 19015 14912 19064 14940
rect 19015 14909 19027 14912
rect 18969 14903 19027 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 16853 14875 16911 14881
rect 16853 14872 16865 14875
rect 8076 14844 11284 14872
rect 11716 14844 16865 14872
rect 8076 14832 8082 14844
rect 2682 14764 2688 14816
rect 2740 14804 2746 14816
rect 2774 14804 2780 14816
rect 2740 14776 2780 14804
rect 2740 14764 2746 14776
rect 2774 14764 2780 14776
rect 2832 14764 2838 14816
rect 3418 14764 3424 14816
rect 3476 14764 3482 14816
rect 4065 14807 4123 14813
rect 4065 14773 4077 14807
rect 4111 14804 4123 14807
rect 5074 14804 5080 14816
rect 4111 14776 5080 14804
rect 4111 14773 4123 14776
rect 4065 14767 4123 14773
rect 5074 14764 5080 14776
rect 5132 14764 5138 14816
rect 5258 14764 5264 14816
rect 5316 14764 5322 14816
rect 5534 14764 5540 14816
rect 5592 14804 5598 14816
rect 5994 14804 6000 14816
rect 5592 14776 6000 14804
rect 5592 14764 5598 14776
rect 5994 14764 6000 14776
rect 6052 14764 6058 14816
rect 6730 14764 6736 14816
rect 6788 14804 6794 14816
rect 7190 14804 7196 14816
rect 6788 14776 7196 14804
rect 6788 14764 6794 14776
rect 7190 14764 7196 14776
rect 7248 14764 7254 14816
rect 7282 14764 7288 14816
rect 7340 14804 7346 14816
rect 7561 14807 7619 14813
rect 7561 14804 7573 14807
rect 7340 14776 7573 14804
rect 7340 14764 7346 14776
rect 7561 14773 7573 14776
rect 7607 14773 7619 14807
rect 7561 14767 7619 14773
rect 8754 14764 8760 14816
rect 8812 14804 8818 14816
rect 9030 14804 9036 14816
rect 8812 14776 9036 14804
rect 8812 14764 8818 14776
rect 9030 14764 9036 14776
rect 9088 14764 9094 14816
rect 9217 14807 9275 14813
rect 9217 14773 9229 14807
rect 9263 14804 9275 14807
rect 9766 14804 9772 14816
rect 9263 14776 9772 14804
rect 9263 14773 9275 14776
rect 9217 14767 9275 14773
rect 9766 14764 9772 14776
rect 9824 14764 9830 14816
rect 9858 14764 9864 14816
rect 9916 14804 9922 14816
rect 10413 14807 10471 14813
rect 10413 14804 10425 14807
rect 9916 14776 10425 14804
rect 9916 14764 9922 14776
rect 10413 14773 10425 14776
rect 10459 14773 10471 14807
rect 10413 14767 10471 14773
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 11716 14804 11744 14844
rect 16853 14841 16865 14844
rect 16899 14841 16911 14875
rect 16853 14835 16911 14841
rect 17126 14832 17132 14884
rect 17184 14872 17190 14884
rect 18046 14872 18052 14884
rect 17184 14844 18052 14872
rect 17184 14832 17190 14844
rect 18046 14832 18052 14844
rect 18104 14832 18110 14884
rect 18230 14832 18236 14884
rect 18288 14872 18294 14884
rect 18506 14872 18512 14884
rect 18288 14844 18512 14872
rect 18288 14832 18294 14844
rect 18506 14832 18512 14844
rect 18564 14832 18570 14884
rect 10652 14776 11744 14804
rect 10652 14764 10658 14776
rect 11790 14764 11796 14816
rect 11848 14764 11854 14816
rect 11977 14807 12035 14813
rect 11977 14773 11989 14807
rect 12023 14804 12035 14807
rect 13262 14804 13268 14816
rect 12023 14776 13268 14804
rect 12023 14773 12035 14776
rect 11977 14767 12035 14773
rect 13262 14764 13268 14776
rect 13320 14764 13326 14816
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 14366 14804 14372 14816
rect 13688 14776 14372 14804
rect 13688 14764 13694 14776
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 18690 14804 18696 14816
rect 14700 14776 18696 14804
rect 14700 14764 14706 14776
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19352 14813 19380 14980
rect 22278 14968 22284 15020
rect 22336 14968 22342 15020
rect 24210 14968 24216 15020
rect 24268 15008 24274 15020
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 24268 14980 24409 15008
rect 24268 14968 24274 14980
rect 24397 14977 24409 14980
rect 24443 14977 24455 15011
rect 24504 15008 24532 15048
rect 24581 15045 24593 15079
rect 24627 15076 24639 15079
rect 24762 15076 24768 15088
rect 24627 15048 24768 15076
rect 24627 15045 24639 15048
rect 24581 15039 24639 15045
rect 24762 15036 24768 15048
rect 24820 15036 24826 15088
rect 24872 15048 25622 15076
rect 24872 15008 24900 15048
rect 27706 15036 27712 15088
rect 27764 15076 27770 15088
rect 27764 15048 31064 15076
rect 27764 15036 27770 15048
rect 24504 14980 24900 15008
rect 24397 14971 24455 14977
rect 27614 14968 27620 15020
rect 27672 14968 27678 15020
rect 28718 14968 28724 15020
rect 28776 14968 28782 15020
rect 29454 14968 29460 15020
rect 29512 15008 29518 15020
rect 29825 15011 29883 15017
rect 29825 15008 29837 15011
rect 29512 14980 29837 15008
rect 29512 14968 29518 14980
rect 29825 14977 29837 14980
rect 29871 14977 29883 15011
rect 29825 14971 29883 14977
rect 30926 14968 30932 15020
rect 30984 14968 30990 15020
rect 31036 15008 31064 15048
rect 31110 15036 31116 15088
rect 31168 15076 31174 15088
rect 41414 15076 41420 15088
rect 31168 15048 41420 15076
rect 31168 15036 31174 15048
rect 41414 15036 41420 15048
rect 41472 15036 41478 15088
rect 33594 15008 33600 15020
rect 31036 14980 33600 15008
rect 33594 14968 33600 14980
rect 33652 14968 33658 15020
rect 19702 14900 19708 14952
rect 19760 14900 19766 14952
rect 19978 14900 19984 14952
rect 20036 14940 20042 14952
rect 20036 14912 22094 14940
rect 20036 14900 20042 14912
rect 21082 14832 21088 14884
rect 21140 14872 21146 14884
rect 21910 14872 21916 14884
rect 21140 14844 21916 14872
rect 21140 14832 21146 14844
rect 21910 14832 21916 14844
rect 21968 14832 21974 14884
rect 19337 14807 19395 14813
rect 19337 14773 19349 14807
rect 19383 14804 19395 14807
rect 20622 14804 20628 14816
rect 19383 14776 20628 14804
rect 19383 14773 19395 14776
rect 19337 14767 19395 14773
rect 20622 14764 20628 14776
rect 20680 14764 20686 14816
rect 21726 14764 21732 14816
rect 21784 14804 21790 14816
rect 21821 14807 21879 14813
rect 21821 14804 21833 14807
rect 21784 14776 21833 14804
rect 21784 14764 21790 14776
rect 21821 14773 21833 14776
rect 21867 14773 21879 14807
rect 22066 14804 22094 14912
rect 22554 14900 22560 14952
rect 22612 14900 22618 14952
rect 23290 14900 23296 14952
rect 23348 14940 23354 14952
rect 24857 14943 24915 14949
rect 24857 14940 24869 14943
rect 23348 14912 24869 14940
rect 23348 14900 23354 14912
rect 24857 14909 24869 14912
rect 24903 14909 24915 14943
rect 24857 14903 24915 14909
rect 25133 14943 25191 14949
rect 25133 14909 25145 14943
rect 25179 14940 25191 14943
rect 28261 14943 28319 14949
rect 28261 14940 28273 14943
rect 25179 14912 28273 14940
rect 25179 14909 25191 14912
rect 25133 14903 25191 14909
rect 28261 14909 28273 14912
rect 28307 14909 28319 14943
rect 28261 14903 28319 14909
rect 28442 14900 28448 14952
rect 28500 14940 28506 14952
rect 31294 14940 31300 14952
rect 28500 14912 31300 14940
rect 28500 14900 28506 14912
rect 31294 14900 31300 14912
rect 31352 14900 31358 14952
rect 31772 14912 38654 14940
rect 24029 14875 24087 14881
rect 24029 14841 24041 14875
rect 24075 14872 24087 14875
rect 24075 14844 24992 14872
rect 24075 14841 24087 14844
rect 24029 14835 24087 14841
rect 24854 14804 24860 14816
rect 22066 14776 24860 14804
rect 21821 14767 21879 14773
rect 24854 14764 24860 14776
rect 24912 14764 24918 14816
rect 24964 14804 24992 14844
rect 26878 14832 26884 14884
rect 26936 14872 26942 14884
rect 27157 14875 27215 14881
rect 27157 14872 27169 14875
rect 26936 14844 27169 14872
rect 26936 14832 26942 14844
rect 27157 14841 27169 14844
rect 27203 14841 27215 14875
rect 27157 14835 27215 14841
rect 27246 14832 27252 14884
rect 27304 14872 27310 14884
rect 31772 14872 31800 14912
rect 27304 14844 31800 14872
rect 38626 14872 38654 14912
rect 44818 14872 44824 14884
rect 38626 14844 44824 14872
rect 27304 14832 27310 14844
rect 44818 14832 44824 14844
rect 44876 14832 44882 14884
rect 25314 14804 25320 14816
rect 24964 14776 25320 14804
rect 25314 14764 25320 14776
rect 25372 14804 25378 14816
rect 25866 14804 25872 14816
rect 25372 14776 25872 14804
rect 25372 14764 25378 14776
rect 25866 14764 25872 14776
rect 25924 14764 25930 14816
rect 26602 14764 26608 14816
rect 26660 14764 26666 14816
rect 27062 14764 27068 14816
rect 27120 14764 27126 14816
rect 29362 14764 29368 14816
rect 29420 14764 29426 14816
rect 30374 14764 30380 14816
rect 30432 14804 30438 14816
rect 30469 14807 30527 14813
rect 30469 14804 30481 14807
rect 30432 14776 30481 14804
rect 30432 14764 30438 14776
rect 30469 14773 30481 14776
rect 30515 14773 30527 14807
rect 30469 14767 30527 14773
rect 31570 14764 31576 14816
rect 31628 14764 31634 14816
rect 31662 14764 31668 14816
rect 31720 14804 31726 14816
rect 31849 14807 31907 14813
rect 31849 14804 31861 14807
rect 31720 14776 31861 14804
rect 31720 14764 31726 14776
rect 31849 14773 31861 14776
rect 31895 14773 31907 14807
rect 31849 14767 31907 14773
rect 33594 14764 33600 14816
rect 33652 14804 33658 14816
rect 40402 14804 40408 14816
rect 33652 14776 40408 14804
rect 33652 14764 33658 14776
rect 40402 14764 40408 14776
rect 40460 14764 40466 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 2130 14600 2136 14612
rect 1820 14572 2136 14600
rect 1820 14560 1826 14572
rect 2130 14560 2136 14572
rect 2188 14560 2194 14612
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3510 14600 3516 14612
rect 3467 14572 3516 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 3881 14603 3939 14609
rect 3881 14569 3893 14603
rect 3927 14600 3939 14603
rect 6270 14600 6276 14612
rect 3927 14572 6276 14600
rect 3927 14569 3939 14572
rect 3881 14563 3939 14569
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 3988 14473 4016 14572
rect 6270 14560 6276 14572
rect 6328 14560 6334 14612
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 6696 14572 7328 14600
rect 6696 14560 6702 14572
rect 7190 14492 7196 14544
rect 7248 14492 7254 14544
rect 7300 14532 7328 14572
rect 7834 14560 7840 14612
rect 7892 14600 7898 14612
rect 9398 14600 9404 14612
rect 7892 14572 9404 14600
rect 7892 14560 7898 14572
rect 9398 14560 9404 14572
rect 9456 14560 9462 14612
rect 10226 14560 10232 14612
rect 10284 14600 10290 14612
rect 12434 14600 12440 14612
rect 10284 14572 12440 14600
rect 10284 14560 10290 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 12526 14560 12532 14612
rect 12584 14600 12590 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 12584 14572 13553 14600
rect 12584 14560 12590 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 13541 14563 13599 14569
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 13964 14572 18736 14600
rect 13964 14560 13970 14572
rect 8573 14535 8631 14541
rect 8573 14532 8585 14535
rect 7300 14504 8585 14532
rect 8573 14501 8585 14504
rect 8619 14501 8631 14535
rect 8573 14495 8631 14501
rect 8662 14492 8668 14544
rect 8720 14532 8726 14544
rect 10413 14535 10471 14541
rect 10413 14532 10425 14535
rect 8720 14504 10425 14532
rect 8720 14492 8726 14504
rect 10413 14501 10425 14504
rect 10459 14501 10471 14535
rect 18708 14532 18736 14572
rect 18782 14560 18788 14612
rect 18840 14600 18846 14612
rect 18877 14603 18935 14609
rect 18877 14600 18889 14603
rect 18840 14572 18889 14600
rect 18840 14560 18846 14572
rect 18877 14569 18889 14572
rect 18923 14569 18935 14603
rect 18877 14563 18935 14569
rect 22554 14560 22560 14612
rect 22612 14600 22618 14612
rect 28905 14603 28963 14609
rect 28905 14600 28917 14603
rect 22612 14572 28917 14600
rect 22612 14560 22618 14572
rect 28905 14569 28917 14572
rect 28951 14569 28963 14603
rect 28905 14563 28963 14569
rect 28994 14560 29000 14612
rect 29052 14600 29058 14612
rect 29730 14600 29736 14612
rect 29052 14572 29736 14600
rect 29052 14560 29058 14572
rect 29730 14560 29736 14572
rect 29788 14560 29794 14612
rect 30377 14603 30435 14609
rect 30377 14569 30389 14603
rect 30423 14600 30435 14603
rect 30926 14600 30932 14612
rect 30423 14572 30932 14600
rect 30423 14569 30435 14572
rect 30377 14563 30435 14569
rect 30926 14560 30932 14572
rect 30984 14560 30990 14612
rect 42518 14600 42524 14612
rect 31726 14572 42524 14600
rect 21542 14532 21548 14544
rect 18708 14504 21548 14532
rect 10413 14495 10471 14501
rect 21542 14492 21548 14504
rect 21600 14492 21606 14544
rect 24210 14532 24216 14544
rect 21836 14504 24216 14532
rect 2041 14467 2099 14473
rect 2041 14464 2053 14467
rect 1360 14436 2053 14464
rect 1360 14424 1366 14436
rect 2041 14433 2053 14436
rect 2087 14433 2099 14467
rect 2041 14427 2099 14433
rect 3973 14467 4031 14473
rect 3973 14433 3985 14467
rect 4019 14433 4031 14467
rect 3973 14427 4031 14433
rect 5074 14424 5080 14476
rect 5132 14424 5138 14476
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5718 14464 5724 14476
rect 5307 14436 5724 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 7208 14464 7236 14492
rect 10873 14467 10931 14473
rect 10873 14464 10885 14467
rect 7208 14436 10885 14464
rect 10873 14433 10885 14436
rect 10919 14433 10931 14467
rect 10873 14427 10931 14433
rect 1765 14399 1823 14405
rect 1765 14365 1777 14399
rect 1811 14396 1823 14399
rect 3602 14396 3608 14408
rect 1811 14368 3608 14396
rect 1811 14365 1823 14368
rect 1765 14359 1823 14365
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 4798 14356 4804 14408
rect 4856 14396 4862 14408
rect 5813 14399 5871 14405
rect 5813 14396 5825 14399
rect 4856 14368 5825 14396
rect 4856 14356 4862 14368
rect 5813 14365 5825 14368
rect 5859 14365 5871 14399
rect 8389 14399 8447 14405
rect 5813 14359 5871 14365
rect 7484 14368 8340 14396
rect 4982 14288 4988 14340
rect 5040 14288 5046 14340
rect 5626 14288 5632 14340
rect 5684 14328 5690 14340
rect 6089 14331 6147 14337
rect 6089 14328 6101 14331
rect 5684 14300 6101 14328
rect 5684 14288 5690 14300
rect 6089 14297 6101 14300
rect 6135 14297 6147 14331
rect 6546 14328 6552 14340
rect 6089 14291 6147 14297
rect 6288 14300 6552 14328
rect 3602 14220 3608 14272
rect 3660 14220 3666 14272
rect 4617 14263 4675 14269
rect 4617 14229 4629 14263
rect 4663 14260 4675 14263
rect 5442 14260 5448 14272
rect 4663 14232 5448 14260
rect 4663 14229 4675 14232
rect 4617 14223 4675 14229
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 5534 14220 5540 14272
rect 5592 14260 5598 14272
rect 6288 14260 6316 14300
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 5592 14232 6316 14260
rect 5592 14220 5598 14232
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 7484 14260 7512 14368
rect 7837 14331 7895 14337
rect 7837 14297 7849 14331
rect 7883 14328 7895 14331
rect 7926 14328 7932 14340
rect 7883 14300 7932 14328
rect 7883 14297 7895 14300
rect 7837 14291 7895 14297
rect 7926 14288 7932 14300
rect 7984 14288 7990 14340
rect 8312 14328 8340 14368
rect 8389 14365 8401 14399
rect 8435 14396 8447 14399
rect 8478 14396 8484 14408
rect 8435 14368 8484 14396
rect 8435 14365 8447 14368
rect 8389 14359 8447 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 8938 14356 8944 14408
rect 8996 14396 9002 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8996 14368 9137 14396
rect 8996 14356 9002 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9401 14399 9459 14405
rect 9401 14365 9413 14399
rect 9447 14396 9459 14399
rect 9582 14396 9588 14408
rect 9447 14368 9588 14396
rect 9447 14365 9459 14368
rect 9401 14359 9459 14365
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10686 14356 10692 14408
rect 10744 14396 10750 14408
rect 10781 14399 10839 14405
rect 10781 14396 10793 14399
rect 10744 14368 10793 14396
rect 10744 14356 10750 14368
rect 10781 14365 10793 14368
rect 10827 14365 10839 14399
rect 10888 14396 10916 14427
rect 10962 14424 10968 14476
rect 11020 14424 11026 14476
rect 14182 14464 14188 14476
rect 11072 14436 14188 14464
rect 11072 14396 11100 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14550 14424 14556 14476
rect 14608 14464 14614 14476
rect 15378 14464 15384 14476
rect 14608 14436 15384 14464
rect 14608 14424 14614 14436
rect 15378 14424 15384 14436
rect 15436 14424 15442 14476
rect 16942 14424 16948 14476
rect 17000 14464 17006 14476
rect 17129 14467 17187 14473
rect 17129 14464 17141 14467
rect 17000 14436 17141 14464
rect 17000 14424 17006 14436
rect 17129 14433 17141 14436
rect 17175 14464 17187 14467
rect 19702 14464 19708 14476
rect 17175 14436 19708 14464
rect 17175 14433 17187 14436
rect 17129 14427 17187 14433
rect 19702 14424 19708 14436
rect 19760 14464 19766 14476
rect 20165 14467 20223 14473
rect 20165 14464 20177 14467
rect 19760 14436 20177 14464
rect 19760 14424 19766 14436
rect 20165 14433 20177 14436
rect 20211 14433 20223 14467
rect 20165 14427 20223 14433
rect 20254 14424 20260 14476
rect 20312 14464 20318 14476
rect 20901 14467 20959 14473
rect 20901 14464 20913 14467
rect 20312 14436 20913 14464
rect 20312 14424 20318 14436
rect 20901 14433 20913 14436
rect 20947 14464 20959 14467
rect 21358 14464 21364 14476
rect 20947 14436 21364 14464
rect 20947 14433 20959 14436
rect 20901 14427 20959 14433
rect 21358 14424 21364 14436
rect 21416 14424 21422 14476
rect 21450 14424 21456 14476
rect 21508 14464 21514 14476
rect 21836 14464 21864 14504
rect 24210 14492 24216 14504
rect 24268 14492 24274 14544
rect 24397 14535 24455 14541
rect 24397 14501 24409 14535
rect 24443 14532 24455 14535
rect 24578 14532 24584 14544
rect 24443 14504 24584 14532
rect 24443 14501 24455 14504
rect 24397 14495 24455 14501
rect 24578 14492 24584 14504
rect 24636 14492 24642 14544
rect 26237 14535 26295 14541
rect 26237 14532 26249 14535
rect 25608 14504 26249 14532
rect 21508 14436 21864 14464
rect 21508 14424 21514 14436
rect 10888 14368 11100 14396
rect 10781 14359 10839 14365
rect 10594 14328 10600 14340
rect 8312 14300 10600 14328
rect 10594 14288 10600 14300
rect 10652 14288 10658 14340
rect 10796 14328 10824 14359
rect 11790 14356 11796 14408
rect 11848 14356 11854 14408
rect 13354 14356 13360 14408
rect 13412 14396 13418 14408
rect 13906 14396 13912 14408
rect 13412 14368 13912 14396
rect 13412 14356 13418 14368
rect 13906 14356 13912 14368
rect 13964 14356 13970 14408
rect 14642 14356 14648 14408
rect 14700 14356 14706 14408
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 19518 14396 19524 14408
rect 18748 14368 19524 14396
rect 18748 14356 18754 14368
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 19852 14368 20637 14396
rect 19852 14356 19858 14368
rect 20625 14365 20637 14368
rect 20671 14396 20683 14399
rect 21729 14399 21787 14405
rect 20671 14368 21680 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 11422 14328 11428 14340
rect 10796 14300 11428 14328
rect 11422 14288 11428 14300
rect 11480 14288 11486 14340
rect 12069 14331 12127 14337
rect 12069 14297 12081 14331
rect 12115 14297 12127 14331
rect 12069 14291 12127 14297
rect 6420 14232 7512 14260
rect 6420 14220 6426 14232
rect 7558 14220 7564 14272
rect 7616 14260 7622 14272
rect 10686 14260 10692 14272
rect 7616 14232 10692 14260
rect 7616 14220 7622 14232
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 12084 14260 12112 14291
rect 12618 14288 12624 14340
rect 12676 14288 12682 14340
rect 13814 14288 13820 14340
rect 13872 14328 13878 14340
rect 14921 14331 14979 14337
rect 14921 14328 14933 14331
rect 13872 14300 14933 14328
rect 13872 14288 13878 14300
rect 14921 14297 14933 14300
rect 14967 14297 14979 14331
rect 14921 14291 14979 14297
rect 15654 14288 15660 14340
rect 15712 14288 15718 14340
rect 16942 14288 16948 14340
rect 17000 14328 17006 14340
rect 17310 14328 17316 14340
rect 17000 14300 17316 14328
rect 17000 14288 17006 14300
rect 17310 14288 17316 14300
rect 17368 14288 17374 14340
rect 17402 14288 17408 14340
rect 17460 14288 17466 14340
rect 17678 14288 17684 14340
rect 17736 14328 17742 14340
rect 17736 14300 17894 14328
rect 17736 14288 17742 14300
rect 19058 14288 19064 14340
rect 19116 14328 19122 14340
rect 19426 14328 19432 14340
rect 19116 14300 19432 14328
rect 19116 14288 19122 14300
rect 19426 14288 19432 14300
rect 19484 14328 19490 14340
rect 21085 14331 21143 14337
rect 21085 14328 21097 14331
rect 19484 14300 21097 14328
rect 19484 14288 19490 14300
rect 21085 14297 21097 14300
rect 21131 14328 21143 14331
rect 21652 14328 21680 14368
rect 21729 14365 21741 14399
rect 21775 14396 21787 14399
rect 21836 14396 21864 14436
rect 21910 14424 21916 14476
rect 21968 14424 21974 14476
rect 22278 14424 22284 14476
rect 22336 14464 22342 14476
rect 23290 14464 23296 14476
rect 22336 14436 23296 14464
rect 22336 14424 22342 14436
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 23474 14424 23480 14476
rect 23532 14464 23538 14476
rect 24029 14467 24087 14473
rect 24029 14464 24041 14467
rect 23532 14436 24041 14464
rect 23532 14424 23538 14436
rect 24029 14433 24041 14436
rect 24075 14464 24087 14467
rect 24486 14464 24492 14476
rect 24075 14436 24492 14464
rect 24075 14433 24087 14436
rect 24029 14427 24087 14433
rect 24486 14424 24492 14436
rect 24544 14424 24550 14476
rect 21775 14368 21864 14396
rect 21775 14365 21787 14368
rect 21729 14359 21787 14365
rect 22094 14356 22100 14408
rect 22152 14396 22158 14408
rect 24578 14396 24584 14408
rect 22152 14368 24584 14396
rect 22152 14356 22158 14368
rect 24578 14356 24584 14368
rect 24636 14356 24642 14408
rect 25498 14356 25504 14408
rect 25556 14396 25562 14408
rect 25608 14405 25636 14504
rect 26237 14501 26249 14504
rect 26283 14532 26295 14535
rect 26421 14535 26479 14541
rect 26421 14532 26433 14535
rect 26283 14504 26433 14532
rect 26283 14501 26295 14504
rect 26237 14495 26295 14501
rect 26421 14501 26433 14504
rect 26467 14501 26479 14535
rect 26421 14495 26479 14501
rect 26786 14492 26792 14544
rect 26844 14532 26850 14544
rect 28442 14532 28448 14544
rect 26844 14504 28448 14532
rect 26844 14492 26850 14504
rect 28442 14492 28448 14504
rect 28500 14492 28506 14544
rect 28810 14492 28816 14544
rect 28868 14532 28874 14544
rect 31726 14532 31754 14572
rect 42518 14560 42524 14572
rect 42576 14560 42582 14612
rect 28868 14504 31754 14532
rect 28868 14492 28874 14504
rect 31846 14492 31852 14544
rect 31904 14532 31910 14544
rect 37642 14532 37648 14544
rect 31904 14504 37648 14532
rect 31904 14492 31910 14504
rect 37642 14492 37648 14504
rect 37700 14492 37706 14544
rect 25866 14424 25872 14476
rect 25924 14424 25930 14476
rect 26694 14424 26700 14476
rect 26752 14464 26758 14476
rect 30282 14464 30288 14476
rect 26752 14436 30288 14464
rect 26752 14424 26758 14436
rect 30282 14424 30288 14436
rect 30340 14424 30346 14476
rect 30742 14424 30748 14476
rect 30800 14464 30806 14476
rect 31113 14467 31171 14473
rect 31113 14464 31125 14467
rect 30800 14436 31125 14464
rect 30800 14424 30806 14436
rect 31113 14433 31125 14436
rect 31159 14433 31171 14467
rect 31113 14427 31171 14433
rect 25593 14399 25651 14405
rect 25593 14396 25605 14399
rect 25556 14368 25605 14396
rect 25556 14356 25562 14368
rect 25593 14365 25605 14368
rect 25639 14365 25651 14399
rect 25884 14396 25912 14424
rect 27157 14399 27215 14405
rect 27157 14396 27169 14399
rect 25884 14368 27169 14396
rect 25593 14359 25651 14365
rect 27157 14365 27169 14368
rect 27203 14365 27215 14399
rect 27157 14359 27215 14365
rect 28261 14399 28319 14405
rect 28261 14365 28273 14399
rect 28307 14396 28319 14399
rect 29362 14396 29368 14408
rect 28307 14368 29368 14396
rect 28307 14365 28319 14368
rect 28261 14359 28319 14365
rect 29362 14356 29368 14368
rect 29420 14356 29426 14408
rect 29472 14368 29684 14396
rect 21131 14300 21496 14328
rect 21652 14300 21864 14328
rect 21131 14297 21143 14300
rect 21085 14291 21143 14297
rect 12802 14260 12808 14272
rect 12084 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13078 14220 13084 14272
rect 13136 14260 13142 14272
rect 15838 14260 15844 14272
rect 13136 14232 15844 14260
rect 13136 14220 13142 14232
rect 15838 14220 15844 14232
rect 15896 14220 15902 14272
rect 16390 14220 16396 14272
rect 16448 14220 16454 14272
rect 16761 14263 16819 14269
rect 16761 14229 16773 14263
rect 16807 14260 16819 14263
rect 17494 14260 17500 14272
rect 16807 14232 17500 14260
rect 16807 14229 16819 14232
rect 16761 14223 16819 14229
rect 17494 14220 17500 14232
rect 17552 14220 17558 14272
rect 18046 14220 18052 14272
rect 18104 14260 18110 14272
rect 19886 14260 19892 14272
rect 18104 14232 19892 14260
rect 18104 14220 18110 14232
rect 19886 14220 19892 14232
rect 19944 14220 19950 14272
rect 21358 14220 21364 14272
rect 21416 14220 21422 14272
rect 21468 14260 21496 14300
rect 21726 14260 21732 14272
rect 21468 14232 21732 14260
rect 21726 14220 21732 14232
rect 21784 14220 21790 14272
rect 21836 14269 21864 14300
rect 22278 14288 22284 14340
rect 22336 14328 22342 14340
rect 22557 14331 22615 14337
rect 22557 14328 22569 14331
rect 22336 14300 22569 14328
rect 22336 14288 22342 14300
rect 22557 14297 22569 14300
rect 22603 14328 22615 14331
rect 23290 14328 23296 14340
rect 22603 14300 23296 14328
rect 22603 14297 22615 14300
rect 22557 14291 22615 14297
rect 23290 14288 23296 14300
rect 23348 14288 23354 14340
rect 23845 14331 23903 14337
rect 23845 14297 23857 14331
rect 23891 14328 23903 14331
rect 24210 14328 24216 14340
rect 23891 14300 24216 14328
rect 23891 14297 23903 14300
rect 23845 14291 23903 14297
rect 24210 14288 24216 14300
rect 24268 14328 24274 14340
rect 24857 14331 24915 14337
rect 24857 14328 24869 14331
rect 24268 14300 24869 14328
rect 24268 14288 24274 14300
rect 24857 14297 24869 14300
rect 24903 14328 24915 14331
rect 29472 14328 29500 14368
rect 24903 14300 29500 14328
rect 29656 14328 29684 14368
rect 29730 14356 29736 14408
rect 29788 14356 29794 14408
rect 30834 14356 30840 14408
rect 30892 14356 30898 14408
rect 46198 14328 46204 14340
rect 29656 14300 46204 14328
rect 24903 14297 24915 14300
rect 24857 14291 24915 14297
rect 46198 14288 46204 14300
rect 46256 14288 46262 14340
rect 21821 14263 21879 14269
rect 21821 14229 21833 14263
rect 21867 14260 21879 14263
rect 21910 14260 21916 14272
rect 21867 14232 21916 14260
rect 21867 14229 21879 14232
rect 21821 14223 21879 14229
rect 21910 14220 21916 14232
rect 21968 14220 21974 14272
rect 22462 14220 22468 14272
rect 22520 14260 22526 14272
rect 22922 14260 22928 14272
rect 22520 14232 22928 14260
rect 22520 14220 22526 14232
rect 22922 14220 22928 14232
rect 22980 14220 22986 14272
rect 23106 14220 23112 14272
rect 23164 14260 23170 14272
rect 23750 14260 23756 14272
rect 23164 14232 23756 14260
rect 23164 14220 23170 14232
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 24121 14263 24179 14269
rect 24121 14229 24133 14263
rect 24167 14260 24179 14263
rect 24302 14260 24308 14272
rect 24167 14232 24308 14260
rect 24167 14229 24179 14232
rect 24121 14223 24179 14229
rect 24302 14220 24308 14232
rect 24360 14220 24366 14272
rect 24762 14220 24768 14272
rect 24820 14220 24826 14272
rect 24946 14220 24952 14272
rect 25004 14260 25010 14272
rect 25225 14263 25283 14269
rect 25225 14260 25237 14263
rect 25004 14232 25237 14260
rect 25004 14220 25010 14232
rect 25225 14229 25237 14232
rect 25271 14229 25283 14263
rect 25225 14223 25283 14229
rect 25682 14220 25688 14272
rect 25740 14260 25746 14272
rect 26510 14260 26516 14272
rect 25740 14232 26516 14260
rect 25740 14220 25746 14232
rect 26510 14220 26516 14232
rect 26568 14260 26574 14272
rect 26605 14263 26663 14269
rect 26605 14260 26617 14263
rect 26568 14232 26617 14260
rect 26568 14220 26574 14232
rect 26605 14229 26617 14232
rect 26651 14260 26663 14263
rect 26694 14260 26700 14272
rect 26651 14232 26700 14260
rect 26651 14229 26663 14232
rect 26605 14223 26663 14229
rect 26694 14220 26700 14232
rect 26752 14220 26758 14272
rect 27706 14220 27712 14272
rect 27764 14260 27770 14272
rect 27801 14263 27859 14269
rect 27801 14260 27813 14263
rect 27764 14232 27813 14260
rect 27764 14220 27770 14232
rect 27801 14229 27813 14232
rect 27847 14229 27859 14263
rect 27801 14223 27859 14229
rect 28810 14220 28816 14272
rect 28868 14260 28874 14272
rect 29270 14260 29276 14272
rect 28868 14232 29276 14260
rect 28868 14220 28874 14232
rect 29270 14220 29276 14232
rect 29328 14220 29334 14272
rect 29362 14220 29368 14272
rect 29420 14220 29426 14272
rect 30282 14220 30288 14272
rect 30340 14260 30346 14272
rect 47854 14260 47860 14272
rect 30340 14232 47860 14260
rect 30340 14220 30346 14232
rect 47854 14220 47860 14232
rect 47912 14220 47918 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 4522 14056 4528 14068
rect 3660 14028 4528 14056
rect 3660 14016 3666 14028
rect 4522 14016 4528 14028
rect 4580 14016 4586 14068
rect 4982 14016 4988 14068
rect 5040 14056 5046 14068
rect 5040 14028 6040 14056
rect 5040 14016 5046 14028
rect 3697 13991 3755 13997
rect 3697 13957 3709 13991
rect 3743 13988 3755 13991
rect 3878 13988 3884 14000
rect 3743 13960 3884 13988
rect 3743 13957 3755 13960
rect 3697 13951 3755 13957
rect 3878 13948 3884 13960
rect 3936 13948 3942 14000
rect 4154 13988 4160 14000
rect 3988 13960 4160 13988
rect 290 13880 296 13932
rect 348 13920 354 13932
rect 1486 13920 1492 13932
rect 348 13892 1492 13920
rect 348 13880 354 13892
rect 1486 13880 1492 13892
rect 1544 13880 1550 13932
rect 1578 13880 1584 13932
rect 1636 13880 1642 13932
rect 2130 13880 2136 13932
rect 2188 13920 2194 13932
rect 3988 13929 4016 13960
rect 4154 13948 4160 13960
rect 4212 13948 4218 14000
rect 5534 13988 5540 14000
rect 5474 13960 5540 13988
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 6012 13997 6040 14028
rect 6914 14016 6920 14068
rect 6972 14056 6978 14068
rect 7377 14059 7435 14065
rect 7377 14056 7389 14059
rect 6972 14028 7389 14056
rect 6972 14016 6978 14028
rect 7377 14025 7389 14028
rect 7423 14025 7435 14059
rect 7377 14019 7435 14025
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 8018 14056 8024 14068
rect 7800 14028 8024 14056
rect 7800 14016 7806 14028
rect 8018 14016 8024 14028
rect 8076 14016 8082 14068
rect 8113 14059 8171 14065
rect 8113 14025 8125 14059
rect 8159 14056 8171 14059
rect 8386 14056 8392 14068
rect 8159 14028 8392 14056
rect 8159 14025 8171 14028
rect 8113 14019 8171 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 8573 14059 8631 14065
rect 8573 14025 8585 14059
rect 8619 14056 8631 14059
rect 9674 14056 9680 14068
rect 8619 14028 9680 14056
rect 8619 14025 8631 14028
rect 8573 14019 8631 14025
rect 9674 14016 9680 14028
rect 9732 14016 9738 14068
rect 12161 14059 12219 14065
rect 12161 14056 12173 14059
rect 9784 14028 12173 14056
rect 5997 13991 6055 13997
rect 5997 13957 6009 13991
rect 6043 13957 6055 13991
rect 5997 13951 6055 13957
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 6549 13991 6607 13997
rect 6549 13988 6561 13991
rect 6420 13960 6561 13988
rect 6420 13948 6426 13960
rect 6549 13957 6561 13960
rect 6595 13957 6607 13991
rect 6549 13951 6607 13957
rect 6638 13948 6644 14000
rect 6696 13988 6702 14000
rect 7285 13991 7343 13997
rect 7285 13988 7297 13991
rect 6696 13960 7297 13988
rect 6696 13948 6702 13960
rect 7285 13957 7297 13960
rect 7331 13957 7343 13991
rect 9784 13988 9812 14028
rect 12161 14025 12173 14028
rect 12207 14025 12219 14059
rect 12161 14019 12219 14025
rect 13262 14016 13268 14068
rect 13320 14056 13326 14068
rect 15565 14059 15623 14065
rect 15565 14056 15577 14059
rect 13320 14028 15577 14056
rect 13320 14016 13326 14028
rect 15565 14025 15577 14028
rect 15611 14056 15623 14059
rect 16393 14059 16451 14065
rect 16393 14056 16405 14059
rect 15611 14028 16405 14056
rect 15611 14025 15623 14028
rect 15565 14019 15623 14025
rect 16393 14025 16405 14028
rect 16439 14025 16451 14059
rect 16393 14019 16451 14025
rect 16666 14016 16672 14068
rect 16724 14056 16730 14068
rect 17126 14056 17132 14068
rect 16724 14028 17132 14056
rect 16724 14016 16730 14028
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 18046 14016 18052 14068
rect 18104 14056 18110 14068
rect 19521 14059 19579 14065
rect 19521 14056 19533 14059
rect 18104 14028 19533 14056
rect 18104 14016 18110 14028
rect 19521 14025 19533 14028
rect 19567 14025 19579 14059
rect 19521 14019 19579 14025
rect 19794 14016 19800 14068
rect 19852 14056 19858 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19852 14028 19901 14056
rect 19852 14016 19858 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 19889 14019 19947 14025
rect 19981 14059 20039 14065
rect 19981 14025 19993 14059
rect 20027 14056 20039 14059
rect 20254 14056 20260 14068
rect 20027 14028 20260 14056
rect 20027 14025 20039 14028
rect 19981 14019 20039 14025
rect 20254 14016 20260 14028
rect 20312 14016 20318 14068
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 20806 14056 20812 14068
rect 20763 14028 20812 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 20898 14016 20904 14068
rect 20956 14056 20962 14068
rect 21542 14056 21548 14068
rect 20956 14028 21548 14056
rect 20956 14016 20962 14028
rect 21542 14016 21548 14028
rect 21600 14016 21606 14068
rect 21726 14016 21732 14068
rect 21784 14056 21790 14068
rect 22189 14059 22247 14065
rect 22189 14056 22201 14059
rect 21784 14028 22201 14056
rect 21784 14016 21790 14028
rect 22189 14025 22201 14028
rect 22235 14056 22247 14059
rect 22278 14056 22284 14068
rect 22235 14028 22284 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 22462 14016 22468 14068
rect 22520 14056 22526 14068
rect 22738 14056 22744 14068
rect 22520 14028 22744 14056
rect 22520 14016 22526 14028
rect 22738 14016 22744 14028
rect 22796 14016 22802 14068
rect 23017 14059 23075 14065
rect 23017 14025 23029 14059
rect 23063 14056 23075 14059
rect 23474 14056 23480 14068
rect 23063 14028 23480 14056
rect 23063 14025 23075 14028
rect 23017 14019 23075 14025
rect 23474 14016 23480 14028
rect 23532 14016 23538 14068
rect 23566 14016 23572 14068
rect 23624 14056 23630 14068
rect 23845 14059 23903 14065
rect 23845 14056 23857 14059
rect 23624 14028 23857 14056
rect 23624 14016 23630 14028
rect 23845 14025 23857 14028
rect 23891 14025 23903 14059
rect 23845 14019 23903 14025
rect 24210 14016 24216 14068
rect 24268 14016 24274 14068
rect 25498 14016 25504 14068
rect 25556 14016 25562 14068
rect 25593 14059 25651 14065
rect 25593 14025 25605 14059
rect 25639 14056 25651 14059
rect 25682 14056 25688 14068
rect 25639 14028 25688 14056
rect 25639 14025 25651 14028
rect 25593 14019 25651 14025
rect 25682 14016 25688 14028
rect 25740 14016 25746 14068
rect 26237 14059 26295 14065
rect 26237 14025 26249 14059
rect 26283 14056 26295 14059
rect 26329 14059 26387 14065
rect 26329 14056 26341 14059
rect 26283 14028 26341 14056
rect 26283 14025 26295 14028
rect 26237 14019 26295 14025
rect 26329 14025 26341 14028
rect 26375 14056 26387 14059
rect 26418 14056 26424 14068
rect 26375 14028 26424 14056
rect 26375 14025 26387 14028
rect 26329 14019 26387 14025
rect 26418 14016 26424 14028
rect 26476 14016 26482 14068
rect 29270 14016 29276 14068
rect 29328 14056 29334 14068
rect 29641 14059 29699 14065
rect 29641 14056 29653 14059
rect 29328 14028 29653 14056
rect 29328 14016 29334 14028
rect 29641 14025 29653 14028
rect 29687 14025 29699 14059
rect 30285 14059 30343 14065
rect 30285 14056 30297 14059
rect 29641 14019 29699 14025
rect 29932 14028 30297 14056
rect 7285 13951 7343 13957
rect 8680 13960 9812 13988
rect 3973 13923 4031 13929
rect 2188 13892 3924 13920
rect 2188 13880 2194 13892
rect 1302 13812 1308 13864
rect 1360 13852 1366 13864
rect 2041 13855 2099 13861
rect 2041 13852 2053 13855
rect 1360 13824 2053 13852
rect 1360 13812 1366 13824
rect 2041 13821 2053 13824
rect 2087 13821 2099 13855
rect 2041 13815 2099 13821
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 3896 13852 3924 13892
rect 3973 13889 3985 13923
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 7558 13920 7564 13932
rect 6328 13892 7564 13920
rect 6328 13880 6334 13892
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 3896 13824 6377 13852
rect 6365 13821 6377 13824
rect 6411 13852 6423 13855
rect 7190 13852 7196 13864
rect 6411 13824 7196 13852
rect 6411 13821 6423 13824
rect 6365 13815 6423 13821
rect 7190 13812 7196 13824
rect 7248 13812 7254 13864
rect 7484 13861 7512 13892
rect 7558 13880 7564 13892
rect 7616 13920 7622 13932
rect 8386 13920 8392 13932
rect 7616 13892 8392 13920
rect 7616 13880 7622 13892
rect 8386 13880 8392 13892
rect 8444 13880 8450 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 7469 13855 7527 13861
rect 7469 13821 7481 13855
rect 7515 13821 7527 13855
rect 7469 13815 7527 13821
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 8496 13852 8524 13883
rect 8570 13880 8576 13932
rect 8628 13920 8634 13932
rect 8680 13920 8708 13960
rect 11146 13948 11152 14000
rect 11204 13988 11210 14000
rect 13541 13991 13599 13997
rect 13541 13988 13553 13991
rect 11204 13960 13553 13988
rect 11204 13948 11210 13960
rect 13541 13957 13553 13960
rect 13587 13988 13599 13991
rect 14369 13991 14427 13997
rect 14369 13988 14381 13991
rect 13587 13960 14381 13988
rect 13587 13957 13599 13960
rect 13541 13951 13599 13957
rect 14369 13957 14381 13960
rect 14415 13957 14427 13991
rect 14369 13951 14427 13957
rect 14642 13948 14648 14000
rect 14700 13988 14706 14000
rect 14700 13960 17172 13988
rect 14700 13948 14706 13960
rect 8628 13892 8708 13920
rect 8628 13880 8634 13892
rect 8665 13855 8723 13861
rect 8665 13852 8677 13855
rect 7708 13824 8524 13852
rect 8588 13824 8677 13852
rect 7708 13812 7714 13824
rect 3329 13787 3387 13793
rect 3329 13753 3341 13787
rect 3375 13784 3387 13787
rect 3786 13784 3792 13796
rect 3375 13756 3792 13784
rect 3375 13753 3387 13756
rect 3329 13747 3387 13753
rect 3786 13744 3792 13756
rect 3844 13744 3850 13796
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 6604 13756 7512 13784
rect 6604 13744 6610 13756
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4230 13719 4288 13725
rect 4230 13716 4242 13719
rect 4028 13688 4242 13716
rect 4028 13676 4034 13688
rect 4230 13685 4242 13688
rect 4276 13685 4288 13719
rect 4230 13679 4288 13685
rect 4706 13676 4712 13728
rect 4764 13716 4770 13728
rect 5350 13716 5356 13728
rect 4764 13688 5356 13716
rect 4764 13676 4770 13688
rect 5350 13676 5356 13688
rect 5408 13716 5414 13728
rect 6270 13716 6276 13728
rect 5408 13688 6276 13716
rect 5408 13676 5414 13688
rect 6270 13676 6276 13688
rect 6328 13676 6334 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 6917 13719 6975 13725
rect 6917 13716 6929 13719
rect 6696 13688 6929 13716
rect 6696 13676 6702 13688
rect 6917 13685 6929 13688
rect 6963 13685 6975 13719
rect 7484 13716 7512 13756
rect 8588 13716 8616 13824
rect 8665 13821 8677 13824
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 9306 13812 9312 13864
rect 9364 13812 9370 13864
rect 10134 13812 10140 13864
rect 10192 13852 10198 13864
rect 10704 13852 10732 13906
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 11793 13923 11851 13929
rect 11793 13920 11805 13923
rect 11296 13892 11805 13920
rect 11296 13880 11302 13892
rect 11793 13889 11805 13892
rect 11839 13920 11851 13923
rect 12529 13923 12587 13929
rect 11839 13892 12480 13920
rect 11839 13889 11851 13892
rect 11793 13883 11851 13889
rect 12452 13852 12480 13892
rect 12529 13889 12541 13923
rect 12575 13920 12587 13923
rect 13265 13923 13323 13929
rect 13265 13920 13277 13923
rect 12575 13892 13277 13920
rect 12575 13889 12587 13892
rect 12529 13883 12587 13889
rect 13265 13889 13277 13892
rect 13311 13920 13323 13923
rect 13630 13920 13636 13932
rect 13311 13892 13636 13920
rect 13311 13889 13323 13892
rect 13265 13883 13323 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13832 13892 14289 13920
rect 12621 13855 12679 13861
rect 12621 13852 12633 13855
rect 10192 13824 10640 13852
rect 10704 13824 11652 13852
rect 12452 13824 12633 13852
rect 10192 13812 10198 13824
rect 10612 13784 10640 13824
rect 10962 13784 10968 13796
rect 10612 13756 10968 13784
rect 10962 13744 10968 13756
rect 11020 13744 11026 13796
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11517 13787 11575 13793
rect 11517 13784 11529 13787
rect 11388 13756 11529 13784
rect 11388 13744 11394 13756
rect 11517 13753 11529 13756
rect 11563 13753 11575 13787
rect 11624 13784 11652 13824
rect 12621 13821 12633 13824
rect 12667 13821 12679 13855
rect 12621 13815 12679 13821
rect 12805 13855 12863 13861
rect 12805 13821 12817 13855
rect 12851 13852 12863 13855
rect 12894 13852 12900 13864
rect 12851 13824 12900 13852
rect 12851 13821 12863 13824
rect 12805 13815 12863 13821
rect 12526 13784 12532 13796
rect 11624 13756 12532 13784
rect 11517 13747 11575 13753
rect 12526 13744 12532 13756
rect 12584 13744 12590 13796
rect 12636 13784 12664 13815
rect 12894 13812 12900 13824
rect 12952 13852 12958 13864
rect 13357 13855 13415 13861
rect 13357 13852 13369 13855
rect 12952 13824 13369 13852
rect 12952 13812 12958 13824
rect 13357 13821 13369 13824
rect 13403 13821 13415 13855
rect 13357 13815 13415 13821
rect 13262 13784 13268 13796
rect 12636 13756 13268 13784
rect 13262 13744 13268 13756
rect 13320 13744 13326 13796
rect 13832 13784 13860 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14918 13920 14924 13932
rect 14277 13883 14335 13889
rect 14476 13892 14924 13920
rect 14476 13852 14504 13892
rect 14918 13880 14924 13892
rect 14976 13880 14982 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 15657 13923 15715 13929
rect 15657 13889 15669 13923
rect 15703 13920 15715 13923
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15703 13892 16221 13920
rect 15703 13889 15715 13892
rect 15657 13883 15715 13889
rect 16209 13889 16221 13892
rect 16255 13920 16267 13923
rect 17034 13920 17040 13932
rect 16255 13892 17040 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 17034 13880 17040 13892
rect 17092 13880 17098 13932
rect 17144 13929 17172 13960
rect 17310 13948 17316 14000
rect 17368 13988 17374 14000
rect 17405 13991 17463 13997
rect 17405 13988 17417 13991
rect 17368 13960 17417 13988
rect 17368 13948 17374 13960
rect 17405 13957 17417 13960
rect 17451 13957 17463 13991
rect 17405 13951 17463 13957
rect 17678 13948 17684 14000
rect 17736 13988 17742 14000
rect 20622 13988 20628 14000
rect 17736 13960 17894 13988
rect 18708 13960 20628 13988
rect 17736 13948 17742 13960
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 13924 13824 14504 13852
rect 14553 13855 14611 13861
rect 13924 13793 13952 13824
rect 14553 13821 14565 13855
rect 14599 13852 14611 13855
rect 15010 13852 15016 13864
rect 14599 13824 15016 13852
rect 14599 13821 14611 13824
rect 14553 13815 14611 13821
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 15212 13793 15240 13880
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16390 13852 16396 13864
rect 15804 13824 16396 13852
rect 15804 13812 15810 13824
rect 16390 13812 16396 13824
rect 16448 13812 16454 13864
rect 18708 13852 18736 13960
rect 20622 13948 20628 13960
rect 20680 13948 20686 14000
rect 22554 13948 22560 14000
rect 22612 13988 22618 14000
rect 24946 13988 24952 14000
rect 22612 13960 24952 13988
rect 22612 13948 22618 13960
rect 24946 13948 24952 13960
rect 25004 13948 25010 14000
rect 29181 13991 29239 13997
rect 29181 13988 29193 13991
rect 25608 13960 29193 13988
rect 21082 13880 21088 13932
rect 21140 13880 21146 13932
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13920 21235 13923
rect 21450 13920 21456 13932
rect 21223 13892 21456 13920
rect 21223 13889 21235 13892
rect 21177 13883 21235 13889
rect 21450 13880 21456 13892
rect 21508 13880 21514 13932
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 24305 13923 24363 13929
rect 24305 13920 24317 13923
rect 21968 13892 24317 13920
rect 21968 13880 21974 13892
rect 24305 13889 24317 13892
rect 24351 13920 24363 13923
rect 24351 13892 24532 13920
rect 24351 13889 24363 13892
rect 24305 13883 24363 13889
rect 16500 13824 18736 13852
rect 13740 13756 13860 13784
rect 13909 13787 13967 13793
rect 7484 13688 8616 13716
rect 9572 13719 9630 13725
rect 6917 13679 6975 13685
rect 9572 13685 9584 13719
rect 9618 13716 9630 13719
rect 10134 13716 10140 13728
rect 9618 13688 10140 13716
rect 9618 13685 9630 13688
rect 9572 13679 9630 13685
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 10594 13676 10600 13728
rect 10652 13716 10658 13728
rect 11054 13716 11060 13728
rect 10652 13688 11060 13716
rect 10652 13676 10658 13688
rect 11054 13676 11060 13688
rect 11112 13676 11118 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 11882 13716 11888 13728
rect 11664 13688 11888 13716
rect 11664 13676 11670 13688
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12066 13676 12072 13728
rect 12124 13716 12130 13728
rect 13078 13716 13084 13728
rect 12124 13688 13084 13716
rect 12124 13676 12130 13688
rect 13078 13676 13084 13688
rect 13136 13676 13142 13728
rect 13630 13676 13636 13728
rect 13688 13716 13694 13728
rect 13740 13725 13768 13756
rect 13909 13753 13921 13787
rect 13955 13753 13967 13787
rect 13909 13747 13967 13753
rect 15197 13787 15255 13793
rect 15197 13753 15209 13787
rect 15243 13753 15255 13787
rect 15197 13747 15255 13753
rect 15562 13744 15568 13796
rect 15620 13784 15626 13796
rect 16500 13784 16528 13824
rect 18874 13812 18880 13864
rect 18932 13812 18938 13864
rect 19518 13812 19524 13864
rect 19576 13852 19582 13864
rect 19978 13852 19984 13864
rect 19576 13824 19984 13852
rect 19576 13812 19582 13824
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 20070 13812 20076 13864
rect 20128 13812 20134 13864
rect 21269 13855 21327 13861
rect 21269 13821 21281 13855
rect 21315 13821 21327 13855
rect 22281 13855 22339 13861
rect 22281 13852 22293 13855
rect 21269 13815 21327 13821
rect 21928 13824 22293 13852
rect 15620 13756 16528 13784
rect 15620 13744 15626 13756
rect 18598 13744 18604 13796
rect 18656 13784 18662 13796
rect 20254 13784 20260 13796
rect 18656 13756 20260 13784
rect 18656 13744 18662 13756
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 20806 13744 20812 13796
rect 20864 13784 20870 13796
rect 21284 13784 21312 13815
rect 20864 13756 21312 13784
rect 20864 13744 20870 13756
rect 13725 13719 13783 13725
rect 13725 13716 13737 13719
rect 13688 13688 13737 13716
rect 13688 13676 13694 13688
rect 13725 13685 13737 13688
rect 13771 13685 13783 13719
rect 13725 13679 13783 13685
rect 14090 13676 14096 13728
rect 14148 13716 14154 13728
rect 18138 13716 18144 13728
rect 14148 13688 18144 13716
rect 14148 13676 14154 13688
rect 18138 13676 18144 13688
rect 18196 13676 18202 13728
rect 18690 13676 18696 13728
rect 18748 13716 18754 13728
rect 19245 13719 19303 13725
rect 19245 13716 19257 13719
rect 18748 13688 19257 13716
rect 18748 13676 18754 13688
rect 19245 13685 19257 13688
rect 19291 13716 19303 13719
rect 21928 13716 21956 13824
rect 22281 13821 22293 13824
rect 22327 13852 22339 13855
rect 23106 13852 23112 13864
rect 22327 13824 23112 13852
rect 22327 13821 22339 13824
rect 22281 13815 22339 13821
rect 23106 13812 23112 13824
rect 23164 13812 23170 13864
rect 23201 13855 23259 13861
rect 23201 13821 23213 13855
rect 23247 13821 23259 13855
rect 23201 13815 23259 13821
rect 22002 13744 22008 13796
rect 22060 13784 22066 13796
rect 22738 13784 22744 13796
rect 22060 13756 22744 13784
rect 22060 13744 22066 13756
rect 22738 13744 22744 13756
rect 22796 13784 22802 13796
rect 23216 13784 23244 13815
rect 23934 13812 23940 13864
rect 23992 13852 23998 13864
rect 24397 13855 24455 13861
rect 24397 13852 24409 13855
rect 23992 13824 24409 13852
rect 23992 13812 23998 13824
rect 24397 13821 24409 13824
rect 24443 13821 24455 13855
rect 24504 13852 24532 13892
rect 24578 13880 24584 13932
rect 24636 13920 24642 13932
rect 25608 13920 25636 13960
rect 29181 13957 29193 13960
rect 29227 13957 29239 13991
rect 29181 13951 29239 13957
rect 26602 13920 26608 13932
rect 24636 13892 25636 13920
rect 26252 13892 26608 13920
rect 24636 13880 24642 13892
rect 24762 13852 24768 13864
rect 24504 13824 24768 13852
rect 24397 13815 24455 13821
rect 24762 13812 24768 13824
rect 24820 13812 24826 13864
rect 24854 13812 24860 13864
rect 24912 13852 24918 13864
rect 25590 13852 25596 13864
rect 24912 13824 25596 13852
rect 24912 13812 24918 13824
rect 25590 13812 25596 13824
rect 25648 13812 25654 13864
rect 25777 13855 25835 13861
rect 25777 13821 25789 13855
rect 25823 13852 25835 13855
rect 26252 13852 26280 13892
rect 26602 13880 26608 13892
rect 26660 13920 26666 13932
rect 27157 13923 27215 13929
rect 27157 13920 27169 13923
rect 26660 13892 27169 13920
rect 26660 13880 26666 13892
rect 27157 13889 27169 13892
rect 27203 13889 27215 13923
rect 27157 13883 27215 13889
rect 28534 13880 28540 13932
rect 28592 13880 28598 13932
rect 29822 13880 29828 13932
rect 29880 13880 29886 13932
rect 29932 13852 29960 14028
rect 30285 14025 30297 14028
rect 30331 14025 30343 14059
rect 30285 14019 30343 14025
rect 40034 13948 40040 14000
rect 40092 13988 40098 14000
rect 42794 13988 42800 14000
rect 40092 13960 42800 13988
rect 40092 13948 40098 13960
rect 42794 13948 42800 13960
rect 42852 13948 42858 14000
rect 30466 13880 30472 13932
rect 30524 13920 30530 13932
rect 30745 13923 30803 13929
rect 30745 13920 30757 13923
rect 30524 13892 30757 13920
rect 30524 13880 30530 13892
rect 30745 13889 30757 13892
rect 30791 13889 30803 13923
rect 30745 13883 30803 13889
rect 25823 13824 26280 13852
rect 26344 13824 29960 13852
rect 25823 13821 25835 13824
rect 25777 13815 25835 13821
rect 22796 13756 23244 13784
rect 22796 13744 22802 13756
rect 23290 13744 23296 13796
rect 23348 13784 23354 13796
rect 25222 13784 25228 13796
rect 23348 13756 25228 13784
rect 23348 13744 23354 13756
rect 25222 13744 25228 13756
rect 25280 13744 25286 13796
rect 25958 13744 25964 13796
rect 26016 13784 26022 13796
rect 26344 13784 26372 13824
rect 26016 13756 26372 13784
rect 26016 13744 26022 13756
rect 28902 13744 28908 13796
rect 28960 13784 28966 13796
rect 36538 13784 36544 13796
rect 28960 13756 36544 13784
rect 28960 13744 28966 13756
rect 36538 13744 36544 13756
rect 36596 13744 36602 13796
rect 19291 13688 21956 13716
rect 19291 13685 19303 13688
rect 19245 13679 19303 13685
rect 22646 13676 22652 13728
rect 22704 13676 22710 13728
rect 22922 13676 22928 13728
rect 22980 13716 22986 13728
rect 23474 13716 23480 13728
rect 22980 13688 23480 13716
rect 22980 13676 22986 13688
rect 23474 13676 23480 13688
rect 23532 13676 23538 13728
rect 23750 13676 23756 13728
rect 23808 13716 23814 13728
rect 24026 13716 24032 13728
rect 23808 13688 24032 13716
rect 23808 13676 23814 13688
rect 24026 13676 24032 13688
rect 24084 13676 24090 13728
rect 24946 13676 24952 13728
rect 25004 13716 25010 13728
rect 25133 13719 25191 13725
rect 25133 13716 25145 13719
rect 25004 13688 25145 13716
rect 25004 13676 25010 13688
rect 25133 13685 25145 13688
rect 25179 13685 25191 13719
rect 25133 13679 25191 13685
rect 27798 13676 27804 13728
rect 27856 13676 27862 13728
rect 29914 13676 29920 13728
rect 29972 13716 29978 13728
rect 39666 13716 39672 13728
rect 29972 13688 39672 13716
rect 29972 13676 29978 13688
rect 39666 13676 39672 13688
rect 39724 13676 39730 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 3605 13515 3663 13521
rect 3605 13481 3617 13515
rect 3651 13512 3663 13515
rect 3786 13512 3792 13524
rect 3651 13484 3792 13512
rect 3651 13481 3663 13484
rect 3605 13475 3663 13481
rect 3786 13472 3792 13484
rect 3844 13472 3850 13524
rect 3973 13515 4031 13521
rect 3973 13481 3985 13515
rect 4019 13512 4031 13515
rect 4246 13512 4252 13524
rect 4019 13484 4252 13512
rect 4019 13481 4031 13484
rect 3973 13475 4031 13481
rect 4246 13472 4252 13484
rect 4304 13472 4310 13524
rect 4338 13472 4344 13524
rect 4396 13512 4402 13524
rect 6086 13512 6092 13524
rect 4396 13484 6092 13512
rect 4396 13472 4402 13484
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 6288 13484 8585 13512
rect 4433 13447 4491 13453
rect 4433 13413 4445 13447
rect 4479 13444 4491 13447
rect 5166 13444 5172 13456
rect 4479 13416 5172 13444
rect 4479 13413 4491 13416
rect 4433 13407 4491 13413
rect 5166 13404 5172 13416
rect 5224 13404 5230 13456
rect 6288 13388 6316 13484
rect 8573 13481 8585 13484
rect 8619 13512 8631 13515
rect 8619 13484 10824 13512
rect 8619 13481 8631 13484
rect 8573 13475 8631 13481
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13444 9183 13447
rect 9950 13444 9956 13456
rect 9171 13416 9956 13444
rect 9171 13413 9183 13416
rect 9125 13407 9183 13413
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 2038 13336 2044 13388
rect 2096 13336 2102 13388
rect 3418 13336 3424 13388
rect 3476 13376 3482 13388
rect 3878 13376 3884 13388
rect 3476 13348 3884 13376
rect 3476 13336 3482 13348
rect 3878 13336 3884 13348
rect 3936 13376 3942 13388
rect 4893 13379 4951 13385
rect 4893 13376 4905 13379
rect 3936 13348 4905 13376
rect 3936 13336 3942 13348
rect 4893 13345 4905 13348
rect 4939 13345 4951 13379
rect 4893 13339 4951 13345
rect 4982 13336 4988 13388
rect 5040 13336 5046 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5316 13348 6101 13376
rect 5316 13336 5322 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 6270 13336 6276 13388
rect 6328 13336 6334 13388
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 9272 13348 9781 13376
rect 9272 13336 9278 13348
rect 9769 13345 9781 13348
rect 9815 13376 9827 13379
rect 10594 13376 10600 13388
rect 9815 13348 10600 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 10594 13336 10600 13348
rect 10652 13336 10658 13388
rect 10796 13376 10824 13484
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 12710 13512 12716 13524
rect 11664 13484 12716 13512
rect 11664 13472 11670 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 14292 13484 15608 13512
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 14292 13444 14320 13484
rect 13320 13416 14320 13444
rect 15580 13444 15608 13484
rect 16298 13472 16304 13524
rect 16356 13472 16362 13524
rect 16482 13472 16488 13524
rect 16540 13472 16546 13524
rect 16666 13472 16672 13524
rect 16724 13512 16730 13524
rect 16945 13515 17003 13521
rect 16945 13512 16957 13515
rect 16724 13484 16957 13512
rect 16724 13472 16730 13484
rect 16945 13481 16957 13484
rect 16991 13512 17003 13515
rect 17034 13512 17040 13524
rect 16991 13484 17040 13512
rect 16991 13481 17003 13484
rect 16945 13475 17003 13481
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 17310 13472 17316 13524
rect 17368 13512 17374 13524
rect 17368 13484 19012 13512
rect 17368 13472 17374 13484
rect 16758 13444 16764 13456
rect 15580 13416 16764 13444
rect 13320 13404 13326 13416
rect 16758 13404 16764 13416
rect 16816 13404 16822 13456
rect 18141 13447 18199 13453
rect 18141 13413 18153 13447
rect 18187 13413 18199 13447
rect 18141 13407 18199 13413
rect 10873 13379 10931 13385
rect 10873 13376 10885 13379
rect 10796 13348 10885 13376
rect 10873 13345 10885 13348
rect 10919 13345 10931 13379
rect 10873 13339 10931 13345
rect 11790 13336 11796 13388
rect 11848 13376 11854 13388
rect 11885 13379 11943 13385
rect 11885 13376 11897 13379
rect 11848 13348 11897 13376
rect 11848 13336 11854 13348
rect 11885 13345 11897 13348
rect 11931 13376 11943 13379
rect 12250 13376 12256 13388
rect 11931 13348 12256 13376
rect 11931 13345 11943 13348
rect 11885 13339 11943 13345
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 12308 13348 14289 13376
rect 12308 13336 12314 13348
rect 14277 13345 14289 13348
rect 14323 13376 14335 13379
rect 14642 13376 14648 13388
rect 14323 13348 14648 13376
rect 14323 13345 14335 13348
rect 14277 13339 14335 13345
rect 14642 13336 14648 13348
rect 14700 13376 14706 13388
rect 14918 13376 14924 13388
rect 14700 13348 14924 13376
rect 14700 13336 14706 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 15010 13336 15016 13388
rect 15068 13376 15074 13388
rect 16666 13376 16672 13388
rect 15068 13348 16672 13376
rect 15068 13336 15074 13348
rect 16666 13336 16672 13348
rect 16724 13336 16730 13388
rect 16850 13336 16856 13388
rect 16908 13376 16914 13388
rect 17405 13379 17463 13385
rect 17405 13376 17417 13379
rect 16908 13348 17417 13376
rect 16908 13336 16914 13348
rect 17405 13345 17417 13348
rect 17451 13345 17463 13379
rect 17405 13339 17463 13345
rect 17586 13336 17592 13388
rect 17644 13336 17650 13388
rect 566 13268 572 13320
rect 624 13308 630 13320
rect 1578 13308 1584 13320
rect 624 13280 1584 13308
rect 624 13268 630 13280
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 3234 13268 3240 13320
rect 3292 13308 3298 13320
rect 4065 13311 4123 13317
rect 4065 13308 4077 13311
rect 3292 13280 4077 13308
rect 3292 13268 3298 13280
rect 4065 13277 4077 13280
rect 4111 13277 4123 13311
rect 4065 13271 4123 13277
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 4212 13280 6837 13308
rect 4212 13268 4218 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 9490 13268 9496 13320
rect 9548 13268 9554 13320
rect 9585 13311 9643 13317
rect 9585 13277 9597 13311
rect 9631 13308 9643 13311
rect 10042 13308 10048 13320
rect 9631 13280 10048 13308
rect 9631 13277 9643 13280
rect 9585 13271 9643 13277
rect 10042 13268 10048 13280
rect 10100 13268 10106 13320
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13308 10747 13311
rect 11514 13308 11520 13320
rect 10735 13280 11520 13308
rect 10735 13277 10747 13280
rect 10689 13271 10747 13277
rect 11514 13268 11520 13280
rect 11572 13268 11578 13320
rect 15654 13268 15660 13320
rect 15712 13268 15718 13320
rect 17310 13308 17316 13320
rect 15948 13280 17316 13308
rect 382 13200 388 13252
rect 440 13240 446 13252
rect 4801 13243 4859 13249
rect 440 13212 3740 13240
rect 440 13200 446 13212
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 1946 13172 1952 13184
rect 1820 13144 1952 13172
rect 1820 13132 1826 13144
rect 1946 13132 1952 13144
rect 2004 13172 2010 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 2004 13144 3433 13172
rect 2004 13132 2010 13144
rect 3421 13141 3433 13144
rect 3467 13172 3479 13175
rect 3510 13172 3516 13184
rect 3467 13144 3516 13172
rect 3467 13141 3479 13144
rect 3421 13135 3479 13141
rect 3510 13132 3516 13144
rect 3568 13132 3574 13184
rect 3712 13172 3740 13212
rect 4801 13209 4813 13243
rect 4847 13240 4859 13243
rect 5074 13240 5080 13252
rect 4847 13212 5080 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5997 13243 6055 13249
rect 5997 13209 6009 13243
rect 6043 13240 6055 13243
rect 6638 13240 6644 13252
rect 6043 13212 6644 13240
rect 6043 13209 6055 13212
rect 5997 13203 6055 13209
rect 6638 13200 6644 13212
rect 6696 13200 6702 13252
rect 7006 13200 7012 13252
rect 7064 13240 7070 13252
rect 7101 13243 7159 13249
rect 7101 13240 7113 13243
rect 7064 13212 7113 13240
rect 7064 13200 7070 13212
rect 7101 13209 7113 13212
rect 7147 13209 7159 13243
rect 7101 13203 7159 13209
rect 7650 13200 7656 13252
rect 7708 13200 7714 13252
rect 9508 13240 9536 13268
rect 10781 13243 10839 13249
rect 10781 13240 10793 13243
rect 9508 13212 10793 13240
rect 10781 13209 10793 13212
rect 10827 13209 10839 13243
rect 10781 13203 10839 13209
rect 10870 13200 10876 13252
rect 10928 13240 10934 13252
rect 11609 13243 11667 13249
rect 11609 13240 11621 13243
rect 10928 13212 11621 13240
rect 10928 13200 10934 13212
rect 11609 13209 11621 13212
rect 11655 13209 11667 13243
rect 11609 13203 11667 13209
rect 11882 13200 11888 13252
rect 11940 13240 11946 13252
rect 12066 13240 12072 13252
rect 11940 13212 12072 13240
rect 11940 13200 11946 13212
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 12161 13243 12219 13249
rect 12161 13209 12173 13243
rect 12207 13240 12219 13243
rect 12207 13212 12434 13240
rect 12207 13209 12219 13212
rect 12161 13203 12219 13209
rect 5442 13172 5448 13184
rect 3712 13144 5448 13172
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 7742 13172 7748 13184
rect 5675 13144 7748 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 10042 13132 10048 13184
rect 10100 13172 10106 13184
rect 10321 13175 10379 13181
rect 10321 13172 10333 13175
rect 10100 13144 10333 13172
rect 10100 13132 10106 13144
rect 10321 13141 10333 13144
rect 10367 13141 10379 13175
rect 10321 13135 10379 13141
rect 10410 13132 10416 13184
rect 10468 13172 10474 13184
rect 11333 13175 11391 13181
rect 11333 13172 11345 13175
rect 10468 13144 11345 13172
rect 10468 13132 10474 13144
rect 11333 13141 11345 13144
rect 11379 13141 11391 13175
rect 12406 13172 12434 13212
rect 12618 13200 12624 13252
rect 12676 13200 12682 13252
rect 14553 13243 14611 13249
rect 14553 13209 14565 13243
rect 14599 13240 14611 13243
rect 14642 13240 14648 13252
rect 14599 13212 14648 13240
rect 14599 13209 14611 13212
rect 14553 13203 14611 13209
rect 14642 13200 14648 13212
rect 14700 13200 14706 13252
rect 12526 13172 12532 13184
rect 12406 13144 12532 13172
rect 11333 13135 11391 13141
rect 12526 13132 12532 13144
rect 12584 13132 12590 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 13136 13144 13645 13172
rect 13136 13132 13142 13144
rect 13633 13141 13645 13144
rect 13679 13172 13691 13175
rect 13998 13172 14004 13184
rect 13679 13144 14004 13172
rect 13679 13141 13691 13144
rect 13633 13135 13691 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14458 13132 14464 13184
rect 14516 13172 14522 13184
rect 15948 13172 15976 13280
rect 17310 13268 17316 13280
rect 17368 13268 17374 13320
rect 17770 13268 17776 13320
rect 17828 13308 17834 13320
rect 18156 13308 18184 13407
rect 18506 13404 18512 13456
rect 18564 13444 18570 13456
rect 18564 13416 18828 13444
rect 18564 13404 18570 13416
rect 18230 13336 18236 13388
rect 18288 13376 18294 13388
rect 18601 13379 18659 13385
rect 18288 13348 18460 13376
rect 18288 13336 18294 13348
rect 17828 13280 18184 13308
rect 18432 13304 18460 13348
rect 18601 13345 18613 13379
rect 18647 13376 18659 13379
rect 18690 13376 18696 13388
rect 18647 13348 18696 13376
rect 18647 13345 18659 13348
rect 18601 13339 18659 13345
rect 18690 13336 18696 13348
rect 18748 13336 18754 13388
rect 18800 13385 18828 13416
rect 18785 13379 18843 13385
rect 18785 13345 18797 13379
rect 18831 13345 18843 13379
rect 18984 13376 19012 13484
rect 19150 13472 19156 13524
rect 19208 13512 19214 13524
rect 21910 13512 21916 13524
rect 19208 13484 21916 13512
rect 19208 13472 19214 13484
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 23845 13515 23903 13521
rect 23845 13481 23857 13515
rect 23891 13512 23903 13515
rect 30834 13512 30840 13524
rect 23891 13484 30840 13512
rect 23891 13481 23903 13484
rect 23845 13475 23903 13481
rect 30834 13472 30840 13484
rect 30892 13472 30898 13524
rect 42702 13512 42708 13524
rect 31726 13484 42708 13512
rect 19337 13447 19395 13453
rect 19337 13413 19349 13447
rect 19383 13444 19395 13447
rect 19383 13416 20392 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 19150 13376 19156 13388
rect 18984 13348 19156 13376
rect 18785 13339 18843 13345
rect 19150 13336 19156 13348
rect 19208 13336 19214 13388
rect 18509 13311 18567 13317
rect 18509 13304 18521 13311
rect 17828 13268 17834 13280
rect 18432 13277 18521 13304
rect 18555 13308 18567 13311
rect 19352 13308 19380 13407
rect 19610 13336 19616 13388
rect 19668 13336 19674 13388
rect 20364 13376 20392 13416
rect 21542 13404 21548 13456
rect 21600 13444 21606 13456
rect 22554 13444 22560 13456
rect 21600 13416 22560 13444
rect 21600 13404 21606 13416
rect 22554 13404 22560 13416
rect 22612 13404 22618 13456
rect 26050 13444 26056 13456
rect 22756 13416 26056 13444
rect 20530 13376 20536 13388
rect 20364 13348 20536 13376
rect 20530 13336 20536 13348
rect 20588 13336 20594 13388
rect 22005 13379 22063 13385
rect 22005 13345 22017 13379
rect 22051 13376 22063 13379
rect 22094 13376 22100 13388
rect 22051 13348 22100 13376
rect 22051 13345 22063 13348
rect 22005 13339 22063 13345
rect 22094 13336 22100 13348
rect 22152 13336 22158 13388
rect 18555 13280 19380 13308
rect 18555 13277 18567 13280
rect 18432 13276 18567 13277
rect 18509 13271 18567 13276
rect 19702 13268 19708 13320
rect 19760 13308 19766 13320
rect 20257 13311 20315 13317
rect 20257 13308 20269 13311
rect 19760 13280 20269 13308
rect 19760 13268 19766 13280
rect 20257 13277 20269 13280
rect 20303 13277 20315 13311
rect 20257 13271 20315 13277
rect 22186 13268 22192 13320
rect 22244 13308 22250 13320
rect 22465 13311 22523 13317
rect 22465 13308 22477 13311
rect 22244 13280 22477 13308
rect 22244 13268 22250 13280
rect 22465 13277 22477 13280
rect 22511 13277 22523 13311
rect 22465 13271 22523 13277
rect 16482 13200 16488 13252
rect 16540 13200 16546 13252
rect 16574 13200 16580 13252
rect 16632 13240 16638 13252
rect 18690 13240 18696 13252
rect 16632 13212 18696 13240
rect 16632 13200 16638 13212
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 19334 13200 19340 13252
rect 19392 13200 19398 13252
rect 20530 13200 20536 13252
rect 20588 13200 20594 13252
rect 20990 13200 20996 13252
rect 21048 13200 21054 13252
rect 14516 13144 15976 13172
rect 14516 13132 14522 13144
rect 16022 13132 16028 13184
rect 16080 13132 16086 13184
rect 16500 13172 16528 13200
rect 17313 13175 17371 13181
rect 17313 13172 17325 13175
rect 16500 13144 17325 13172
rect 17313 13141 17325 13144
rect 17359 13141 17371 13175
rect 17313 13135 17371 13141
rect 17862 13132 17868 13184
rect 17920 13172 17926 13184
rect 19352 13172 19380 13200
rect 17920 13144 19380 13172
rect 17920 13132 17926 13144
rect 19518 13132 19524 13184
rect 19576 13172 19582 13184
rect 22756 13172 22784 13416
rect 26050 13404 26056 13416
rect 26108 13404 26114 13456
rect 29641 13447 29699 13453
rect 29641 13413 29653 13447
rect 29687 13444 29699 13447
rect 29730 13444 29736 13456
rect 29687 13416 29736 13444
rect 29687 13413 29699 13416
rect 29641 13407 29699 13413
rect 29730 13404 29736 13416
rect 29788 13404 29794 13456
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 24118 13376 24124 13388
rect 23532 13348 24124 13376
rect 23532 13336 23538 13348
rect 24118 13336 24124 13348
rect 24176 13336 24182 13388
rect 24210 13336 24216 13388
rect 24268 13376 24274 13388
rect 24578 13376 24584 13388
rect 24268 13348 24584 13376
rect 24268 13336 24274 13348
rect 24578 13336 24584 13348
rect 24636 13336 24642 13388
rect 25130 13336 25136 13388
rect 25188 13336 25194 13388
rect 27798 13376 27804 13388
rect 25792 13348 27804 13376
rect 23106 13268 23112 13320
rect 23164 13308 23170 13320
rect 24029 13311 24087 13317
rect 24029 13308 24041 13311
rect 23164 13280 24041 13308
rect 23164 13268 23170 13280
rect 24029 13277 24041 13280
rect 24075 13277 24087 13311
rect 24029 13271 24087 13277
rect 24946 13268 24952 13320
rect 25004 13268 25010 13320
rect 25792 13317 25820 13348
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 28626 13336 28632 13388
rect 28684 13376 28690 13388
rect 31726 13376 31754 13484
rect 42702 13472 42708 13484
rect 42760 13472 42766 13524
rect 28684 13348 31754 13376
rect 28684 13336 28690 13348
rect 25777 13311 25835 13317
rect 25777 13277 25789 13311
rect 25823 13277 25835 13311
rect 25777 13271 25835 13277
rect 26694 13268 26700 13320
rect 26752 13308 26758 13320
rect 27157 13311 27215 13317
rect 27157 13308 27169 13311
rect 26752 13280 27169 13308
rect 26752 13268 26758 13280
rect 27157 13277 27169 13280
rect 27203 13277 27215 13311
rect 27157 13271 27215 13277
rect 28261 13311 28319 13317
rect 28261 13277 28273 13311
rect 28307 13308 28319 13311
rect 37550 13308 37556 13320
rect 28307 13280 37556 13308
rect 28307 13277 28319 13280
rect 28261 13271 28319 13277
rect 37550 13268 37556 13280
rect 37608 13268 37614 13320
rect 22830 13200 22836 13252
rect 22888 13240 22894 13252
rect 23201 13243 23259 13249
rect 23201 13240 23213 13243
rect 22888 13212 23213 13240
rect 22888 13200 22894 13212
rect 23201 13209 23213 13212
rect 23247 13209 23259 13243
rect 23201 13203 23259 13209
rect 23290 13200 23296 13252
rect 23348 13240 23354 13252
rect 27801 13243 27859 13249
rect 27801 13240 27813 13243
rect 23348 13212 27813 13240
rect 23348 13200 23354 13212
rect 27801 13209 27813 13212
rect 27847 13209 27859 13243
rect 27801 13203 27859 13209
rect 28902 13200 28908 13252
rect 28960 13200 28966 13252
rect 19576 13144 22784 13172
rect 19576 13132 19582 13144
rect 23474 13132 23480 13184
rect 23532 13172 23538 13184
rect 23658 13172 23664 13184
rect 23532 13144 23664 13172
rect 23532 13132 23538 13144
rect 23658 13132 23664 13144
rect 23716 13132 23722 13184
rect 24026 13132 24032 13184
rect 24084 13172 24090 13184
rect 24581 13175 24639 13181
rect 24581 13172 24593 13175
rect 24084 13144 24593 13172
rect 24084 13132 24090 13144
rect 24581 13141 24593 13144
rect 24627 13141 24639 13175
rect 24581 13135 24639 13141
rect 25041 13175 25099 13181
rect 25041 13141 25053 13175
rect 25087 13172 25099 13175
rect 26142 13172 26148 13184
rect 25087 13144 26148 13172
rect 25087 13141 25099 13144
rect 25041 13135 25099 13141
rect 26142 13132 26148 13144
rect 26200 13132 26206 13184
rect 26234 13132 26240 13184
rect 26292 13172 26298 13184
rect 26421 13175 26479 13181
rect 26421 13172 26433 13175
rect 26292 13144 26433 13172
rect 26292 13132 26298 13144
rect 26421 13141 26433 13144
rect 26467 13141 26479 13175
rect 26421 13135 26479 13141
rect 26510 13132 26516 13184
rect 26568 13172 26574 13184
rect 26697 13175 26755 13181
rect 26697 13172 26709 13175
rect 26568 13144 26709 13172
rect 26568 13132 26574 13144
rect 26697 13141 26709 13144
rect 26743 13141 26755 13175
rect 26697 13135 26755 13141
rect 27706 13132 27712 13184
rect 27764 13172 27770 13184
rect 27890 13172 27896 13184
rect 27764 13144 27896 13172
rect 27764 13132 27770 13144
rect 27890 13132 27896 13144
rect 27948 13132 27954 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 2961 12971 3019 12977
rect 2961 12937 2973 12971
rect 3007 12968 3019 12971
rect 3694 12968 3700 12980
rect 3007 12940 3700 12968
rect 3007 12937 3019 12940
rect 2961 12931 3019 12937
rect 3694 12928 3700 12940
rect 3752 12928 3758 12980
rect 4154 12928 4160 12980
rect 4212 12968 4218 12980
rect 4798 12968 4804 12980
rect 4212 12940 4804 12968
rect 4212 12928 4218 12940
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 5258 12928 5264 12980
rect 5316 12968 5322 12980
rect 5718 12968 5724 12980
rect 5316 12940 5724 12968
rect 5316 12928 5322 12940
rect 5718 12928 5724 12940
rect 5776 12968 5782 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5776 12940 5917 12968
rect 5776 12928 5782 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 6822 12928 6828 12980
rect 6880 12968 6886 12980
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 6880 12940 10885 12968
rect 6880 12928 6886 12940
rect 10873 12937 10885 12940
rect 10919 12968 10931 12971
rect 11790 12968 11796 12980
rect 10919 12940 11796 12968
rect 10919 12937 10931 12940
rect 10873 12931 10931 12937
rect 11790 12928 11796 12940
rect 11848 12928 11854 12980
rect 11974 12928 11980 12980
rect 12032 12928 12038 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12437 12971 12495 12977
rect 12437 12968 12449 12971
rect 12124 12940 12449 12968
rect 12124 12928 12130 12940
rect 12437 12937 12449 12940
rect 12483 12968 12495 12971
rect 13633 12971 13691 12977
rect 12483 12940 13584 12968
rect 12483 12937 12495 12940
rect 12437 12931 12495 12937
rect 3234 12900 3240 12912
rect 1872 12872 3240 12900
rect 1872 12841 1900 12872
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 4430 12860 4436 12912
rect 4488 12860 4494 12912
rect 6178 12900 6184 12912
rect 5658 12872 6184 12900
rect 6178 12860 6184 12872
rect 6236 12900 6242 12912
rect 7650 12900 7656 12912
rect 6236 12872 7656 12900
rect 6236 12860 6242 12872
rect 7650 12860 7656 12872
rect 7708 12900 7714 12912
rect 8018 12900 8024 12912
rect 7708 12872 8024 12900
rect 7708 12860 7714 12872
rect 8018 12860 8024 12872
rect 8076 12900 8082 12912
rect 8076 12872 8418 12900
rect 8076 12860 8082 12872
rect 9398 12860 9404 12912
rect 9456 12900 9462 12912
rect 9674 12900 9680 12912
rect 9456 12872 9680 12900
rect 9456 12860 9462 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 10045 12903 10103 12909
rect 10045 12869 10057 12903
rect 10091 12900 10103 12903
rect 10226 12900 10232 12912
rect 10091 12872 10232 12900
rect 10091 12869 10103 12872
rect 10045 12863 10103 12869
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10778 12860 10784 12912
rect 10836 12860 10842 12912
rect 11698 12860 11704 12912
rect 11756 12900 11762 12912
rect 13354 12900 13360 12912
rect 11756 12872 13360 12900
rect 11756 12860 11762 12872
rect 13354 12860 13360 12872
rect 13412 12860 13418 12912
rect 13556 12900 13584 12940
rect 13633 12937 13645 12971
rect 13679 12968 13691 12971
rect 16482 12968 16488 12980
rect 13679 12940 16488 12968
rect 13679 12937 13691 12940
rect 13633 12931 13691 12937
rect 16482 12928 16488 12940
rect 16540 12928 16546 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17681 12971 17739 12977
rect 17681 12968 17693 12971
rect 17000 12940 17693 12968
rect 17000 12928 17006 12940
rect 17681 12937 17693 12940
rect 17727 12937 17739 12971
rect 17681 12931 17739 12937
rect 17770 12928 17776 12980
rect 17828 12968 17834 12980
rect 17828 12940 18368 12968
rect 17828 12928 17834 12940
rect 14458 12900 14464 12912
rect 13556 12872 14464 12900
rect 14458 12860 14464 12872
rect 14516 12860 14522 12912
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 16669 12903 16727 12909
rect 16669 12900 16681 12903
rect 14884 12872 16681 12900
rect 14884 12860 14890 12872
rect 16669 12869 16681 12872
rect 16715 12869 16727 12903
rect 16669 12863 16727 12869
rect 16758 12860 16764 12912
rect 16816 12900 16822 12912
rect 18340 12900 18368 12940
rect 18874 12928 18880 12980
rect 18932 12968 18938 12980
rect 22186 12968 22192 12980
rect 18932 12940 22192 12968
rect 18932 12928 18938 12940
rect 22186 12928 22192 12940
rect 22244 12968 22250 12980
rect 22557 12971 22615 12977
rect 22557 12968 22569 12971
rect 22244 12940 22569 12968
rect 22244 12928 22250 12940
rect 22557 12937 22569 12940
rect 22603 12937 22615 12971
rect 22557 12931 22615 12937
rect 22940 12940 25912 12968
rect 19610 12900 19616 12912
rect 16816 12872 18276 12900
rect 18340 12872 19616 12900
rect 16816 12860 16822 12872
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 1857 12795 1915 12801
rect 2746 12804 3341 12832
rect 1118 12724 1124 12776
rect 1176 12764 1182 12776
rect 1581 12767 1639 12773
rect 1581 12764 1593 12767
rect 1176 12736 1593 12764
rect 1176 12724 1182 12736
rect 1581 12733 1593 12736
rect 1627 12733 1639 12767
rect 1581 12727 1639 12733
rect 1670 12724 1676 12776
rect 1728 12764 1734 12776
rect 2746 12764 2774 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3694 12832 3700 12844
rect 3329 12795 3387 12801
rect 3528 12804 3700 12832
rect 3528 12773 3556 12804
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 4154 12792 4160 12844
rect 4212 12792 4218 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6270 12832 6276 12844
rect 5776 12804 6276 12832
rect 5776 12792 5782 12804
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 6457 12835 6515 12841
rect 6457 12801 6469 12835
rect 6503 12832 6515 12835
rect 6546 12832 6552 12844
rect 6503 12804 6552 12832
rect 6503 12801 6515 12804
rect 6457 12795 6515 12801
rect 1728 12736 2774 12764
rect 3421 12767 3479 12773
rect 1728 12724 1734 12736
rect 3421 12733 3433 12767
rect 3467 12733 3479 12767
rect 3421 12727 3479 12733
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 3620 12736 5488 12764
rect 3326 12656 3332 12708
rect 3384 12696 3390 12708
rect 3436 12696 3464 12727
rect 3384 12668 3464 12696
rect 3384 12656 3390 12668
rect 3510 12588 3516 12640
rect 3568 12628 3574 12640
rect 3620 12628 3648 12736
rect 4062 12656 4068 12708
rect 4120 12696 4126 12708
rect 5460 12696 5488 12736
rect 6086 12724 6092 12776
rect 6144 12764 6150 12776
rect 6472 12764 6500 12795
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 7190 12792 7196 12844
rect 7248 12792 7254 12844
rect 10134 12792 10140 12844
rect 10192 12832 10198 12844
rect 11330 12832 11336 12844
rect 10192 12804 11336 12832
rect 10192 12792 10198 12804
rect 11330 12792 11336 12804
rect 11388 12792 11394 12844
rect 11514 12792 11520 12844
rect 11572 12832 11578 12844
rect 11609 12835 11667 12841
rect 11609 12832 11621 12835
rect 11572 12804 11621 12832
rect 11572 12792 11578 12804
rect 11609 12801 11621 12804
rect 11655 12832 11667 12835
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 11655 12804 12357 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 12345 12801 12357 12804
rect 12391 12832 12403 12835
rect 12391 12804 12664 12832
rect 12391 12801 12403 12804
rect 12345 12795 12403 12801
rect 6144 12736 6500 12764
rect 6144 12724 6150 12736
rect 7650 12724 7656 12776
rect 7708 12724 7714 12776
rect 7929 12767 7987 12773
rect 7929 12764 7941 12767
rect 7760 12736 7941 12764
rect 7760 12696 7788 12736
rect 7929 12733 7941 12736
rect 7975 12733 7987 12767
rect 7929 12727 7987 12733
rect 8938 12724 8944 12776
rect 8996 12764 9002 12776
rect 9677 12767 9735 12773
rect 9677 12764 9689 12767
rect 8996 12736 9689 12764
rect 8996 12724 9002 12736
rect 9677 12733 9689 12736
rect 9723 12733 9735 12767
rect 9677 12727 9735 12733
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10594 12764 10600 12776
rect 9916 12736 10600 12764
rect 9916 12724 9922 12736
rect 10594 12724 10600 12736
rect 10652 12724 10658 12776
rect 11054 12724 11060 12776
rect 11112 12724 11118 12776
rect 11698 12724 11704 12776
rect 11756 12764 11762 12776
rect 12529 12767 12587 12773
rect 12529 12764 12541 12767
rect 11756 12736 12541 12764
rect 11756 12724 11762 12736
rect 12529 12733 12541 12736
rect 12575 12733 12587 12767
rect 12636 12764 12664 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13541 12835 13599 12841
rect 13541 12832 13553 12835
rect 12768 12804 13553 12832
rect 12768 12792 12774 12804
rect 13541 12801 13553 12804
rect 13587 12801 13599 12835
rect 13541 12795 13599 12801
rect 14277 12835 14335 12841
rect 14277 12801 14289 12835
rect 14323 12832 14335 12835
rect 14737 12835 14795 12841
rect 14737 12832 14749 12835
rect 14323 12804 14749 12832
rect 14323 12801 14335 12804
rect 14277 12795 14335 12801
rect 14737 12801 14749 12804
rect 14783 12832 14795 12835
rect 15194 12832 15200 12844
rect 14783 12804 15200 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 15194 12792 15200 12804
rect 15252 12792 15258 12844
rect 15930 12792 15936 12844
rect 15988 12792 15994 12844
rect 16025 12835 16083 12841
rect 16025 12801 16037 12835
rect 16071 12832 16083 12835
rect 16071 12804 16443 12832
rect 16071 12801 16083 12804
rect 16025 12795 16083 12801
rect 13262 12764 13268 12776
rect 12636 12736 13268 12764
rect 12529 12727 12587 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13817 12767 13875 12773
rect 13817 12733 13829 12767
rect 13863 12764 13875 12767
rect 14550 12764 14556 12776
rect 13863 12736 14556 12764
rect 13863 12733 13875 12736
rect 13817 12727 13875 12733
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12764 15071 12767
rect 15059 12736 16068 12764
rect 15059 12733 15071 12736
rect 15013 12727 15071 12733
rect 4120 12668 4292 12696
rect 5460 12668 7788 12696
rect 4120 12656 4126 12668
rect 3568 12600 3648 12628
rect 3568 12588 3574 12600
rect 3878 12588 3884 12640
rect 3936 12628 3942 12640
rect 4154 12628 4160 12640
rect 3936 12600 4160 12628
rect 3936 12588 3942 12600
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 4264 12628 4292 12668
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 9640 12668 12296 12696
rect 9640 12656 9646 12668
rect 4614 12628 4620 12640
rect 4264 12600 4620 12628
rect 4614 12588 4620 12600
rect 4672 12588 4678 12640
rect 5166 12588 5172 12640
rect 5224 12628 5230 12640
rect 5626 12628 5632 12640
rect 5224 12600 5632 12628
rect 5224 12588 5230 12600
rect 5626 12588 5632 12600
rect 5684 12588 5690 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 9214 12628 9220 12640
rect 6604 12600 9220 12628
rect 6604 12588 6610 12600
rect 9214 12588 9220 12600
rect 9272 12588 9278 12640
rect 9950 12588 9956 12640
rect 10008 12628 10014 12640
rect 10134 12628 10140 12640
rect 10008 12600 10140 12628
rect 10008 12588 10014 12600
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10318 12588 10324 12640
rect 10376 12628 10382 12640
rect 10413 12631 10471 12637
rect 10413 12628 10425 12631
rect 10376 12600 10425 12628
rect 10376 12588 10382 12600
rect 10413 12597 10425 12600
rect 10459 12597 10471 12631
rect 10413 12591 10471 12597
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 11514 12628 11520 12640
rect 10744 12600 11520 12628
rect 10744 12588 10750 12600
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 12268 12628 12296 12668
rect 12618 12656 12624 12708
rect 12676 12696 12682 12708
rect 13078 12696 13084 12708
rect 12676 12668 13084 12696
rect 12676 12656 12682 12668
rect 13078 12656 13084 12668
rect 13136 12656 13142 12708
rect 13170 12656 13176 12708
rect 13228 12656 13234 12708
rect 13354 12656 13360 12708
rect 13412 12696 13418 12708
rect 15838 12696 15844 12708
rect 13412 12668 15844 12696
rect 13412 12656 13418 12668
rect 15838 12656 15844 12668
rect 15896 12656 15902 12708
rect 13814 12628 13820 12640
rect 12268 12600 13820 12628
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 14366 12588 14372 12640
rect 14424 12588 14430 12640
rect 15562 12588 15568 12640
rect 15620 12588 15626 12640
rect 16040 12628 16068 12736
rect 16206 12724 16212 12776
rect 16264 12724 16270 12776
rect 16415 12696 16443 12804
rect 17310 12792 17316 12844
rect 17368 12832 17374 12844
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 17368 12804 17601 12832
rect 17368 12792 17374 12804
rect 17589 12801 17601 12804
rect 17635 12832 17647 12835
rect 17635 12804 17816 12832
rect 17635 12801 17647 12804
rect 17589 12795 17647 12801
rect 16482 12724 16488 12776
rect 16540 12764 16546 12776
rect 16540 12736 17724 12764
rect 16540 12724 16546 12736
rect 17586 12696 17592 12708
rect 16415 12668 17592 12696
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 16482 12628 16488 12640
rect 16040 12600 16488 12628
rect 16482 12588 16488 12600
rect 16540 12588 16546 12640
rect 16942 12588 16948 12640
rect 17000 12628 17006 12640
rect 17221 12631 17279 12637
rect 17221 12628 17233 12631
rect 17000 12600 17233 12628
rect 17000 12588 17006 12600
rect 17221 12597 17233 12600
rect 17267 12597 17279 12631
rect 17696 12628 17724 12736
rect 17788 12696 17816 12804
rect 17862 12724 17868 12776
rect 17920 12724 17926 12776
rect 18248 12764 18276 12872
rect 19610 12860 19616 12872
rect 19668 12860 19674 12912
rect 21542 12900 21548 12912
rect 21206 12872 21548 12900
rect 21542 12860 21548 12872
rect 21600 12860 21606 12912
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12832 18475 12835
rect 18598 12832 18604 12844
rect 18463 12804 18604 12832
rect 18463 12801 18475 12804
rect 18417 12795 18475 12801
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18693 12835 18751 12841
rect 18693 12801 18705 12835
rect 18739 12832 18751 12835
rect 19518 12832 19524 12844
rect 18739 12804 19524 12832
rect 18739 12801 18751 12804
rect 18693 12795 18751 12801
rect 19518 12792 19524 12804
rect 19576 12792 19582 12844
rect 19702 12792 19708 12844
rect 19760 12792 19766 12844
rect 22002 12792 22008 12844
rect 22060 12832 22066 12844
rect 22097 12835 22155 12841
rect 22097 12832 22109 12835
rect 22060 12804 22109 12832
rect 22060 12792 22066 12804
rect 22097 12801 22109 12804
rect 22143 12801 22155 12835
rect 22097 12795 22155 12801
rect 19150 12764 19156 12776
rect 18248 12736 19156 12764
rect 19150 12724 19156 12736
rect 19208 12724 19214 12776
rect 19981 12767 20039 12773
rect 19981 12733 19993 12767
rect 20027 12764 20039 12767
rect 22370 12764 22376 12776
rect 20027 12736 22376 12764
rect 20027 12733 20039 12736
rect 19981 12727 20039 12733
rect 22370 12724 22376 12736
rect 22428 12724 22434 12776
rect 22940 12773 22968 12940
rect 23201 12903 23259 12909
rect 23201 12869 23213 12903
rect 23247 12900 23259 12903
rect 23290 12900 23296 12912
rect 23247 12872 23296 12900
rect 23247 12869 23259 12872
rect 23201 12863 23259 12869
rect 23290 12860 23296 12872
rect 23348 12860 23354 12912
rect 25133 12903 25191 12909
rect 25133 12869 25145 12903
rect 25179 12900 25191 12903
rect 25222 12900 25228 12912
rect 25179 12872 25228 12900
rect 25179 12869 25191 12872
rect 25133 12863 25191 12869
rect 25222 12860 25228 12872
rect 25280 12860 25286 12912
rect 25884 12909 25912 12940
rect 26050 12928 26056 12980
rect 26108 12968 26114 12980
rect 36722 12968 36728 12980
rect 26108 12940 36728 12968
rect 26108 12928 26114 12940
rect 36722 12928 36728 12940
rect 36780 12928 36786 12980
rect 25869 12903 25927 12909
rect 25869 12869 25881 12903
rect 25915 12900 25927 12903
rect 25958 12900 25964 12912
rect 25915 12872 25964 12900
rect 25915 12869 25927 12872
rect 25869 12863 25927 12869
rect 25958 12860 25964 12872
rect 26016 12860 26022 12912
rect 24302 12792 24308 12844
rect 24360 12792 24366 12844
rect 25240 12832 25268 12860
rect 26329 12835 26387 12841
rect 26329 12832 26341 12835
rect 25240 12804 26341 12832
rect 26329 12801 26341 12804
rect 26375 12801 26387 12835
rect 26329 12795 26387 12801
rect 27157 12835 27215 12841
rect 27157 12801 27169 12835
rect 27203 12801 27215 12835
rect 27157 12795 27215 12801
rect 28353 12835 28411 12841
rect 28353 12801 28365 12835
rect 28399 12832 28411 12835
rect 31570 12832 31576 12844
rect 28399 12804 31576 12832
rect 28399 12801 28411 12804
rect 28353 12795 28411 12801
rect 22925 12767 22983 12773
rect 22925 12733 22937 12767
rect 22971 12733 22983 12767
rect 22925 12727 22983 12733
rect 18874 12696 18880 12708
rect 17788 12668 18880 12696
rect 18874 12656 18880 12668
rect 18932 12656 18938 12708
rect 22278 12656 22284 12708
rect 22336 12656 22342 12708
rect 22462 12656 22468 12708
rect 22520 12696 22526 12708
rect 22940 12696 22968 12727
rect 23290 12724 23296 12776
rect 23348 12764 23354 12776
rect 24673 12767 24731 12773
rect 24673 12764 24685 12767
rect 23348 12736 24685 12764
rect 23348 12724 23354 12736
rect 24673 12733 24685 12736
rect 24719 12764 24731 12767
rect 27172 12764 27200 12795
rect 31570 12792 31576 12804
rect 31628 12792 31634 12844
rect 24719 12736 27200 12764
rect 24719 12733 24731 12736
rect 24673 12727 24731 12733
rect 28902 12724 28908 12776
rect 28960 12724 28966 12776
rect 24854 12696 24860 12708
rect 22520 12668 22968 12696
rect 24228 12668 24860 12696
rect 22520 12656 22526 12668
rect 20070 12628 20076 12640
rect 17696 12600 20076 12628
rect 17221 12591 17279 12597
rect 20070 12588 20076 12600
rect 20128 12588 20134 12640
rect 20162 12588 20168 12640
rect 20220 12628 20226 12640
rect 21450 12628 21456 12640
rect 20220 12600 21456 12628
rect 20220 12588 20226 12600
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 22554 12588 22560 12640
rect 22612 12628 22618 12640
rect 24228 12628 24256 12668
rect 24854 12656 24860 12668
rect 24912 12656 24918 12708
rect 22612 12600 24256 12628
rect 22612 12588 22618 12600
rect 24302 12588 24308 12640
rect 24360 12628 24366 12640
rect 26513 12631 26571 12637
rect 26513 12628 26525 12631
rect 24360 12600 26525 12628
rect 24360 12588 24366 12600
rect 26513 12597 26525 12600
rect 26559 12628 26571 12631
rect 27062 12628 27068 12640
rect 26559 12600 27068 12628
rect 26559 12597 26571 12600
rect 26513 12591 26571 12597
rect 27062 12588 27068 12600
rect 27120 12588 27126 12640
rect 27801 12631 27859 12637
rect 27801 12597 27813 12631
rect 27847 12628 27859 12631
rect 28350 12628 28356 12640
rect 27847 12600 28356 12628
rect 27847 12597 27859 12600
rect 27801 12591 27859 12597
rect 28350 12588 28356 12600
rect 28408 12588 28414 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 2222 12384 2228 12436
rect 2280 12384 2286 12436
rect 4065 12427 4123 12433
rect 4065 12393 4077 12427
rect 4111 12424 4123 12427
rect 4246 12424 4252 12436
rect 4111 12396 4252 12424
rect 4111 12393 4123 12396
rect 4065 12387 4123 12393
rect 4246 12384 4252 12396
rect 4304 12384 4310 12436
rect 6270 12424 6276 12436
rect 5000 12396 6276 12424
rect 2406 12316 2412 12368
rect 2464 12316 2470 12368
rect 5000 12365 5028 12396
rect 6270 12384 6276 12396
rect 6328 12384 6334 12436
rect 8570 12424 8576 12436
rect 6748 12396 8576 12424
rect 6748 12368 6776 12396
rect 8570 12384 8576 12396
rect 8628 12424 8634 12436
rect 9030 12424 9036 12436
rect 8628 12396 9036 12424
rect 8628 12384 8634 12396
rect 9030 12384 9036 12396
rect 9088 12384 9094 12436
rect 9401 12427 9459 12433
rect 9401 12393 9413 12427
rect 9447 12424 9459 12427
rect 9490 12424 9496 12436
rect 9447 12396 9496 12424
rect 9447 12393 9459 12396
rect 9401 12387 9459 12393
rect 9490 12384 9496 12396
rect 9548 12384 9554 12436
rect 11606 12424 11612 12436
rect 9600 12396 11612 12424
rect 4985 12359 5043 12365
rect 4985 12325 4997 12359
rect 5031 12325 5043 12359
rect 4985 12319 5043 12325
rect 5166 12316 5172 12368
rect 5224 12356 5230 12368
rect 5442 12356 5448 12368
rect 5224 12328 5448 12356
rect 5224 12316 5230 12328
rect 5442 12316 5448 12328
rect 5500 12316 5506 12368
rect 6730 12316 6736 12368
rect 6788 12316 6794 12368
rect 7282 12316 7288 12368
rect 7340 12356 7346 12368
rect 7834 12356 7840 12368
rect 7340 12328 7840 12356
rect 7340 12316 7346 12328
rect 7834 12316 7840 12328
rect 7892 12316 7898 12368
rect 2424 12288 2452 12316
rect 8573 12291 8631 12297
rect 2424 12260 2544 12288
rect 1854 12180 1860 12232
rect 1912 12220 1918 12232
rect 2406 12220 2412 12232
rect 1912 12192 2412 12220
rect 1912 12180 1918 12192
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 2133 12155 2191 12161
rect 2133 12121 2145 12155
rect 2179 12152 2191 12155
rect 2222 12152 2228 12164
rect 2179 12124 2228 12152
rect 2179 12121 2191 12124
rect 2133 12115 2191 12121
rect 2222 12112 2228 12124
rect 2280 12152 2286 12164
rect 2516 12152 2544 12260
rect 2792 12260 8064 12288
rect 2792 12229 2820 12260
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 4338 12180 4344 12232
rect 4396 12180 4402 12232
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5442 12220 5448 12232
rect 4856 12192 5448 12220
rect 4856 12180 4862 12192
rect 5442 12180 5448 12192
rect 5500 12180 5506 12232
rect 7466 12180 7472 12232
rect 7524 12180 7530 12232
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 7929 12223 7987 12229
rect 7929 12220 7941 12223
rect 7892 12192 7941 12220
rect 7892 12180 7898 12192
rect 7929 12189 7941 12192
rect 7975 12189 7987 12223
rect 8036 12220 8064 12260
rect 8573 12257 8585 12291
rect 8619 12288 8631 12291
rect 9600 12288 9628 12396
rect 11606 12384 11612 12396
rect 11664 12384 11670 12436
rect 12989 12427 13047 12433
rect 12989 12424 13001 12427
rect 11716 12396 13001 12424
rect 10870 12316 10876 12368
rect 10928 12356 10934 12368
rect 11716 12356 11744 12396
rect 12989 12393 13001 12396
rect 13035 12393 13047 12427
rect 12989 12387 13047 12393
rect 13538 12384 13544 12436
rect 13596 12424 13602 12436
rect 14734 12424 14740 12436
rect 13596 12396 14740 12424
rect 13596 12384 13602 12396
rect 14734 12384 14740 12396
rect 14792 12384 14798 12436
rect 16942 12424 16948 12436
rect 14844 12396 16948 12424
rect 10928 12328 11744 12356
rect 11793 12359 11851 12365
rect 10928 12316 10934 12328
rect 11793 12325 11805 12359
rect 11839 12325 11851 12359
rect 14093 12359 14151 12365
rect 14093 12356 14105 12359
rect 11793 12319 11851 12325
rect 12452 12328 14105 12356
rect 8619 12260 9628 12288
rect 8619 12257 8631 12260
rect 8573 12251 8631 12257
rect 9950 12248 9956 12300
rect 10008 12248 10014 12300
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 11149 12291 11207 12297
rect 11149 12288 11161 12291
rect 10468 12260 11161 12288
rect 10468 12248 10474 12260
rect 11149 12257 11161 12260
rect 11195 12257 11207 12291
rect 11149 12251 11207 12257
rect 9398 12220 9404 12232
rect 8036 12192 9404 12220
rect 7929 12183 7987 12189
rect 9398 12180 9404 12192
rect 9456 12180 9462 12232
rect 10594 12220 10600 12232
rect 10336 12192 10600 12220
rect 2280 12124 2544 12152
rect 3421 12155 3479 12161
rect 2280 12112 2286 12124
rect 3421 12121 3433 12155
rect 3467 12152 3479 12155
rect 4522 12152 4528 12164
rect 3467 12124 4528 12152
rect 3467 12121 3479 12124
rect 3421 12115 3479 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 5721 12155 5779 12161
rect 5721 12121 5733 12155
rect 5767 12121 5779 12155
rect 5721 12115 5779 12121
rect 1578 12044 1584 12096
rect 1636 12044 1642 12096
rect 1765 12087 1823 12093
rect 1765 12053 1777 12087
rect 1811 12084 1823 12087
rect 1854 12084 1860 12096
rect 1811 12056 1860 12084
rect 1811 12053 1823 12056
rect 1765 12047 1823 12053
rect 1854 12044 1860 12056
rect 1912 12084 1918 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 1912 12056 3801 12084
rect 1912 12044 1918 12056
rect 3789 12053 3801 12056
rect 3835 12084 3847 12087
rect 4614 12084 4620 12096
rect 3835 12056 4620 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 4614 12044 4620 12056
rect 4672 12084 4678 12096
rect 4982 12084 4988 12096
rect 4672 12056 4988 12084
rect 4672 12044 4678 12056
rect 4982 12044 4988 12056
rect 5040 12044 5046 12096
rect 5736 12084 5764 12115
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 10042 12152 10048 12164
rect 9692 12124 10048 12152
rect 6362 12084 6368 12096
rect 5736 12056 6368 12084
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 8018 12044 8024 12096
rect 8076 12084 8082 12096
rect 8478 12084 8484 12096
rect 8076 12056 8484 12084
rect 8076 12044 8082 12056
rect 8478 12044 8484 12056
rect 8536 12084 8542 12096
rect 9030 12084 9036 12096
rect 8536 12056 9036 12084
rect 8536 12044 8542 12056
rect 9030 12044 9036 12056
rect 9088 12044 9094 12096
rect 9398 12044 9404 12096
rect 9456 12084 9462 12096
rect 9692 12084 9720 12124
rect 10042 12112 10048 12124
rect 10100 12112 10106 12164
rect 9456 12056 9720 12084
rect 9456 12044 9462 12056
rect 9766 12044 9772 12096
rect 9824 12044 9830 12096
rect 9861 12087 9919 12093
rect 9861 12053 9873 12087
rect 9907 12084 9919 12087
rect 10336 12084 10364 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11514 12180 11520 12232
rect 11572 12220 11578 12232
rect 11808 12220 11836 12319
rect 12342 12248 12348 12300
rect 12400 12248 12406 12300
rect 11572 12192 11836 12220
rect 11572 12180 11578 12192
rect 11974 12180 11980 12232
rect 12032 12220 12038 12232
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 12032 12192 12265 12220
rect 12032 12180 12038 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12452 12220 12480 12328
rect 14093 12325 14105 12328
rect 14139 12325 14151 12359
rect 14093 12319 14151 12325
rect 12618 12248 12624 12300
rect 12676 12288 12682 12300
rect 12894 12288 12900 12300
rect 12676 12260 12900 12288
rect 12676 12248 12682 12260
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13538 12248 13544 12300
rect 13596 12248 13602 12300
rect 12253 12183 12311 12189
rect 12360 12192 12480 12220
rect 13449 12223 13507 12229
rect 10965 12155 11023 12161
rect 10965 12121 10977 12155
rect 11011 12152 11023 12155
rect 11011 12124 11836 12152
rect 11011 12121 11023 12124
rect 10965 12115 11023 12121
rect 9907 12056 10364 12084
rect 9907 12053 9919 12056
rect 9861 12047 9919 12053
rect 10594 12044 10600 12096
rect 10652 12044 10658 12096
rect 10686 12044 10692 12096
rect 10744 12084 10750 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10744 12056 11069 12084
rect 10744 12044 10750 12056
rect 11057 12053 11069 12056
rect 11103 12053 11115 12087
rect 11808 12084 11836 12124
rect 11882 12112 11888 12164
rect 11940 12152 11946 12164
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 11940 12124 12173 12152
rect 11940 12112 11946 12124
rect 12161 12121 12173 12124
rect 12207 12152 12219 12155
rect 12360 12152 12388 12192
rect 13449 12189 13461 12223
rect 13495 12220 13507 12223
rect 14844 12220 14872 12396
rect 16942 12384 16948 12396
rect 17000 12384 17006 12436
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17092 12396 18276 12424
rect 17092 12384 17098 12396
rect 15194 12316 15200 12368
rect 15252 12356 15258 12368
rect 15654 12356 15660 12368
rect 15252 12328 15660 12356
rect 15252 12316 15258 12328
rect 15654 12316 15660 12328
rect 15712 12316 15718 12368
rect 18046 12356 18052 12368
rect 17972 12328 18052 12356
rect 14918 12248 14924 12300
rect 14976 12288 14982 12300
rect 15473 12291 15531 12297
rect 15473 12288 15485 12291
rect 14976 12260 15485 12288
rect 14976 12248 14982 12260
rect 15473 12257 15485 12260
rect 15519 12288 15531 12291
rect 16117 12291 16175 12297
rect 16117 12288 16129 12291
rect 15519 12260 16129 12288
rect 15519 12257 15531 12260
rect 15473 12251 15531 12257
rect 16117 12257 16129 12260
rect 16163 12257 16175 12291
rect 16117 12251 16175 12257
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17972 12288 18000 12328
rect 18046 12316 18052 12328
rect 18104 12316 18110 12368
rect 18248 12356 18276 12396
rect 18874 12384 18880 12436
rect 18932 12384 18938 12436
rect 20346 12424 20352 12436
rect 19444 12396 20352 12424
rect 18969 12359 19027 12365
rect 18969 12356 18981 12359
rect 18248 12328 18981 12356
rect 18969 12325 18981 12328
rect 19015 12325 19027 12359
rect 18969 12319 19027 12325
rect 16908 12260 18000 12288
rect 18325 12291 18383 12297
rect 16908 12248 16914 12260
rect 18325 12257 18337 12291
rect 18371 12288 18383 12291
rect 18598 12288 18604 12300
rect 18371 12260 18604 12288
rect 18371 12257 18383 12260
rect 18325 12251 18383 12257
rect 18598 12248 18604 12260
rect 18656 12248 18662 12300
rect 19444 12297 19472 12396
rect 20346 12384 20352 12396
rect 20404 12384 20410 12436
rect 20714 12384 20720 12436
rect 20772 12424 20778 12436
rect 21634 12424 21640 12436
rect 20772 12396 21640 12424
rect 20772 12384 20778 12396
rect 21634 12384 21640 12396
rect 21692 12384 21698 12436
rect 21726 12384 21732 12436
rect 21784 12424 21790 12436
rect 25222 12424 25228 12436
rect 21784 12396 25228 12424
rect 21784 12384 21790 12396
rect 25222 12384 25228 12396
rect 25280 12384 25286 12436
rect 25685 12427 25743 12433
rect 25685 12393 25697 12427
rect 25731 12424 25743 12427
rect 27614 12424 27620 12436
rect 25731 12396 27620 12424
rect 25731 12393 25743 12396
rect 25685 12387 25743 12393
rect 27614 12384 27620 12396
rect 27672 12384 27678 12436
rect 28442 12384 28448 12436
rect 28500 12384 28506 12436
rect 29270 12384 29276 12436
rect 29328 12424 29334 12436
rect 29730 12424 29736 12436
rect 29328 12396 29736 12424
rect 29328 12384 29334 12396
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 24118 12316 24124 12368
rect 24176 12356 24182 12368
rect 24176 12328 27292 12356
rect 24176 12316 24182 12328
rect 19429 12291 19487 12297
rect 19429 12257 19441 12291
rect 19475 12257 19487 12291
rect 19429 12251 19487 12257
rect 20073 12291 20131 12297
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 22281 12291 22339 12297
rect 22281 12288 22293 12291
rect 20119 12260 22293 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 22281 12257 22293 12260
rect 22327 12288 22339 12291
rect 22554 12288 22560 12300
rect 22327 12260 22560 12288
rect 22327 12257 22339 12260
rect 22281 12251 22339 12257
rect 22554 12248 22560 12260
rect 22612 12248 22618 12300
rect 24302 12248 24308 12300
rect 24360 12288 24366 12300
rect 24578 12288 24584 12300
rect 24360 12260 24584 12288
rect 24360 12248 24366 12260
rect 24578 12248 24584 12260
rect 24636 12248 24642 12300
rect 13495 12192 14872 12220
rect 13495 12189 13507 12192
rect 13449 12183 13507 12189
rect 18506 12180 18512 12232
rect 18564 12220 18570 12232
rect 19978 12220 19984 12232
rect 18564 12192 19984 12220
rect 18564 12180 18570 12192
rect 19978 12180 19984 12192
rect 20036 12180 20042 12232
rect 24394 12180 24400 12232
rect 24452 12220 24458 12232
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 24452 12192 25053 12220
rect 24452 12180 24458 12192
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 26786 12180 26792 12232
rect 26844 12220 26850 12232
rect 27157 12223 27215 12229
rect 27157 12220 27169 12223
rect 26844 12192 27169 12220
rect 26844 12180 26850 12192
rect 27157 12189 27169 12192
rect 27203 12189 27215 12223
rect 27264 12220 27292 12328
rect 27706 12316 27712 12368
rect 27764 12356 27770 12368
rect 35986 12356 35992 12368
rect 27764 12328 35992 12356
rect 27764 12316 27770 12328
rect 35986 12316 35992 12328
rect 36044 12316 36050 12368
rect 27338 12248 27344 12300
rect 27396 12288 27402 12300
rect 29638 12288 29644 12300
rect 27396 12260 29644 12288
rect 27396 12248 27402 12260
rect 29638 12248 29644 12260
rect 29696 12248 29702 12300
rect 31662 12220 31668 12232
rect 27264 12192 31668 12220
rect 27157 12183 27215 12189
rect 31662 12180 31668 12192
rect 31720 12180 31726 12232
rect 14461 12155 14519 12161
rect 12207 12124 12388 12152
rect 12544 12124 14412 12152
rect 12207 12121 12219 12124
rect 12161 12115 12219 12121
rect 12544 12084 12572 12124
rect 11808 12056 12572 12084
rect 11057 12047 11115 12053
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 12802 12084 12808 12096
rect 12676 12056 12808 12084
rect 12676 12044 12682 12056
rect 12802 12044 12808 12056
rect 12860 12044 12866 12096
rect 13357 12087 13415 12093
rect 13357 12053 13369 12087
rect 13403 12084 13415 12087
rect 13630 12084 13636 12096
rect 13403 12056 13636 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 14384 12084 14412 12124
rect 14461 12121 14473 12155
rect 14507 12152 14519 12155
rect 14737 12155 14795 12161
rect 14737 12152 14749 12155
rect 14507 12124 14749 12152
rect 14507 12121 14519 12124
rect 14461 12115 14519 12121
rect 14737 12121 14749 12124
rect 14783 12152 14795 12155
rect 15194 12152 15200 12164
rect 14783 12124 15200 12152
rect 14783 12121 14795 12124
rect 14737 12115 14795 12121
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 16397 12161 16403 12164
rect 16393 12115 16403 12161
rect 16397 12112 16403 12115
rect 16455 12112 16461 12164
rect 16850 12112 16856 12164
rect 16908 12112 16914 12164
rect 20349 12155 20407 12161
rect 18156 12124 20300 12152
rect 15010 12084 15016 12096
rect 14384 12056 15016 12084
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15838 12044 15844 12096
rect 15896 12084 15902 12096
rect 16574 12084 16580 12096
rect 15896 12056 16580 12084
rect 15896 12044 15902 12056
rect 16574 12044 16580 12056
rect 16632 12044 16638 12096
rect 16666 12044 16672 12096
rect 16724 12084 16730 12096
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 16724 12056 17877 12084
rect 16724 12044 16730 12056
rect 17865 12053 17877 12056
rect 17911 12084 17923 12087
rect 18156 12084 18184 12124
rect 20272 12096 20300 12124
rect 20349 12121 20361 12155
rect 20395 12121 20407 12155
rect 21726 12152 21732 12164
rect 21574 12124 21732 12152
rect 20349 12115 20407 12121
rect 17911 12056 18184 12084
rect 17911 12053 17923 12056
rect 17865 12047 17923 12053
rect 18230 12044 18236 12096
rect 18288 12084 18294 12096
rect 19518 12084 19524 12096
rect 18288 12056 19524 12084
rect 18288 12044 18294 12056
rect 19518 12044 19524 12056
rect 19576 12044 19582 12096
rect 19610 12044 19616 12096
rect 19668 12084 19674 12096
rect 19794 12084 19800 12096
rect 19668 12056 19800 12084
rect 19668 12044 19674 12056
rect 19794 12044 19800 12056
rect 19852 12044 19858 12096
rect 20254 12044 20260 12096
rect 20312 12044 20318 12096
rect 20364 12084 20392 12115
rect 21726 12112 21732 12124
rect 21784 12152 21790 12164
rect 21784 12124 21956 12152
rect 21784 12112 21790 12124
rect 21634 12084 21640 12096
rect 20364 12056 21640 12084
rect 21634 12044 21640 12056
rect 21692 12044 21698 12096
rect 21818 12044 21824 12096
rect 21876 12044 21882 12096
rect 21928 12084 21956 12124
rect 22554 12112 22560 12164
rect 22612 12112 22618 12164
rect 23782 12124 24532 12152
rect 22830 12084 22836 12096
rect 21928 12056 22836 12084
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 24026 12044 24032 12096
rect 24084 12044 24090 12096
rect 24504 12093 24532 12124
rect 24670 12112 24676 12164
rect 24728 12152 24734 12164
rect 28353 12155 28411 12161
rect 28353 12152 28365 12155
rect 24728 12124 28365 12152
rect 24728 12112 24734 12124
rect 28353 12121 28365 12124
rect 28399 12152 28411 12155
rect 28813 12155 28871 12161
rect 28813 12152 28825 12155
rect 28399 12124 28825 12152
rect 28399 12121 28411 12124
rect 28353 12115 28411 12121
rect 28813 12121 28825 12124
rect 28859 12121 28871 12155
rect 28813 12115 28871 12121
rect 24489 12087 24547 12093
rect 24489 12053 24501 12087
rect 24535 12084 24547 12087
rect 24578 12084 24584 12096
rect 24535 12056 24584 12084
rect 24535 12053 24547 12056
rect 24489 12047 24547 12053
rect 24578 12044 24584 12056
rect 24636 12044 24642 12096
rect 27614 12044 27620 12096
rect 27672 12084 27678 12096
rect 27801 12087 27859 12093
rect 27801 12084 27813 12087
rect 27672 12056 27813 12084
rect 27672 12044 27678 12056
rect 27801 12053 27813 12056
rect 27847 12053 27859 12087
rect 27801 12047 27859 12053
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 934 11840 940 11892
rect 992 11880 998 11892
rect 1397 11883 1455 11889
rect 1397 11880 1409 11883
rect 992 11852 1409 11880
rect 992 11840 998 11852
rect 1397 11849 1409 11852
rect 1443 11849 1455 11883
rect 1397 11843 1455 11849
rect 2590 11840 2596 11892
rect 2648 11840 2654 11892
rect 5442 11840 5448 11892
rect 5500 11880 5506 11892
rect 5500 11852 9352 11880
rect 5500 11840 5506 11852
rect 1302 11772 1308 11824
rect 1360 11812 1366 11824
rect 5258 11812 5264 11824
rect 1360 11784 5264 11812
rect 1360 11772 1366 11784
rect 5258 11772 5264 11784
rect 5316 11812 5322 11824
rect 5316 11784 5580 11812
rect 5316 11772 5322 11784
rect 1946 11704 1952 11756
rect 2004 11704 2010 11756
rect 2774 11704 2780 11756
rect 2832 11744 2838 11756
rect 3053 11747 3111 11753
rect 3053 11744 3065 11747
rect 2832 11716 3065 11744
rect 2832 11704 2838 11716
rect 3053 11713 3065 11716
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3326 11704 3332 11756
rect 3384 11744 3390 11756
rect 3602 11744 3608 11756
rect 3384 11716 3608 11744
rect 3384 11704 3390 11716
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 4157 11747 4215 11753
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 5166 11744 5172 11756
rect 4203 11716 5172 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 5166 11704 5172 11716
rect 5224 11704 5230 11756
rect 5552 11744 5580 11784
rect 5626 11772 5632 11824
rect 5684 11772 5690 11824
rect 5718 11772 5724 11824
rect 5776 11812 5782 11824
rect 5994 11812 6000 11824
rect 5776 11784 6000 11812
rect 5776 11772 5782 11784
rect 5994 11772 6000 11784
rect 6052 11772 6058 11824
rect 6457 11815 6515 11821
rect 6457 11781 6469 11815
rect 6503 11812 6515 11815
rect 6549 11815 6607 11821
rect 6549 11812 6561 11815
rect 6503 11784 6561 11812
rect 6503 11781 6515 11784
rect 6457 11775 6515 11781
rect 6549 11781 6561 11784
rect 6595 11812 6607 11815
rect 6822 11812 6828 11824
rect 6595 11784 6828 11812
rect 6595 11781 6607 11784
rect 6549 11775 6607 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7208 11753 7236 11852
rect 9324 11824 9352 11852
rect 9582 11840 9588 11892
rect 9640 11880 9646 11892
rect 11422 11880 11428 11892
rect 9640 11852 11428 11880
rect 9640 11840 9646 11852
rect 11422 11840 11428 11852
rect 11480 11840 11486 11892
rect 11514 11840 11520 11892
rect 11572 11880 11578 11892
rect 11882 11880 11888 11892
rect 11572 11852 11888 11880
rect 11572 11840 11578 11852
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 11974 11840 11980 11892
rect 12032 11840 12038 11892
rect 12342 11880 12348 11892
rect 12176 11852 12348 11880
rect 7466 11772 7472 11824
rect 7524 11772 7530 11824
rect 8478 11772 8484 11824
rect 8536 11772 8542 11824
rect 9306 11772 9312 11824
rect 9364 11812 9370 11824
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 9364 11784 10149 11812
rect 9364 11772 9370 11784
rect 10137 11781 10149 11784
rect 10183 11781 10195 11815
rect 10137 11775 10195 11781
rect 10962 11772 10968 11824
rect 11020 11772 11026 11824
rect 11701 11815 11759 11821
rect 11701 11781 11713 11815
rect 11747 11812 11759 11815
rect 12066 11812 12072 11824
rect 11747 11784 12072 11812
rect 11747 11781 11759 11784
rect 11701 11775 11759 11781
rect 12066 11772 12072 11784
rect 12124 11772 12130 11824
rect 7193 11747 7251 11753
rect 5552 11716 5856 11744
rect 3234 11636 3240 11688
rect 3292 11676 3298 11688
rect 4614 11676 4620 11688
rect 3292 11648 4620 11676
rect 3292 11636 3298 11648
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5258 11676 5264 11688
rect 5040 11648 5264 11676
rect 5040 11636 5046 11648
rect 5258 11636 5264 11648
rect 5316 11636 5322 11688
rect 5718 11636 5724 11688
rect 5776 11636 5782 11688
rect 5828 11685 5856 11716
rect 7193 11713 7205 11747
rect 7239 11713 7251 11747
rect 7193 11707 7251 11713
rect 9122 11704 9128 11756
rect 9180 11744 9186 11756
rect 9401 11747 9459 11753
rect 9401 11744 9413 11747
rect 9180 11716 9413 11744
rect 9180 11704 9186 11716
rect 9401 11713 9413 11716
rect 9447 11744 9459 11747
rect 9674 11744 9680 11756
rect 9447 11716 9680 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9674 11704 9680 11716
rect 9732 11704 9738 11756
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11744 11207 11747
rect 11238 11744 11244 11756
rect 11195 11716 11244 11744
rect 11195 11713 11207 11716
rect 11149 11707 11207 11713
rect 11238 11704 11244 11716
rect 11296 11704 11302 11756
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12176 11744 12204 11852
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 14182 11880 14188 11892
rect 12492 11852 14188 11880
rect 12492 11840 12498 11852
rect 14182 11840 14188 11852
rect 14240 11840 14246 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 14424 11852 15424 11880
rect 14424 11840 14430 11852
rect 12250 11772 12256 11824
rect 12308 11812 12314 11824
rect 12308 11784 13216 11812
rect 12308 11772 12314 11784
rect 11940 11716 12204 11744
rect 11940 11704 11946 11716
rect 12342 11704 12348 11756
rect 12400 11704 12406 11756
rect 12437 11747 12495 11753
rect 12437 11713 12449 11747
rect 12483 11744 12495 11747
rect 12802 11744 12808 11756
rect 12483 11716 12808 11744
rect 12483 11713 12495 11716
rect 12437 11707 12495 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13188 11753 13216 11784
rect 13446 11772 13452 11824
rect 13504 11772 13510 11824
rect 15286 11812 15292 11824
rect 14674 11784 15292 11812
rect 15286 11772 15292 11784
rect 15344 11772 15350 11824
rect 15396 11812 15424 11852
rect 15470 11840 15476 11892
rect 15528 11840 15534 11892
rect 16022 11840 16028 11892
rect 16080 11880 16086 11892
rect 16206 11880 16212 11892
rect 16080 11852 16212 11880
rect 16080 11840 16086 11852
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 16298 11840 16304 11892
rect 16356 11880 16362 11892
rect 16574 11880 16580 11892
rect 16356 11852 16580 11880
rect 16356 11840 16362 11852
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 17313 11883 17371 11889
rect 17313 11880 17325 11883
rect 16684 11852 17325 11880
rect 16684 11812 16712 11852
rect 17313 11849 17325 11852
rect 17359 11849 17371 11883
rect 17313 11843 17371 11849
rect 17405 11883 17463 11889
rect 17405 11849 17417 11883
rect 17451 11880 17463 11883
rect 17678 11880 17684 11892
rect 17451 11852 17684 11880
rect 17451 11849 17463 11852
rect 17405 11843 17463 11849
rect 17678 11840 17684 11852
rect 17736 11840 17742 11892
rect 18322 11880 18328 11892
rect 17972 11852 18328 11880
rect 15396 11784 16712 11812
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 17972 11812 18000 11852
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18874 11840 18880 11892
rect 18932 11880 18938 11892
rect 18932 11852 19840 11880
rect 18932 11840 18938 11852
rect 17552 11784 18000 11812
rect 17552 11772 17558 11784
rect 13173 11747 13231 11753
rect 13173 11713 13185 11747
rect 13219 11713 13231 11747
rect 14918 11744 14924 11756
rect 13173 11707 13231 11713
rect 14660 11716 14924 11744
rect 5813 11679 5871 11685
rect 5813 11645 5825 11679
rect 5859 11645 5871 11679
rect 5813 11639 5871 11645
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 6880 11648 11652 11676
rect 6880 11636 6886 11648
rect 382 11568 388 11620
rect 440 11608 446 11620
rect 4801 11611 4859 11617
rect 4801 11608 4813 11611
rect 440 11580 4813 11608
rect 440 11568 446 11580
rect 4801 11577 4813 11580
rect 4847 11577 4859 11611
rect 6730 11608 6736 11620
rect 4801 11571 4859 11577
rect 5184 11580 6736 11608
rect 566 11500 572 11552
rect 624 11540 630 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 624 11512 1593 11540
rect 624 11500 630 11512
rect 1581 11509 1593 11512
rect 1627 11540 1639 11543
rect 2590 11540 2596 11552
rect 1627 11512 2596 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 2590 11500 2596 11512
rect 2648 11500 2654 11552
rect 3694 11500 3700 11552
rect 3752 11500 3758 11552
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 5184 11540 5212 11580
rect 6730 11568 6736 11580
rect 6788 11568 6794 11620
rect 8570 11568 8576 11620
rect 8628 11608 8634 11620
rect 9122 11608 9128 11620
rect 8628 11580 9128 11608
rect 8628 11568 8634 11580
rect 9122 11568 9128 11580
rect 9180 11568 9186 11620
rect 11624 11608 11652 11648
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 12250 11676 12256 11688
rect 11756 11648 12256 11676
rect 11756 11636 11762 11648
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11676 12679 11679
rect 13906 11676 13912 11688
rect 12667 11648 13912 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 13906 11636 13912 11648
rect 13964 11676 13970 11688
rect 14660 11676 14688 11716
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 15838 11704 15844 11756
rect 15896 11704 15902 11756
rect 16390 11704 16396 11756
rect 16448 11744 16454 11756
rect 16448 11716 16896 11744
rect 16448 11704 16454 11716
rect 15930 11676 15936 11688
rect 13964 11648 14688 11676
rect 14844 11648 15936 11676
rect 13964 11636 13970 11648
rect 12894 11608 12900 11620
rect 11624 11580 12900 11608
rect 12894 11568 12900 11580
rect 12952 11568 12958 11620
rect 4304 11512 5212 11540
rect 5261 11543 5319 11549
rect 4304 11500 4310 11512
rect 5261 11509 5273 11543
rect 5307 11540 5319 11543
rect 6914 11540 6920 11552
rect 5307 11512 6920 11540
rect 5307 11509 5319 11512
rect 5261 11503 5319 11509
rect 6914 11500 6920 11512
rect 6972 11500 6978 11552
rect 7834 11500 7840 11552
rect 7892 11540 7898 11552
rect 8941 11543 8999 11549
rect 8941 11540 8953 11543
rect 7892 11512 8953 11540
rect 7892 11500 7898 11512
rect 8941 11509 8953 11512
rect 8987 11509 8999 11543
rect 8941 11503 8999 11509
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 14844 11540 14872 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11676 16175 11679
rect 16758 11676 16764 11688
rect 16163 11648 16764 11676
rect 16163 11645 16175 11648
rect 16117 11639 16175 11645
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 16868 11676 16896 11716
rect 19610 11704 19616 11756
rect 19668 11704 19674 11756
rect 19812 11744 19840 11852
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20990 11880 20996 11892
rect 20312 11852 20996 11880
rect 20312 11840 20318 11852
rect 20990 11840 20996 11852
rect 21048 11840 21054 11892
rect 21542 11840 21548 11892
rect 21600 11880 21606 11892
rect 21637 11883 21695 11889
rect 21637 11880 21649 11883
rect 21600 11852 21649 11880
rect 21600 11840 21606 11852
rect 21637 11849 21649 11852
rect 21683 11880 21695 11883
rect 21683 11852 24072 11880
rect 21683 11849 21695 11852
rect 21637 11843 21695 11849
rect 20346 11772 20352 11824
rect 20404 11812 20410 11824
rect 21821 11815 21879 11821
rect 21821 11812 21833 11815
rect 20404 11784 21833 11812
rect 20404 11772 20410 11784
rect 21821 11781 21833 11784
rect 21867 11812 21879 11815
rect 22002 11812 22008 11824
rect 21867 11784 22008 11812
rect 21867 11781 21879 11784
rect 21821 11775 21879 11781
rect 22002 11772 22008 11784
rect 22060 11772 22066 11824
rect 22094 11772 22100 11824
rect 22152 11812 22158 11824
rect 23014 11812 23020 11824
rect 22152 11784 23020 11812
rect 22152 11772 22158 11784
rect 23014 11772 23020 11784
rect 23072 11772 23078 11824
rect 24044 11812 24072 11852
rect 24578 11840 24584 11892
rect 24636 11880 24642 11892
rect 25866 11880 25872 11892
rect 24636 11852 25872 11880
rect 24636 11840 24642 11852
rect 25866 11840 25872 11852
rect 25924 11840 25930 11892
rect 27798 11840 27804 11892
rect 27856 11880 27862 11892
rect 28261 11883 28319 11889
rect 28261 11880 28273 11883
rect 27856 11852 28273 11880
rect 27856 11840 27862 11852
rect 28261 11849 28273 11852
rect 28307 11849 28319 11883
rect 28261 11843 28319 11849
rect 30374 11840 30380 11892
rect 30432 11880 30438 11892
rect 34514 11880 34520 11892
rect 30432 11852 34520 11880
rect 30432 11840 30438 11852
rect 34514 11840 34520 11852
rect 34572 11840 34578 11892
rect 24210 11812 24216 11824
rect 23966 11784 24216 11812
rect 24210 11772 24216 11784
rect 24268 11812 24274 11824
rect 24596 11812 24624 11840
rect 24268 11784 24624 11812
rect 24268 11772 24274 11784
rect 24946 11772 24952 11824
rect 25004 11812 25010 11824
rect 25130 11812 25136 11824
rect 25004 11784 25136 11812
rect 25004 11772 25010 11784
rect 25130 11772 25136 11784
rect 25188 11772 25194 11824
rect 25222 11772 25228 11824
rect 25280 11812 25286 11824
rect 33410 11812 33416 11824
rect 25280 11784 33416 11812
rect 25280 11772 25286 11784
rect 33410 11772 33416 11784
rect 33468 11772 33474 11824
rect 20441 11747 20499 11753
rect 20441 11744 20453 11747
rect 19812 11716 20453 11744
rect 20441 11713 20453 11716
rect 20487 11744 20499 11747
rect 20622 11744 20628 11756
rect 20487 11716 20628 11744
rect 20487 11713 20499 11716
rect 20441 11707 20499 11713
rect 20622 11704 20628 11716
rect 20680 11704 20686 11756
rect 20717 11747 20775 11753
rect 20717 11713 20729 11747
rect 20763 11744 20775 11747
rect 21174 11744 21180 11756
rect 20763 11716 21180 11744
rect 20763 11713 20775 11716
rect 20717 11707 20775 11713
rect 21174 11704 21180 11716
rect 21232 11704 21238 11756
rect 22462 11704 22468 11756
rect 22520 11704 22526 11756
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11744 25743 11747
rect 26234 11744 26240 11756
rect 25731 11716 26240 11744
rect 25731 11713 25743 11716
rect 25685 11707 25743 11713
rect 26234 11704 26240 11716
rect 26292 11704 26298 11756
rect 27154 11704 27160 11756
rect 27212 11704 27218 11756
rect 32398 11704 32404 11756
rect 32456 11744 32462 11756
rect 40034 11744 40040 11756
rect 32456 11716 40040 11744
rect 32456 11704 32462 11716
rect 40034 11704 40040 11716
rect 40092 11704 40098 11756
rect 16868 11648 17540 11676
rect 14918 11568 14924 11620
rect 14976 11568 14982 11620
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 17034 11608 17040 11620
rect 15712 11580 17040 11608
rect 15712 11568 15718 11580
rect 17034 11568 17040 11580
rect 17092 11568 17098 11620
rect 17512 11608 17540 11648
rect 17586 11636 17592 11688
rect 17644 11636 17650 11688
rect 18233 11679 18291 11685
rect 18233 11645 18245 11679
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 18509 11679 18567 11685
rect 18509 11645 18521 11679
rect 18555 11676 18567 11679
rect 19242 11676 19248 11688
rect 18555 11648 19248 11676
rect 18555 11645 18567 11648
rect 18509 11639 18567 11645
rect 17862 11608 17868 11620
rect 17512 11580 17868 11608
rect 17862 11568 17868 11580
rect 17920 11568 17926 11620
rect 12492 11512 14872 11540
rect 12492 11500 12498 11512
rect 16666 11500 16672 11552
rect 16724 11540 16730 11552
rect 16945 11543 17003 11549
rect 16945 11540 16957 11543
rect 16724 11512 16957 11540
rect 16724 11500 16730 11512
rect 16945 11509 16957 11512
rect 16991 11509 17003 11543
rect 16945 11503 17003 11509
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 18248 11540 18276 11639
rect 19242 11636 19248 11648
rect 19300 11636 19306 11688
rect 19518 11636 19524 11688
rect 19576 11676 19582 11688
rect 21082 11676 21088 11688
rect 19576 11648 21088 11676
rect 19576 11636 19582 11648
rect 21082 11636 21088 11648
rect 21140 11636 21146 11688
rect 21818 11636 21824 11688
rect 21876 11676 21882 11688
rect 22278 11676 22284 11688
rect 21876 11648 22284 11676
rect 21876 11636 21882 11648
rect 22278 11636 22284 11648
rect 22336 11636 22342 11688
rect 22741 11679 22799 11685
rect 22741 11645 22753 11679
rect 22787 11676 22799 11679
rect 26329 11679 26387 11685
rect 26329 11676 26341 11679
rect 22787 11648 26341 11676
rect 22787 11645 22799 11648
rect 22741 11639 22799 11645
rect 26329 11645 26341 11648
rect 26375 11645 26387 11679
rect 26329 11639 26387 11645
rect 19610 11568 19616 11620
rect 19668 11608 19674 11620
rect 21726 11608 21732 11620
rect 19668 11580 21732 11608
rect 19668 11568 19674 11580
rect 21726 11568 21732 11580
rect 21784 11568 21790 11620
rect 22094 11568 22100 11620
rect 22152 11568 22158 11620
rect 24946 11608 24952 11620
rect 24228 11580 24952 11608
rect 19702 11540 19708 11552
rect 17460 11512 19708 11540
rect 17460 11500 17466 11512
rect 19702 11500 19708 11512
rect 19760 11500 19766 11552
rect 19794 11500 19800 11552
rect 19852 11540 19858 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 19852 11512 19993 11540
rect 19852 11500 19858 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 20714 11500 20720 11552
rect 20772 11540 20778 11552
rect 23842 11540 23848 11552
rect 20772 11512 23848 11540
rect 20772 11500 20778 11512
rect 23842 11500 23848 11512
rect 23900 11500 23906 11552
rect 23934 11500 23940 11552
rect 23992 11540 23998 11552
rect 24228 11549 24256 11580
rect 24946 11568 24952 11580
rect 25004 11568 25010 11620
rect 25866 11568 25872 11620
rect 25924 11608 25930 11620
rect 32214 11608 32220 11620
rect 25924 11580 32220 11608
rect 25924 11568 25930 11580
rect 32214 11568 32220 11580
rect 32272 11568 32278 11620
rect 24213 11543 24271 11549
rect 24213 11540 24225 11543
rect 23992 11512 24225 11540
rect 23992 11500 23998 11512
rect 24213 11509 24225 11512
rect 24259 11509 24271 11543
rect 24213 11503 24271 11509
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 27706 11540 27712 11552
rect 24636 11512 27712 11540
rect 24636 11500 24642 11512
rect 27706 11500 27712 11512
rect 27764 11500 27770 11552
rect 27798 11500 27804 11552
rect 27856 11500 27862 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 2314 11296 2320 11348
rect 2372 11296 2378 11348
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 3510 11336 3516 11348
rect 3467 11308 3516 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 5810 11296 5816 11348
rect 5868 11336 5874 11348
rect 7193 11339 7251 11345
rect 7193 11336 7205 11339
rect 5868 11308 7205 11336
rect 5868 11296 5874 11308
rect 7193 11305 7205 11308
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7374 11296 7380 11348
rect 7432 11336 7438 11348
rect 7558 11336 7564 11348
rect 7432 11308 7564 11336
rect 7432 11296 7438 11308
rect 7558 11296 7564 11308
rect 7616 11336 7622 11348
rect 12434 11336 12440 11348
rect 7616 11308 12440 11336
rect 7616 11296 7622 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13538 11336 13544 11348
rect 13320 11308 13544 11336
rect 13320 11296 13326 11308
rect 13538 11296 13544 11308
rect 13596 11296 13602 11348
rect 13814 11296 13820 11348
rect 13872 11296 13878 11348
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 14516 11308 16160 11336
rect 14516 11296 14522 11308
rect 2406 11228 2412 11280
rect 2464 11268 2470 11280
rect 4249 11271 4307 11277
rect 4249 11268 4261 11271
rect 2464 11240 4261 11268
rect 2464 11228 2470 11240
rect 4249 11237 4261 11240
rect 4295 11237 4307 11271
rect 4249 11231 4307 11237
rect 4724 11240 4936 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 1452 11172 2452 11200
rect 1452 11160 1458 11172
rect 2424 11144 2452 11172
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 4724 11200 4752 11240
rect 2648 11172 4752 11200
rect 2648 11160 2654 11172
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 4908 11200 4936 11240
rect 7098 11228 7104 11280
rect 7156 11268 7162 11280
rect 7156 11240 9260 11268
rect 7156 11228 7162 11240
rect 6549 11203 6607 11209
rect 4908 11172 6500 11200
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11132 1731 11135
rect 2130 11132 2136 11144
rect 1719 11104 2136 11132
rect 1719 11101 1731 11104
rect 1673 11095 1731 11101
rect 2130 11092 2136 11104
rect 2188 11092 2194 11144
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 3510 11132 3516 11144
rect 2823 11104 3516 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 3510 11092 3516 11104
rect 3568 11092 3574 11144
rect 4062 11092 4068 11144
rect 4120 11092 4126 11144
rect 6178 11092 6184 11144
rect 6236 11092 6242 11144
rect 6472 11132 6500 11172
rect 6549 11169 6561 11203
rect 6595 11200 6607 11203
rect 7190 11200 7196 11212
rect 6595 11172 7196 11200
rect 6595 11169 6607 11172
rect 6549 11163 6607 11169
rect 7190 11160 7196 11172
rect 7248 11160 7254 11212
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 7800 11172 8309 11200
rect 7800 11160 7806 11172
rect 8297 11169 8309 11172
rect 8343 11169 8355 11203
rect 8297 11163 8355 11169
rect 8389 11203 8447 11209
rect 8389 11169 8401 11203
rect 8435 11169 8447 11203
rect 8389 11163 8447 11169
rect 7374 11132 7380 11144
rect 6472 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 8404 11132 8432 11163
rect 8570 11160 8576 11212
rect 8628 11200 8634 11212
rect 9125 11203 9183 11209
rect 9125 11200 9137 11203
rect 8628 11172 9137 11200
rect 8628 11160 8634 11172
rect 9125 11169 9137 11172
rect 9171 11169 9183 11203
rect 9125 11163 9183 11169
rect 9232 11144 9260 11240
rect 9306 11228 9312 11280
rect 9364 11268 9370 11280
rect 10778 11268 10784 11280
rect 9364 11240 10784 11268
rect 9364 11228 9370 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 11057 11271 11115 11277
rect 11057 11237 11069 11271
rect 11103 11268 11115 11271
rect 11146 11268 11152 11280
rect 11103 11240 11152 11268
rect 11103 11237 11115 11240
rect 11057 11231 11115 11237
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 12860 11240 13676 11268
rect 12860 11228 12866 11240
rect 9950 11160 9956 11212
rect 10008 11160 10014 11212
rect 10137 11203 10195 11209
rect 10137 11169 10149 11203
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 7892 11104 8432 11132
rect 7892 11092 7898 11104
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8938 11132 8944 11144
rect 8536 11104 8944 11132
rect 8536 11092 8542 11104
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9214 11092 9220 11144
rect 9272 11092 9278 11144
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 10042 11132 10048 11144
rect 9907 11104 10048 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 10042 11092 10048 11104
rect 10100 11092 10106 11144
rect 10152 11132 10180 11163
rect 11422 11160 11428 11212
rect 11480 11200 11486 11212
rect 12158 11200 12164 11212
rect 11480 11172 12164 11200
rect 11480 11160 11486 11172
rect 12158 11160 12164 11172
rect 12216 11160 12222 11212
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 13648 11209 13676 11240
rect 14182 11228 14188 11280
rect 14240 11268 14246 11280
rect 14369 11271 14427 11277
rect 14369 11268 14381 11271
rect 14240 11240 14381 11268
rect 14240 11228 14246 11240
rect 14369 11237 14381 11240
rect 14415 11268 14427 11271
rect 14550 11268 14556 11280
rect 14415 11240 14556 11268
rect 14415 11237 14427 11240
rect 14369 11231 14427 11237
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 16132 11212 16160 11308
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17386 11339 17444 11345
rect 17386 11336 17398 11339
rect 17000 11308 17398 11336
rect 17000 11296 17006 11308
rect 17386 11305 17398 11308
rect 17432 11305 17444 11339
rect 17386 11299 17444 11305
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 23201 11339 23259 11345
rect 23201 11336 23213 11339
rect 17828 11308 23213 11336
rect 17828 11296 17834 11308
rect 23201 11305 23213 11308
rect 23247 11305 23259 11339
rect 23201 11299 23259 11305
rect 25130 11296 25136 11348
rect 25188 11336 25194 11348
rect 25498 11336 25504 11348
rect 25188 11308 25504 11336
rect 25188 11296 25194 11308
rect 25498 11296 25504 11308
rect 25556 11296 25562 11348
rect 26329 11339 26387 11345
rect 26329 11305 26341 11339
rect 26375 11336 26387 11339
rect 27154 11336 27160 11348
rect 26375 11308 27160 11336
rect 26375 11305 26387 11308
rect 26329 11299 26387 11305
rect 27154 11296 27160 11308
rect 27212 11296 27218 11348
rect 32125 11339 32183 11345
rect 32125 11305 32137 11339
rect 32171 11336 32183 11339
rect 32214 11336 32220 11348
rect 32171 11308 32220 11336
rect 32171 11305 32183 11308
rect 32125 11299 32183 11305
rect 18598 11268 18604 11280
rect 18432 11240 18604 11268
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12308 11172 13277 11200
rect 12308 11160 12314 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 13814 11200 13820 11212
rect 13679 11172 13820 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 16114 11160 16120 11212
rect 16172 11200 16178 11212
rect 16393 11203 16451 11209
rect 16393 11200 16405 11203
rect 16172 11172 16405 11200
rect 16172 11160 16178 11172
rect 16393 11169 16405 11172
rect 16439 11169 16451 11203
rect 16393 11163 16451 11169
rect 17129 11203 17187 11209
rect 17129 11169 17141 11203
rect 17175 11200 17187 11203
rect 17402 11200 17408 11212
rect 17175 11172 17408 11200
rect 17175 11169 17187 11172
rect 17129 11163 17187 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18432 11200 18460 11240
rect 18598 11228 18604 11240
rect 18656 11268 18662 11280
rect 18877 11271 18935 11277
rect 18877 11268 18889 11271
rect 18656 11240 18889 11268
rect 18656 11228 18662 11240
rect 18877 11237 18889 11240
rect 18923 11237 18935 11271
rect 18877 11231 18935 11237
rect 20622 11228 20628 11280
rect 20680 11228 20686 11280
rect 22278 11228 22284 11280
rect 22336 11268 22342 11280
rect 25225 11271 25283 11277
rect 22336 11240 23796 11268
rect 22336 11228 22342 11240
rect 19610 11200 19616 11212
rect 17920 11172 18460 11200
rect 19306 11172 19616 11200
rect 17920 11160 17926 11172
rect 10778 11132 10784 11144
rect 10152 11104 10784 11132
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 10962 11092 10968 11144
rect 11020 11132 11026 11144
rect 11517 11135 11575 11141
rect 11517 11132 11529 11135
rect 11020 11104 11529 11132
rect 11020 11092 11026 11104
rect 11517 11101 11529 11104
rect 11563 11101 11575 11135
rect 11517 11095 11575 11101
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 14645 11135 14703 11141
rect 14645 11132 14657 11135
rect 14516 11104 14657 11132
rect 14516 11092 14522 11104
rect 14645 11101 14657 11104
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 18874 11092 18880 11144
rect 18932 11132 18938 11144
rect 19306 11132 19334 11172
rect 19610 11160 19616 11172
rect 19668 11160 19674 11212
rect 19702 11160 19708 11212
rect 19760 11200 19766 11212
rect 20165 11203 20223 11209
rect 20165 11200 20177 11203
rect 19760 11172 20177 11200
rect 19760 11160 19766 11172
rect 20165 11169 20177 11172
rect 20211 11169 20223 11203
rect 20165 11163 20223 11169
rect 20254 11160 20260 11212
rect 20312 11200 20318 11212
rect 20993 11203 21051 11209
rect 20993 11200 21005 11203
rect 20312 11172 21005 11200
rect 20312 11160 20318 11172
rect 20993 11169 21005 11172
rect 21039 11200 21051 11203
rect 21910 11200 21916 11212
rect 21039 11172 21916 11200
rect 21039 11169 21051 11172
rect 20993 11163 21051 11169
rect 21910 11160 21916 11172
rect 21968 11200 21974 11212
rect 22462 11200 22468 11212
rect 21968 11172 22468 11200
rect 21968 11160 21974 11172
rect 22462 11160 22468 11172
rect 22520 11160 22526 11212
rect 22738 11160 22744 11212
rect 22796 11160 22802 11212
rect 23382 11160 23388 11212
rect 23440 11200 23446 11212
rect 23768 11209 23796 11240
rect 25225 11237 25237 11271
rect 25271 11268 25283 11271
rect 26694 11268 26700 11280
rect 25271 11240 26700 11268
rect 25271 11237 25283 11240
rect 25225 11231 25283 11237
rect 26694 11228 26700 11240
rect 26752 11228 26758 11280
rect 27430 11228 27436 11280
rect 27488 11228 27494 11280
rect 28718 11228 28724 11280
rect 28776 11268 28782 11280
rect 29638 11268 29644 11280
rect 28776 11240 29644 11268
rect 28776 11228 28782 11240
rect 29638 11228 29644 11240
rect 29696 11228 29702 11280
rect 23661 11203 23719 11209
rect 23661 11200 23673 11203
rect 23440 11172 23673 11200
rect 23440 11160 23446 11172
rect 23661 11169 23673 11172
rect 23707 11169 23719 11203
rect 23661 11163 23719 11169
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11200 23811 11203
rect 23799 11172 25728 11200
rect 23799 11169 23811 11172
rect 23753 11163 23811 11169
rect 18932 11104 19334 11132
rect 18932 11092 18938 11104
rect 19426 11092 19432 11144
rect 19484 11092 19490 11144
rect 23566 11092 23572 11144
rect 23624 11092 23630 11144
rect 24578 11092 24584 11144
rect 24636 11092 24642 11144
rect 25700 11141 25728 11172
rect 25958 11160 25964 11212
rect 26016 11200 26022 11212
rect 29733 11203 29791 11209
rect 29733 11200 29745 11203
rect 26016 11172 29745 11200
rect 26016 11160 26022 11172
rect 29733 11169 29745 11172
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 25685 11135 25743 11141
rect 25685 11101 25697 11135
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 26789 11135 26847 11141
rect 26789 11101 26801 11135
rect 26835 11132 26847 11135
rect 27062 11132 27068 11144
rect 26835 11104 27068 11132
rect 26835 11101 26847 11104
rect 26789 11095 26847 11101
rect 27062 11092 27068 11104
rect 27120 11092 27126 11144
rect 27154 11092 27160 11144
rect 27212 11132 27218 11144
rect 28905 11135 28963 11141
rect 28905 11132 28917 11135
rect 27212 11104 28917 11132
rect 27212 11092 27218 11104
rect 28905 11101 28917 11104
rect 28951 11101 28963 11135
rect 32140 11132 32168 11299
rect 32214 11296 32220 11308
rect 32272 11296 32278 11348
rect 31142 11104 32168 11132
rect 28905 11095 28963 11101
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 5077 11067 5135 11073
rect 5077 11064 5089 11067
rect 4212 11036 5089 11064
rect 4212 11024 4218 11036
rect 5077 11033 5089 11036
rect 5123 11033 5135 11067
rect 5077 11027 5135 11033
rect 7098 11024 7104 11076
rect 7156 11024 7162 11076
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 9398 11064 9404 11076
rect 8251 11036 9404 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 9398 11024 9404 11036
rect 9456 11024 9462 11076
rect 10873 11067 10931 11073
rect 10873 11033 10885 11067
rect 10919 11064 10931 11067
rect 10919 11036 11008 11064
rect 10919 11033 10931 11036
rect 10873 11027 10931 11033
rect 2774 10956 2780 11008
rect 2832 10996 2838 11008
rect 6546 10996 6552 11008
rect 2832 10968 6552 10996
rect 2832 10956 2838 10968
rect 6546 10956 6552 10968
rect 6604 10996 6610 11008
rect 7558 10996 7564 11008
rect 6604 10968 7564 10996
rect 6604 10956 6610 10968
rect 7558 10956 7564 10968
rect 7616 10956 7622 11008
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7800 10968 7849 10996
rect 7800 10956 7806 10968
rect 7837 10965 7849 10968
rect 7883 10965 7895 10999
rect 7837 10959 7895 10965
rect 9490 10956 9496 11008
rect 9548 10956 9554 11008
rect 10980 10996 11008 11036
rect 11790 11024 11796 11076
rect 11848 11024 11854 11076
rect 12802 11024 12808 11076
rect 12860 11024 12866 11076
rect 14185 11067 14243 11073
rect 14185 11033 14197 11067
rect 14231 11064 14243 11067
rect 14366 11064 14372 11076
rect 14231 11036 14372 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 14366 11024 14372 11036
rect 14424 11024 14430 11076
rect 14918 11024 14924 11076
rect 14976 11024 14982 11076
rect 15378 11064 15384 11076
rect 15304 11036 15384 11064
rect 11974 10996 11980 11008
rect 10980 10968 11980 10996
rect 11974 10956 11980 10968
rect 12032 10956 12038 11008
rect 12434 10956 12440 11008
rect 12492 10996 12498 11008
rect 12710 10996 12716 11008
rect 12492 10968 12716 10996
rect 12492 10956 12498 10968
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14826 10996 14832 11008
rect 13872 10968 14832 10996
rect 13872 10956 13878 10968
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 15304 10996 15332 11036
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 16758 11024 16764 11076
rect 16816 11064 16822 11076
rect 18690 11064 18696 11076
rect 16816 11036 17356 11064
rect 18630 11036 18696 11064
rect 16816 11024 16822 11036
rect 16850 10996 16856 11008
rect 15304 10968 16856 10996
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 17328 10996 17356 11036
rect 18690 11024 18696 11036
rect 18748 11064 18754 11076
rect 19518 11064 19524 11076
rect 18748 11036 19524 11064
rect 18748 11024 18754 11036
rect 19518 11024 19524 11036
rect 19576 11024 19582 11076
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 21174 11064 21180 11076
rect 19668 11036 21180 11064
rect 19668 11024 19674 11036
rect 21174 11024 21180 11036
rect 21232 11024 21238 11076
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21358 11064 21364 11076
rect 21315 11036 21364 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 23106 11064 23112 11076
rect 22494 11036 23112 11064
rect 23106 11024 23112 11036
rect 23164 11064 23170 11076
rect 24210 11064 24216 11076
rect 23164 11036 24216 11064
rect 23164 11024 23170 11036
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 24854 11024 24860 11076
rect 24912 11064 24918 11076
rect 26694 11064 26700 11076
rect 24912 11036 26700 11064
rect 24912 11024 24918 11036
rect 26694 11024 26700 11036
rect 26752 11024 26758 11076
rect 27798 11064 27804 11076
rect 27356 11036 27804 11064
rect 20714 10996 20720 11008
rect 17328 10968 20720 10996
rect 20714 10956 20720 10968
rect 20772 10956 20778 11008
rect 23566 10956 23572 11008
rect 23624 10996 23630 11008
rect 24118 10996 24124 11008
rect 23624 10968 24124 10996
rect 23624 10956 23630 10968
rect 24118 10956 24124 10968
rect 24176 10956 24182 11008
rect 25406 10956 25412 11008
rect 25464 10996 25470 11008
rect 27356 10996 27384 11036
rect 27798 11024 27804 11036
rect 27856 11024 27862 11076
rect 27985 11067 28043 11073
rect 27985 11033 27997 11067
rect 28031 11033 28043 11067
rect 27985 11027 28043 11033
rect 28169 11067 28227 11073
rect 28169 11033 28181 11067
rect 28215 11064 28227 11067
rect 28626 11064 28632 11076
rect 28215 11036 28632 11064
rect 28215 11033 28227 11036
rect 28169 11027 28227 11033
rect 25464 10968 27384 10996
rect 25464 10956 25470 10968
rect 27706 10956 27712 11008
rect 27764 10996 27770 11008
rect 28000 10996 28028 11027
rect 28626 11024 28632 11036
rect 28684 11024 28690 11076
rect 28718 11024 28724 11076
rect 28776 11064 28782 11076
rect 29181 11067 29239 11073
rect 29181 11064 29193 11067
rect 28776 11036 29193 11064
rect 28776 11024 28782 11036
rect 29181 11033 29193 11036
rect 29227 11033 29239 11067
rect 29181 11027 29239 11033
rect 30006 11024 30012 11076
rect 30064 11024 30070 11076
rect 31294 11024 31300 11076
rect 31352 11064 31358 11076
rect 31757 11067 31815 11073
rect 31757 11064 31769 11067
rect 31352 11036 31769 11064
rect 31352 11024 31358 11036
rect 31757 11033 31769 11036
rect 31803 11064 31815 11067
rect 47762 11064 47768 11076
rect 31803 11036 47768 11064
rect 31803 11033 31815 11036
rect 31757 11027 31815 11033
rect 47762 11024 47768 11036
rect 47820 11024 47826 11076
rect 27764 10968 28028 10996
rect 27764 10956 27770 10968
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 1578 10752 1584 10804
rect 1636 10752 1642 10804
rect 6822 10792 6828 10804
rect 4172 10764 6828 10792
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1912 10628 1961 10656
rect 1912 10616 1918 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 3050 10616 3056 10668
rect 3108 10616 3114 10668
rect 4172 10665 4200 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 6914 10752 6920 10804
rect 6972 10752 6978 10804
rect 11514 10792 11520 10804
rect 8404 10764 11520 10792
rect 5997 10727 6055 10733
rect 5997 10693 6009 10727
rect 6043 10724 6055 10727
rect 8404 10724 8432 10764
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11698 10752 11704 10804
rect 11756 10752 11762 10804
rect 14458 10792 14464 10804
rect 12406 10764 14464 10792
rect 6043 10696 8432 10724
rect 6043 10693 6055 10696
rect 5997 10687 6055 10693
rect 9030 10684 9036 10736
rect 9088 10684 9094 10736
rect 9674 10684 9680 10736
rect 9732 10724 9738 10736
rect 10226 10724 10232 10736
rect 9732 10696 10232 10724
rect 9732 10684 9738 10696
rect 10226 10684 10232 10696
rect 10284 10684 10290 10736
rect 11054 10684 11060 10736
rect 11112 10724 11118 10736
rect 12406 10724 12434 10764
rect 14458 10752 14464 10764
rect 14516 10752 14522 10804
rect 14550 10752 14556 10804
rect 14608 10752 14614 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 15212 10764 16313 10792
rect 15212 10736 15240 10764
rect 16301 10761 16313 10764
rect 16347 10792 16359 10795
rect 18138 10792 18144 10804
rect 16347 10764 18144 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 19518 10792 19524 10804
rect 19444 10764 19524 10792
rect 11112 10696 11284 10724
rect 11112 10684 11118 10696
rect 4157 10659 4215 10665
rect 4157 10625 4169 10659
rect 4203 10625 4215 10659
rect 4157 10619 4215 10625
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5353 10659 5411 10665
rect 5353 10656 5365 10659
rect 5040 10628 5365 10656
rect 5040 10616 5046 10628
rect 5353 10625 5365 10628
rect 5399 10625 5411 10659
rect 5353 10619 5411 10625
rect 5442 10616 5448 10668
rect 5500 10656 5506 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 5500 10628 7021 10656
rect 5500 10616 5506 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 7009 10619 7067 10625
rect 9398 10616 9404 10668
rect 9456 10656 9462 10668
rect 9456 10628 9904 10656
rect 9456 10616 9462 10628
rect 1578 10548 1584 10600
rect 1636 10588 1642 10600
rect 4798 10588 4804 10600
rect 1636 10560 4804 10588
rect 1636 10548 1642 10560
rect 4798 10548 4804 10560
rect 4856 10548 4862 10600
rect 6730 10548 6736 10600
rect 6788 10588 6794 10600
rect 7098 10588 7104 10600
rect 6788 10560 7104 10588
rect 6788 10548 6794 10560
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 7190 10548 7196 10600
rect 7248 10548 7254 10600
rect 7650 10548 7656 10600
rect 7708 10588 7714 10600
rect 7745 10591 7803 10597
rect 7745 10588 7757 10591
rect 7708 10560 7757 10588
rect 7708 10548 7714 10560
rect 7745 10557 7757 10560
rect 7791 10557 7803 10591
rect 7745 10551 7803 10557
rect 1489 10523 1547 10529
rect 1489 10489 1501 10523
rect 1535 10520 1547 10523
rect 2958 10520 2964 10532
rect 1535 10492 2964 10520
rect 1535 10489 1547 10492
rect 1489 10483 1547 10489
rect 2958 10480 2964 10492
rect 3016 10480 3022 10532
rect 5166 10480 5172 10532
rect 5224 10520 5230 10532
rect 6914 10520 6920 10532
rect 5224 10492 6920 10520
rect 5224 10480 5230 10492
rect 6914 10480 6920 10492
rect 6972 10480 6978 10532
rect 2590 10412 2596 10464
rect 2648 10412 2654 10464
rect 2774 10412 2780 10464
rect 2832 10452 2838 10464
rect 3697 10455 3755 10461
rect 3697 10452 3709 10455
rect 2832 10424 3709 10452
rect 2832 10412 2838 10424
rect 3697 10421 3709 10424
rect 3743 10421 3755 10455
rect 3697 10415 3755 10421
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5902 10452 5908 10464
rect 4847 10424 5908 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6549 10455 6607 10461
rect 6549 10421 6561 10455
rect 6595 10452 6607 10455
rect 6822 10452 6828 10464
rect 6595 10424 6828 10452
rect 6595 10421 6607 10424
rect 6549 10415 6607 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 7760 10452 7788 10551
rect 8018 10548 8024 10600
rect 8076 10548 8082 10600
rect 9769 10591 9827 10597
rect 9769 10588 9781 10591
rect 9646 10560 9781 10588
rect 9122 10480 9128 10532
rect 9180 10520 9186 10532
rect 9646 10520 9674 10560
rect 9769 10557 9781 10560
rect 9815 10557 9827 10591
rect 9769 10551 9827 10557
rect 9180 10492 9674 10520
rect 9180 10480 9186 10492
rect 8478 10452 8484 10464
rect 7760 10424 8484 10452
rect 8478 10412 8484 10424
rect 8536 10452 8542 10464
rect 9766 10452 9772 10464
rect 8536 10424 9772 10452
rect 8536 10412 8542 10424
rect 9766 10412 9772 10424
rect 9824 10412 9830 10464
rect 9876 10452 9904 10628
rect 10594 10548 10600 10600
rect 10652 10588 10658 10600
rect 10962 10588 10968 10600
rect 10652 10560 10968 10588
rect 10652 10548 10658 10560
rect 10962 10548 10968 10560
rect 11020 10548 11026 10600
rect 11256 10588 11284 10696
rect 12268 10696 12434 10724
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 12268 10665 12296 10696
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 12860 10696 13018 10724
rect 12860 10684 12866 10696
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14921 10727 14979 10733
rect 14921 10724 14933 10727
rect 14148 10696 14933 10724
rect 14148 10684 14154 10696
rect 14921 10693 14933 10696
rect 14967 10724 14979 10727
rect 15194 10724 15200 10736
rect 14967 10696 15200 10724
rect 14967 10693 14979 10696
rect 14921 10687 14979 10693
rect 15194 10684 15200 10696
rect 15252 10684 15258 10736
rect 15749 10727 15807 10733
rect 15749 10693 15761 10727
rect 15795 10724 15807 10727
rect 16850 10724 16856 10736
rect 15795 10696 16856 10724
rect 15795 10693 15807 10696
rect 15749 10687 15807 10693
rect 16850 10684 16856 10696
rect 16908 10684 16914 10736
rect 17402 10684 17408 10736
rect 17460 10724 17466 10736
rect 17773 10727 17831 10733
rect 17773 10724 17785 10727
rect 17460 10696 17785 10724
rect 17460 10684 17466 10696
rect 17773 10693 17785 10696
rect 17819 10693 17831 10727
rect 19444 10724 19472 10764
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 21266 10752 21272 10804
rect 21324 10792 21330 10804
rect 22373 10795 22431 10801
rect 22373 10792 22385 10795
rect 21324 10764 22385 10792
rect 21324 10752 21330 10764
rect 22373 10761 22385 10764
rect 22419 10761 22431 10795
rect 22373 10755 22431 10761
rect 22465 10795 22523 10801
rect 22465 10761 22477 10795
rect 22511 10792 22523 10795
rect 22646 10792 22652 10804
rect 22511 10764 22652 10792
rect 22511 10761 22523 10764
rect 22465 10755 22523 10761
rect 22646 10752 22652 10764
rect 22704 10752 22710 10804
rect 22830 10752 22836 10804
rect 22888 10792 22894 10804
rect 29362 10792 29368 10804
rect 22888 10764 29368 10792
rect 22888 10752 22894 10764
rect 29362 10752 29368 10764
rect 29420 10752 29426 10804
rect 29457 10795 29515 10801
rect 29457 10761 29469 10795
rect 29503 10792 29515 10795
rect 30006 10792 30012 10804
rect 29503 10764 30012 10792
rect 29503 10761 29515 10764
rect 29457 10755 29515 10761
rect 30006 10752 30012 10764
rect 30064 10752 30070 10804
rect 20254 10724 20260 10736
rect 18998 10696 19472 10724
rect 19720 10696 20260 10724
rect 17773 10687 17831 10693
rect 12253 10659 12311 10665
rect 12253 10656 12265 10659
rect 11572 10628 12265 10656
rect 11572 10616 11578 10628
rect 12253 10625 12265 10628
rect 12299 10625 12311 10659
rect 12253 10619 12311 10625
rect 15930 10616 15936 10668
rect 15988 10656 15994 10668
rect 16117 10659 16175 10665
rect 16117 10656 16129 10659
rect 15988 10628 16129 10656
rect 15988 10616 15994 10628
rect 16117 10625 16129 10628
rect 16163 10625 16175 10659
rect 16117 10619 16175 10625
rect 17494 10616 17500 10668
rect 17552 10616 17558 10668
rect 19720 10665 19748 10696
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 21726 10724 21732 10736
rect 21206 10696 21732 10724
rect 21726 10684 21732 10696
rect 21784 10684 21790 10736
rect 22094 10684 22100 10736
rect 22152 10724 22158 10736
rect 24118 10724 24124 10736
rect 22152 10696 24124 10724
rect 22152 10684 22158 10696
rect 24118 10684 24124 10696
rect 24176 10684 24182 10736
rect 25590 10684 25596 10736
rect 25648 10724 25654 10736
rect 27249 10727 27307 10733
rect 25648 10696 25820 10724
rect 25648 10684 25654 10696
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10625 19763 10659
rect 19705 10619 19763 10625
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 23106 10656 23112 10668
rect 22888 10628 23112 10656
rect 22888 10616 22894 10628
rect 23106 10616 23112 10628
rect 23164 10616 23170 10668
rect 23477 10659 23535 10665
rect 23477 10625 23489 10659
rect 23523 10656 23535 10659
rect 23934 10656 23940 10668
rect 23523 10628 23940 10656
rect 23523 10625 23535 10628
rect 23477 10619 23535 10625
rect 23934 10616 23940 10628
rect 23992 10616 23998 10668
rect 24026 10616 24032 10668
rect 24084 10656 24090 10668
rect 24581 10659 24639 10665
rect 24581 10656 24593 10659
rect 24084 10628 24593 10656
rect 24084 10616 24090 10628
rect 24581 10625 24593 10628
rect 24627 10625 24639 10659
rect 24581 10619 24639 10625
rect 25222 10616 25228 10668
rect 25280 10616 25286 10668
rect 25685 10659 25743 10665
rect 25685 10625 25697 10659
rect 25731 10625 25743 10659
rect 25685 10619 25743 10625
rect 12066 10588 12072 10600
rect 11256 10560 12072 10588
rect 12066 10548 12072 10560
rect 12124 10548 12130 10600
rect 12529 10591 12587 10597
rect 12529 10557 12541 10591
rect 12575 10588 12587 10591
rect 14366 10588 14372 10600
rect 12575 10560 14372 10588
rect 12575 10557 12587 10560
rect 12529 10551 12587 10557
rect 14366 10548 14372 10560
rect 14424 10548 14430 10600
rect 14734 10548 14740 10600
rect 14792 10588 14798 10600
rect 16853 10591 16911 10597
rect 16853 10588 16865 10591
rect 14792 10560 16865 10588
rect 14792 10548 14798 10560
rect 16853 10557 16865 10560
rect 16899 10557 16911 10591
rect 18414 10588 18420 10600
rect 16853 10551 16911 10557
rect 16960 10560 18420 10588
rect 11882 10520 11888 10532
rect 11256 10492 11888 10520
rect 10870 10452 10876 10464
rect 9876 10424 10876 10452
rect 10870 10412 10876 10424
rect 10928 10412 10934 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11256 10452 11284 10492
rect 11882 10480 11888 10492
rect 11940 10520 11946 10532
rect 11940 10492 12112 10520
rect 11940 10480 11946 10492
rect 11112 10424 11284 10452
rect 11609 10455 11667 10461
rect 11112 10412 11118 10424
rect 11609 10421 11621 10455
rect 11655 10452 11667 10455
rect 11698 10452 11704 10464
rect 11655 10424 11704 10452
rect 11655 10421 11667 10424
rect 11609 10415 11667 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 11974 10412 11980 10464
rect 12032 10412 12038 10464
rect 12084 10452 12112 10492
rect 13538 10480 13544 10532
rect 13596 10520 13602 10532
rect 13596 10492 14780 10520
rect 13596 10480 13602 10492
rect 14752 10464 14780 10492
rect 15930 10480 15936 10532
rect 15988 10520 15994 10532
rect 16960 10520 16988 10560
rect 18414 10548 18420 10560
rect 18472 10548 18478 10600
rect 19981 10591 20039 10597
rect 19076 10560 19380 10588
rect 15988 10492 16988 10520
rect 15988 10480 15994 10492
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 12084 10424 14013 10452
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 14369 10455 14427 10461
rect 14369 10421 14381 10455
rect 14415 10452 14427 10455
rect 14550 10452 14556 10464
rect 14415 10424 14556 10452
rect 14415 10421 14427 10424
rect 14369 10415 14427 10421
rect 14550 10412 14556 10424
rect 14608 10412 14614 10464
rect 14734 10412 14740 10464
rect 14792 10412 14798 10464
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 16758 10452 16764 10464
rect 15160 10424 16764 10452
rect 15160 10412 15166 10424
rect 16758 10412 16764 10424
rect 16816 10412 16822 10464
rect 17034 10412 17040 10464
rect 17092 10452 17098 10464
rect 19076 10452 19104 10560
rect 19352 10520 19380 10560
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 22462 10588 22468 10600
rect 20027 10560 22468 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 22462 10548 22468 10560
rect 22520 10548 22526 10600
rect 22557 10591 22615 10597
rect 22557 10557 22569 10591
rect 22603 10557 22615 10591
rect 22557 10551 22615 10557
rect 24121 10591 24179 10597
rect 24121 10557 24133 10591
rect 24167 10588 24179 10591
rect 25700 10588 25728 10619
rect 24167 10560 25728 10588
rect 25792 10588 25820 10696
rect 27249 10693 27261 10727
rect 27295 10724 27307 10727
rect 27295 10696 35894 10724
rect 27295 10693 27307 10696
rect 27249 10687 27307 10693
rect 27430 10616 27436 10668
rect 27488 10616 27494 10668
rect 28810 10616 28816 10668
rect 28868 10616 28874 10668
rect 35866 10656 35894 10696
rect 36078 10656 36084 10668
rect 35866 10628 36084 10656
rect 36078 10616 36084 10628
rect 36136 10616 36142 10668
rect 32582 10588 32588 10600
rect 25792 10560 32588 10588
rect 24167 10557 24179 10560
rect 24121 10551 24179 10557
rect 19610 10520 19616 10532
rect 19352 10492 19616 10520
rect 19610 10480 19616 10492
rect 19668 10480 19674 10532
rect 21174 10480 21180 10532
rect 21232 10520 21238 10532
rect 22005 10523 22063 10529
rect 22005 10520 22017 10523
rect 21232 10492 22017 10520
rect 21232 10480 21238 10492
rect 22005 10489 22017 10492
rect 22051 10489 22063 10523
rect 22005 10483 22063 10489
rect 17092 10424 19104 10452
rect 19245 10455 19303 10461
rect 17092 10412 17098 10424
rect 19245 10421 19257 10455
rect 19291 10452 19303 10455
rect 20070 10452 20076 10464
rect 19291 10424 20076 10452
rect 19291 10421 19303 10424
rect 19245 10415 19303 10421
rect 20070 10412 20076 10424
rect 20128 10452 20134 10464
rect 20714 10452 20720 10464
rect 20128 10424 20720 10452
rect 20128 10412 20134 10424
rect 20714 10412 20720 10424
rect 20772 10412 20778 10464
rect 20990 10412 20996 10464
rect 21048 10452 21054 10464
rect 21453 10455 21511 10461
rect 21453 10452 21465 10455
rect 21048 10424 21465 10452
rect 21048 10412 21054 10424
rect 21453 10421 21465 10424
rect 21499 10452 21511 10455
rect 22572 10452 22600 10551
rect 32582 10548 32588 10560
rect 32640 10548 32646 10600
rect 24210 10480 24216 10532
rect 24268 10520 24274 10532
rect 26329 10523 26387 10529
rect 26329 10520 26341 10523
rect 24268 10492 26341 10520
rect 24268 10480 24274 10492
rect 26329 10489 26341 10492
rect 26375 10489 26387 10523
rect 28534 10520 28540 10532
rect 26329 10483 26387 10489
rect 26436 10492 28540 10520
rect 21499 10424 22600 10452
rect 21499 10421 21511 10424
rect 21453 10415 21511 10421
rect 23842 10412 23848 10464
rect 23900 10452 23906 10464
rect 26436 10452 26464 10492
rect 28534 10480 28540 10492
rect 28592 10480 28598 10532
rect 23900 10424 26464 10452
rect 23900 10412 23906 10424
rect 27706 10412 27712 10464
rect 27764 10412 27770 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 2314 10208 2320 10260
rect 2372 10248 2378 10260
rect 3142 10248 3148 10260
rect 2372 10220 3148 10248
rect 2372 10208 2378 10220
rect 3142 10208 3148 10220
rect 3200 10208 3206 10260
rect 3421 10251 3479 10257
rect 3421 10217 3433 10251
rect 3467 10248 3479 10251
rect 8018 10248 8024 10260
rect 3467 10220 8024 10248
rect 3467 10217 3479 10220
rect 3421 10211 3479 10217
rect 8018 10208 8024 10220
rect 8076 10208 8082 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 11054 10248 11060 10260
rect 8168 10220 11060 10248
rect 8168 10208 8174 10220
rect 11054 10208 11060 10220
rect 11112 10208 11118 10260
rect 11238 10208 11244 10260
rect 11296 10208 11302 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 15286 10248 15292 10260
rect 11388 10220 15292 10248
rect 11388 10208 11394 10220
rect 15286 10208 15292 10220
rect 15344 10208 15350 10260
rect 15838 10208 15844 10260
rect 15896 10248 15902 10260
rect 17954 10248 17960 10260
rect 15896 10220 17960 10248
rect 15896 10208 15902 10220
rect 17954 10208 17960 10220
rect 18012 10208 18018 10260
rect 18138 10208 18144 10260
rect 18196 10248 18202 10260
rect 19061 10251 19119 10257
rect 19061 10248 19073 10251
rect 18196 10220 19073 10248
rect 18196 10208 18202 10220
rect 19061 10217 19073 10220
rect 19107 10248 19119 10251
rect 19426 10248 19432 10260
rect 19107 10220 19432 10248
rect 19107 10217 19119 10220
rect 19061 10211 19119 10217
rect 19426 10208 19432 10220
rect 19484 10208 19490 10260
rect 19610 10208 19616 10260
rect 19668 10248 19674 10260
rect 20162 10248 20168 10260
rect 19668 10220 20168 10248
rect 19668 10208 19674 10220
rect 20162 10208 20168 10220
rect 20220 10208 20226 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 20864 10220 24348 10248
rect 20864 10208 20870 10220
rect 2222 10140 2228 10192
rect 2280 10180 2286 10192
rect 2958 10180 2964 10192
rect 2280 10152 2964 10180
rect 2280 10140 2286 10152
rect 2958 10140 2964 10152
rect 3016 10140 3022 10192
rect 3234 10140 3240 10192
rect 3292 10180 3298 10192
rect 3786 10180 3792 10192
rect 3292 10152 3792 10180
rect 3292 10140 3298 10152
rect 3786 10140 3792 10152
rect 3844 10140 3850 10192
rect 3973 10183 4031 10189
rect 3973 10149 3985 10183
rect 4019 10180 4031 10183
rect 4062 10180 4068 10192
rect 4019 10152 4068 10180
rect 4019 10149 4031 10152
rect 3973 10143 4031 10149
rect 4062 10140 4068 10152
rect 4120 10140 4126 10192
rect 4338 10140 4344 10192
rect 4396 10180 4402 10192
rect 7193 10183 7251 10189
rect 7193 10180 7205 10183
rect 4396 10152 7205 10180
rect 4396 10140 4402 10152
rect 7193 10149 7205 10152
rect 7239 10149 7251 10183
rect 7193 10143 7251 10149
rect 7300 10152 9260 10180
rect 6089 10115 6147 10121
rect 2792 10084 6040 10112
rect 2792 10053 2820 10084
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 2777 10047 2835 10053
rect 2777 10013 2789 10047
rect 2823 10013 2835 10047
rect 2777 10007 2835 10013
rect 4249 10047 4307 10053
rect 4249 10013 4261 10047
rect 4295 10013 4307 10047
rect 4249 10007 4307 10013
rect 1688 9976 1716 10007
rect 4062 9976 4068 9988
rect 1688 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 4264 9976 4292 10007
rect 5350 10004 5356 10056
rect 5408 10044 5414 10056
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 5408 10016 5457 10044
rect 5408 10004 5414 10016
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 6012 10044 6040 10084
rect 6089 10081 6101 10115
rect 6135 10112 6147 10115
rect 6730 10112 6736 10124
rect 6135 10084 6736 10112
rect 6135 10081 6147 10084
rect 6089 10075 6147 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 6270 10044 6276 10056
rect 6012 10016 6276 10044
rect 5445 10007 5503 10013
rect 6270 10004 6276 10016
rect 6328 10004 6334 10056
rect 6549 10047 6607 10053
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 7300 10044 7328 10152
rect 8202 10072 8208 10124
rect 8260 10112 8266 10124
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 8260 10084 8309 10112
rect 8260 10072 8266 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 8297 10075 8355 10081
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 6595 10016 7328 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 7558 10004 7564 10056
rect 7616 10044 7622 10056
rect 8404 10044 8432 10075
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 9030 10112 9036 10124
rect 8904 10084 9036 10112
rect 8904 10072 8910 10084
rect 9030 10072 9036 10084
rect 9088 10072 9094 10124
rect 9232 10112 9260 10152
rect 10778 10140 10784 10192
rect 10836 10180 10842 10192
rect 10873 10183 10931 10189
rect 10873 10180 10885 10183
rect 10836 10152 10885 10180
rect 10836 10140 10842 10152
rect 10873 10149 10885 10152
rect 10919 10149 10931 10183
rect 10873 10143 10931 10149
rect 11348 10152 11652 10180
rect 11348 10124 11376 10152
rect 11054 10112 11060 10124
rect 9232 10084 11060 10112
rect 11054 10072 11060 10084
rect 11112 10072 11118 10124
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 11624 10112 11652 10152
rect 13814 10140 13820 10192
rect 13872 10140 13878 10192
rect 15930 10140 15936 10192
rect 15988 10180 15994 10192
rect 16209 10183 16267 10189
rect 16209 10180 16221 10183
rect 15988 10152 16221 10180
rect 15988 10140 15994 10152
rect 16209 10149 16221 10152
rect 16255 10149 16267 10183
rect 16209 10143 16267 10149
rect 18230 10140 18236 10192
rect 18288 10180 18294 10192
rect 18693 10183 18751 10189
rect 18693 10180 18705 10183
rect 18288 10152 18705 10180
rect 18288 10140 18294 10152
rect 18693 10149 18705 10152
rect 18739 10149 18751 10183
rect 18693 10143 18751 10149
rect 23842 10140 23848 10192
rect 23900 10140 23906 10192
rect 13541 10115 13599 10121
rect 13541 10112 13553 10115
rect 11624 10084 13553 10112
rect 13541 10081 13553 10084
rect 13587 10112 13599 10115
rect 14090 10112 14096 10124
rect 13587 10084 14096 10112
rect 13587 10081 13599 10084
rect 13541 10075 13599 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 16669 10115 16727 10121
rect 16669 10081 16681 10115
rect 16715 10112 16727 10115
rect 17494 10112 17500 10124
rect 16715 10084 17500 10112
rect 16715 10081 16727 10084
rect 16669 10075 16727 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 17586 10072 17592 10124
rect 17644 10112 17650 10124
rect 18417 10115 18475 10121
rect 18417 10112 18429 10115
rect 17644 10084 18429 10112
rect 17644 10072 17650 10084
rect 18417 10081 18429 10084
rect 18463 10112 18475 10115
rect 19426 10112 19432 10124
rect 18463 10084 19432 10112
rect 18463 10081 18475 10084
rect 18417 10075 18475 10081
rect 19426 10072 19432 10084
rect 19484 10072 19490 10124
rect 19797 10115 19855 10121
rect 19797 10081 19809 10115
rect 19843 10112 19855 10115
rect 24210 10112 24216 10124
rect 19843 10084 24216 10112
rect 19843 10081 19855 10084
rect 19797 10075 19855 10081
rect 24210 10072 24216 10084
rect 24268 10072 24274 10124
rect 24320 10112 24348 10220
rect 24670 10140 24676 10192
rect 24728 10180 24734 10192
rect 27203 10183 27261 10189
rect 27203 10180 27215 10183
rect 24728 10152 27215 10180
rect 24728 10140 24734 10152
rect 27203 10149 27215 10152
rect 27249 10149 27261 10183
rect 27203 10143 27261 10149
rect 30374 10112 30380 10124
rect 24320 10084 25452 10112
rect 7616 10016 8432 10044
rect 7616 10004 7622 10016
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8536 10016 9137 10044
rect 8536 10004 8542 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 14458 10004 14464 10056
rect 14516 10004 14522 10056
rect 19521 10047 19579 10053
rect 19521 10013 19533 10047
rect 19567 10013 19579 10047
rect 19521 10007 19579 10013
rect 22097 10047 22155 10053
rect 22097 10013 22109 10047
rect 22143 10044 22155 10047
rect 22738 10044 22744 10056
rect 22143 10016 22744 10044
rect 22143 10013 22155 10016
rect 22097 10007 22155 10013
rect 8110 9976 8116 9988
rect 4264 9948 8116 9976
rect 8110 9936 8116 9948
rect 8168 9936 8174 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9401 9979 9459 9985
rect 9401 9976 9413 9979
rect 8444 9948 9413 9976
rect 8444 9936 8450 9948
rect 9401 9945 9413 9948
rect 9447 9945 9459 9979
rect 11793 9979 11851 9985
rect 11793 9976 11805 9979
rect 9401 9939 9459 9945
rect 9600 9948 9890 9976
rect 10704 9948 11805 9976
rect 2314 9868 2320 9920
rect 2372 9868 2378 9920
rect 4893 9911 4951 9917
rect 4893 9877 4905 9911
rect 4939 9908 4951 9911
rect 5442 9908 5448 9920
rect 4939 9880 5448 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5442 9868 5448 9880
rect 5500 9868 5506 9920
rect 7374 9868 7380 9920
rect 7432 9908 7438 9920
rect 7469 9911 7527 9917
rect 7469 9908 7481 9911
rect 7432 9880 7481 9908
rect 7432 9868 7438 9880
rect 7469 9877 7481 9880
rect 7515 9877 7527 9911
rect 7469 9871 7527 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 7837 9911 7895 9917
rect 7837 9908 7849 9911
rect 7800 9880 7849 9908
rect 7800 9868 7806 9880
rect 7837 9877 7849 9880
rect 7883 9877 7895 9911
rect 7837 9871 7895 9877
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 8570 9908 8576 9920
rect 8251 9880 8576 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8570 9868 8576 9880
rect 8628 9868 8634 9920
rect 8846 9868 8852 9920
rect 8904 9908 8910 9920
rect 9600 9908 9628 9948
rect 8904 9880 9628 9908
rect 8904 9868 8910 9880
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10704 9908 10732 9948
rect 11793 9945 11805 9948
rect 11839 9945 11851 9979
rect 11793 9939 11851 9945
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 11940 9948 12282 9976
rect 13648 9948 14136 9976
rect 11940 9936 11946 9948
rect 9732 9880 10732 9908
rect 12176 9908 12204 9948
rect 12710 9908 12716 9920
rect 12176 9880 12716 9908
rect 9732 9868 9738 9880
rect 12710 9868 12716 9880
rect 12768 9868 12774 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13265 9911 13323 9917
rect 13265 9908 13277 9911
rect 13228 9880 13277 9908
rect 13228 9868 13234 9880
rect 13265 9877 13277 9880
rect 13311 9877 13323 9911
rect 13265 9871 13323 9877
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 13648 9908 13676 9948
rect 14108 9920 14136 9948
rect 14734 9936 14740 9988
rect 14792 9936 14798 9988
rect 15378 9936 15384 9988
rect 15436 9936 15442 9988
rect 16942 9936 16948 9988
rect 17000 9936 17006 9988
rect 18690 9976 18696 9988
rect 18170 9948 18696 9976
rect 18690 9936 18696 9948
rect 18748 9936 18754 9988
rect 19536 9976 19564 10007
rect 22738 10004 22744 10016
rect 22796 10004 22802 10056
rect 23201 10047 23259 10053
rect 23201 10013 23213 10047
rect 23247 10044 23259 10047
rect 23290 10044 23296 10056
rect 23247 10016 23296 10044
rect 23247 10013 23259 10016
rect 23201 10007 23259 10013
rect 23290 10004 23296 10016
rect 23348 10004 23354 10056
rect 24026 10004 24032 10056
rect 24084 10004 24090 10056
rect 24949 10047 25007 10053
rect 24949 10013 24961 10047
rect 24995 10044 25007 10047
rect 25314 10044 25320 10056
rect 24995 10016 25320 10044
rect 24995 10013 25007 10016
rect 24949 10007 25007 10013
rect 25314 10004 25320 10016
rect 25372 10004 25378 10056
rect 25424 10053 25452 10084
rect 26528 10084 30380 10112
rect 25409 10047 25467 10053
rect 25409 10013 25421 10047
rect 25455 10013 25467 10047
rect 25409 10007 25467 10013
rect 19702 9976 19708 9988
rect 19536 9948 19708 9976
rect 19702 9936 19708 9948
rect 19760 9936 19766 9988
rect 21726 9976 21732 9988
rect 21022 9948 21732 9976
rect 21726 9936 21732 9948
rect 21784 9936 21790 9988
rect 22278 9936 22284 9988
rect 22336 9976 22342 9988
rect 24044 9976 24072 10004
rect 26528 9976 26556 10084
rect 30374 10072 30380 10084
rect 30432 10072 30438 10124
rect 26973 10047 27031 10053
rect 26973 10044 26985 10047
rect 22336 9948 24072 9976
rect 24780 9948 26556 9976
rect 26620 10016 26985 10044
rect 22336 9936 22342 9948
rect 13596 9880 13676 9908
rect 13596 9868 13602 9880
rect 14090 9868 14096 9920
rect 14148 9868 14154 9920
rect 14185 9911 14243 9917
rect 14185 9877 14197 9911
rect 14231 9908 14243 9911
rect 14826 9908 14832 9920
rect 14231 9880 14832 9908
rect 14231 9877 14243 9880
rect 14185 9871 14243 9877
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 15470 9868 15476 9920
rect 15528 9908 15534 9920
rect 17678 9908 17684 9920
rect 15528 9880 17684 9908
rect 15528 9868 15534 9880
rect 17678 9868 17684 9880
rect 17736 9868 17742 9920
rect 17954 9868 17960 9920
rect 18012 9908 18018 9920
rect 19518 9908 19524 9920
rect 18012 9880 19524 9908
rect 18012 9868 18018 9880
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 19886 9868 19892 9920
rect 19944 9908 19950 9920
rect 20714 9908 20720 9920
rect 19944 9880 20720 9908
rect 19944 9868 19950 9880
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 21266 9868 21272 9920
rect 21324 9868 21330 9920
rect 22738 9868 22744 9920
rect 22796 9868 22802 9920
rect 24780 9917 24808 9948
rect 26620 9920 26648 10016
rect 26973 10013 26985 10016
rect 27019 10013 27031 10047
rect 26973 10007 27031 10013
rect 26694 9936 26700 9988
rect 26752 9976 26758 9988
rect 33318 9976 33324 9988
rect 26752 9948 33324 9976
rect 26752 9936 26758 9948
rect 33318 9936 33324 9948
rect 33376 9936 33382 9988
rect 24765 9911 24823 9917
rect 24765 9877 24777 9911
rect 24811 9877 24823 9911
rect 24765 9871 24823 9877
rect 26050 9868 26056 9920
rect 26108 9868 26114 9920
rect 26602 9868 26608 9920
rect 26660 9868 26666 9920
rect 28261 9911 28319 9917
rect 28261 9877 28273 9911
rect 28307 9908 28319 9911
rect 28442 9908 28448 9920
rect 28307 9880 28448 9908
rect 28307 9877 28319 9880
rect 28261 9871 28319 9877
rect 28442 9868 28448 9880
rect 28500 9868 28506 9920
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 1486 9664 1492 9716
rect 1544 9704 1550 9716
rect 2682 9704 2688 9716
rect 1544 9676 2688 9704
rect 1544 9664 1550 9676
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 3694 9664 3700 9716
rect 3752 9704 3758 9716
rect 6549 9707 6607 9713
rect 3752 9676 4568 9704
rect 3752 9664 3758 9676
rect 1946 9596 1952 9648
rect 2004 9636 2010 9648
rect 2866 9636 2872 9648
rect 2004 9608 2872 9636
rect 2004 9596 2010 9608
rect 2866 9596 2872 9608
rect 2924 9596 2930 9648
rect 658 9528 664 9580
rect 716 9568 722 9580
rect 842 9568 848 9580
rect 716 9540 848 9568
rect 716 9528 722 9540
rect 842 9528 848 9540
rect 900 9528 906 9580
rect 2041 9571 2099 9577
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2222 9568 2228 9580
rect 2087 9540 2228 9568
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9568 3203 9571
rect 3694 9568 3700 9580
rect 3191 9540 3700 9568
rect 3191 9537 3203 9540
rect 3145 9531 3203 9537
rect 3694 9528 3700 9540
rect 3752 9528 3758 9580
rect 4246 9528 4252 9580
rect 4304 9528 4310 9580
rect 4540 9568 4568 9676
rect 6549 9673 6561 9707
rect 6595 9674 6607 9707
rect 6595 9673 6629 9674
rect 6549 9667 6629 9673
rect 5626 9596 5632 9648
rect 5684 9636 5690 9648
rect 5684 9608 6040 9636
rect 5684 9596 5690 9608
rect 6012 9577 6040 9608
rect 6454 9596 6460 9648
rect 6512 9636 6518 9648
rect 6564 9646 6629 9667
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 9398 9704 9404 9716
rect 6972 9676 9404 9704
rect 6972 9664 6978 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 12066 9704 12072 9716
rect 9548 9676 12072 9704
rect 9548 9664 9554 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 12158 9664 12164 9716
rect 12216 9704 12222 9716
rect 12216 9676 13308 9704
rect 12216 9664 12222 9676
rect 6564 9636 6592 9646
rect 8662 9636 8668 9648
rect 6512 9608 6592 9636
rect 8496 9608 8668 9636
rect 6512 9596 6518 9608
rect 5353 9571 5411 9577
rect 5353 9568 5365 9571
rect 4540 9540 5365 9568
rect 5353 9537 5365 9540
rect 5399 9537 5411 9571
rect 5353 9531 5411 9537
rect 5997 9571 6055 9577
rect 5997 9537 6009 9571
rect 6043 9537 6055 9571
rect 5997 9531 6055 9537
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9568 6791 9571
rect 7374 9568 7380 9580
rect 6779 9540 7380 9568
rect 6779 9537 6791 9540
rect 6733 9531 6791 9537
rect 7374 9528 7380 9540
rect 7432 9528 7438 9580
rect 7558 9528 7564 9580
rect 7616 9528 7622 9580
rect 7653 9571 7711 9577
rect 7653 9537 7665 9571
rect 7699 9568 7711 9571
rect 8496 9568 8524 9608
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 8904 9608 9246 9636
rect 8904 9596 8910 9608
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 11241 9639 11299 9645
rect 11241 9636 11253 9639
rect 10284 9608 11253 9636
rect 10284 9596 10290 9608
rect 11241 9605 11253 9608
rect 11287 9636 11299 9639
rect 11330 9636 11336 9648
rect 11287 9608 11336 9636
rect 11287 9605 11299 9608
rect 11241 9599 11299 9605
rect 11330 9596 11336 9608
rect 11388 9596 11394 9648
rect 11882 9596 11888 9648
rect 11940 9636 11946 9648
rect 11940 9608 12466 9636
rect 11940 9596 11946 9608
rect 7699 9540 8524 9568
rect 7699 9537 7711 9540
rect 7653 9531 7711 9537
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11701 9571 11759 9577
rect 11701 9568 11713 9571
rect 11572 9540 11713 9568
rect 11572 9528 11578 9540
rect 11701 9537 11713 9540
rect 11747 9537 11759 9571
rect 11701 9531 11759 9537
rect 474 9460 480 9512
rect 532 9500 538 9512
rect 3789 9503 3847 9509
rect 3789 9500 3801 9503
rect 532 9472 3801 9500
rect 532 9460 538 9472
rect 3789 9469 3801 9472
rect 3835 9469 3847 9503
rect 3789 9463 3847 9469
rect 4893 9503 4951 9509
rect 4893 9469 4905 9503
rect 4939 9500 4951 9503
rect 5626 9500 5632 9512
rect 4939 9472 5632 9500
rect 4939 9469 4951 9472
rect 4893 9463 4951 9469
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 6822 9460 6828 9512
rect 6880 9500 6886 9512
rect 7745 9503 7803 9509
rect 7745 9500 7757 9503
rect 6880 9472 7757 9500
rect 6880 9460 6886 9472
rect 7745 9469 7757 9472
rect 7791 9469 7803 9503
rect 7745 9463 7803 9469
rect 8478 9460 8484 9512
rect 8536 9460 8542 9512
rect 8757 9503 8815 9509
rect 8757 9500 8769 9503
rect 8588 9472 8769 9500
rect 1394 9392 1400 9444
rect 1452 9392 1458 9444
rect 1581 9435 1639 9441
rect 1581 9401 1593 9435
rect 1627 9432 1639 9435
rect 3234 9432 3240 9444
rect 1627 9404 3240 9432
rect 1627 9401 1639 9404
rect 1581 9395 1639 9401
rect 3234 9392 3240 9404
rect 3292 9392 3298 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 5074 9432 5080 9444
rect 4120 9404 5080 9432
rect 4120 9392 4126 9404
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 7098 9392 7104 9444
rect 7156 9432 7162 9444
rect 8588 9432 8616 9472
rect 8757 9469 8769 9472
rect 8803 9469 8815 9503
rect 8757 9463 8815 9469
rect 9214 9460 9220 9512
rect 9272 9500 9278 9512
rect 10965 9503 11023 9509
rect 10965 9500 10977 9503
rect 9272 9472 10977 9500
rect 9272 9460 9278 9472
rect 10965 9469 10977 9472
rect 11011 9469 11023 9503
rect 10965 9463 11023 9469
rect 11146 9460 11152 9512
rect 11204 9500 11210 9512
rect 12066 9500 12072 9512
rect 11204 9472 12072 9500
rect 11204 9460 11210 9472
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12526 9460 12532 9512
rect 12584 9500 12590 9512
rect 13170 9500 13176 9512
rect 12584 9472 13176 9500
rect 12584 9460 12590 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13280 9500 13308 9676
rect 13354 9664 13360 9716
rect 13412 9704 13418 9716
rect 13538 9704 13544 9716
rect 13412 9676 13544 9704
rect 13412 9664 13418 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 14458 9664 14464 9716
rect 14516 9704 14522 9716
rect 16850 9704 16856 9716
rect 14516 9676 16856 9704
rect 14516 9664 14522 9676
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 18690 9704 18696 9716
rect 17368 9676 18696 9704
rect 17368 9664 17374 9676
rect 14476 9577 14504 9664
rect 14734 9596 14740 9648
rect 14792 9596 14798 9648
rect 15378 9596 15384 9648
rect 15436 9596 15442 9648
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 17512 9636 17540 9676
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 27801 9707 27859 9713
rect 22612 9676 23888 9704
rect 22612 9664 22618 9676
rect 17092 9608 17618 9636
rect 17092 9596 17098 9608
rect 18598 9596 18604 9648
rect 18656 9636 18662 9648
rect 19058 9636 19064 9648
rect 18656 9608 19064 9636
rect 18656 9596 18662 9608
rect 19058 9596 19064 9608
rect 19116 9596 19122 9648
rect 19889 9639 19947 9645
rect 19889 9605 19901 9639
rect 19935 9636 19947 9639
rect 23566 9636 23572 9648
rect 19935 9608 23572 9636
rect 19935 9605 19947 9608
rect 19889 9599 19947 9605
rect 23566 9596 23572 9608
rect 23624 9596 23630 9648
rect 23860 9645 23888 9676
rect 27801 9673 27813 9707
rect 27847 9704 27859 9707
rect 28810 9704 28816 9716
rect 27847 9676 28816 9704
rect 27847 9673 27859 9676
rect 27801 9667 27859 9673
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 23845 9639 23903 9645
rect 23845 9605 23857 9639
rect 23891 9605 23903 9639
rect 27614 9636 27620 9648
rect 23845 9599 23903 9605
rect 24504 9608 27620 9636
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 14461 9531 14519 9537
rect 18414 9528 18420 9580
rect 18472 9568 18478 9580
rect 19797 9571 19855 9577
rect 19797 9568 19809 9571
rect 18472 9540 19809 9568
rect 18472 9528 18478 9540
rect 19797 9537 19809 9540
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 20622 9528 20628 9580
rect 20680 9528 20686 9580
rect 21450 9528 21456 9580
rect 21508 9568 21514 9580
rect 22005 9571 22063 9577
rect 22005 9568 22017 9571
rect 21508 9540 22017 9568
rect 21508 9528 21514 9540
rect 22005 9537 22017 9540
rect 22051 9537 22063 9571
rect 22005 9531 22063 9537
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9568 23259 9571
rect 24504 9568 24532 9608
rect 27614 9596 27620 9608
rect 27672 9596 27678 9648
rect 27706 9596 27712 9648
rect 27764 9636 27770 9648
rect 32030 9636 32036 9648
rect 27764 9608 32036 9636
rect 27764 9596 27770 9608
rect 32030 9596 32036 9608
rect 32088 9596 32094 9648
rect 23247 9540 24532 9568
rect 24581 9571 24639 9577
rect 23247 9537 23259 9540
rect 23201 9531 23259 9537
rect 24581 9537 24593 9571
rect 24627 9568 24639 9571
rect 25222 9568 25228 9580
rect 24627 9540 25228 9568
rect 24627 9537 24639 9540
rect 24581 9531 24639 9537
rect 25222 9528 25228 9540
rect 25280 9528 25286 9580
rect 25314 9528 25320 9580
rect 25372 9568 25378 9580
rect 25685 9571 25743 9577
rect 25685 9568 25697 9571
rect 25372 9540 25697 9568
rect 25372 9528 25378 9540
rect 25685 9537 25697 9540
rect 25731 9537 25743 9571
rect 25685 9531 25743 9537
rect 26326 9528 26332 9580
rect 26384 9568 26390 9580
rect 27157 9571 27215 9577
rect 27157 9568 27169 9571
rect 26384 9540 27169 9568
rect 26384 9528 26390 9540
rect 27157 9537 27169 9540
rect 27203 9537 27215 9571
rect 27157 9531 27215 9537
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 13280 9472 16221 9500
rect 16209 9469 16221 9472
rect 16255 9469 16267 9503
rect 16209 9463 16267 9469
rect 16850 9460 16856 9512
rect 16908 9460 16914 9512
rect 17129 9503 17187 9509
rect 17129 9469 17141 9503
rect 17175 9500 17187 9503
rect 20073 9503 20131 9509
rect 17175 9472 19656 9500
rect 17175 9469 17187 9472
rect 17129 9463 17187 9469
rect 7156 9404 8616 9432
rect 7156 9392 7162 9404
rect 11514 9392 11520 9444
rect 11572 9432 11578 9444
rect 11572 9404 11836 9432
rect 11572 9392 11578 9404
rect 934 9324 940 9376
rect 992 9364 998 9376
rect 1412 9364 1440 9392
rect 1673 9367 1731 9373
rect 1673 9364 1685 9367
rect 992 9336 1685 9364
rect 992 9324 998 9336
rect 1673 9333 1685 9336
rect 1719 9333 1731 9367
rect 1673 9327 1731 9333
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 2406 9364 2412 9376
rect 1912 9336 2412 9364
rect 1912 9324 1918 9336
rect 2406 9324 2412 9336
rect 2464 9324 2470 9376
rect 2682 9324 2688 9376
rect 2740 9324 2746 9376
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 5258 9364 5264 9376
rect 4856 9336 5264 9364
rect 4856 9324 4862 9336
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 5776 9336 7205 9364
rect 5776 9324 5782 9336
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 7193 9327 7251 9333
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 10042 9364 10048 9376
rect 9824 9336 10048 9364
rect 9824 9324 9830 9336
rect 10042 9324 10048 9336
rect 10100 9324 10106 9376
rect 10134 9324 10140 9376
rect 10192 9364 10198 9376
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 10192 9336 10241 9364
rect 10192 9324 10198 9336
rect 10229 9333 10241 9336
rect 10275 9333 10287 9367
rect 11808 9364 11836 9404
rect 13078 9392 13084 9444
rect 13136 9432 13142 9444
rect 13725 9435 13783 9441
rect 13725 9432 13737 9435
rect 13136 9404 13737 9432
rect 13136 9392 13142 9404
rect 13725 9401 13737 9404
rect 13771 9432 13783 9435
rect 13771 9404 14596 9432
rect 13771 9401 13783 9404
rect 13725 9395 13783 9401
rect 14568 9376 14596 9404
rect 15838 9392 15844 9444
rect 15896 9432 15902 9444
rect 16022 9432 16028 9444
rect 15896 9404 16028 9432
rect 15896 9392 15902 9404
rect 16022 9392 16028 9404
rect 16080 9392 16086 9444
rect 19334 9392 19340 9444
rect 19392 9432 19398 9444
rect 19429 9435 19487 9441
rect 19429 9432 19441 9435
rect 19392 9404 19441 9432
rect 19392 9392 19398 9404
rect 19429 9401 19441 9404
rect 19475 9401 19487 9435
rect 19628 9432 19656 9472
rect 20073 9469 20085 9503
rect 20119 9500 20131 9503
rect 21266 9500 21272 9512
rect 20119 9472 21272 9500
rect 20119 9469 20131 9472
rect 20073 9463 20131 9469
rect 21266 9460 21272 9472
rect 21324 9460 21330 9512
rect 21634 9460 21640 9512
rect 21692 9500 21698 9512
rect 21692 9472 25268 9500
rect 21692 9460 21698 9472
rect 23750 9432 23756 9444
rect 19628 9404 23756 9432
rect 19429 9395 19487 9401
rect 23750 9392 23756 9404
rect 23808 9392 23814 9444
rect 25240 9441 25268 9472
rect 26142 9460 26148 9512
rect 26200 9500 26206 9512
rect 31846 9500 31852 9512
rect 26200 9472 31852 9500
rect 26200 9460 26206 9472
rect 31846 9460 31852 9472
rect 31904 9460 31910 9512
rect 25225 9435 25283 9441
rect 25225 9401 25237 9435
rect 25271 9401 25283 9435
rect 25225 9395 25283 9401
rect 26234 9392 26240 9444
rect 26292 9432 26298 9444
rect 26329 9435 26387 9441
rect 26329 9432 26341 9435
rect 26292 9404 26341 9432
rect 26292 9392 26298 9404
rect 26329 9401 26341 9404
rect 26375 9401 26387 9435
rect 26329 9395 26387 9401
rect 11958 9367 12016 9373
rect 11958 9364 11970 9367
rect 11808 9336 11970 9364
rect 10229 9327 10287 9333
rect 11958 9333 11970 9336
rect 12004 9333 12016 9367
rect 11958 9327 12016 9333
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 13449 9367 13507 9373
rect 13449 9364 13461 9367
rect 12124 9336 13461 9364
rect 12124 9324 12130 9336
rect 13449 9333 13461 9336
rect 13495 9333 13507 9367
rect 13449 9327 13507 9333
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 13909 9367 13967 9373
rect 13909 9364 13921 9367
rect 13872 9336 13921 9364
rect 13872 9324 13878 9336
rect 13909 9333 13921 9336
rect 13955 9333 13967 9367
rect 13909 9327 13967 9333
rect 14182 9324 14188 9376
rect 14240 9324 14246 9376
rect 14550 9324 14556 9376
rect 14608 9324 14614 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 18138 9364 18144 9376
rect 17276 9336 18144 9364
rect 17276 9324 17282 9336
rect 18138 9324 18144 9336
rect 18196 9364 18202 9376
rect 18601 9367 18659 9373
rect 18601 9364 18613 9367
rect 18196 9336 18613 9364
rect 18196 9324 18202 9336
rect 18601 9333 18613 9336
rect 18647 9333 18659 9367
rect 18601 9327 18659 9333
rect 20530 9324 20536 9376
rect 20588 9364 20594 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20588 9336 21281 9364
rect 20588 9324 20594 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 22649 9367 22707 9373
rect 22649 9333 22661 9367
rect 22695 9364 22707 9367
rect 26786 9364 26792 9376
rect 22695 9336 26792 9364
rect 22695 9333 22707 9336
rect 22649 9327 22707 9333
rect 26786 9324 26792 9336
rect 26844 9324 26850 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 1210 9120 1216 9172
rect 1268 9160 1274 9172
rect 2222 9160 2228 9172
rect 1268 9132 2228 9160
rect 1268 9120 1274 9132
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 3786 9120 3792 9172
rect 3844 9120 3850 9172
rect 6362 9160 6368 9172
rect 4264 9132 6368 9160
rect 2317 9095 2375 9101
rect 2317 9061 2329 9095
rect 2363 9092 2375 9095
rect 4264 9092 4292 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 10042 9160 10048 9172
rect 7616 9132 10048 9160
rect 7616 9120 7622 9132
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 11054 9120 11060 9172
rect 11112 9160 11118 9172
rect 13725 9163 13783 9169
rect 13725 9160 13737 9163
rect 11112 9132 13737 9160
rect 11112 9120 11118 9132
rect 13725 9129 13737 9132
rect 13771 9129 13783 9163
rect 13725 9123 13783 9129
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9160 14335 9163
rect 15838 9160 15844 9172
rect 14323 9132 15844 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 15838 9120 15844 9132
rect 15896 9120 15902 9172
rect 17862 9160 17868 9172
rect 15948 9132 17868 9160
rect 2363 9064 4292 9092
rect 6273 9095 6331 9101
rect 2363 9061 2375 9064
rect 2317 9055 2375 9061
rect 6273 9061 6285 9095
rect 6319 9092 6331 9095
rect 9766 9092 9772 9104
rect 6319 9064 9772 9092
rect 6319 9061 6331 9064
rect 6273 9055 6331 9061
rect 9766 9052 9772 9064
rect 9824 9052 9830 9104
rect 10502 9052 10508 9104
rect 10560 9052 10566 9104
rect 12713 9095 12771 9101
rect 11072 9064 12204 9092
rect 290 8984 296 9036
rect 348 9024 354 9036
rect 1210 9024 1216 9036
rect 348 8996 1216 9024
rect 348 8984 354 8996
rect 1210 8984 1216 8996
rect 1268 8984 1274 9036
rect 3786 8984 3792 9036
rect 3844 9024 3850 9036
rect 7190 9024 7196 9036
rect 3844 8996 7196 9024
rect 3844 8984 3850 8996
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 10520 9024 10548 9052
rect 9140 8996 10548 9024
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2406 8956 2412 8968
rect 1719 8928 2412 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 2774 8916 2780 8968
rect 2832 8916 2838 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4706 8956 4712 8968
rect 4295 8928 4712 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4706 8916 4712 8928
rect 4764 8916 4770 8968
rect 5626 8916 5632 8968
rect 5684 8916 5690 8968
rect 5902 8916 5908 8968
rect 5960 8956 5966 8968
rect 9140 8965 9168 8996
rect 6733 8959 6791 8965
rect 6733 8956 6745 8959
rect 5960 8928 6745 8956
rect 5960 8916 5966 8928
rect 6733 8925 6745 8928
rect 6779 8925 6791 8959
rect 6733 8919 6791 8925
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8925 7987 8959
rect 7929 8919 7987 8925
rect 9125 8959 9183 8965
rect 9125 8925 9137 8959
rect 9171 8925 9183 8959
rect 9125 8919 9183 8925
rect 4338 8848 4344 8900
rect 4396 8888 4402 8900
rect 7190 8888 7196 8900
rect 4396 8860 7196 8888
rect 4396 8848 4402 8860
rect 7190 8848 7196 8860
rect 7248 8848 7254 8900
rect 7944 8888 7972 8919
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9456 8928 9812 8956
rect 9456 8916 9462 8928
rect 9784 8897 9812 8928
rect 10134 8916 10140 8968
rect 10192 8956 10198 8968
rect 11072 8956 11100 9064
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 12176 9033 12204 9064
rect 12713 9061 12725 9095
rect 12759 9092 12771 9095
rect 14090 9092 14096 9104
rect 12759 9064 14096 9092
rect 12759 9061 12771 9064
rect 12713 9055 12771 9061
rect 12161 9027 12219 9033
rect 11388 8996 12112 9024
rect 11388 8984 11394 8996
rect 10192 8928 11100 8956
rect 10192 8916 10198 8928
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11977 8959 12035 8965
rect 11977 8956 11989 8959
rect 11204 8928 11989 8956
rect 11204 8916 11210 8928
rect 11977 8925 11989 8928
rect 12023 8925 12035 8959
rect 12084 8956 12112 8996
rect 12161 8993 12173 9027
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 12728 8956 12756 9055
rect 14090 9052 14096 9064
rect 14148 9052 14154 9104
rect 14550 9052 14556 9104
rect 14608 9092 14614 9104
rect 15948 9092 15976 9132
rect 17862 9120 17868 9132
rect 17920 9120 17926 9172
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 18782 9160 18788 9172
rect 18564 9132 18788 9160
rect 18564 9120 18570 9132
rect 18782 9120 18788 9132
rect 18840 9120 18846 9172
rect 20073 9163 20131 9169
rect 20073 9129 20085 9163
rect 20119 9160 20131 9163
rect 20254 9160 20260 9172
rect 20119 9132 20260 9160
rect 20119 9129 20131 9132
rect 20073 9123 20131 9129
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 21358 9120 21364 9172
rect 21416 9160 21422 9172
rect 23753 9163 23811 9169
rect 23753 9160 23765 9163
rect 21416 9132 23765 9160
rect 21416 9120 21422 9132
rect 23753 9129 23765 9132
rect 23799 9129 23811 9163
rect 23753 9123 23811 9129
rect 26326 9120 26332 9172
rect 26384 9120 26390 9172
rect 27433 9163 27491 9169
rect 27433 9129 27445 9163
rect 27479 9160 27491 9163
rect 28261 9163 28319 9169
rect 28261 9160 28273 9163
rect 27479 9132 28273 9160
rect 27479 9129 27491 9132
rect 27433 9123 27491 9129
rect 28261 9129 28273 9132
rect 28307 9160 28319 9163
rect 31294 9160 31300 9172
rect 28307 9132 31300 9160
rect 28307 9129 28319 9132
rect 28261 9123 28319 9129
rect 31294 9120 31300 9132
rect 31352 9120 31358 9172
rect 20898 9092 20904 9104
rect 14608 9064 15976 9092
rect 16224 9064 20904 9092
rect 14608 9052 14614 9064
rect 12894 8984 12900 9036
rect 12952 9024 12958 9036
rect 12952 8996 13492 9024
rect 12952 8984 12958 8996
rect 12084 8928 12756 8956
rect 13081 8959 13139 8965
rect 11977 8919 12035 8925
rect 13081 8925 13093 8959
rect 13127 8956 13139 8959
rect 13354 8956 13360 8968
rect 13127 8928 13360 8956
rect 13127 8925 13139 8928
rect 13081 8919 13139 8925
rect 13354 8916 13360 8928
rect 13412 8916 13418 8968
rect 13464 8956 13492 8996
rect 14918 8984 14924 9036
rect 14976 8984 14982 9036
rect 16224 9033 16252 9064
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 21818 9092 21824 9104
rect 21468 9064 21824 9092
rect 16209 9027 16267 9033
rect 16209 8993 16221 9027
rect 16255 8993 16267 9027
rect 16209 8987 16267 8993
rect 16482 8984 16488 9036
rect 16540 9024 16546 9036
rect 21468 9024 21496 9064
rect 21818 9052 21824 9064
rect 21876 9052 21882 9104
rect 22370 9052 22376 9104
rect 22428 9092 22434 9104
rect 22649 9095 22707 9101
rect 22649 9092 22661 9095
rect 22428 9064 22661 9092
rect 22428 9052 22434 9064
rect 22649 9061 22661 9064
rect 22695 9061 22707 9095
rect 22649 9055 22707 9061
rect 25038 9052 25044 9104
rect 25096 9092 25102 9104
rect 27706 9092 27712 9104
rect 25096 9064 27712 9092
rect 25096 9052 25102 9064
rect 27706 9052 27712 9064
rect 27764 9052 27770 9104
rect 32766 9052 32772 9104
rect 32824 9092 32830 9104
rect 40586 9092 40592 9104
rect 32824 9064 40592 9092
rect 32824 9052 32830 9064
rect 40586 9052 40592 9064
rect 40644 9052 40650 9104
rect 16540 8996 21496 9024
rect 21545 9027 21603 9033
rect 16540 8984 16546 8996
rect 21545 8993 21557 9027
rect 21591 9024 21603 9027
rect 21591 8996 22692 9024
rect 21591 8993 21603 8996
rect 21545 8987 21603 8993
rect 16022 8956 16028 8968
rect 13464 8928 16028 8956
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 17126 8916 17132 8968
rect 17184 8916 17190 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18782 8956 18788 8968
rect 18279 8928 18788 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 18877 8959 18935 8965
rect 18877 8925 18889 8959
rect 18923 8956 18935 8959
rect 19429 8959 19487 8965
rect 19429 8956 19441 8959
rect 18923 8928 19441 8956
rect 18923 8925 18935 8928
rect 18877 8919 18935 8925
rect 19429 8925 19441 8928
rect 19475 8925 19487 8959
rect 19429 8919 19487 8925
rect 20898 8916 20904 8968
rect 20956 8916 20962 8968
rect 22002 8916 22008 8968
rect 22060 8965 22066 8968
rect 22060 8959 22074 8965
rect 22062 8925 22074 8959
rect 22664 8956 22692 8996
rect 28994 8984 29000 9036
rect 29052 9024 29058 9036
rect 38470 9024 38476 9036
rect 29052 8996 38476 9024
rect 29052 8984 29058 8996
rect 38470 8984 38476 8996
rect 38528 8984 38534 9036
rect 23109 8959 23167 8965
rect 23109 8956 23121 8959
rect 22664 8928 23121 8956
rect 22060 8919 22074 8925
rect 23109 8925 23121 8928
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 24581 8959 24639 8965
rect 24581 8925 24593 8959
rect 24627 8925 24639 8959
rect 24581 8919 24639 8925
rect 22060 8916 22066 8919
rect 9769 8891 9827 8897
rect 7944 8860 9674 8888
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 4706 8820 4712 8832
rect 3467 8792 4712 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 4706 8780 4712 8792
rect 4764 8780 4770 8832
rect 4890 8780 4896 8832
rect 4948 8780 4954 8832
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 5350 8780 5356 8832
rect 5408 8820 5414 8832
rect 6454 8820 6460 8832
rect 5408 8792 6460 8820
rect 5408 8780 5414 8792
rect 6454 8780 6460 8792
rect 6512 8780 6518 8832
rect 7377 8823 7435 8829
rect 7377 8789 7389 8823
rect 7423 8820 7435 8823
rect 8386 8820 8392 8832
rect 7423 8792 8392 8820
rect 7423 8789 7435 8792
rect 7377 8783 7435 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8754 8820 8760 8832
rect 8619 8792 8760 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9646 8820 9674 8860
rect 9769 8857 9781 8891
rect 9815 8857 9827 8891
rect 9769 8851 9827 8857
rect 10226 8848 10232 8900
rect 10284 8848 10290 8900
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 10965 8891 11023 8897
rect 10965 8888 10977 8891
rect 10468 8860 10977 8888
rect 10468 8848 10474 8860
rect 10965 8857 10977 8860
rect 11011 8857 11023 8891
rect 10965 8851 11023 8857
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 14645 8891 14703 8897
rect 11112 8860 12204 8888
rect 11112 8848 11118 8860
rect 11330 8820 11336 8832
rect 9646 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 11882 8820 11888 8832
rect 11655 8792 11888 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 12176 8820 12204 8860
rect 14645 8857 14657 8891
rect 14691 8888 14703 8891
rect 15102 8888 15108 8900
rect 14691 8860 15108 8888
rect 14691 8857 14703 8860
rect 14645 8851 14703 8857
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 17773 8891 17831 8897
rect 15580 8860 17724 8888
rect 12894 8820 12900 8832
rect 12176 8792 12900 8820
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 13906 8820 13912 8832
rect 13412 8792 13912 8820
rect 13412 8780 13418 8792
rect 13906 8780 13912 8792
rect 13964 8780 13970 8832
rect 14737 8823 14795 8829
rect 14737 8789 14749 8823
rect 14783 8820 14795 8823
rect 14918 8820 14924 8832
rect 14783 8792 14924 8820
rect 14783 8789 14795 8792
rect 14737 8783 14795 8789
rect 14918 8780 14924 8792
rect 14976 8780 14982 8832
rect 15580 8829 15608 8860
rect 15565 8823 15623 8829
rect 15565 8789 15577 8823
rect 15611 8789 15623 8823
rect 15565 8783 15623 8789
rect 15930 8780 15936 8832
rect 15988 8780 15994 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16577 8823 16635 8829
rect 16577 8820 16589 8823
rect 16080 8792 16589 8820
rect 16080 8780 16086 8792
rect 16577 8789 16589 8792
rect 16623 8789 16635 8823
rect 16577 8783 16635 8789
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 17494 8820 17500 8832
rect 16899 8792 17500 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 17494 8780 17500 8792
rect 17552 8780 17558 8832
rect 17696 8820 17724 8860
rect 17773 8857 17785 8891
rect 17819 8888 17831 8891
rect 17862 8888 17868 8900
rect 17819 8860 17868 8888
rect 17819 8857 17831 8860
rect 17773 8851 17831 8857
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 19058 8848 19064 8900
rect 19116 8888 19122 8900
rect 24596 8888 24624 8919
rect 25682 8916 25688 8968
rect 25740 8916 25746 8968
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 19116 8860 20576 8888
rect 19116 8848 19122 8860
rect 20438 8820 20444 8832
rect 17696 8792 20444 8820
rect 20438 8780 20444 8792
rect 20496 8780 20502 8832
rect 20548 8820 20576 8860
rect 22572 8860 24624 8888
rect 22572 8820 22600 8860
rect 26234 8848 26240 8900
rect 26292 8888 26298 8900
rect 27172 8888 27200 8919
rect 27614 8916 27620 8968
rect 27672 8956 27678 8968
rect 41322 8956 41328 8968
rect 27672 8928 41328 8956
rect 27672 8916 27678 8928
rect 41322 8916 41328 8928
rect 41380 8916 41386 8968
rect 26292 8860 28120 8888
rect 26292 8848 26298 8860
rect 20548 8792 22600 8820
rect 25222 8780 25228 8832
rect 25280 8780 25286 8832
rect 27617 8823 27675 8829
rect 27617 8789 27629 8823
rect 27663 8820 27675 8823
rect 27706 8820 27712 8832
rect 27663 8792 27712 8820
rect 27663 8789 27675 8792
rect 27617 8783 27675 8789
rect 27706 8780 27712 8792
rect 27764 8780 27770 8832
rect 28092 8829 28120 8860
rect 28077 8823 28135 8829
rect 28077 8789 28089 8823
rect 28123 8820 28135 8823
rect 28350 8820 28356 8832
rect 28123 8792 28356 8820
rect 28123 8789 28135 8792
rect 28077 8783 28135 8789
rect 28350 8780 28356 8792
rect 28408 8780 28414 8832
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 1578 8576 1584 8628
rect 1636 8576 1642 8628
rect 1670 8576 1676 8628
rect 1728 8576 1734 8628
rect 3789 8619 3847 8625
rect 3789 8585 3801 8619
rect 3835 8616 3847 8619
rect 3970 8616 3976 8628
rect 3835 8588 3976 8616
rect 3835 8585 3847 8588
rect 3789 8579 3847 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4893 8619 4951 8625
rect 4893 8585 4905 8619
rect 4939 8616 4951 8619
rect 5534 8616 5540 8628
rect 4939 8588 5540 8616
rect 4939 8585 4951 8588
rect 4893 8579 4951 8585
rect 5534 8576 5540 8588
rect 5592 8576 5598 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 7006 8616 7012 8628
rect 6043 8588 7012 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 12158 8616 12164 8628
rect 8220 8588 12164 8616
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 7193 8551 7251 8557
rect 2648 8520 4292 8548
rect 2648 8508 2654 8520
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 4264 8489 4292 8520
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 7558 8548 7564 8560
rect 7239 8520 7564 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 7558 8508 7564 8520
rect 7616 8508 7622 8560
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1636 8452 2053 8480
rect 1636 8440 1642 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 4249 8483 4307 8489
rect 4249 8449 4261 8483
rect 4295 8449 4307 8483
rect 4249 8443 4307 8449
rect 1946 8372 1952 8424
rect 2004 8412 2010 8424
rect 2590 8412 2596 8424
rect 2004 8384 2596 8412
rect 2004 8372 2010 8384
rect 2590 8372 2596 8384
rect 2648 8372 2654 8424
rect 3160 8412 3188 8443
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5353 8483 5411 8489
rect 5353 8480 5365 8483
rect 4948 8452 5365 8480
rect 4948 8440 4954 8452
rect 5353 8449 5365 8452
rect 5399 8449 5411 8483
rect 5353 8443 5411 8449
rect 6546 8440 6552 8492
rect 6604 8440 6610 8492
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 8220 8480 8248 8588
rect 12158 8576 12164 8588
rect 12216 8576 12222 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 18414 8616 18420 8628
rect 13219 8588 18420 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 18782 8576 18788 8628
rect 18840 8616 18846 8628
rect 19521 8619 19579 8625
rect 19521 8616 19533 8619
rect 18840 8588 19533 8616
rect 18840 8576 18846 8588
rect 19521 8585 19533 8588
rect 19567 8585 19579 8619
rect 19521 8579 19579 8585
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 22462 8576 22468 8628
rect 22520 8616 22526 8628
rect 22649 8619 22707 8625
rect 22649 8616 22661 8619
rect 22520 8588 22661 8616
rect 22520 8576 22526 8588
rect 22649 8585 22661 8588
rect 22695 8585 22707 8619
rect 22649 8579 22707 8585
rect 23750 8576 23756 8628
rect 23808 8576 23814 8628
rect 24118 8576 24124 8628
rect 24176 8616 24182 8628
rect 24213 8619 24271 8625
rect 24213 8616 24225 8619
rect 24176 8588 24225 8616
rect 24176 8576 24182 8588
rect 24213 8585 24225 8588
rect 24259 8585 24271 8619
rect 24213 8579 24271 8585
rect 9769 8551 9827 8557
rect 9769 8517 9781 8551
rect 9815 8548 9827 8551
rect 10042 8548 10048 8560
rect 9815 8520 10048 8548
rect 9815 8517 9827 8520
rect 9769 8511 9827 8517
rect 10042 8508 10048 8520
rect 10100 8508 10106 8560
rect 12526 8548 12532 8560
rect 10980 8520 12532 8548
rect 7699 8452 8248 8480
rect 8297 8483 8355 8489
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8343 8452 8708 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 6362 8412 6368 8424
rect 3160 8384 6368 8412
rect 6362 8372 6368 8384
rect 6420 8372 6426 8424
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 8570 8412 8576 8424
rect 7524 8384 8576 8412
rect 7524 8372 7530 8384
rect 8570 8372 8576 8384
rect 8628 8372 8634 8424
rect 8680 8412 8708 8452
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 9214 8440 9220 8492
rect 9272 8480 9278 8492
rect 10226 8480 10232 8492
rect 9272 8452 10232 8480
rect 9272 8440 9278 8452
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10980 8424 11008 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 16761 8551 16819 8557
rect 16761 8548 16773 8551
rect 13464 8520 15516 8548
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11112 8452 11192 8480
rect 11112 8440 11118 8452
rect 9490 8412 9496 8424
rect 8680 8384 9496 8412
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 10042 8372 10048 8424
rect 10100 8372 10106 8424
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8381 10931 8415
rect 10873 8375 10931 8381
rect 2314 8304 2320 8356
rect 2372 8344 2378 8356
rect 4062 8344 4068 8356
rect 2372 8316 4068 8344
rect 2372 8304 2378 8316
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 7006 8344 7012 8356
rect 5644 8316 7012 8344
rect 1026 8236 1032 8288
rect 1084 8276 1090 8288
rect 1946 8276 1952 8288
rect 1084 8248 1952 8276
rect 1084 8236 1090 8248
rect 1946 8236 1952 8248
rect 2004 8236 2010 8288
rect 2685 8279 2743 8285
rect 2685 8245 2697 8279
rect 2731 8276 2743 8279
rect 5644 8276 5672 8316
rect 7006 8304 7012 8316
rect 7064 8304 7070 8356
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 10226 8344 10232 8356
rect 7800 8316 10232 8344
rect 7800 8304 7806 8316
rect 10226 8304 10232 8316
rect 10284 8304 10290 8356
rect 10413 8347 10471 8353
rect 10413 8313 10425 8347
rect 10459 8344 10471 8347
rect 10686 8344 10692 8356
rect 10459 8316 10692 8344
rect 10459 8313 10471 8316
rect 10413 8307 10471 8313
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 10888 8344 10916 8375
rect 10962 8372 10968 8424
rect 11020 8372 11026 8424
rect 11054 8344 11060 8356
rect 10888 8316 11060 8344
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 2731 8248 5672 8276
rect 2731 8245 2743 8248
rect 2685 8239 2743 8245
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6822 8276 6828 8288
rect 5776 8248 6828 8276
rect 5776 8236 5782 8248
rect 6822 8236 6828 8248
rect 6880 8236 6886 8288
rect 9398 8236 9404 8288
rect 9456 8236 9462 8288
rect 9674 8236 9680 8288
rect 9732 8276 9738 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9732 8248 9965 8276
rect 9732 8236 9738 8248
rect 9953 8245 9965 8248
rect 9999 8276 10011 8279
rect 11164 8276 11192 8452
rect 11514 8440 11520 8492
rect 11572 8440 11578 8492
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12345 8483 12403 8489
rect 12345 8480 12357 8483
rect 12124 8452 12357 8480
rect 12124 8440 12130 8452
rect 12345 8449 12357 8452
rect 12391 8449 12403 8483
rect 13464 8480 13492 8520
rect 12345 8443 12403 8449
rect 12636 8452 13492 8480
rect 13541 8483 13599 8489
rect 11532 8412 11560 8440
rect 12250 8412 12256 8424
rect 11532 8384 12256 8412
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12636 8421 12664 8452
rect 13541 8449 13553 8483
rect 13587 8480 13599 8483
rect 14550 8480 14556 8492
rect 13587 8452 14556 8480
rect 13587 8449 13599 8452
rect 13541 8443 13599 8449
rect 14550 8440 14556 8452
rect 14608 8440 14614 8492
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 15488 8480 15516 8520
rect 15672 8520 16773 8548
rect 15672 8489 15700 8520
rect 16761 8517 16773 8520
rect 16807 8548 16819 8551
rect 16807 8520 21220 8548
rect 16807 8517 16819 8520
rect 16761 8511 16819 8517
rect 15657 8483 15715 8489
rect 15488 8452 15608 8480
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8381 12495 8415
rect 12437 8375 12495 8381
rect 12621 8415 12679 8421
rect 12621 8381 12633 8415
rect 12667 8381 12679 8415
rect 12621 8375 12679 8381
rect 13633 8415 13691 8421
rect 13633 8381 13645 8415
rect 13679 8381 13691 8415
rect 13633 8375 13691 8381
rect 13725 8415 13783 8421
rect 13725 8381 13737 8415
rect 13771 8381 13783 8415
rect 13725 8375 13783 8381
rect 14369 8415 14427 8421
rect 14369 8381 14381 8415
rect 14415 8412 14427 8415
rect 15378 8412 15384 8424
rect 14415 8384 15384 8412
rect 14415 8381 14427 8384
rect 14369 8375 14427 8381
rect 11974 8304 11980 8356
rect 12032 8304 12038 8356
rect 9999 8248 11192 8276
rect 9999 8245 10011 8248
rect 9953 8239 10011 8245
rect 11330 8236 11336 8288
rect 11388 8276 11394 8288
rect 12158 8276 12164 8288
rect 11388 8248 12164 8276
rect 11388 8236 11394 8248
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 12452 8276 12480 8375
rect 13538 8304 13544 8356
rect 13596 8344 13602 8356
rect 13648 8344 13676 8375
rect 13596 8316 13676 8344
rect 13740 8344 13768 8375
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15580 8412 15608 8452
rect 15657 8449 15669 8483
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 18877 8483 18935 8489
rect 17972 8452 18828 8480
rect 17972 8412 18000 8452
rect 15580 8384 18000 8412
rect 18046 8372 18052 8424
rect 18104 8372 18110 8424
rect 18800 8412 18828 8452
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18966 8480 18972 8492
rect 18923 8452 18972 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19978 8440 19984 8492
rect 20036 8440 20042 8492
rect 19334 8412 19340 8424
rect 18800 8384 19340 8412
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 19518 8372 19524 8424
rect 19576 8412 19582 8424
rect 21085 8415 21143 8421
rect 21085 8412 21097 8415
rect 19576 8384 21097 8412
rect 19576 8372 19582 8384
rect 21085 8381 21097 8384
rect 21131 8381 21143 8415
rect 21192 8412 21220 8520
rect 21726 8508 21732 8560
rect 21784 8548 21790 8560
rect 24228 8548 24256 8579
rect 25958 8576 25964 8628
rect 26016 8616 26022 8628
rect 26053 8619 26111 8625
rect 26053 8616 26065 8619
rect 26016 8588 26065 8616
rect 26016 8576 26022 8588
rect 26053 8585 26065 8588
rect 26099 8585 26111 8619
rect 26053 8579 26111 8585
rect 28350 8576 28356 8628
rect 28408 8616 28414 8628
rect 36354 8616 36360 8628
rect 28408 8588 36360 8616
rect 28408 8576 28414 8588
rect 36354 8576 36360 8588
rect 36412 8576 36418 8628
rect 24673 8551 24731 8557
rect 24673 8548 24685 8551
rect 21784 8520 23520 8548
rect 24228 8520 24685 8548
rect 21784 8508 21790 8520
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8480 22063 8483
rect 22738 8480 22744 8492
rect 22051 8452 22744 8480
rect 22051 8449 22063 8452
rect 22005 8443 22063 8449
rect 22738 8440 22744 8452
rect 22796 8440 22802 8492
rect 23109 8483 23167 8489
rect 23109 8449 23121 8483
rect 23155 8480 23167 8483
rect 23382 8480 23388 8492
rect 23155 8452 23388 8480
rect 23155 8449 23167 8452
rect 23109 8443 23167 8449
rect 23382 8440 23388 8452
rect 23440 8440 23446 8492
rect 23492 8480 23520 8520
rect 24673 8517 24685 8520
rect 24719 8517 24731 8551
rect 24673 8511 24731 8517
rect 25593 8551 25651 8557
rect 25593 8517 25605 8551
rect 25639 8548 25651 8551
rect 26510 8548 26516 8560
rect 25639 8520 26516 8548
rect 25639 8517 25651 8520
rect 25593 8511 25651 8517
rect 26510 8508 26516 8520
rect 26568 8508 26574 8560
rect 24857 8483 24915 8489
rect 24857 8480 24869 8483
rect 23492 8452 24869 8480
rect 24857 8449 24869 8452
rect 24903 8449 24915 8483
rect 24857 8443 24915 8449
rect 25409 8483 25467 8489
rect 25409 8449 25421 8483
rect 25455 8480 25467 8483
rect 29730 8480 29736 8492
rect 25455 8452 29736 8480
rect 25455 8449 25467 8452
rect 25409 8443 25467 8449
rect 29730 8440 29736 8452
rect 29788 8440 29794 8492
rect 21192 8384 22094 8412
rect 21085 8375 21143 8381
rect 19352 8344 19380 8372
rect 20990 8344 20996 8356
rect 13740 8316 16804 8344
rect 13596 8304 13602 8316
rect 12710 8276 12716 8288
rect 12452 8248 12716 8276
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 12802 8236 12808 8288
rect 12860 8276 12866 8288
rect 14274 8276 14280 8288
rect 12860 8248 14280 8276
rect 12860 8236 12866 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 16301 8279 16359 8285
rect 16301 8245 16313 8279
rect 16347 8276 16359 8279
rect 16390 8276 16396 8288
rect 16347 8248 16396 8276
rect 16347 8245 16359 8248
rect 16301 8239 16359 8245
rect 16390 8236 16396 8248
rect 16448 8236 16454 8288
rect 16776 8276 16804 8316
rect 17972 8316 18184 8344
rect 19352 8316 20996 8344
rect 17972 8276 18000 8316
rect 16776 8248 18000 8276
rect 18156 8276 18184 8316
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 22066 8344 22094 8384
rect 27798 8372 27804 8424
rect 27856 8412 27862 8424
rect 31018 8412 31024 8424
rect 27856 8384 31024 8412
rect 27856 8372 27862 8384
rect 31018 8372 31024 8384
rect 31076 8372 31082 8424
rect 32306 8344 32312 8356
rect 22066 8316 32312 8344
rect 32306 8304 32312 8316
rect 32364 8304 32370 8356
rect 23934 8276 23940 8288
rect 18156 8248 23940 8276
rect 23934 8236 23940 8248
rect 23992 8236 23998 8288
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 2314 8032 2320 8084
rect 2372 8032 2378 8084
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 3421 8075 3479 8081
rect 3421 8072 3433 8075
rect 2464 8044 3433 8072
rect 2464 8032 2470 8044
rect 3421 8041 3433 8044
rect 3467 8041 3479 8075
rect 3421 8035 3479 8041
rect 4709 8075 4767 8081
rect 4709 8041 4721 8075
rect 4755 8072 4767 8075
rect 4798 8072 4804 8084
rect 4755 8044 4804 8072
rect 4755 8041 4767 8044
rect 4709 8035 4767 8041
rect 4798 8032 4804 8044
rect 4856 8032 4862 8084
rect 5074 8032 5080 8084
rect 5132 8072 5138 8084
rect 5810 8072 5816 8084
rect 5132 8044 5816 8072
rect 5132 8032 5138 8044
rect 5810 8032 5816 8044
rect 5868 8032 5874 8084
rect 6086 8032 6092 8084
rect 6144 8072 6150 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 6144 8044 6193 8072
rect 6144 8032 6150 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7469 8075 7527 8081
rect 7469 8072 7481 8075
rect 7248 8044 7481 8072
rect 7248 8032 7254 8044
rect 7469 8041 7481 8044
rect 7515 8041 7527 8075
rect 7469 8035 7527 8041
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 8352 8044 8585 8072
rect 8352 8032 8358 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 8754 8032 8760 8084
rect 8812 8072 8818 8084
rect 9674 8072 9680 8084
rect 8812 8044 9680 8072
rect 8812 8032 8818 8044
rect 9674 8032 9680 8044
rect 9732 8032 9738 8084
rect 9858 8032 9864 8084
rect 9916 8032 9922 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 11514 8072 11520 8084
rect 10100 8044 11520 8072
rect 10100 8032 10106 8044
rect 11514 8032 11520 8044
rect 11572 8032 11578 8084
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 13170 8072 13176 8084
rect 11756 8044 13176 8072
rect 11756 8032 11762 8044
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 13722 8032 13728 8084
rect 13780 8032 13786 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 17037 8075 17095 8081
rect 17037 8072 17049 8075
rect 16816 8044 17049 8072
rect 16816 8032 16822 8044
rect 17037 8041 17049 8044
rect 17083 8041 17095 8075
rect 17037 8035 17095 8041
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 17184 8044 18153 8072
rect 17184 8032 17190 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 20898 8032 20904 8084
rect 20956 8072 20962 8084
rect 22649 8075 22707 8081
rect 22649 8072 22661 8075
rect 20956 8044 22661 8072
rect 20956 8032 20962 8044
rect 22649 8041 22661 8044
rect 22695 8041 22707 8075
rect 22649 8035 22707 8041
rect 23382 8032 23388 8084
rect 23440 8072 23446 8084
rect 23753 8075 23811 8081
rect 23753 8072 23765 8075
rect 23440 8044 23765 8072
rect 23440 8032 23446 8044
rect 23753 8041 23765 8044
rect 23799 8041 23811 8075
rect 23753 8035 23811 8041
rect 24394 8032 24400 8084
rect 24452 8072 24458 8084
rect 24452 8044 25452 8072
rect 24452 8032 24458 8044
rect 1302 7964 1308 8016
rect 1360 8004 1366 8016
rect 4338 8004 4344 8016
rect 1360 7976 4344 8004
rect 1360 7964 1366 7976
rect 4338 7964 4344 7976
rect 4396 7964 4402 8016
rect 10962 8004 10968 8016
rect 6564 7976 10968 8004
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 4080 7908 5825 7936
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 2222 7868 2228 7880
rect 1719 7840 2228 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7837 2835 7871
rect 2777 7831 2835 7837
rect 2792 7800 2820 7831
rect 3510 7828 3516 7880
rect 3568 7868 3574 7880
rect 3970 7868 3976 7880
rect 3568 7840 3976 7868
rect 3568 7828 3574 7840
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4080 7877 4108 7908
rect 5813 7905 5825 7908
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6564 7877 6592 7976
rect 10962 7964 10968 7976
rect 11020 7964 11026 8016
rect 11146 7964 11152 8016
rect 11204 8004 11210 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 11204 7976 14105 8004
rect 11204 7964 11210 7976
rect 14093 7973 14105 7976
rect 14139 7973 14151 8007
rect 14093 7967 14151 7973
rect 15194 7964 15200 8016
rect 15252 8004 15258 8016
rect 21545 8007 21603 8013
rect 15252 7976 18644 8004
rect 15252 7964 15258 7976
rect 9217 7939 9275 7945
rect 6656 7908 8064 7936
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 5169 7871 5227 7877
rect 5169 7837 5181 7871
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 4890 7800 4896 7812
rect 2792 7772 4896 7800
rect 4890 7760 4896 7772
rect 4948 7760 4954 7812
rect 5184 7800 5212 7831
rect 5258 7800 5264 7812
rect 5184 7772 5264 7800
rect 5258 7760 5264 7772
rect 5316 7800 5322 7812
rect 6656 7800 6684 7908
rect 6822 7828 6828 7880
rect 6880 7868 6886 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 6880 7840 7941 7868
rect 6880 7828 6886 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 8036 7868 8064 7908
rect 9217 7905 9229 7939
rect 9263 7936 9275 7939
rect 9582 7936 9588 7948
rect 9263 7908 9588 7936
rect 9263 7905 9275 7908
rect 9217 7899 9275 7905
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 10413 7939 10471 7945
rect 10413 7905 10425 7939
rect 10459 7936 10471 7939
rect 10870 7936 10876 7948
rect 10459 7908 10876 7936
rect 10459 7905 10471 7908
rect 10413 7899 10471 7905
rect 10042 7868 10048 7880
rect 8036 7840 10048 7868
rect 7929 7831 7987 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10318 7868 10324 7880
rect 10275 7840 10324 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 10428 7800 10456 7899
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11054 7896 11060 7948
rect 11112 7936 11118 7948
rect 13906 7936 13912 7948
rect 11112 7908 13912 7936
rect 11112 7896 11118 7908
rect 13906 7896 13912 7908
rect 13964 7896 13970 7948
rect 14645 7939 14703 7945
rect 14645 7905 14657 7939
rect 14691 7936 14703 7939
rect 15930 7936 15936 7948
rect 14691 7908 15936 7936
rect 14691 7905 14703 7908
rect 14645 7899 14703 7905
rect 15930 7896 15936 7908
rect 15988 7896 15994 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 17862 7936 17868 7948
rect 16172 7908 17868 7936
rect 16172 7896 16178 7908
rect 17862 7896 17868 7908
rect 17920 7896 17926 7948
rect 18616 7945 18644 7976
rect 19444 7976 19932 8004
rect 19444 7945 19472 7976
rect 18601 7939 18659 7945
rect 18601 7905 18613 7939
rect 18647 7905 18659 7939
rect 18601 7899 18659 7905
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7905 19487 7939
rect 19904 7936 19932 7976
rect 21545 7973 21557 8007
rect 21591 8004 21603 8007
rect 25314 8004 25320 8016
rect 21591 7976 25320 8004
rect 21591 7973 21603 7976
rect 21545 7967 21603 7973
rect 25314 7964 25320 7976
rect 25372 7964 25378 8016
rect 25424 8004 25452 8044
rect 25498 8032 25504 8084
rect 25556 8072 25562 8084
rect 39390 8072 39396 8084
rect 25556 8044 39396 8072
rect 25556 8032 25562 8044
rect 39390 8032 39396 8044
rect 39448 8032 39454 8084
rect 49050 8004 49056 8016
rect 25424 7976 49056 8004
rect 49050 7964 49056 7976
rect 49108 7964 49114 8016
rect 22186 7936 22192 7948
rect 19429 7899 19487 7905
rect 19628 7908 19840 7936
rect 19904 7908 22192 7936
rect 11238 7828 11244 7880
rect 11296 7868 11302 7880
rect 11517 7871 11575 7877
rect 11517 7868 11529 7871
rect 11296 7840 11529 7868
rect 11296 7828 11302 7840
rect 11517 7837 11529 7840
rect 11563 7837 11575 7871
rect 11517 7831 11575 7837
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7868 12035 7871
rect 12158 7868 12164 7880
rect 12023 7840 12164 7868
rect 12023 7837 12035 7840
rect 11977 7831 12035 7837
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12621 7871 12679 7877
rect 12621 7837 12633 7871
rect 12667 7868 12679 7871
rect 13081 7871 13139 7877
rect 13081 7868 13093 7871
rect 12667 7840 13093 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 13081 7837 13093 7840
rect 13127 7837 13139 7871
rect 13081 7831 13139 7837
rect 13170 7828 13176 7880
rect 13228 7868 13234 7880
rect 14918 7868 14924 7880
rect 13228 7840 14924 7868
rect 13228 7828 13234 7840
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7868 15347 7871
rect 15746 7868 15752 7880
rect 15335 7840 15752 7868
rect 15335 7837 15347 7840
rect 15289 7831 15347 7837
rect 15746 7828 15752 7840
rect 15804 7828 15810 7880
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 17497 7871 17555 7877
rect 17497 7837 17509 7871
rect 17543 7868 17555 7871
rect 18874 7868 18880 7880
rect 17543 7840 18880 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 18874 7828 18880 7840
rect 18932 7828 18938 7880
rect 18966 7828 18972 7880
rect 19024 7868 19030 7880
rect 19628 7868 19656 7908
rect 19024 7840 19656 7868
rect 19024 7828 19030 7840
rect 19702 7828 19708 7880
rect 19760 7828 19766 7880
rect 19812 7868 19840 7908
rect 22186 7896 22192 7908
rect 22244 7896 22250 7948
rect 24854 7896 24860 7948
rect 24912 7896 24918 7948
rect 25225 7939 25283 7945
rect 25225 7905 25237 7939
rect 25271 7936 25283 7939
rect 25590 7936 25596 7948
rect 25271 7908 25596 7936
rect 25271 7905 25283 7908
rect 25225 7899 25283 7905
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 20901 7871 20959 7877
rect 20901 7868 20913 7871
rect 19812 7840 20913 7868
rect 20901 7837 20913 7840
rect 20947 7837 20959 7871
rect 20901 7831 20959 7837
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 22005 7871 22063 7877
rect 22005 7868 22017 7871
rect 21324 7840 22017 7868
rect 21324 7828 21330 7840
rect 22005 7837 22017 7840
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 23106 7828 23112 7880
rect 23164 7828 23170 7880
rect 24762 7828 24768 7880
rect 24820 7868 24826 7880
rect 24820 7840 35894 7868
rect 24820 7828 24826 7840
rect 5316 7772 6684 7800
rect 7116 7772 10456 7800
rect 11333 7803 11391 7809
rect 5316 7760 5322 7772
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 7116 7732 7144 7772
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 12066 7800 12072 7812
rect 11379 7772 12072 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 16482 7800 16488 7812
rect 15252 7772 16488 7800
rect 15252 7760 15258 7772
rect 16482 7760 16488 7772
rect 16540 7800 16546 7812
rect 24673 7803 24731 7809
rect 16540 7772 24624 7800
rect 16540 7760 16546 7772
rect 2832 7704 7144 7732
rect 7193 7735 7251 7741
rect 2832 7692 2838 7704
rect 7193 7701 7205 7735
rect 7239 7732 7251 7735
rect 7558 7732 7564 7744
rect 7239 7704 7564 7732
rect 7239 7701 7251 7704
rect 7193 7695 7251 7701
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 10226 7692 10232 7744
rect 10284 7732 10290 7744
rect 10321 7735 10379 7741
rect 10321 7732 10333 7735
rect 10284 7704 10333 7732
rect 10284 7692 10290 7704
rect 10321 7701 10333 7704
rect 10367 7701 10379 7735
rect 10321 7695 10379 7701
rect 10594 7692 10600 7744
rect 10652 7732 10658 7744
rect 10873 7735 10931 7741
rect 10873 7732 10885 7735
rect 10652 7704 10885 7732
rect 10652 7692 10658 7704
rect 10873 7701 10885 7704
rect 10919 7701 10931 7735
rect 10873 7695 10931 7701
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 12342 7732 12348 7744
rect 11020 7704 12348 7732
rect 11020 7692 11026 7704
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 14274 7692 14280 7744
rect 14332 7692 14338 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15712 7704 15945 7732
rect 15712 7692 15718 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 24118 7732 24124 7744
rect 18564 7704 24124 7732
rect 18564 7692 18570 7704
rect 24118 7692 24124 7704
rect 24176 7692 24182 7744
rect 24596 7732 24624 7772
rect 24673 7769 24685 7803
rect 24719 7800 24731 7803
rect 24854 7800 24860 7812
rect 24719 7772 24860 7800
rect 24719 7769 24731 7772
rect 24673 7763 24731 7769
rect 24854 7760 24860 7772
rect 24912 7800 24918 7812
rect 25590 7800 25596 7812
rect 24912 7772 25596 7800
rect 24912 7760 24918 7772
rect 25590 7760 25596 7772
rect 25648 7760 25654 7812
rect 27798 7732 27804 7744
rect 24596 7704 27804 7732
rect 27798 7692 27804 7704
rect 27856 7692 27862 7744
rect 35866 7732 35894 7840
rect 38746 7732 38752 7744
rect 35866 7704 38752 7732
rect 38746 7692 38752 7704
rect 38804 7692 38810 7744
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 1486 7488 1492 7540
rect 1544 7488 1550 7540
rect 2498 7488 2504 7540
rect 2556 7488 2562 7540
rect 3605 7531 3663 7537
rect 3605 7497 3617 7531
rect 3651 7528 3663 7531
rect 4154 7528 4160 7540
rect 3651 7500 4160 7528
rect 3651 7497 3663 7500
rect 3605 7491 3663 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4709 7531 4767 7537
rect 4709 7528 4721 7531
rect 4488 7500 4721 7528
rect 4488 7488 4494 7500
rect 4709 7497 4721 7500
rect 4755 7497 4767 7531
rect 4709 7491 4767 7497
rect 4982 7488 4988 7540
rect 5040 7488 5046 7540
rect 6546 7488 6552 7540
rect 6604 7528 6610 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 6604 7500 9597 7528
rect 6604 7488 6610 7500
rect 9585 7497 9597 7500
rect 9631 7497 9643 7531
rect 9585 7491 9643 7497
rect 10045 7531 10103 7537
rect 10045 7497 10057 7531
rect 10091 7528 10103 7531
rect 10962 7528 10968 7540
rect 10091 7500 10968 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11054 7488 11060 7540
rect 11112 7528 11118 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11112 7500 11529 7528
rect 11112 7488 11118 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12434 7528 12440 7540
rect 12308 7500 12440 7528
rect 12308 7488 12314 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 15197 7531 15255 7537
rect 12544 7500 14136 7528
rect 1210 7420 1216 7472
rect 1268 7460 1274 7472
rect 1578 7460 1584 7472
rect 1268 7432 1584 7460
rect 1268 7420 1274 7432
rect 1578 7420 1584 7432
rect 1636 7420 1642 7472
rect 2130 7420 2136 7472
rect 2188 7460 2194 7472
rect 7377 7463 7435 7469
rect 7377 7460 7389 7463
rect 2188 7432 7389 7460
rect 2188 7420 2194 7432
rect 7377 7429 7389 7432
rect 7423 7429 7435 7463
rect 7377 7423 7435 7429
rect 8386 7420 8392 7472
rect 8444 7460 8450 7472
rect 8444 7432 11100 7460
rect 8444 7420 8450 7432
rect 1854 7352 1860 7404
rect 1912 7352 1918 7404
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 2976 7324 3004 7355
rect 4062 7352 4068 7404
rect 4120 7352 4126 7404
rect 4706 7352 4712 7404
rect 4764 7392 4770 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 4764 7364 5365 7392
rect 4764 7352 4770 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6779 7364 7788 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 5258 7324 5264 7336
rect 2976 7296 5264 7324
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5997 7327 6055 7333
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 7098 7324 7104 7336
rect 6043 7296 7104 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 7098 7284 7104 7296
rect 7156 7284 7162 7336
rect 7760 7324 7788 7364
rect 7834 7352 7840 7404
rect 7892 7352 7898 7404
rect 7926 7352 7932 7404
rect 7984 7392 7990 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 7984 7364 8953 7392
rect 7984 7352 7990 7364
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 7760 7296 8616 7324
rect 3510 7216 3516 7268
rect 3568 7256 3574 7268
rect 4706 7256 4712 7268
rect 3568 7228 4712 7256
rect 3568 7216 3574 7228
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 7926 7256 7932 7268
rect 5500 7228 7932 7256
rect 5500 7216 5506 7228
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 4614 7148 4620 7200
rect 4672 7188 4678 7200
rect 5534 7188 5540 7200
rect 4672 7160 5540 7188
rect 4672 7148 4678 7160
rect 5534 7148 5540 7160
rect 5592 7148 5598 7200
rect 6457 7191 6515 7197
rect 6457 7157 6469 7191
rect 6503 7188 6515 7191
rect 6730 7188 6736 7200
rect 6503 7160 6736 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8481 7191 8539 7197
rect 8481 7188 8493 7191
rect 8352 7160 8493 7188
rect 8352 7148 8358 7160
rect 8481 7157 8493 7160
rect 8527 7157 8539 7191
rect 8588 7188 8616 7296
rect 10318 7284 10324 7336
rect 10376 7324 10382 7336
rect 10505 7327 10563 7333
rect 10505 7324 10517 7327
rect 10376 7296 10517 7324
rect 10376 7284 10382 7296
rect 10505 7293 10517 7296
rect 10551 7293 10563 7327
rect 10505 7287 10563 7293
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 11072 7324 11100 7432
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 12544 7460 12572 7500
rect 11204 7432 12572 7460
rect 11204 7420 11210 7432
rect 12618 7420 12624 7472
rect 12676 7460 12682 7472
rect 14001 7463 14059 7469
rect 14001 7460 14013 7463
rect 12676 7432 14013 7460
rect 12676 7420 12682 7432
rect 14001 7429 14013 7432
rect 14047 7429 14059 7463
rect 14001 7423 14059 7429
rect 11238 7352 11244 7404
rect 11296 7392 11302 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 11296 7364 12265 7392
rect 11296 7352 11302 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 12253 7355 12311 7361
rect 12728 7364 13369 7392
rect 12728 7324 12756 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 11072 7296 12756 7324
rect 12894 7284 12900 7336
rect 12952 7284 12958 7336
rect 14108 7324 14136 7500
rect 15197 7497 15209 7531
rect 15243 7528 15255 7531
rect 15286 7528 15292 7540
rect 15243 7500 15292 7528
rect 15243 7497 15255 7500
rect 15197 7491 15255 7497
rect 15286 7488 15292 7500
rect 15344 7488 15350 7540
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 16853 7531 16911 7537
rect 16853 7528 16865 7531
rect 16816 7500 16865 7528
rect 16816 7488 16822 7500
rect 16853 7497 16865 7500
rect 16899 7497 16911 7531
rect 16853 7491 16911 7497
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 19978 7488 19984 7540
rect 20036 7528 20042 7540
rect 20073 7531 20131 7537
rect 20073 7528 20085 7531
rect 20036 7500 20085 7528
rect 20036 7488 20042 7500
rect 20073 7497 20085 7500
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 21450 7488 21456 7540
rect 21508 7488 21514 7540
rect 21542 7488 21548 7540
rect 21600 7528 21606 7540
rect 23106 7528 23112 7540
rect 21600 7500 23112 7528
rect 21600 7488 21606 7500
rect 23106 7488 23112 7500
rect 23164 7488 23170 7540
rect 23750 7488 23756 7540
rect 23808 7528 23814 7540
rect 25682 7528 25688 7540
rect 23808 7500 25688 7528
rect 23808 7488 23814 7500
rect 25682 7488 25688 7500
rect 25740 7488 25746 7540
rect 15102 7420 15108 7472
rect 15160 7460 15166 7472
rect 18785 7463 18843 7469
rect 18785 7460 18797 7463
rect 15160 7432 18797 7460
rect 15160 7420 15166 7432
rect 18785 7429 18797 7432
rect 18831 7429 18843 7463
rect 18785 7423 18843 7429
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 21177 7463 21235 7469
rect 21177 7460 21189 7463
rect 19300 7432 21189 7460
rect 19300 7420 19306 7432
rect 21177 7429 21189 7432
rect 21223 7429 21235 7463
rect 21177 7423 21235 7429
rect 22278 7420 22284 7472
rect 22336 7420 22342 7472
rect 22830 7420 22836 7472
rect 22888 7420 22894 7472
rect 24857 7463 24915 7469
rect 24857 7460 24869 7463
rect 24228 7432 24869 7460
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7392 14611 7395
rect 15194 7392 15200 7404
rect 14599 7364 15200 7392
rect 14599 7361 14611 7364
rect 14553 7355 14611 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 16666 7392 16672 7404
rect 15764 7364 16672 7392
rect 15378 7324 15384 7336
rect 14108 7296 15384 7324
rect 15378 7284 15384 7296
rect 15436 7284 15442 7336
rect 9398 7216 9404 7268
rect 9456 7256 9462 7268
rect 10962 7256 10968 7268
rect 9456 7228 10968 7256
rect 9456 7216 9462 7228
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 11330 7216 11336 7268
rect 11388 7216 11394 7268
rect 11514 7216 11520 7268
rect 11572 7256 11578 7268
rect 11885 7259 11943 7265
rect 11885 7256 11897 7259
rect 11572 7228 11897 7256
rect 11572 7216 11578 7228
rect 11885 7225 11897 7228
rect 11931 7225 11943 7259
rect 15764 7256 15792 7364
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 17037 7395 17095 7401
rect 17037 7361 17049 7395
rect 17083 7392 17095 7395
rect 17126 7392 17132 7404
rect 17083 7364 17132 7392
rect 17083 7361 17095 7364
rect 17037 7355 17095 7361
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18506 7392 18512 7404
rect 17727 7364 18512 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 19429 7395 19487 7401
rect 19429 7361 19441 7395
rect 19475 7392 19487 7395
rect 19794 7392 19800 7404
rect 19475 7364 19800 7392
rect 19475 7361 19487 7364
rect 19429 7355 19487 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 20530 7352 20536 7404
rect 20588 7352 20594 7404
rect 21910 7352 21916 7404
rect 21968 7392 21974 7404
rect 24228 7401 24256 7432
rect 24857 7429 24869 7432
rect 24903 7460 24915 7463
rect 28994 7460 29000 7472
rect 24903 7432 29000 7460
rect 24903 7429 24915 7432
rect 24857 7423 24915 7429
rect 28994 7420 29000 7432
rect 29052 7420 29058 7472
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21968 7364 22017 7392
rect 21968 7352 21974 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 24213 7395 24271 7401
rect 24213 7361 24225 7395
rect 24259 7361 24271 7395
rect 24213 7355 24271 7361
rect 16114 7284 16120 7336
rect 16172 7324 16178 7336
rect 24854 7324 24860 7336
rect 16172 7296 24860 7324
rect 16172 7284 16178 7296
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 11885 7219 11943 7225
rect 15488 7228 15792 7256
rect 8938 7188 8944 7200
rect 8588 7160 8944 7188
rect 8481 7151 8539 7157
rect 8938 7148 8944 7160
rect 8996 7188 9002 7200
rect 11701 7191 11759 7197
rect 11701 7188 11713 7191
rect 8996 7160 11713 7188
rect 8996 7148 9002 7160
rect 11701 7157 11713 7160
rect 11747 7157 11759 7191
rect 11701 7151 11759 7157
rect 12066 7148 12072 7200
rect 12124 7188 12130 7200
rect 15488 7188 15516 7228
rect 16666 7216 16672 7268
rect 16724 7256 16730 7268
rect 17218 7256 17224 7268
rect 16724 7228 17224 7256
rect 16724 7216 16730 7228
rect 17218 7216 17224 7228
rect 17276 7256 17282 7268
rect 18966 7256 18972 7268
rect 17276 7228 18972 7256
rect 17276 7216 17282 7228
rect 18966 7216 18972 7228
rect 19024 7216 19030 7268
rect 24394 7216 24400 7268
rect 24452 7216 24458 7268
rect 12124 7160 15516 7188
rect 12124 7148 12130 7160
rect 15654 7148 15660 7200
rect 15712 7188 15718 7200
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 15712 7160 16313 7188
rect 15712 7148 15718 7160
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 17126 7148 17132 7200
rect 17184 7188 17190 7200
rect 17313 7191 17371 7197
rect 17313 7188 17325 7191
rect 17184 7160 17325 7188
rect 17184 7148 17190 7160
rect 17313 7157 17325 7160
rect 17359 7188 17371 7191
rect 25774 7188 25780 7200
rect 17359 7160 25780 7188
rect 17359 7157 17371 7160
rect 17313 7151 17371 7157
rect 25774 7148 25780 7160
rect 25832 7148 25838 7200
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 5350 6984 5356 6996
rect 2648 6956 5356 6984
rect 2648 6944 2654 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 6362 6944 6368 6996
rect 6420 6944 6426 6996
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 9214 6984 9220 6996
rect 7340 6956 9220 6984
rect 7340 6944 7346 6956
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9861 6987 9919 6993
rect 9861 6953 9873 6987
rect 9907 6984 9919 6987
rect 13722 6984 13728 6996
rect 9907 6956 13728 6984
rect 9907 6953 9919 6956
rect 9861 6947 9919 6953
rect 13722 6944 13728 6956
rect 13780 6944 13786 6996
rect 15838 6984 15844 6996
rect 14016 6956 15844 6984
rect 1118 6876 1124 6928
rect 1176 6916 1182 6928
rect 2682 6916 2688 6928
rect 1176 6888 2688 6916
rect 1176 6876 1182 6888
rect 2682 6876 2688 6888
rect 2740 6876 2746 6928
rect 3694 6876 3700 6928
rect 3752 6916 3758 6928
rect 3752 6888 6914 6916
rect 3752 6876 3758 6888
rect 1762 6808 1768 6860
rect 1820 6808 1826 6860
rect 6886 6848 6914 6888
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 10594 6916 10600 6928
rect 7248 6888 10600 6916
rect 7248 6876 7254 6888
rect 10594 6876 10600 6888
rect 10652 6876 10658 6928
rect 10686 6876 10692 6928
rect 10744 6916 10750 6928
rect 14016 6916 14044 6956
rect 15838 6944 15844 6956
rect 15896 6944 15902 6996
rect 15930 6944 15936 6996
rect 15988 6984 15994 6996
rect 20165 6987 20223 6993
rect 15988 6956 19334 6984
rect 15988 6944 15994 6956
rect 10744 6888 14044 6916
rect 10744 6876 10750 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 16298 6916 16304 6928
rect 14792 6888 16304 6916
rect 14792 6876 14798 6888
rect 16298 6876 16304 6888
rect 16356 6876 16362 6928
rect 7374 6848 7380 6860
rect 6886 6820 7380 6848
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 7800 6820 8524 6848
rect 7800 6808 7806 6820
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1780 6780 1808 6808
rect 2130 6780 2136 6792
rect 1719 6752 2136 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2590 6780 2596 6792
rect 2547 6752 2596 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6780 3479 6783
rect 3510 6780 3516 6792
rect 3467 6752 3516 6780
rect 3467 6749 3479 6752
rect 3421 6743 3479 6749
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 4157 6783 4215 6789
rect 3927 6776 4108 6780
rect 4157 6776 4169 6783
rect 3927 6752 4169 6776
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 4080 6749 4169 6752
rect 4203 6780 4215 6783
rect 4246 6780 4252 6792
rect 4203 6752 4252 6780
rect 4203 6749 4215 6752
rect 4080 6748 4215 6749
rect 4157 6743 4215 6748
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 4617 6783 4675 6789
rect 4617 6780 4629 6783
rect 4396 6752 4629 6780
rect 4396 6740 4402 6752
rect 4617 6749 4629 6752
rect 4663 6749 4675 6783
rect 4617 6743 4675 6749
rect 5258 6740 5264 6792
rect 5316 6740 5322 6792
rect 5718 6740 5724 6792
rect 5776 6740 5782 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6825 6783 6883 6789
rect 6825 6780 6837 6783
rect 6052 6752 6837 6780
rect 6052 6740 6058 6752
rect 6825 6749 6837 6752
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7469 6783 7527 6789
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7929 6783 7987 6789
rect 7929 6780 7941 6783
rect 7515 6752 7941 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 7929 6749 7941 6752
rect 7975 6749 7987 6783
rect 8496 6780 8524 6820
rect 8570 6808 8576 6860
rect 8628 6808 8634 6860
rect 10226 6848 10232 6860
rect 8680 6820 10232 6848
rect 8680 6780 8708 6820
rect 10226 6808 10232 6820
rect 10284 6808 10290 6860
rect 10778 6808 10784 6860
rect 10836 6808 10842 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11020 6820 12020 6848
rect 11020 6808 11026 6820
rect 8496 6752 8708 6780
rect 7929 6743 7987 6749
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 9088 6752 9137 6780
rect 9088 6740 9094 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 11517 6783 11575 6789
rect 11517 6749 11529 6783
rect 11563 6780 11575 6783
rect 11698 6780 11704 6792
rect 11563 6752 11704 6780
rect 11563 6749 11575 6752
rect 11517 6743 11575 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 11992 6789 12020 6820
rect 12526 6808 12532 6860
rect 12584 6848 12590 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12584 6820 12633 6848
rect 12584 6808 12590 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12728 6820 13216 6848
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6749 12035 6783
rect 11977 6743 12035 6749
rect 12066 6740 12072 6792
rect 12124 6780 12130 6792
rect 12728 6780 12756 6820
rect 12124 6752 12756 6780
rect 13081 6783 13139 6789
rect 12124 6740 12130 6752
rect 13081 6749 13093 6783
rect 13127 6749 13139 6783
rect 13188 6780 13216 6820
rect 13446 6808 13452 6860
rect 13504 6848 13510 6860
rect 13725 6851 13783 6857
rect 13725 6848 13737 6851
rect 13504 6820 13737 6848
rect 13504 6808 13510 6820
rect 13725 6817 13737 6820
rect 13771 6817 13783 6851
rect 13725 6811 13783 6817
rect 14550 6808 14556 6860
rect 14608 6808 14614 6860
rect 15930 6848 15936 6860
rect 14660 6820 15936 6848
rect 14660 6780 14688 6820
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6848 16451 6851
rect 16482 6848 16488 6860
rect 16439 6820 16488 6848
rect 16439 6817 16451 6820
rect 16393 6811 16451 6817
rect 16482 6808 16488 6820
rect 16540 6808 16546 6860
rect 16574 6808 16580 6860
rect 16632 6848 16638 6860
rect 17405 6851 17463 6857
rect 17405 6848 17417 6851
rect 16632 6820 17417 6848
rect 16632 6808 16638 6820
rect 17405 6817 17417 6820
rect 17451 6817 17463 6851
rect 17405 6811 17463 6817
rect 17494 6808 17500 6860
rect 17552 6848 17558 6860
rect 17552 6820 18000 6848
rect 17552 6808 17558 6820
rect 13188 6752 14688 6780
rect 13081 6743 13139 6749
rect 3234 6672 3240 6724
rect 3292 6672 3298 6724
rect 7834 6672 7840 6724
rect 7892 6712 7898 6724
rect 9674 6712 9680 6724
rect 7892 6684 9680 6712
rect 7892 6672 7898 6684
rect 9674 6672 9680 6684
rect 9732 6672 9738 6724
rect 1762 6604 1768 6656
rect 1820 6604 1826 6656
rect 1946 6604 1952 6656
rect 2004 6644 2010 6656
rect 2593 6647 2651 6653
rect 2593 6644 2605 6647
rect 2004 6616 2605 6644
rect 2004 6604 2010 6616
rect 2593 6613 2605 6616
rect 2639 6613 2651 6647
rect 2593 6607 2651 6613
rect 3694 6604 3700 6656
rect 3752 6644 3758 6656
rect 3973 6647 4031 6653
rect 3973 6644 3985 6647
rect 3752 6616 3985 6644
rect 3752 6604 3758 6616
rect 3973 6613 3985 6616
rect 4019 6613 4031 6647
rect 3973 6607 4031 6613
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 9030 6644 9036 6656
rect 6512 6616 9036 6644
rect 6512 6604 6518 6616
rect 9030 6604 9036 6616
rect 9088 6604 9094 6656
rect 10137 6647 10195 6653
rect 10137 6613 10149 6647
rect 10183 6644 10195 6647
rect 10226 6644 10232 6656
rect 10183 6616 10232 6644
rect 10183 6613 10195 6616
rect 10137 6607 10195 6613
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 10502 6604 10508 6656
rect 10560 6604 10566 6656
rect 10597 6647 10655 6653
rect 10597 6613 10609 6647
rect 10643 6644 10655 6647
rect 10686 6644 10692 6656
rect 10643 6616 10692 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 10686 6604 10692 6616
rect 10744 6604 10750 6656
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 10928 6616 11345 6644
rect 10928 6604 10934 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 13096 6644 13124 6743
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 15470 6740 15476 6792
rect 15528 6740 15534 6792
rect 16758 6740 16764 6792
rect 16816 6740 16822 6792
rect 17865 6783 17923 6789
rect 17865 6749 17877 6783
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 13906 6672 13912 6724
rect 13964 6712 13970 6724
rect 16022 6712 16028 6724
rect 13964 6684 16028 6712
rect 13964 6672 13970 6684
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 16390 6672 16396 6724
rect 16448 6712 16454 6724
rect 17880 6712 17908 6743
rect 16448 6684 17908 6712
rect 17972 6712 18000 6820
rect 18506 6808 18512 6860
rect 18564 6808 18570 6860
rect 19306 6848 19334 6956
rect 20165 6953 20177 6987
rect 20211 6984 20223 6987
rect 20530 6984 20536 6996
rect 20211 6956 20536 6984
rect 20211 6953 20223 6956
rect 20165 6947 20223 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 22278 6944 22284 6996
rect 22336 6984 22342 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 22336 6956 22477 6984
rect 22336 6944 22342 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22465 6947 22523 6953
rect 22830 6944 22836 6996
rect 22888 6984 22894 6996
rect 23845 6987 23903 6993
rect 23845 6984 23857 6987
rect 22888 6956 23857 6984
rect 22888 6944 22894 6956
rect 23845 6953 23857 6956
rect 23891 6953 23903 6987
rect 23845 6947 23903 6953
rect 25314 6944 25320 6996
rect 25372 6984 25378 6996
rect 26878 6984 26884 6996
rect 25372 6956 26884 6984
rect 25372 6944 25378 6956
rect 26878 6944 26884 6956
rect 26936 6944 26942 6996
rect 26878 6848 26884 6860
rect 19306 6820 26884 6848
rect 26878 6808 26884 6820
rect 26936 6808 26942 6860
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19521 6783 19579 6789
rect 19521 6780 19533 6783
rect 19392 6752 19533 6780
rect 19392 6740 19398 6752
rect 19521 6749 19533 6752
rect 19567 6749 19579 6783
rect 19521 6743 19579 6749
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6780 20683 6783
rect 20806 6780 20812 6792
rect 20671 6752 20812 6780
rect 20671 6749 20683 6752
rect 20625 6743 20683 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21269 6783 21327 6789
rect 21269 6749 21281 6783
rect 21315 6780 21327 6783
rect 21821 6783 21879 6789
rect 21821 6780 21833 6783
rect 21315 6752 21833 6780
rect 21315 6749 21327 6752
rect 21269 6743 21327 6749
rect 21821 6749 21833 6752
rect 21867 6749 21879 6783
rect 21821 6743 21879 6749
rect 21726 6712 21732 6724
rect 17972 6684 21732 6712
rect 16448 6672 16454 6684
rect 21726 6672 21732 6684
rect 21784 6672 21790 6724
rect 23014 6672 23020 6724
rect 23072 6672 23078 6724
rect 23198 6672 23204 6724
rect 23256 6672 23262 6724
rect 15194 6644 15200 6656
rect 13096 6616 15200 6644
rect 11333 6607 11391 6613
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 17586 6604 17592 6656
rect 17644 6644 17650 6656
rect 21174 6644 21180 6656
rect 17644 6616 21180 6644
rect 17644 6604 17650 6616
rect 21174 6604 21180 6616
rect 21232 6604 21238 6656
rect 24118 6604 24124 6656
rect 24176 6644 24182 6656
rect 30466 6644 30472 6656
rect 24176 6616 30472 6644
rect 24176 6604 24182 6616
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3970 6440 3976 6452
rect 3384 6412 3976 6440
rect 3384 6400 3390 6412
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 4062 6400 4068 6452
rect 4120 6440 4126 6452
rect 4120 6412 4844 6440
rect 4120 6400 4126 6412
rect 3786 6332 3792 6384
rect 3844 6372 3850 6384
rect 4816 6372 4844 6412
rect 4890 6400 4896 6452
rect 4948 6400 4954 6452
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 10045 6443 10103 6449
rect 10045 6440 10057 6443
rect 5684 6412 10057 6440
rect 5684 6400 5690 6412
rect 10045 6409 10057 6412
rect 10091 6409 10103 6443
rect 12621 6443 12679 6449
rect 12621 6440 12633 6443
rect 10045 6403 10103 6409
rect 10152 6412 12633 6440
rect 3844 6344 4292 6372
rect 4816 6344 7328 6372
rect 3844 6332 3850 6344
rect 1302 6264 1308 6316
rect 1360 6304 1366 6316
rect 1581 6307 1639 6313
rect 1581 6304 1593 6307
rect 1360 6276 1593 6304
rect 1360 6264 1366 6276
rect 1581 6273 1593 6276
rect 1627 6304 1639 6307
rect 1946 6304 1952 6316
rect 1627 6276 1952 6304
rect 1627 6273 1639 6276
rect 1581 6267 1639 6273
rect 1946 6264 1952 6276
rect 2004 6264 2010 6316
rect 3053 6307 3111 6313
rect 3053 6273 3065 6307
rect 3099 6273 3111 6307
rect 3053 6267 3111 6273
rect 3605 6308 3663 6313
rect 3605 6307 3740 6308
rect 3605 6273 3617 6307
rect 3651 6304 3740 6307
rect 4062 6304 4068 6316
rect 3651 6280 4068 6304
rect 3651 6273 3663 6280
rect 3712 6276 4068 6280
rect 3605 6267 3663 6273
rect 1857 6239 1915 6245
rect 1857 6205 1869 6239
rect 1903 6236 1915 6239
rect 2682 6236 2688 6248
rect 1903 6208 2688 6236
rect 1903 6205 1915 6208
rect 1857 6199 1915 6205
rect 2682 6196 2688 6208
rect 2740 6196 2746 6248
rect 3068 6236 3096 6267
rect 4062 6264 4068 6276
rect 4120 6264 4126 6316
rect 4264 6313 4292 6344
rect 4249 6307 4307 6313
rect 4249 6273 4261 6307
rect 4295 6273 4307 6307
rect 4249 6267 4307 6273
rect 5350 6264 5356 6316
rect 5408 6264 5414 6316
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 7300 6304 7328 6344
rect 7742 6332 7748 6384
rect 7800 6372 7806 6384
rect 7837 6375 7895 6381
rect 7837 6372 7849 6375
rect 7800 6344 7849 6372
rect 7800 6332 7806 6344
rect 7837 6341 7849 6344
rect 7883 6341 7895 6375
rect 8941 6375 8999 6381
rect 8941 6372 8953 6375
rect 7837 6335 7895 6341
rect 7944 6344 8953 6372
rect 7944 6304 7972 6344
rect 8941 6341 8953 6344
rect 8987 6341 8999 6375
rect 8941 6335 8999 6341
rect 9030 6332 9036 6384
rect 9088 6372 9094 6384
rect 10152 6372 10180 6412
rect 12621 6409 12633 6412
rect 12667 6409 12679 6443
rect 12621 6403 12679 6409
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 16758 6440 16764 6452
rect 15243 6412 16764 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 17497 6443 17555 6449
rect 17497 6409 17509 6443
rect 17543 6440 17555 6443
rect 17770 6440 17776 6452
rect 17543 6412 17776 6440
rect 17543 6409 17555 6412
rect 17497 6403 17555 6409
rect 17770 6400 17776 6412
rect 17828 6400 17834 6452
rect 19705 6443 19763 6449
rect 19705 6440 19717 6443
rect 18340 6412 19717 6440
rect 9088 6344 10180 6372
rect 9088 6332 9094 6344
rect 10686 6332 10692 6384
rect 10744 6372 10750 6384
rect 16206 6372 16212 6384
rect 10744 6344 13400 6372
rect 10744 6332 10750 6344
rect 7300 6276 7972 6304
rect 7193 6267 7251 6273
rect 3068 6208 3648 6236
rect 2869 6171 2927 6177
rect 2869 6137 2881 6171
rect 2915 6168 2927 6171
rect 3510 6168 3516 6180
rect 2915 6140 3516 6168
rect 2915 6137 2927 6140
rect 2869 6131 2927 6137
rect 3510 6128 3516 6140
rect 3568 6128 3574 6180
rect 3620 6168 3648 6208
rect 3970 6196 3976 6248
rect 4028 6236 4034 6248
rect 5997 6239 6055 6245
rect 5997 6236 6009 6239
rect 4028 6208 6009 6236
rect 4028 6196 4034 6208
rect 5997 6205 6009 6208
rect 6043 6205 6055 6239
rect 5997 6199 6055 6205
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 6512 6208 6561 6236
rect 6512 6196 6518 6208
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 7208 6236 7236 6267
rect 8294 6264 8300 6316
rect 8352 6264 8358 6316
rect 9401 6307 9459 6313
rect 9401 6273 9413 6307
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 10505 6307 10563 6313
rect 10505 6273 10517 6307
rect 10551 6304 10563 6307
rect 10962 6304 10968 6316
rect 10551 6276 10968 6304
rect 10551 6273 10563 6276
rect 10505 6267 10563 6273
rect 8938 6236 8944 6248
rect 7208 6208 8944 6236
rect 6549 6199 6607 6205
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 9416 6236 9444 6267
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12158 6304 12164 6316
rect 12023 6276 12164 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 11054 6236 11060 6248
rect 9416 6208 11060 6236
rect 11054 6196 11060 6208
rect 11112 6196 11118 6248
rect 13372 6236 13400 6344
rect 13464 6344 16212 6372
rect 13464 6313 13492 6344
rect 16206 6332 16212 6344
rect 16264 6332 16270 6384
rect 16298 6332 16304 6384
rect 16356 6332 16362 6384
rect 16942 6332 16948 6384
rect 17000 6372 17006 6384
rect 18340 6372 18368 6412
rect 19705 6409 19717 6412
rect 19751 6409 19763 6443
rect 19705 6403 19763 6409
rect 20806 6400 20812 6452
rect 20864 6400 20870 6452
rect 21269 6443 21327 6449
rect 21269 6409 21281 6443
rect 21315 6440 21327 6443
rect 23014 6440 23020 6452
rect 21315 6412 23020 6440
rect 21315 6409 21327 6412
rect 21269 6403 21327 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23290 6400 23296 6452
rect 23348 6440 23354 6452
rect 23753 6443 23811 6449
rect 23753 6440 23765 6443
rect 23348 6412 23765 6440
rect 23348 6400 23354 6412
rect 23753 6409 23765 6412
rect 23799 6440 23811 6443
rect 26234 6440 26240 6452
rect 23799 6412 26240 6440
rect 23799 6409 23811 6412
rect 23753 6403 23811 6409
rect 26234 6400 26240 6412
rect 26292 6400 26298 6452
rect 26878 6400 26884 6452
rect 26936 6440 26942 6452
rect 33870 6440 33876 6452
rect 26936 6412 33876 6440
rect 26936 6400 26942 6412
rect 33870 6400 33876 6412
rect 33928 6400 33934 6452
rect 26050 6372 26056 6384
rect 17000 6344 18368 6372
rect 19076 6344 26056 6372
rect 17000 6332 17006 6344
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6273 13507 6307
rect 13449 6267 13507 6273
rect 13722 6264 13728 6316
rect 13780 6304 13786 6316
rect 14553 6307 14611 6313
rect 14553 6304 14565 6307
rect 13780 6276 14565 6304
rect 13780 6264 13786 6276
rect 14553 6273 14565 6276
rect 14599 6273 14611 6307
rect 14553 6267 14611 6273
rect 15654 6264 15660 6316
rect 15712 6264 15718 6316
rect 19076 6313 19104 6344
rect 26050 6332 26056 6344
rect 26108 6332 26114 6384
rect 16853 6307 16911 6313
rect 16853 6273 16865 6307
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6304 18015 6307
rect 19061 6307 19119 6313
rect 18003 6276 19012 6304
rect 18003 6273 18015 6276
rect 17957 6267 18015 6273
rect 16758 6236 16764 6248
rect 13372 6208 16764 6236
rect 16758 6196 16764 6208
rect 16816 6196 16822 6248
rect 16868 6236 16896 6267
rect 18601 6239 18659 6245
rect 18601 6236 18613 6239
rect 16868 6208 18613 6236
rect 18601 6205 18613 6208
rect 18647 6205 18659 6239
rect 18984 6236 19012 6276
rect 19061 6273 19073 6307
rect 19107 6273 19119 6307
rect 19061 6267 19119 6273
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 20990 6304 20996 6316
rect 20211 6276 20996 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 21450 6264 21456 6316
rect 21508 6264 21514 6316
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 22465 6307 22523 6313
rect 22465 6304 22477 6307
rect 22244 6276 22477 6304
rect 22244 6264 22250 6276
rect 22465 6273 22477 6276
rect 22511 6273 22523 6307
rect 22465 6267 22523 6273
rect 22830 6264 22836 6316
rect 22888 6304 22894 6316
rect 23290 6304 23296 6316
rect 22888 6276 23296 6304
rect 22888 6264 22894 6276
rect 23290 6264 23296 6276
rect 23348 6264 23354 6316
rect 25222 6236 25228 6248
rect 18984 6208 25228 6236
rect 18601 6199 18659 6205
rect 25222 6196 25228 6208
rect 25280 6196 25286 6248
rect 27614 6196 27620 6248
rect 27672 6236 27678 6248
rect 43622 6236 43628 6248
rect 27672 6208 43628 6236
rect 27672 6196 27678 6208
rect 43622 6196 43628 6208
rect 43680 6196 43686 6248
rect 3620 6140 4108 6168
rect 3326 6060 3332 6112
rect 3384 6100 3390 6112
rect 3697 6103 3755 6109
rect 3697 6100 3709 6103
rect 3384 6072 3709 6100
rect 3384 6060 3390 6072
rect 3697 6069 3709 6072
rect 3743 6069 3755 6103
rect 4080 6100 4108 6140
rect 4154 6128 4160 6180
rect 4212 6168 4218 6180
rect 4212 6140 6592 6168
rect 4212 6128 4218 6140
rect 6362 6100 6368 6112
rect 4080 6072 6368 6100
rect 3697 6063 3755 6069
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6454 6060 6460 6112
rect 6512 6060 6518 6112
rect 6564 6100 6592 6140
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 13081 6171 13139 6177
rect 13081 6168 13093 6171
rect 6788 6140 13093 6168
rect 6788 6128 6794 6140
rect 13081 6137 13093 6140
rect 13127 6137 13139 6171
rect 13081 6131 13139 6137
rect 14182 6128 14188 6180
rect 14240 6168 14246 6180
rect 14240 6140 17264 6168
rect 14240 6128 14246 6140
rect 9858 6100 9864 6112
rect 6564 6072 9864 6100
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 11146 6060 11152 6112
rect 11204 6060 11210 6112
rect 11698 6060 11704 6112
rect 11756 6060 11762 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 12897 6103 12955 6109
rect 12897 6100 12909 6103
rect 12768 6072 12909 6100
rect 12768 6060 12774 6072
rect 12897 6069 12909 6072
rect 12943 6069 12955 6103
rect 12897 6063 12955 6069
rect 14093 6103 14151 6109
rect 14093 6069 14105 6103
rect 14139 6100 14151 6103
rect 14550 6100 14556 6112
rect 14139 6072 14556 6100
rect 14139 6069 14151 6072
rect 14093 6063 14151 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 17126 6100 17132 6112
rect 14884 6072 17132 6100
rect 14884 6060 14890 6072
rect 17126 6060 17132 6072
rect 17184 6060 17190 6112
rect 17236 6100 17264 6140
rect 18322 6128 18328 6180
rect 18380 6168 18386 6180
rect 21542 6168 21548 6180
rect 18380 6140 21548 6168
rect 18380 6128 18386 6140
rect 21542 6128 21548 6140
rect 21600 6128 21606 6180
rect 23750 6168 23756 6180
rect 23124 6140 23756 6168
rect 23124 6109 23152 6140
rect 23750 6128 23756 6140
rect 23808 6128 23814 6180
rect 26142 6128 26148 6180
rect 26200 6168 26206 6180
rect 42058 6168 42064 6180
rect 26200 6140 42064 6168
rect 26200 6128 26206 6140
rect 42058 6128 42064 6140
rect 42116 6128 42122 6180
rect 22005 6103 22063 6109
rect 22005 6100 22017 6103
rect 17236 6072 22017 6100
rect 22005 6069 22017 6072
rect 22051 6069 22063 6103
rect 22005 6063 22063 6069
rect 23109 6103 23167 6109
rect 23109 6069 23121 6103
rect 23155 6069 23167 6103
rect 23109 6063 23167 6069
rect 23290 6060 23296 6112
rect 23348 6060 23354 6112
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 2777 5899 2835 5905
rect 2777 5865 2789 5899
rect 2823 5896 2835 5899
rect 4430 5896 4436 5908
rect 2823 5868 4436 5896
rect 2823 5865 2835 5868
rect 2777 5859 2835 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 5442 5856 5448 5908
rect 5500 5856 5506 5908
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7469 5899 7527 5905
rect 7469 5896 7481 5899
rect 7432 5868 7481 5896
rect 7432 5856 7438 5868
rect 7469 5865 7481 5868
rect 7515 5865 7527 5899
rect 7469 5859 7527 5865
rect 10226 5856 10232 5908
rect 10284 5896 10290 5908
rect 10413 5899 10471 5905
rect 10413 5896 10425 5899
rect 10284 5868 10425 5896
rect 10284 5856 10290 5868
rect 10413 5865 10425 5868
rect 10459 5865 10471 5899
rect 10413 5859 10471 5865
rect 11517 5899 11575 5905
rect 11517 5865 11529 5899
rect 11563 5896 11575 5899
rect 11606 5896 11612 5908
rect 11563 5868 11612 5896
rect 11563 5865 11575 5868
rect 11517 5859 11575 5865
rect 11606 5856 11612 5868
rect 11664 5856 11670 5908
rect 12621 5899 12679 5905
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12802 5896 12808 5908
rect 12667 5868 12808 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13722 5856 13728 5908
rect 13780 5856 13786 5908
rect 19337 5899 19395 5905
rect 19337 5896 19349 5899
rect 13924 5868 19349 5896
rect 750 5788 756 5840
rect 808 5828 814 5840
rect 3326 5828 3332 5840
rect 808 5800 3332 5828
rect 808 5788 814 5800
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 3418 5788 3424 5840
rect 3476 5788 3482 5840
rect 3694 5788 3700 5840
rect 3752 5828 3758 5840
rect 13924 5828 13952 5868
rect 3752 5800 13952 5828
rect 3752 5788 3758 5800
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5760 1915 5763
rect 2038 5760 2044 5772
rect 1903 5732 2044 5760
rect 1903 5729 1915 5732
rect 1857 5723 1915 5729
rect 2038 5720 2044 5732
rect 2096 5720 2102 5772
rect 4893 5763 4951 5769
rect 4893 5760 4905 5763
rect 2746 5732 4905 5760
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1578 5692 1584 5704
rect 1360 5664 1584 5692
rect 1360 5652 1366 5664
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 2746 5556 2774 5732
rect 4893 5729 4905 5732
rect 4939 5729 4951 5763
rect 6365 5763 6423 5769
rect 6365 5760 6377 5763
rect 4893 5723 4951 5729
rect 5276 5732 6377 5760
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3786 5692 3792 5704
rect 3283 5664 3792 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5692 4307 5695
rect 5276 5692 5304 5732
rect 6365 5729 6377 5732
rect 6411 5729 6423 5763
rect 6365 5723 6423 5729
rect 9125 5763 9183 5769
rect 9125 5729 9137 5763
rect 9171 5760 9183 5763
rect 9306 5760 9312 5772
rect 9171 5732 9312 5760
rect 9171 5729 9183 5732
rect 9125 5723 9183 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 9950 5720 9956 5772
rect 10008 5760 10014 5772
rect 10008 5732 12020 5760
rect 10008 5720 10014 5732
rect 4295 5664 5304 5692
rect 4295 5661 4307 5664
rect 4249 5655 4307 5661
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5721 5695 5779 5701
rect 5721 5692 5733 5695
rect 5592 5664 5733 5692
rect 5592 5652 5598 5664
rect 5721 5661 5733 5664
rect 5767 5661 5779 5695
rect 5721 5655 5779 5661
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 7466 5692 7472 5704
rect 6871 5664 7472 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 7466 5652 7472 5664
rect 7524 5652 7530 5704
rect 7926 5652 7932 5704
rect 7984 5652 7990 5704
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 11992 5701 12020 5732
rect 15286 5720 15292 5772
rect 15344 5720 15350 5772
rect 16850 5720 16856 5772
rect 16908 5760 16914 5772
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16908 5732 17141 5760
rect 16908 5720 16914 5732
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 17405 5763 17463 5769
rect 17405 5729 17417 5763
rect 17451 5760 17463 5763
rect 18598 5760 18604 5772
rect 17451 5732 18604 5760
rect 17451 5729 17463 5732
rect 17405 5723 17463 5729
rect 18598 5720 18604 5732
rect 18656 5720 18662 5772
rect 18800 5760 18828 5868
rect 19337 5865 19349 5868
rect 19383 5865 19395 5899
rect 19337 5859 19395 5865
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 23842 5896 23848 5908
rect 20763 5868 23848 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 23842 5856 23848 5868
rect 23900 5856 23906 5908
rect 18877 5831 18935 5837
rect 18877 5797 18889 5831
rect 18923 5828 18935 5831
rect 20990 5828 20996 5840
rect 18923 5800 20996 5828
rect 18923 5797 18935 5800
rect 18877 5791 18935 5797
rect 20990 5788 20996 5800
rect 21048 5788 21054 5840
rect 21174 5788 21180 5840
rect 21232 5788 21238 5840
rect 30650 5828 30656 5840
rect 23308 5800 30656 5828
rect 19429 5763 19487 5769
rect 19429 5760 19441 5763
rect 18800 5732 19441 5760
rect 19429 5729 19441 5732
rect 19475 5729 19487 5763
rect 19429 5723 19487 5729
rect 19702 5720 19708 5772
rect 19760 5720 19766 5772
rect 23308 5769 23336 5800
rect 30650 5788 30656 5800
rect 30708 5788 30714 5840
rect 21637 5763 21695 5769
rect 21637 5760 21649 5763
rect 19812 5732 21649 5760
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5661 12035 5695
rect 11977 5655 12035 5661
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13081 5695 13139 5701
rect 12492 5664 12940 5692
rect 12492 5652 12498 5664
rect 3881 5627 3939 5633
rect 3881 5593 3893 5627
rect 3927 5624 3939 5627
rect 4614 5624 4620 5636
rect 3927 5596 4620 5624
rect 3927 5593 3939 5596
rect 3881 5587 3939 5593
rect 4614 5584 4620 5596
rect 4672 5584 4678 5636
rect 6546 5584 6552 5636
rect 6604 5624 6610 5636
rect 6604 5596 9674 5624
rect 6604 5584 6610 5596
rect 1912 5528 2774 5556
rect 1912 5516 1918 5528
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5166 5556 5172 5568
rect 4948 5528 5172 5556
rect 4948 5516 4954 5528
rect 5166 5516 5172 5528
rect 5224 5516 5230 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8573 5559 8631 5565
rect 8573 5556 8585 5559
rect 8352 5528 8585 5556
rect 8352 5516 8358 5528
rect 8573 5525 8585 5528
rect 8619 5525 8631 5559
rect 9646 5556 9674 5596
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 12802 5624 12808 5636
rect 11848 5596 12808 5624
rect 11848 5584 11854 5596
rect 12802 5584 12808 5596
rect 12860 5584 12866 5636
rect 12912 5624 12940 5664
rect 13081 5661 13093 5695
rect 13127 5692 13139 5695
rect 13906 5692 13912 5704
rect 13127 5664 13912 5692
rect 13127 5661 13139 5664
rect 13081 5655 13139 5661
rect 13906 5652 13912 5664
rect 13964 5652 13970 5704
rect 14274 5652 14280 5704
rect 14332 5652 14338 5704
rect 19150 5652 19156 5704
rect 19208 5692 19214 5704
rect 19812 5692 19840 5732
rect 21637 5729 21649 5732
rect 21683 5729 21695 5763
rect 21637 5723 21695 5729
rect 23293 5763 23351 5769
rect 23293 5729 23305 5763
rect 23339 5729 23351 5763
rect 23293 5723 23351 5729
rect 23845 5763 23903 5769
rect 23845 5729 23857 5763
rect 23891 5760 23903 5763
rect 27706 5760 27712 5772
rect 23891 5732 27712 5760
rect 23891 5729 23903 5732
rect 23845 5723 23903 5729
rect 19208 5664 19840 5692
rect 19208 5652 19214 5664
rect 20346 5652 20352 5704
rect 20404 5692 20410 5704
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 20404 5664 20913 5692
rect 20404 5652 20410 5664
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21361 5695 21419 5701
rect 21361 5692 21373 5695
rect 21232 5664 21373 5692
rect 21232 5652 21238 5664
rect 21361 5661 21373 5664
rect 21407 5661 21419 5695
rect 22700 5695 22758 5701
rect 22700 5692 22712 5695
rect 21361 5655 21419 5661
rect 22066 5664 22712 5692
rect 14461 5627 14519 5633
rect 14461 5624 14473 5627
rect 12912 5596 14473 5624
rect 14461 5593 14473 5596
rect 14507 5624 14519 5627
rect 14507 5596 16528 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 12526 5556 12532 5568
rect 9646 5528 12532 5556
rect 8573 5519 8631 5525
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 15102 5556 15108 5568
rect 13596 5528 15108 5556
rect 13596 5516 13602 5528
rect 15102 5516 15108 5528
rect 15160 5516 15166 5568
rect 16500 5565 16528 5596
rect 17310 5584 17316 5636
rect 17368 5624 17374 5636
rect 22066 5624 22094 5664
rect 22700 5661 22712 5664
rect 22746 5692 22758 5695
rect 23860 5692 23888 5723
rect 27706 5720 27712 5732
rect 27764 5720 27770 5772
rect 22746 5664 23888 5692
rect 22746 5661 22758 5664
rect 22700 5655 22758 5661
rect 17368 5596 17894 5624
rect 18708 5596 22094 5624
rect 22787 5627 22845 5633
rect 17368 5584 17374 5596
rect 16485 5559 16543 5565
rect 16485 5525 16497 5559
rect 16531 5556 16543 5559
rect 18708 5556 18736 5596
rect 22787 5593 22799 5627
rect 22833 5624 22845 5627
rect 24946 5624 24952 5636
rect 22833 5596 24952 5624
rect 22833 5593 22845 5596
rect 22787 5587 22845 5593
rect 24946 5584 24952 5596
rect 25004 5584 25010 5636
rect 16531 5528 18736 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 23750 5516 23756 5568
rect 23808 5556 23814 5568
rect 27062 5556 27068 5568
rect 23808 5528 27068 5556
rect 23808 5516 23814 5528
rect 27062 5516 27068 5528
rect 27120 5516 27126 5568
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 2406 5312 2412 5364
rect 2464 5352 2470 5364
rect 3418 5352 3424 5364
rect 2464 5324 3424 5352
rect 2464 5312 2470 5324
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 3878 5312 3884 5364
rect 3936 5312 3942 5364
rect 4157 5355 4215 5361
rect 4157 5321 4169 5355
rect 4203 5352 4215 5355
rect 5074 5352 5080 5364
rect 4203 5324 5080 5352
rect 4203 5321 4215 5324
rect 4157 5315 4215 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 6549 5355 6607 5361
rect 6549 5321 6561 5355
rect 6595 5352 6607 5355
rect 7190 5352 7196 5364
rect 6595 5324 7196 5352
rect 6595 5321 6607 5324
rect 6549 5315 6607 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 7742 5312 7748 5364
rect 7800 5352 7806 5364
rect 7837 5355 7895 5361
rect 7837 5352 7849 5355
rect 7800 5324 7849 5352
rect 7800 5312 7806 5324
rect 7837 5321 7849 5324
rect 7883 5321 7895 5355
rect 7837 5315 7895 5321
rect 8938 5312 8944 5364
rect 8996 5312 9002 5364
rect 11330 5312 11336 5364
rect 11388 5352 11394 5364
rect 11609 5355 11667 5361
rect 11609 5352 11621 5355
rect 11388 5324 11621 5352
rect 11388 5312 11394 5324
rect 11609 5321 11621 5324
rect 11655 5352 11667 5355
rect 12066 5352 12072 5364
rect 11655 5324 12072 5352
rect 11655 5321 11667 5324
rect 11609 5315 11667 5321
rect 12066 5312 12072 5324
rect 12124 5312 12130 5364
rect 12802 5312 12808 5364
rect 12860 5312 12866 5364
rect 13446 5312 13452 5364
rect 13504 5352 13510 5364
rect 13504 5324 14136 5352
rect 13504 5312 13510 5324
rect 2222 5244 2228 5296
rect 2280 5284 2286 5296
rect 5261 5287 5319 5293
rect 5261 5284 5273 5287
rect 2280 5256 5273 5284
rect 2280 5244 2286 5256
rect 5261 5253 5273 5256
rect 5307 5253 5319 5287
rect 5261 5247 5319 5253
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 8386 5284 8392 5296
rect 5859 5256 8392 5284
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 9122 5244 9128 5296
rect 9180 5284 9186 5296
rect 9180 5256 10548 5284
rect 9180 5244 9186 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 4522 5216 4528 5228
rect 1719 5188 4528 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 4522 5176 4528 5188
rect 4580 5176 4586 5228
rect 4617 5219 4675 5225
rect 4617 5185 4629 5219
rect 4663 5216 4675 5219
rect 5718 5216 5724 5228
rect 4663 5188 5724 5216
rect 4663 5185 4675 5188
rect 4617 5179 4675 5185
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 7193 5219 7251 5225
rect 7193 5185 7205 5219
rect 7239 5216 7251 5219
rect 8202 5216 8208 5228
rect 7239 5188 8208 5216
rect 7239 5185 7251 5188
rect 7193 5179 7251 5185
rect 8202 5176 8208 5188
rect 8260 5176 8266 5228
rect 8294 5176 8300 5228
rect 8352 5176 8358 5228
rect 9401 5219 9459 5225
rect 9401 5185 9413 5219
rect 9447 5216 9459 5219
rect 10134 5216 10140 5228
rect 9447 5188 10140 5216
rect 9447 5185 9459 5188
rect 9401 5179 9459 5185
rect 10134 5176 10140 5188
rect 10192 5176 10198 5228
rect 10520 5225 10548 5256
rect 10962 5244 10968 5296
rect 11020 5284 11026 5296
rect 14001 5287 14059 5293
rect 14001 5284 14013 5287
rect 11020 5256 14013 5284
rect 11020 5244 11026 5256
rect 14001 5253 14013 5256
rect 14047 5253 14059 5287
rect 14108 5284 14136 5324
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 17402 5352 17408 5364
rect 15304 5324 17408 5352
rect 15304 5284 15332 5324
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 18322 5352 18328 5364
rect 17543 5324 18328 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 18322 5312 18328 5324
rect 18380 5312 18386 5364
rect 21174 5312 21180 5364
rect 21232 5352 21238 5364
rect 21545 5355 21603 5361
rect 21545 5352 21557 5355
rect 21232 5324 21557 5352
rect 21232 5312 21238 5324
rect 21545 5321 21557 5324
rect 21591 5321 21603 5355
rect 29730 5352 29736 5364
rect 21545 5315 21603 5321
rect 22066 5324 29736 5352
rect 19426 5284 19432 5296
rect 14108 5256 15332 5284
rect 16868 5256 19432 5284
rect 14001 5247 14059 5253
rect 10505 5219 10563 5225
rect 10505 5185 10517 5219
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11149 5219 11207 5225
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 12161 5219 12219 5225
rect 12161 5216 12173 5219
rect 11195 5188 12173 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 12161 5185 12173 5188
rect 12207 5185 12219 5219
rect 12161 5179 12219 5185
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 12710 5216 12716 5228
rect 12492 5188 12716 5216
rect 12492 5176 12498 5188
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 13354 5176 13360 5228
rect 13412 5176 13418 5228
rect 14550 5176 14556 5228
rect 14608 5176 14614 5228
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 15838 5216 15844 5228
rect 15703 5188 15844 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 16868 5225 16896 5256
rect 19426 5244 19432 5256
rect 19484 5244 19490 5296
rect 19610 5244 19616 5296
rect 19668 5284 19674 5296
rect 22066 5284 22094 5324
rect 29730 5312 29736 5324
rect 29788 5312 29794 5364
rect 19668 5256 22094 5284
rect 22741 5287 22799 5293
rect 19668 5244 19674 5256
rect 22741 5253 22753 5287
rect 22787 5284 22799 5287
rect 22833 5287 22891 5293
rect 22833 5284 22845 5287
rect 22787 5256 22845 5284
rect 22787 5253 22799 5256
rect 22741 5247 22799 5253
rect 22833 5253 22845 5256
rect 22879 5284 22891 5287
rect 23658 5284 23664 5296
rect 22879 5256 23664 5284
rect 22879 5253 22891 5256
rect 22833 5247 22891 5253
rect 23658 5244 23664 5256
rect 23716 5244 23722 5296
rect 24946 5244 24952 5296
rect 25004 5244 25010 5296
rect 26605 5287 26663 5293
rect 26605 5253 26617 5287
rect 26651 5284 26663 5287
rect 27522 5284 27528 5296
rect 26651 5256 27528 5284
rect 26651 5253 26663 5256
rect 26605 5247 26663 5253
rect 27522 5244 27528 5256
rect 27580 5284 27586 5296
rect 31297 5287 31355 5293
rect 27580 5256 31248 5284
rect 27580 5244 27586 5256
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17000 5188 18644 5216
rect 17000 5176 17006 5188
rect 2777 5151 2835 5157
rect 2777 5117 2789 5151
rect 2823 5148 2835 5151
rect 2958 5148 2964 5160
rect 2823 5120 2964 5148
rect 2823 5117 2835 5120
rect 2777 5111 2835 5117
rect 2958 5108 2964 5120
rect 3016 5108 3022 5160
rect 3053 5151 3111 5157
rect 3053 5117 3065 5151
rect 3099 5117 3111 5151
rect 3053 5111 3111 5117
rect 658 5040 664 5092
rect 716 5080 722 5092
rect 3068 5080 3096 5111
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 10410 5148 10416 5160
rect 9272 5120 10416 5148
rect 9272 5108 9278 5120
rect 10410 5108 10416 5120
rect 10468 5108 10474 5160
rect 11698 5108 11704 5160
rect 11756 5108 11762 5160
rect 13906 5108 13912 5160
rect 13964 5148 13970 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 13964 5120 18061 5148
rect 13964 5108 13970 5120
rect 18049 5117 18061 5120
rect 18095 5148 18107 5151
rect 18417 5151 18475 5157
rect 18417 5148 18429 5151
rect 18095 5120 18429 5148
rect 18095 5117 18107 5120
rect 18049 5111 18107 5117
rect 18417 5117 18429 5120
rect 18463 5117 18475 5151
rect 18616 5148 18644 5188
rect 18690 5176 18696 5228
rect 18748 5176 18754 5228
rect 19794 5216 19800 5228
rect 18800 5188 19800 5216
rect 18800 5148 18828 5188
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 19978 5176 19984 5228
rect 20036 5176 20042 5228
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5216 21143 5219
rect 21266 5216 21272 5228
rect 21131 5188 21272 5216
rect 21131 5185 21143 5188
rect 21085 5179 21143 5185
rect 21266 5176 21272 5188
rect 21324 5216 21330 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21324 5188 21833 5216
rect 21324 5176 21330 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 22186 5176 22192 5228
rect 22244 5224 22250 5228
rect 22244 5218 22282 5224
rect 22270 5216 22282 5218
rect 23290 5216 23296 5228
rect 22270 5188 23296 5216
rect 22270 5187 22299 5188
rect 22270 5184 22282 5187
rect 22244 5178 22282 5184
rect 22244 5176 22250 5178
rect 23290 5176 23296 5188
rect 23348 5176 23354 5228
rect 31220 5216 31248 5256
rect 31297 5253 31309 5287
rect 31343 5284 31355 5287
rect 31754 5284 31760 5296
rect 31343 5256 31760 5284
rect 31343 5253 31355 5256
rect 31297 5247 31355 5253
rect 31754 5244 31760 5256
rect 31812 5244 31818 5296
rect 31220 5188 38654 5216
rect 18616 5120 18828 5148
rect 18417 5111 18475 5117
rect 18874 5108 18880 5160
rect 18932 5148 18938 5160
rect 19705 5151 19763 5157
rect 19705 5148 19717 5151
rect 18932 5120 19717 5148
rect 18932 5108 18938 5120
rect 19705 5117 19717 5120
rect 19751 5117 19763 5151
rect 24302 5148 24308 5160
rect 19705 5111 19763 5117
rect 19812 5120 24308 5148
rect 716 5052 3096 5080
rect 5997 5083 6055 5089
rect 716 5040 722 5052
rect 5997 5049 6009 5083
rect 6043 5080 6055 5083
rect 6362 5080 6368 5092
rect 6043 5052 6368 5080
rect 6043 5049 6055 5052
rect 5997 5043 6055 5049
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 15654 5080 15660 5092
rect 7300 5052 15660 5080
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2317 5015 2375 5021
rect 2317 5012 2329 5015
rect 1728 4984 2329 5012
rect 1728 4972 1734 4984
rect 2317 4981 2329 4984
rect 2363 4981 2375 5015
rect 2317 4975 2375 4981
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 5442 5012 5448 5024
rect 4387 4984 5448 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 6178 4972 6184 5024
rect 6236 5012 6242 5024
rect 7300 5012 7328 5052
rect 15654 5040 15660 5052
rect 15712 5040 15718 5092
rect 19812 5080 19840 5120
rect 24302 5108 24308 5120
rect 24360 5108 24366 5160
rect 24765 5151 24823 5157
rect 24765 5117 24777 5151
rect 24811 5117 24823 5151
rect 24765 5111 24823 5117
rect 27157 5151 27215 5157
rect 27157 5117 27169 5151
rect 27203 5117 27215 5151
rect 27157 5111 27215 5117
rect 24780 5080 24808 5111
rect 25498 5080 25504 5092
rect 15764 5052 19840 5080
rect 19904 5052 24716 5080
rect 24780 5052 25504 5080
rect 6236 4984 7328 5012
rect 6236 4972 6242 4984
rect 9306 4972 9312 5024
rect 9364 5012 9370 5024
rect 10045 5015 10103 5021
rect 10045 5012 10057 5015
rect 9364 4984 10057 5012
rect 9364 4972 9370 4984
rect 10045 4981 10057 4984
rect 10091 4981 10103 5015
rect 10045 4975 10103 4981
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 13814 5012 13820 5024
rect 12124 4984 13820 5012
rect 12124 4972 12130 4984
rect 13814 4972 13820 4984
rect 13872 4972 13878 5024
rect 14090 4972 14096 5024
rect 14148 5012 14154 5024
rect 15764 5012 15792 5052
rect 14148 4984 15792 5012
rect 14148 4972 14154 4984
rect 16298 4972 16304 5024
rect 16356 4972 16362 5024
rect 18414 4972 18420 5024
rect 18472 5012 18478 5024
rect 19904 5012 19932 5052
rect 18472 4984 19932 5012
rect 18472 4972 18478 4984
rect 21174 4972 21180 5024
rect 21232 4972 21238 5024
rect 22327 5015 22385 5021
rect 22327 4981 22339 5015
rect 22373 5012 22385 5015
rect 22554 5012 22560 5024
rect 22373 4984 22560 5012
rect 22373 4981 22385 4984
rect 22327 4975 22385 4981
rect 22554 4972 22560 4984
rect 22612 4972 22618 5024
rect 24688 5012 24716 5052
rect 25498 5040 25504 5052
rect 25556 5040 25562 5092
rect 27062 5012 27068 5024
rect 24688 4984 27068 5012
rect 27062 4972 27068 4984
rect 27120 4972 27126 5024
rect 27172 5012 27200 5111
rect 27338 5108 27344 5160
rect 27396 5108 27402 5160
rect 28902 5108 28908 5160
rect 28960 5108 28966 5160
rect 29457 5151 29515 5157
rect 29457 5117 29469 5151
rect 29503 5117 29515 5151
rect 29457 5111 29515 5117
rect 29472 5080 29500 5111
rect 29638 5108 29644 5160
rect 29696 5108 29702 5160
rect 33502 5080 33508 5092
rect 29472 5052 33508 5080
rect 33502 5040 33508 5052
rect 33560 5040 33566 5092
rect 30834 5012 30840 5024
rect 27172 4984 30840 5012
rect 30834 4972 30840 4984
rect 30892 4972 30898 5024
rect 38626 5012 38654 5188
rect 49418 5012 49424 5024
rect 38626 4984 49424 5012
rect 49418 4972 49424 4984
rect 49476 4972 49482 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 2774 4768 2780 4820
rect 2832 4808 2838 4820
rect 3421 4811 3479 4817
rect 3421 4808 3433 4811
rect 2832 4780 3433 4808
rect 2832 4768 2838 4780
rect 3421 4777 3433 4780
rect 3467 4777 3479 4811
rect 3421 4771 3479 4777
rect 4522 4768 4528 4820
rect 4580 4808 4586 4820
rect 4617 4811 4675 4817
rect 4617 4808 4629 4811
rect 4580 4780 4629 4808
rect 4580 4768 4586 4780
rect 4617 4777 4629 4780
rect 4663 4777 4675 4811
rect 4617 4771 4675 4777
rect 5261 4811 5319 4817
rect 5261 4777 5273 4811
rect 5307 4808 5319 4811
rect 5350 4808 5356 4820
rect 5307 4780 5356 4808
rect 5307 4777 5319 4780
rect 5261 4771 5319 4777
rect 5350 4768 5356 4780
rect 5408 4768 5414 4820
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 7282 4808 7288 4820
rect 6595 4780 7288 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 7466 4768 7472 4820
rect 7524 4768 7530 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8573 4811 8631 4817
rect 8573 4808 8585 4811
rect 8260 4780 8585 4808
rect 8260 4768 8266 4780
rect 8573 4777 8585 4780
rect 8619 4777 8631 4811
rect 8573 4771 8631 4777
rect 9950 4768 9956 4820
rect 10008 4768 10014 4820
rect 11422 4808 11428 4820
rect 10704 4780 11428 4808
rect 1578 4700 1584 4752
rect 1636 4740 1642 4752
rect 10229 4743 10287 4749
rect 10229 4740 10241 4743
rect 1636 4712 10241 4740
rect 1636 4700 1642 4712
rect 10229 4709 10241 4712
rect 10275 4709 10287 4743
rect 10229 4703 10287 4709
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4672 1915 4675
rect 1903 4644 3464 4672
rect 1903 4641 1915 4644
rect 1857 4635 1915 4641
rect 1302 4564 1308 4616
rect 1360 4604 1366 4616
rect 1581 4607 1639 4613
rect 1581 4604 1593 4607
rect 1360 4576 1593 4604
rect 1360 4564 1366 4576
rect 1581 4573 1593 4576
rect 1627 4604 1639 4607
rect 1762 4604 1768 4616
rect 1627 4576 1768 4604
rect 1627 4573 1639 4576
rect 1581 4567 1639 4573
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 2958 4564 2964 4616
rect 3016 4564 3022 4616
rect 3142 4564 3148 4616
rect 3200 4564 3206 4616
rect 3436 4536 3464 4644
rect 5718 4632 5724 4684
rect 5776 4672 5782 4684
rect 7190 4672 7196 4684
rect 5776 4644 7196 4672
rect 5776 4632 5782 4644
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 10704 4681 10732 4780
rect 11422 4768 11428 4780
rect 11480 4808 11486 4820
rect 11793 4811 11851 4817
rect 11793 4808 11805 4811
rect 11480 4780 11805 4808
rect 11480 4768 11486 4780
rect 11793 4777 11805 4780
rect 11839 4777 11851 4811
rect 11793 4771 11851 4777
rect 12066 4768 12072 4820
rect 12124 4768 12130 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12406 4780 13093 4808
rect 10870 4700 10876 4752
rect 10928 4740 10934 4752
rect 12406 4740 12434 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 14366 4768 14372 4820
rect 14424 4808 14430 4820
rect 14921 4811 14979 4817
rect 14921 4808 14933 4811
rect 14424 4780 14933 4808
rect 14424 4768 14430 4780
rect 14921 4777 14933 4780
rect 14967 4777 14979 4811
rect 14921 4771 14979 4777
rect 15102 4768 15108 4820
rect 15160 4808 15166 4820
rect 16942 4808 16948 4820
rect 15160 4780 16948 4808
rect 15160 4768 15166 4780
rect 16942 4768 16948 4780
rect 17000 4768 17006 4820
rect 18598 4768 18604 4820
rect 18656 4768 18662 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 18969 4811 19027 4817
rect 18969 4808 18981 4811
rect 18932 4780 18981 4808
rect 18932 4768 18938 4780
rect 18969 4777 18981 4780
rect 19015 4777 19027 4811
rect 18969 4771 19027 4777
rect 20990 4768 20996 4820
rect 21048 4768 21054 4820
rect 22465 4811 22523 4817
rect 22465 4777 22477 4811
rect 22511 4808 22523 4811
rect 22830 4808 22836 4820
rect 22511 4780 22836 4808
rect 22511 4777 22523 4780
rect 22465 4771 22523 4777
rect 22830 4768 22836 4780
rect 22888 4768 22894 4820
rect 23063 4811 23121 4817
rect 23063 4777 23075 4811
rect 23109 4808 23121 4811
rect 27338 4808 27344 4820
rect 23109 4780 27344 4808
rect 23109 4777 23121 4780
rect 23063 4771 23121 4777
rect 27338 4768 27344 4780
rect 27396 4768 27402 4820
rect 31754 4768 31760 4820
rect 31812 4808 31818 4820
rect 41414 4808 41420 4820
rect 31812 4780 41420 4808
rect 31812 4768 31818 4780
rect 41414 4768 41420 4780
rect 41472 4768 41478 4820
rect 10928 4712 12434 4740
rect 10928 4700 10934 4712
rect 16298 4700 16304 4752
rect 16356 4740 16362 4752
rect 23750 4740 23756 4752
rect 16356 4712 23756 4740
rect 16356 4700 16362 4712
rect 23750 4700 23756 4712
rect 23808 4700 23814 4752
rect 24719 4743 24777 4749
rect 24719 4709 24731 4743
rect 24765 4740 24777 4743
rect 29638 4740 29644 4752
rect 24765 4712 29644 4740
rect 24765 4709 24777 4712
rect 24719 4703 24777 4709
rect 29638 4700 29644 4712
rect 29696 4700 29702 4752
rect 29730 4700 29736 4752
rect 29788 4740 29794 4752
rect 34698 4740 34704 4752
rect 29788 4712 34704 4740
rect 29788 4700 29794 4712
rect 34698 4700 34704 4712
rect 34756 4700 34762 4752
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 10689 4635 10747 4641
rect 10962 4632 10968 4684
rect 11020 4632 11026 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11204 4644 14320 4672
rect 11204 4632 11210 4644
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4604 4031 4607
rect 4614 4604 4620 4616
rect 4019 4576 4620 4604
rect 4019 4573 4031 4576
rect 3973 4567 4031 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 5166 4564 5172 4616
rect 5224 4604 5230 4616
rect 6270 4604 6276 4616
rect 5224 4576 6276 4604
rect 5224 4564 5230 4576
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6822 4564 6828 4616
rect 6880 4564 6886 4616
rect 7006 4564 7012 4616
rect 7064 4604 7070 4616
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7064 4576 7941 4604
rect 7064 4564 7070 4576
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 9306 4564 9312 4616
rect 9364 4564 9370 4616
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 12342 4604 12348 4616
rect 9456 4576 12348 4604
rect 9456 4564 9462 4576
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 12437 4607 12495 4613
rect 12437 4573 12449 4607
rect 12483 4573 12495 4607
rect 12437 4567 12495 4573
rect 3436 4508 5396 4536
rect 3510 4428 3516 4480
rect 3568 4468 3574 4480
rect 5258 4468 5264 4480
rect 3568 4440 5264 4468
rect 3568 4428 3574 4440
rect 5258 4428 5264 4440
rect 5316 4428 5322 4480
rect 5368 4468 5396 4508
rect 5902 4496 5908 4548
rect 5960 4496 5966 4548
rect 6086 4496 6092 4548
rect 6144 4496 6150 4548
rect 7558 4496 7564 4548
rect 7616 4536 7622 4548
rect 7616 4508 9674 4536
rect 7616 4496 7622 4508
rect 5994 4468 6000 4480
rect 5368 4440 6000 4468
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 7524 4440 8953 4468
rect 7524 4428 7530 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 9646 4468 9674 4508
rect 12452 4468 12480 4567
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13722 4604 13728 4616
rect 12768 4576 13728 4604
rect 12768 4564 12774 4576
rect 13722 4564 13728 4576
rect 13780 4564 13786 4616
rect 14292 4613 14320 4644
rect 15654 4632 15660 4684
rect 15712 4632 15718 4684
rect 19242 4632 19248 4684
rect 19300 4672 19306 4684
rect 19429 4675 19487 4681
rect 19429 4672 19441 4675
rect 19300 4644 19441 4672
rect 19300 4632 19306 4644
rect 19429 4641 19441 4644
rect 19475 4641 19487 4675
rect 19429 4635 19487 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 20714 4672 20720 4684
rect 19751 4644 20720 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 20714 4632 20720 4644
rect 20772 4632 20778 4684
rect 21910 4632 21916 4684
rect 21968 4632 21974 4684
rect 22554 4632 22560 4684
rect 22612 4672 22618 4684
rect 25869 4675 25927 4681
rect 25869 4672 25881 4675
rect 22612 4644 25881 4672
rect 22612 4632 22618 4644
rect 25869 4641 25881 4644
rect 25915 4641 25927 4675
rect 25869 4635 25927 4641
rect 27062 4632 27068 4684
rect 27120 4632 27126 4684
rect 27154 4632 27160 4684
rect 27212 4672 27218 4684
rect 30742 4672 30748 4684
rect 27212 4644 30748 4672
rect 27212 4632 27218 4644
rect 30742 4632 30748 4644
rect 30800 4632 30806 4684
rect 14277 4607 14335 4613
rect 14277 4573 14289 4607
rect 14323 4573 14335 4607
rect 14277 4567 14335 4573
rect 17052 4576 17632 4604
rect 12618 4496 12624 4548
rect 12676 4536 12682 4548
rect 14458 4536 14464 4548
rect 12676 4508 14464 4536
rect 12676 4496 12682 4508
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 15841 4539 15899 4545
rect 15841 4536 15853 4539
rect 14568 4508 15853 4536
rect 9646 4440 12480 4468
rect 13449 4471 13507 4477
rect 8941 4431 8999 4437
rect 13449 4437 13461 4471
rect 13495 4468 13507 4471
rect 13541 4471 13599 4477
rect 13541 4468 13553 4471
rect 13495 4440 13553 4468
rect 13495 4437 13507 4440
rect 13449 4431 13507 4437
rect 13541 4437 13553 4440
rect 13587 4468 13599 4471
rect 13630 4468 13636 4480
rect 13587 4440 13636 4468
rect 13587 4437 13599 4440
rect 13541 4431 13599 4437
rect 13630 4428 13636 4440
rect 13688 4428 13694 4480
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 14568 4468 14596 4508
rect 15841 4505 15853 4508
rect 15887 4536 15899 4539
rect 17052 4536 17080 4576
rect 15887 4508 17080 4536
rect 15887 4505 15899 4508
rect 15841 4499 15899 4505
rect 17402 4496 17408 4548
rect 17460 4536 17466 4548
rect 17497 4539 17555 4545
rect 17497 4536 17509 4539
rect 17460 4508 17509 4536
rect 17460 4496 17466 4508
rect 17497 4505 17509 4508
rect 17543 4505 17555 4539
rect 17604 4536 17632 4576
rect 17862 4564 17868 4616
rect 17920 4604 17926 4616
rect 17957 4607 18015 4613
rect 17957 4604 17969 4607
rect 17920 4576 17969 4604
rect 17920 4564 17926 4576
rect 17957 4573 17969 4576
rect 18003 4573 18015 4607
rect 17957 4567 18015 4573
rect 20898 4564 20904 4616
rect 20956 4564 20962 4616
rect 22960 4607 23018 4613
rect 22960 4604 22972 4607
rect 22296 4576 22972 4604
rect 22186 4536 22192 4548
rect 17604 4508 22192 4536
rect 17497 4499 17555 4505
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 13780 4440 14596 4468
rect 13780 4428 13786 4440
rect 20346 4428 20352 4480
rect 20404 4468 20410 4480
rect 20533 4471 20591 4477
rect 20533 4468 20545 4471
rect 20404 4440 20545 4468
rect 20404 4428 20410 4440
rect 20533 4437 20545 4440
rect 20579 4437 20591 4471
rect 20533 4431 20591 4437
rect 21358 4428 21364 4480
rect 21416 4468 21422 4480
rect 22296 4468 22324 4576
rect 22960 4573 22972 4576
rect 23006 4573 23018 4607
rect 22960 4567 23018 4573
rect 23474 4564 23480 4616
rect 23532 4604 23538 4616
rect 24616 4607 24674 4613
rect 24616 4604 24628 4607
rect 23532 4576 24628 4604
rect 23532 4564 23538 4576
rect 24616 4573 24628 4576
rect 24662 4573 24674 4607
rect 24616 4567 24674 4573
rect 25685 4607 25743 4613
rect 25685 4573 25697 4607
rect 25731 4573 25743 4607
rect 25685 4567 25743 4573
rect 21416 4440 22324 4468
rect 25700 4468 25728 4567
rect 27798 4468 27804 4480
rect 25700 4440 27804 4468
rect 21416 4428 21422 4440
rect 27798 4428 27804 4440
rect 27856 4428 27862 4480
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 3142 4224 3148 4276
rect 3200 4264 3206 4276
rect 5813 4267 5871 4273
rect 3200 4236 5764 4264
rect 3200 4224 3206 4236
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 5169 4199 5227 4205
rect 2004 4168 4108 4196
rect 2004 4156 2010 4168
rect 1486 4088 1492 4140
rect 1544 4128 1550 4140
rect 1581 4131 1639 4137
rect 1581 4128 1593 4131
rect 1544 4100 1593 4128
rect 1544 4088 1550 4100
rect 1581 4097 1593 4100
rect 1627 4097 1639 4131
rect 1581 4091 1639 4097
rect 1596 3924 1624 4091
rect 2314 4088 2320 4140
rect 2372 4128 2378 4140
rect 2869 4131 2927 4137
rect 2869 4128 2881 4131
rect 2372 4100 2881 4128
rect 2372 4088 2378 4100
rect 2869 4097 2881 4100
rect 2915 4097 2927 4131
rect 2869 4091 2927 4097
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 1857 4063 1915 4069
rect 1857 4029 1869 4063
rect 1903 4060 1915 4063
rect 2774 4060 2780 4072
rect 1903 4032 2780 4060
rect 1903 4029 1915 4032
rect 1857 4023 1915 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 4080 3992 4108 4168
rect 5169 4165 5181 4199
rect 5215 4196 5227 4199
rect 5534 4196 5540 4208
rect 5215 4168 5540 4196
rect 5215 4165 5227 4168
rect 5169 4159 5227 4165
rect 5534 4156 5540 4168
rect 5592 4156 5598 4208
rect 5736 4196 5764 4236
rect 5813 4233 5825 4267
rect 5859 4264 5871 4267
rect 6178 4264 6184 4276
rect 5859 4236 6184 4264
rect 5859 4233 5871 4236
rect 5813 4227 5871 4233
rect 6178 4224 6184 4236
rect 6236 4224 6242 4276
rect 11514 4264 11520 4276
rect 8404 4236 11520 4264
rect 7466 4196 7472 4208
rect 5736 4168 7472 4196
rect 7466 4156 7472 4168
rect 7524 4156 7530 4208
rect 7561 4199 7619 4205
rect 7561 4165 7573 4199
rect 7607 4196 7619 4199
rect 7653 4199 7711 4205
rect 7653 4196 7665 4199
rect 7607 4168 7665 4196
rect 7607 4165 7619 4168
rect 7561 4159 7619 4165
rect 7653 4165 7665 4168
rect 7699 4196 7711 4199
rect 7699 4168 8248 4196
rect 7699 4165 7711 4168
rect 7653 4159 7711 4165
rect 4614 4088 4620 4140
rect 4672 4088 4678 4140
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 5997 4131 6055 4137
rect 5997 4097 6009 4131
rect 6043 4097 6055 4131
rect 5997 4091 6055 4097
rect 6012 4060 6040 4091
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 7190 4088 7196 4140
rect 7248 4088 7254 4140
rect 7650 4060 7656 4072
rect 6012 4032 7656 4060
rect 7650 4020 7656 4032
rect 7708 4020 7714 4072
rect 8220 4060 8248 4168
rect 8404 4137 8432 4236
rect 11514 4224 11520 4236
rect 11572 4224 11578 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 13722 4264 13728 4276
rect 11756 4236 13728 4264
rect 11756 4224 11762 4236
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 14185 4267 14243 4273
rect 14185 4233 14197 4267
rect 14231 4264 14243 4267
rect 17862 4264 17868 4276
rect 14231 4236 17868 4264
rect 14231 4233 14243 4236
rect 14185 4227 14243 4233
rect 17862 4224 17868 4236
rect 17920 4224 17926 4276
rect 19153 4267 19211 4273
rect 19153 4233 19165 4267
rect 19199 4264 19211 4267
rect 19242 4264 19248 4276
rect 19199 4236 19248 4264
rect 19199 4233 19211 4236
rect 19153 4227 19211 4233
rect 19242 4224 19248 4236
rect 19300 4224 19306 4276
rect 20441 4267 20499 4273
rect 20441 4264 20453 4267
rect 19352 4236 20453 4264
rect 9950 4196 9956 4208
rect 8496 4168 9956 4196
rect 8389 4131 8447 4137
rect 8389 4097 8401 4131
rect 8435 4097 8447 4131
rect 8389 4091 8447 4097
rect 8496 4060 8524 4168
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 10965 4199 11023 4205
rect 10965 4165 10977 4199
rect 11011 4196 11023 4199
rect 12345 4199 12403 4205
rect 12345 4196 12357 4199
rect 11011 4168 12357 4196
rect 11011 4165 11023 4168
rect 10965 4159 11023 4165
rect 12345 4165 12357 4168
rect 12391 4165 12403 4199
rect 14090 4196 14096 4208
rect 12345 4159 12403 4165
rect 12452 4168 14096 4196
rect 8846 4088 8852 4140
rect 8904 4088 8910 4140
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9585 4091 9643 4097
rect 8220 4032 8524 4060
rect 9306 4020 9312 4072
rect 9364 4060 9370 4072
rect 9600 4060 9628 4091
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 11422 4128 11428 4140
rect 10100 4100 11428 4128
rect 10100 4088 10106 4100
rect 11422 4088 11428 4100
rect 11480 4088 11486 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4128 11759 4131
rect 12066 4128 12072 4140
rect 11747 4100 12072 4128
rect 11747 4097 11759 4100
rect 11701 4091 11759 4097
rect 12066 4088 12072 4100
rect 12124 4088 12130 4140
rect 12158 4088 12164 4140
rect 12216 4128 12222 4140
rect 12452 4128 12480 4168
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 14274 4156 14280 4208
rect 14332 4196 14338 4208
rect 14332 4168 18276 4196
rect 14332 4156 14338 4168
rect 12216 4100 12480 4128
rect 13081 4131 13139 4137
rect 12216 4088 12222 4100
rect 13081 4097 13093 4131
rect 13127 4128 13139 4131
rect 13354 4128 13360 4140
rect 13127 4100 13360 4128
rect 13127 4097 13139 4100
rect 13081 4091 13139 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13538 4088 13544 4140
rect 13596 4088 13602 4140
rect 14642 4088 14648 4140
rect 14700 4088 14706 4140
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 15286 4128 15292 4140
rect 14792 4100 15292 4128
rect 14792 4088 14798 4100
rect 15286 4088 15292 4100
rect 15344 4088 15350 4140
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16117 4131 16175 4137
rect 16117 4128 16129 4131
rect 15528 4100 16129 4128
rect 15528 4088 15534 4100
rect 16117 4097 16129 4100
rect 16163 4097 16175 4131
rect 18248 4128 18276 4168
rect 19352 4128 19380 4236
rect 20441 4233 20453 4236
rect 20487 4233 20499 4267
rect 20441 4227 20499 4233
rect 21085 4267 21143 4273
rect 21085 4233 21097 4267
rect 21131 4264 21143 4267
rect 25130 4264 25136 4276
rect 21131 4236 25136 4264
rect 21131 4233 21143 4236
rect 21085 4227 21143 4233
rect 25130 4224 25136 4236
rect 25188 4224 25194 4276
rect 22830 4196 22836 4208
rect 21836 4168 22836 4196
rect 18248 4100 19380 4128
rect 19429 4131 19487 4137
rect 16117 4091 16175 4097
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 19475 4100 20576 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 9364 4032 9628 4060
rect 9692 4032 10517 4060
rect 9364 4020 9370 4032
rect 9692 3992 9720 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 11146 4020 11152 4072
rect 11204 4020 11210 4072
rect 11330 4020 11336 4072
rect 11388 4060 11394 4072
rect 16853 4063 16911 4069
rect 16853 4060 16865 4063
rect 11388 4032 16865 4060
rect 11388 4020 11394 4032
rect 16853 4029 16865 4032
rect 16899 4029 16911 4063
rect 16853 4023 16911 4029
rect 17037 4063 17095 4069
rect 17037 4029 17049 4063
rect 17083 4060 17095 4063
rect 17126 4060 17132 4072
rect 17083 4032 17132 4060
rect 17083 4029 17095 4032
rect 17037 4023 17095 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 18693 4063 18751 4069
rect 18693 4029 18705 4063
rect 18739 4060 18751 4063
rect 20070 4060 20076 4072
rect 18739 4032 20076 4060
rect 18739 4029 18751 4032
rect 18693 4023 18751 4029
rect 20070 4020 20076 4032
rect 20128 4020 20134 4072
rect 20548 4060 20576 4100
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 21545 4131 21603 4137
rect 21545 4128 21557 4131
rect 20680 4100 21557 4128
rect 20680 4088 20686 4100
rect 21545 4097 21557 4100
rect 21591 4097 21603 4131
rect 21545 4091 21603 4097
rect 20898 4060 20904 4072
rect 20548 4032 20904 4060
rect 20898 4020 20904 4032
rect 20956 4060 20962 4072
rect 21836 4069 21864 4168
rect 22830 4156 22836 4168
rect 22888 4156 22894 4208
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 20956 4032 21833 4060
rect 20956 4020 20962 4032
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 21821 4023 21879 4029
rect 4080 3964 9720 3992
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 13446 3992 13452 4004
rect 10008 3964 13452 3992
rect 10008 3952 10014 3964
rect 13446 3952 13452 3964
rect 13504 3952 13510 4004
rect 13722 3952 13728 4004
rect 13780 3992 13786 4004
rect 31202 3992 31208 4004
rect 13780 3964 31208 3992
rect 13780 3952 13786 3964
rect 31202 3952 31208 3964
rect 31260 3952 31266 4004
rect 2866 3924 2872 3936
rect 1596 3896 2872 3924
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3510 3884 3516 3936
rect 3568 3884 3574 3936
rect 8481 3927 8539 3933
rect 8481 3893 8493 3927
rect 8527 3924 8539 3927
rect 8754 3924 8760 3936
rect 8527 3896 8760 3924
rect 8527 3893 8539 3896
rect 8481 3887 8539 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 9122 3884 9128 3936
rect 9180 3884 9186 3936
rect 9490 3884 9496 3936
rect 9548 3924 9554 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 9548 3896 10241 3924
rect 9548 3884 9554 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 10229 3887 10287 3893
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 12584 3896 12909 3924
rect 12584 3884 12590 3896
rect 12897 3893 12909 3896
rect 12943 3893 12955 3927
rect 12897 3887 12955 3893
rect 15286 3884 15292 3936
rect 15344 3884 15350 3936
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15657 3927 15715 3933
rect 15657 3924 15669 3927
rect 15528 3896 15669 3924
rect 15528 3884 15534 3896
rect 15657 3893 15669 3896
rect 15703 3893 15715 3927
rect 15657 3887 15715 3893
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16209 3927 16267 3933
rect 16209 3924 16221 3927
rect 16172 3896 16221 3924
rect 16172 3884 16178 3896
rect 16209 3893 16221 3896
rect 16255 3893 16267 3927
rect 16209 3887 16267 3893
rect 19518 3884 19524 3936
rect 19576 3884 19582 3936
rect 19886 3884 19892 3936
rect 19944 3884 19950 3936
rect 21634 3884 21640 3936
rect 21692 3924 21698 3936
rect 23474 3924 23480 3936
rect 21692 3896 23480 3924
rect 21692 3884 21698 3896
rect 23474 3884 23480 3896
rect 23532 3884 23538 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 2314 3680 2320 3732
rect 2372 3680 2378 3732
rect 3970 3680 3976 3732
rect 4028 3720 4034 3732
rect 5261 3723 5319 3729
rect 5261 3720 5273 3723
rect 4028 3692 5273 3720
rect 4028 3680 4034 3692
rect 5261 3689 5273 3692
rect 5307 3689 5319 3723
rect 8662 3720 8668 3732
rect 5261 3683 5319 3689
rect 5368 3692 8668 3720
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 5368 3652 5396 3692
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9033 3723 9091 3729
rect 9033 3689 9045 3723
rect 9079 3720 9091 3723
rect 9674 3720 9680 3732
rect 9079 3692 9680 3720
rect 9079 3689 9091 3692
rect 9033 3683 9091 3689
rect 9674 3680 9680 3692
rect 9732 3680 9738 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 12158 3720 12164 3732
rect 11287 3692 12164 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 12158 3680 12164 3692
rect 12216 3680 12222 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13538 3720 13544 3732
rect 13035 3692 13544 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 18506 3720 18512 3732
rect 14476 3692 18512 3720
rect 2832 3624 5396 3652
rect 7009 3655 7067 3661
rect 2832 3612 2838 3624
rect 7009 3621 7021 3655
rect 7055 3652 7067 3655
rect 11330 3652 11336 3664
rect 7055 3624 11336 3652
rect 7055 3621 7067 3624
rect 7009 3615 7067 3621
rect 11330 3612 11336 3624
rect 11388 3612 11394 3664
rect 11701 3655 11759 3661
rect 11701 3621 11713 3655
rect 11747 3652 11759 3655
rect 14476 3652 14504 3692
rect 18506 3680 18512 3692
rect 18564 3680 18570 3732
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 21634 3720 21640 3732
rect 19944 3692 21640 3720
rect 19944 3680 19950 3692
rect 21634 3680 21640 3692
rect 21692 3680 21698 3732
rect 11747 3624 14504 3652
rect 11747 3621 11759 3624
rect 11701 3615 11759 3621
rect 14550 3612 14556 3664
rect 14608 3612 14614 3664
rect 15289 3655 15347 3661
rect 15289 3621 15301 3655
rect 15335 3652 15347 3655
rect 15378 3652 15384 3664
rect 15335 3624 15384 3652
rect 15335 3621 15347 3624
rect 15289 3615 15347 3621
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 15746 3612 15752 3664
rect 15804 3612 15810 3664
rect 15930 3612 15936 3664
rect 15988 3612 15994 3664
rect 17126 3612 17132 3664
rect 17184 3652 17190 3664
rect 21358 3652 21364 3664
rect 17184 3624 21364 3652
rect 17184 3612 17190 3624
rect 21358 3612 21364 3624
rect 21416 3612 21422 3664
rect 22094 3612 22100 3664
rect 22152 3652 22158 3664
rect 28718 3652 28724 3664
rect 22152 3624 28724 3652
rect 22152 3612 22158 3624
rect 28718 3612 28724 3624
rect 28776 3612 28782 3664
rect 842 3544 848 3596
rect 900 3584 906 3596
rect 3973 3587 4031 3593
rect 3973 3584 3985 3587
rect 900 3556 3985 3584
rect 900 3544 906 3556
rect 3973 3553 3985 3556
rect 4019 3553 4031 3587
rect 3973 3547 4031 3553
rect 5721 3587 5779 3593
rect 5721 3553 5733 3587
rect 5767 3584 5779 3587
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 5767 3556 9137 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 9125 3553 9137 3556
rect 9171 3584 9183 3587
rect 9398 3584 9404 3596
rect 9171 3556 9404 3584
rect 9171 3553 9183 3556
rect 9125 3547 9183 3553
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 19518 3584 19524 3596
rect 9824 3556 12112 3584
rect 9824 3544 9830 3556
rect 1670 3476 1676 3528
rect 1728 3476 1734 3528
rect 2774 3476 2780 3528
rect 2832 3476 2838 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3485 4675 3519
rect 4617 3479 4675 3485
rect 1394 3408 1400 3460
rect 1452 3448 1458 3460
rect 4632 3448 4660 3479
rect 5994 3476 6000 3528
rect 6052 3476 6058 3528
rect 6914 3476 6920 3528
rect 6972 3516 6978 3528
rect 7193 3519 7251 3525
rect 7193 3516 7205 3519
rect 6972 3488 7205 3516
rect 6972 3476 6978 3488
rect 7193 3485 7205 3488
rect 7239 3485 7251 3519
rect 7193 3479 7251 3485
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 8435 3488 9444 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 8294 3448 8300 3460
rect 1452 3420 8300 3448
rect 1452 3408 1458 3420
rect 8294 3408 8300 3420
rect 8352 3408 8358 3460
rect 8570 3408 8576 3460
rect 8628 3408 8634 3460
rect 9416 3448 9444 3488
rect 9490 3476 9496 3528
rect 9548 3476 9554 3528
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10597 3519 10655 3525
rect 10597 3516 10609 3519
rect 10183 3488 10609 3516
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 10597 3485 10609 3488
rect 10643 3485 10655 3519
rect 10597 3479 10655 3485
rect 11882 3476 11888 3528
rect 11940 3476 11946 3528
rect 9674 3448 9680 3460
rect 9416 3420 9680 3448
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 11974 3448 11980 3460
rect 9968 3420 11980 3448
rect 3421 3383 3479 3389
rect 3421 3349 3433 3383
rect 3467 3380 3479 3383
rect 3878 3380 3884 3392
rect 3467 3352 3884 3380
rect 3467 3349 3479 3352
rect 3421 3343 3479 3349
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 4062 3340 4068 3392
rect 4120 3380 4126 3392
rect 5810 3380 5816 3392
rect 4120 3352 5816 3380
rect 4120 3340 4126 3352
rect 5810 3340 5816 3352
rect 5868 3340 5874 3392
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 9968 3380 9996 3420
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 12084 3448 12112 3556
rect 12360 3556 19524 3584
rect 12360 3528 12388 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 20717 3587 20775 3593
rect 20717 3553 20729 3587
rect 20763 3584 20775 3587
rect 21082 3584 21088 3596
rect 20763 3556 21088 3584
rect 20763 3553 20775 3556
rect 20717 3547 20775 3553
rect 21082 3544 21088 3556
rect 21140 3544 21146 3596
rect 12342 3476 12348 3528
rect 12400 3476 12406 3528
rect 14642 3516 14648 3528
rect 12820 3488 14648 3516
rect 12820 3448 12848 3488
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 15028 3488 15700 3516
rect 13541 3451 13599 3457
rect 13541 3448 13553 3451
rect 12084 3420 12848 3448
rect 12912 3420 13553 3448
rect 7699 3352 9996 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 10502 3340 10508 3392
rect 10560 3380 10566 3392
rect 12912 3380 12940 3420
rect 13541 3417 13553 3420
rect 13587 3417 13599 3451
rect 13541 3411 13599 3417
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3448 14427 3451
rect 15028 3448 15056 3488
rect 14415 3420 15056 3448
rect 14415 3417 14427 3420
rect 14369 3411 14427 3417
rect 15102 3408 15108 3460
rect 15160 3408 15166 3460
rect 15672 3457 15700 3488
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 16301 3519 16359 3525
rect 16301 3516 16313 3519
rect 15804 3488 16313 3516
rect 15804 3476 15810 3488
rect 16301 3485 16313 3488
rect 16347 3485 16359 3519
rect 16301 3479 16359 3485
rect 16577 3519 16635 3525
rect 16577 3485 16589 3519
rect 16623 3516 16635 3519
rect 17034 3516 17040 3528
rect 16623 3488 17040 3516
rect 16623 3485 16635 3488
rect 16577 3479 16635 3485
rect 17034 3476 17040 3488
rect 17092 3476 17098 3528
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 17736 3488 17877 3516
rect 17736 3476 17742 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 19613 3519 19671 3525
rect 19613 3516 19625 3519
rect 17865 3479 17923 3485
rect 18800 3488 19625 3516
rect 15657 3451 15715 3457
rect 15657 3417 15669 3451
rect 15703 3448 15715 3451
rect 18414 3448 18420 3460
rect 15703 3420 18420 3448
rect 15703 3417 15715 3420
rect 15657 3411 15715 3417
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 10560 3352 12940 3380
rect 10560 3340 10566 3352
rect 17218 3340 17224 3392
rect 17276 3380 17282 3392
rect 17678 3380 17684 3392
rect 17276 3352 17684 3380
rect 17276 3340 17282 3352
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 18690 3340 18696 3392
rect 18748 3380 18754 3392
rect 18800 3389 18828 3488
rect 19613 3485 19625 3488
rect 19659 3485 19671 3519
rect 19613 3479 19671 3485
rect 20257 3519 20315 3525
rect 20257 3485 20269 3519
rect 20303 3485 20315 3519
rect 20257 3479 20315 3485
rect 18874 3408 18880 3460
rect 18932 3448 18938 3460
rect 19061 3451 19119 3457
rect 19061 3448 19073 3451
rect 18932 3420 19073 3448
rect 18932 3408 18938 3420
rect 19061 3417 19073 3420
rect 19107 3448 19119 3451
rect 20272 3448 20300 3479
rect 28902 3476 28908 3528
rect 28960 3516 28966 3528
rect 44082 3516 44088 3528
rect 28960 3488 44088 3516
rect 28960 3476 28966 3488
rect 44082 3476 44088 3488
rect 44140 3476 44146 3528
rect 19107 3420 20300 3448
rect 19107 3417 19119 3420
rect 19061 3411 19119 3417
rect 27062 3408 27068 3460
rect 27120 3448 27126 3460
rect 46750 3448 46756 3460
rect 27120 3420 46756 3448
rect 27120 3408 27126 3420
rect 46750 3408 46756 3420
rect 46808 3408 46814 3460
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18748 3352 18797 3380
rect 18748 3340 18754 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 19334 3340 19340 3392
rect 19392 3380 19398 3392
rect 19429 3383 19487 3389
rect 19429 3380 19441 3383
rect 19392 3352 19441 3380
rect 19392 3340 19398 3352
rect 19429 3349 19441 3352
rect 19475 3349 19487 3383
rect 19429 3343 19487 3349
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19852 3352 20085 3380
rect 19852 3340 19858 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 2869 3179 2927 3185
rect 2869 3145 2881 3179
rect 2915 3176 2927 3179
rect 10597 3179 10655 3185
rect 2915 3148 10456 3176
rect 2915 3145 2927 3148
rect 2869 3139 2927 3145
rect 5813 3111 5871 3117
rect 5813 3077 5825 3111
rect 5859 3108 5871 3111
rect 9214 3108 9220 3120
rect 5859 3080 9220 3108
rect 5859 3077 5871 3080
rect 5813 3071 5871 3077
rect 9214 3068 9220 3080
rect 9272 3068 9278 3120
rect 10428 3108 10456 3148
rect 10597 3145 10609 3179
rect 10643 3176 10655 3179
rect 12066 3176 12072 3188
rect 10643 3148 12072 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 15102 3176 15108 3188
rect 12268 3148 15108 3176
rect 12268 3108 12296 3148
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 17586 3136 17592 3188
rect 17644 3176 17650 3188
rect 17862 3176 17868 3188
rect 17644 3148 17868 3176
rect 17644 3136 17650 3148
rect 17862 3136 17868 3148
rect 17920 3176 17926 3188
rect 18049 3179 18107 3185
rect 18049 3176 18061 3179
rect 17920 3148 18061 3176
rect 17920 3136 17926 3148
rect 18049 3145 18061 3148
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 20806 3136 20812 3188
rect 20864 3136 20870 3188
rect 10428 3080 12296 3108
rect 12406 3080 13584 3108
rect 3050 3000 3056 3052
rect 3108 3000 3114 3052
rect 3510 3000 3516 3052
rect 3568 3000 3574 3052
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 4617 3043 4675 3049
rect 4617 3040 4629 3043
rect 3936 3012 4629 3040
rect 3936 3000 3942 3012
rect 4617 3009 4629 3012
rect 4663 3009 4675 3043
rect 4617 3003 4675 3009
rect 5261 3043 5319 3049
rect 5261 3009 5273 3043
rect 5307 3040 5319 3043
rect 6549 3043 6607 3049
rect 6549 3040 6561 3043
rect 5307 3012 6561 3040
rect 5307 3009 5319 3012
rect 5261 3003 5319 3009
rect 6549 3009 6561 3012
rect 6595 3009 6607 3043
rect 6549 3003 6607 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3040 7251 3043
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7239 3012 7757 3040
rect 7239 3009 7251 3012
rect 7193 3003 7251 3009
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 7745 3003 7803 3009
rect 8478 3000 8484 3052
rect 8536 3040 8542 3052
rect 8849 3043 8907 3049
rect 8849 3040 8861 3043
rect 8536 3012 8861 3040
rect 8536 3000 8542 3012
rect 8849 3009 8861 3012
rect 8895 3009 8907 3043
rect 10594 3040 10600 3052
rect 10258 3012 10600 3040
rect 8849 3003 8907 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10870 3000 10876 3052
rect 10928 3000 10934 3052
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11793 3043 11851 3049
rect 11793 3040 11805 3043
rect 11379 3012 11805 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11793 3009 11805 3012
rect 11839 3040 11851 3043
rect 12158 3040 12164 3052
rect 11839 3012 12164 3040
rect 11839 3009 11851 3012
rect 11793 3003 11851 3009
rect 12158 3000 12164 3012
rect 12216 3000 12222 3052
rect 1578 2932 1584 2984
rect 1636 2932 1642 2984
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 8389 2975 8447 2981
rect 1903 2944 8340 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 3326 2864 3332 2916
rect 3384 2904 3390 2916
rect 3878 2904 3884 2916
rect 3384 2876 3884 2904
rect 3384 2864 3390 2876
rect 3878 2864 3884 2876
rect 3936 2864 3942 2916
rect 4062 2864 4068 2916
rect 4120 2904 4126 2916
rect 8312 2904 8340 2944
rect 8389 2941 8401 2975
rect 8435 2972 8447 2975
rect 9125 2975 9183 2981
rect 9125 2972 9137 2975
rect 8435 2944 9137 2972
rect 8435 2941 8447 2944
rect 8389 2935 8447 2941
rect 9125 2941 9137 2944
rect 9171 2941 9183 2975
rect 9125 2935 9183 2941
rect 9858 2932 9864 2984
rect 9916 2972 9922 2984
rect 12406 2972 12434 3080
rect 13556 3052 13584 3080
rect 14826 3068 14832 3120
rect 14884 3068 14890 3120
rect 15010 3068 15016 3120
rect 15068 3068 15074 3120
rect 15841 3111 15899 3117
rect 15841 3077 15853 3111
rect 15887 3108 15899 3111
rect 18693 3111 18751 3117
rect 18693 3108 18705 3111
rect 15887 3080 18705 3108
rect 15887 3077 15899 3080
rect 15841 3071 15899 3077
rect 18693 3077 18705 3080
rect 18739 3108 18751 3111
rect 19886 3108 19892 3120
rect 18739 3080 19892 3108
rect 18739 3077 18751 3080
rect 18693 3071 18751 3077
rect 19886 3068 19892 3080
rect 19944 3068 19950 3120
rect 20349 3111 20407 3117
rect 20349 3077 20361 3111
rect 20395 3108 20407 3111
rect 22738 3108 22744 3120
rect 20395 3080 22744 3108
rect 20395 3077 20407 3080
rect 20349 3071 20407 3077
rect 22738 3068 22744 3080
rect 22796 3068 22802 3120
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 12710 3040 12716 3052
rect 12575 3012 12716 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 13078 3000 13084 3052
rect 13136 3000 13142 3052
rect 13538 3000 13544 3052
rect 13596 3000 13602 3052
rect 14093 3043 14151 3049
rect 14093 3009 14105 3043
rect 14139 3040 14151 3043
rect 17126 3040 17132 3052
rect 14139 3012 17132 3040
rect 14139 3009 14151 3012
rect 14093 3003 14151 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 18414 3040 18420 3052
rect 17267 3012 18420 3040
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 18414 3000 18420 3012
rect 18472 3000 18478 3052
rect 18506 3000 18512 3052
rect 18564 3000 18570 3052
rect 22186 3000 22192 3052
rect 22244 3040 22250 3052
rect 22465 3043 22523 3049
rect 22465 3040 22477 3043
rect 22244 3012 22477 3040
rect 22244 3000 22250 3012
rect 22465 3009 22477 3012
rect 22511 3009 22523 3043
rect 22465 3003 22523 3009
rect 9916 2944 12434 2972
rect 9916 2932 9922 2944
rect 15930 2932 15936 2984
rect 15988 2972 15994 2984
rect 16945 2975 17003 2981
rect 16945 2972 16957 2975
rect 15988 2944 16957 2972
rect 15988 2932 15994 2944
rect 16945 2941 16957 2944
rect 16991 2941 17003 2975
rect 16945 2935 17003 2941
rect 8846 2904 8852 2916
rect 4120 2876 4292 2904
rect 8312 2876 8852 2904
rect 4120 2864 4126 2876
rect 4154 2796 4160 2848
rect 4212 2796 4218 2848
rect 4264 2836 4292 2876
rect 8846 2864 8852 2876
rect 8904 2864 8910 2916
rect 16390 2904 16396 2916
rect 10152 2876 16396 2904
rect 10152 2836 10180 2876
rect 16390 2864 16396 2876
rect 16448 2864 16454 2916
rect 4264 2808 10180 2836
rect 11882 2796 11888 2848
rect 11940 2796 11946 2848
rect 12618 2796 12624 2848
rect 12676 2796 12682 2848
rect 13354 2796 13360 2848
rect 13412 2796 13418 2848
rect 14182 2796 14188 2848
rect 14240 2796 14246 2848
rect 15378 2796 15384 2848
rect 15436 2796 15442 2848
rect 15930 2796 15936 2848
rect 15988 2796 15994 2848
rect 20806 2796 20812 2848
rect 20864 2836 20870 2848
rect 22005 2839 22063 2845
rect 22005 2836 22017 2839
rect 20864 2808 22017 2836
rect 20864 2796 20870 2808
rect 22005 2805 22017 2808
rect 22051 2805 22063 2839
rect 22005 2799 22063 2805
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 2038 2592 2044 2644
rect 2096 2632 2102 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2096 2604 2881 2632
rect 2096 2592 2102 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 5534 2592 5540 2644
rect 5592 2632 5598 2644
rect 6365 2635 6423 2641
rect 6365 2632 6377 2635
rect 5592 2604 6377 2632
rect 5592 2592 5598 2604
rect 6365 2601 6377 2604
rect 6411 2601 6423 2635
rect 6365 2595 6423 2601
rect 8294 2592 8300 2644
rect 8352 2632 8358 2644
rect 9125 2635 9183 2641
rect 9125 2632 9137 2635
rect 8352 2604 9137 2632
rect 8352 2592 8358 2604
rect 9125 2601 9137 2604
rect 9171 2601 9183 2635
rect 9125 2595 9183 2601
rect 13538 2592 13544 2644
rect 13596 2632 13602 2644
rect 13817 2635 13875 2641
rect 13817 2632 13829 2635
rect 13596 2604 13829 2632
rect 13596 2592 13602 2604
rect 13817 2601 13829 2604
rect 13863 2601 13875 2635
rect 13817 2595 13875 2601
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14921 2635 14979 2641
rect 14921 2632 14933 2635
rect 14056 2604 14933 2632
rect 14056 2592 14062 2604
rect 14921 2601 14933 2604
rect 14967 2601 14979 2635
rect 14921 2595 14979 2601
rect 15194 2592 15200 2644
rect 15252 2632 15258 2644
rect 15930 2632 15936 2644
rect 15252 2604 15936 2632
rect 15252 2592 15258 2604
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 16942 2592 16948 2644
rect 17000 2592 17006 2644
rect 17586 2592 17592 2644
rect 17644 2592 17650 2644
rect 17678 2592 17684 2644
rect 17736 2632 17742 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 17736 2604 20085 2632
rect 17736 2592 17742 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 22002 2592 22008 2644
rect 22060 2592 22066 2644
rect 22554 2592 22560 2644
rect 22612 2632 22618 2644
rect 23382 2632 23388 2644
rect 22612 2604 23388 2632
rect 22612 2592 22618 2604
rect 23382 2592 23388 2604
rect 23440 2592 23446 2644
rect 25498 2592 25504 2644
rect 25556 2592 25562 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 27856 2604 28181 2632
rect 27856 2592 27862 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 30834 2592 30840 2644
rect 30892 2592 30898 2644
rect 33502 2592 33508 2644
rect 33560 2592 33566 2644
rect 1118 2524 1124 2576
rect 1176 2564 1182 2576
rect 3789 2567 3847 2573
rect 3789 2564 3801 2567
rect 1176 2536 3801 2564
rect 1176 2524 1182 2536
rect 3789 2533 3801 2536
rect 3835 2533 3847 2567
rect 8665 2567 8723 2573
rect 8665 2564 8677 2567
rect 3789 2527 3847 2533
rect 3896 2536 8677 2564
rect 658 2456 664 2508
rect 716 2496 722 2508
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 716 2468 1869 2496
rect 716 2456 722 2468
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 3237 2499 3295 2505
rect 3237 2465 3249 2499
rect 3283 2496 3295 2499
rect 3326 2496 3332 2508
rect 3283 2468 3332 2496
rect 3283 2465 3295 2468
rect 3237 2459 3295 2465
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 1360 2400 1593 2428
rect 1360 2388 1366 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 1596 2360 1624 2391
rect 1762 2388 1768 2440
rect 1820 2428 1826 2440
rect 3896 2428 3924 2536
rect 8665 2533 8677 2536
rect 8711 2533 8723 2567
rect 14182 2564 14188 2576
rect 8665 2527 8723 2533
rect 11808 2536 14188 2564
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4120 2468 4629 2496
rect 4120 2456 4126 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 4617 2459 4675 2465
rect 5810 2456 5816 2508
rect 5868 2456 5874 2508
rect 6089 2499 6147 2505
rect 6089 2465 6101 2499
rect 6135 2496 6147 2499
rect 6178 2496 6184 2508
rect 6135 2468 6184 2496
rect 6135 2465 6147 2468
rect 6089 2459 6147 2465
rect 6178 2456 6184 2468
rect 6236 2456 6242 2508
rect 6730 2456 6736 2508
rect 6788 2496 6794 2508
rect 7285 2499 7343 2505
rect 7285 2496 7297 2499
rect 6788 2468 7297 2496
rect 6788 2456 6794 2468
rect 7285 2465 7297 2468
rect 7331 2465 7343 2499
rect 7285 2459 7343 2465
rect 9398 2456 9404 2508
rect 9456 2496 9462 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9456 2468 9965 2496
rect 9456 2456 9462 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 9953 2459 10011 2465
rect 1820 2400 3924 2428
rect 1820 2388 1826 2400
rect 4338 2388 4344 2440
rect 4396 2388 4402 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2397 7067 2431
rect 7009 2391 7067 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2428 9643 2431
rect 11808 2428 11836 2536
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 18233 2567 18291 2573
rect 18233 2564 18245 2567
rect 15068 2536 18245 2564
rect 15068 2524 15074 2536
rect 18233 2533 18245 2536
rect 18279 2533 18291 2567
rect 18233 2527 18291 2533
rect 18414 2524 18420 2576
rect 18472 2564 18478 2576
rect 18472 2536 19334 2564
rect 18472 2524 18478 2536
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12124 2468 12633 2496
rect 12124 2456 12130 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 14642 2456 14648 2508
rect 14700 2496 14706 2508
rect 14700 2468 16344 2496
rect 14700 2456 14706 2468
rect 9631 2400 11836 2428
rect 12345 2431 12403 2437
rect 9631 2397 9643 2400
rect 9585 2391 9643 2397
rect 12345 2397 12357 2431
rect 12391 2428 12403 2431
rect 15194 2428 15200 2440
rect 12391 2400 15200 2428
rect 12391 2397 12403 2400
rect 12345 2391 12403 2397
rect 7024 2360 7052 2391
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 12618 2360 12624 2372
rect 1596 2332 6914 2360
rect 7024 2332 12624 2360
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 4890 2292 4896 2304
rect 2823 2264 4896 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 4890 2252 4896 2264
rect 4948 2252 4954 2304
rect 6886 2292 6914 2332
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 14829 2363 14887 2369
rect 14829 2360 14841 2363
rect 14200 2332 14841 2360
rect 14200 2304 14228 2332
rect 14829 2329 14841 2332
rect 14875 2329 14887 2363
rect 14829 2323 14887 2329
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 6886 2264 8493 2292
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8481 2255 8539 2261
rect 9030 2252 9036 2304
rect 9088 2252 9094 2304
rect 11146 2252 11152 2304
rect 11204 2252 11210 2304
rect 11514 2252 11520 2304
rect 11572 2252 11578 2304
rect 14182 2252 14188 2304
rect 14240 2252 14246 2304
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 15488 2292 15516 2391
rect 15746 2388 15752 2440
rect 15804 2388 15810 2440
rect 16316 2360 16344 2468
rect 16390 2456 16396 2508
rect 16448 2496 16454 2508
rect 19306 2496 19334 2536
rect 19426 2524 19432 2576
rect 19484 2524 19490 2576
rect 32398 2564 32404 2576
rect 28966 2536 32404 2564
rect 28966 2496 28994 2536
rect 32398 2524 32404 2536
rect 32456 2524 32462 2576
rect 16448 2468 18460 2496
rect 19306 2468 28994 2496
rect 16448 2456 16454 2468
rect 16482 2388 16488 2440
rect 16540 2428 16546 2440
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 16540 2400 17141 2428
rect 16540 2388 16546 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 18432 2437 18460 2468
rect 36354 2456 36360 2508
rect 36412 2456 36418 2508
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2397 18475 2431
rect 19426 2428 19432 2440
rect 18417 2391 18475 2397
rect 18800 2400 19432 2428
rect 18800 2360 18828 2400
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 22189 2431 22247 2437
rect 22189 2397 22201 2431
rect 22235 2428 22247 2431
rect 22554 2428 22560 2440
rect 22235 2400 22560 2428
rect 22235 2397 22247 2400
rect 22189 2391 22247 2397
rect 20272 2360 20300 2391
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 25406 2388 25412 2440
rect 25464 2428 25470 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25464 2400 25697 2428
rect 25464 2388 25470 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 25961 2431 26019 2437
rect 25961 2428 25973 2431
rect 25731 2400 25973 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 25961 2397 25973 2400
rect 26007 2397 26019 2431
rect 25961 2391 26019 2397
rect 28350 2388 28356 2440
rect 28408 2428 28414 2440
rect 28629 2431 28687 2437
rect 28629 2428 28641 2431
rect 28408 2400 28641 2428
rect 28408 2388 28414 2400
rect 28629 2397 28641 2400
rect 28675 2397 28687 2431
rect 28629 2391 28687 2397
rect 30742 2388 30748 2440
rect 30800 2428 30806 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30800 2400 31033 2428
rect 30800 2388 30806 2400
rect 31021 2397 31033 2400
rect 31067 2428 31079 2431
rect 31297 2431 31355 2437
rect 31297 2428 31309 2431
rect 31067 2400 31309 2428
rect 31067 2397 31079 2400
rect 31021 2391 31079 2397
rect 31297 2397 31309 2400
rect 31343 2397 31355 2431
rect 31297 2391 31355 2397
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 33689 2431 33747 2437
rect 33689 2428 33701 2431
rect 33468 2400 33701 2428
rect 33468 2388 33474 2400
rect 33689 2397 33701 2400
rect 33735 2428 33747 2431
rect 33965 2431 34023 2437
rect 33965 2428 33977 2431
rect 33735 2400 33977 2428
rect 33735 2397 33747 2400
rect 33689 2391 33747 2397
rect 33965 2397 33977 2400
rect 34011 2397 34023 2431
rect 33965 2391 34023 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 37277 2431 37335 2437
rect 37277 2428 37289 2431
rect 36136 2400 37289 2428
rect 36136 2388 36142 2400
rect 37277 2397 37289 2400
rect 37323 2397 37335 2431
rect 37277 2391 37335 2397
rect 16316 2332 18828 2360
rect 19306 2332 20300 2360
rect 14424 2264 15516 2292
rect 14424 2252 14430 2264
rect 18782 2252 18788 2304
rect 18840 2252 18846 2304
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 19306 2292 19334 2332
rect 20714 2320 20720 2372
rect 20772 2320 20778 2372
rect 20898 2320 20904 2372
rect 20956 2360 20962 2372
rect 28718 2360 28724 2372
rect 20956 2332 28724 2360
rect 20956 2320 20962 2332
rect 28718 2320 28724 2332
rect 28776 2320 28782 2372
rect 19024 2264 19334 2292
rect 19024 2252 19030 2264
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 11514 2088 11520 2100
rect 2924 2060 11520 2088
rect 2924 2048 2930 2060
rect 11514 2048 11520 2060
rect 11572 2048 11578 2100
rect 15194 2088 15200 2100
rect 11624 2060 15200 2088
rect 9030 1980 9036 2032
rect 9088 2020 9094 2032
rect 11624 2020 11652 2060
rect 15194 2048 15200 2060
rect 15252 2048 15258 2100
rect 18782 2048 18788 2100
rect 18840 2088 18846 2100
rect 19610 2088 19616 2100
rect 18840 2060 19616 2088
rect 18840 2048 18846 2060
rect 19610 2048 19616 2060
rect 19668 2048 19674 2100
rect 9088 1992 11652 2020
rect 9088 1980 9094 1992
rect 11698 1980 11704 2032
rect 11756 2020 11762 2032
rect 22094 2020 22100 2032
rect 11756 1992 22100 2020
rect 11756 1980 11762 1992
rect 22094 1980 22100 1992
rect 22152 1980 22158 2032
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 17770 1952 17776 1964
rect 4212 1924 17776 1952
rect 4212 1912 4218 1924
rect 17770 1912 17776 1924
rect 17828 1912 17834 1964
rect 3418 1844 3424 1896
rect 3476 1884 3482 1896
rect 15378 1884 15384 1896
rect 3476 1856 15384 1884
rect 3476 1844 3482 1856
rect 15378 1844 15384 1856
rect 15436 1884 15442 1896
rect 16482 1884 16488 1896
rect 15436 1856 16488 1884
rect 15436 1844 15442 1856
rect 16482 1844 16488 1856
rect 16540 1844 16546 1896
rect 17494 1844 17500 1896
rect 17552 1884 17558 1896
rect 20898 1884 20904 1896
rect 17552 1856 20904 1884
rect 17552 1844 17558 1856
rect 20898 1844 20904 1856
rect 20956 1844 20962 1896
rect 3602 1776 3608 1828
rect 3660 1816 3666 1828
rect 3660 1788 12434 1816
rect 3660 1776 3666 1788
rect 11882 1748 11888 1760
rect 6886 1720 11888 1748
rect 4338 1640 4344 1692
rect 4396 1680 4402 1692
rect 6886 1680 6914 1720
rect 11882 1708 11888 1720
rect 11940 1708 11946 1760
rect 12406 1748 12434 1788
rect 18966 1748 18972 1760
rect 12406 1720 18972 1748
rect 18966 1708 18972 1720
rect 19024 1708 19030 1760
rect 4396 1652 6914 1680
rect 4396 1640 4402 1652
rect 10962 1640 10968 1692
rect 11020 1680 11026 1692
rect 20714 1680 20720 1692
rect 11020 1652 20720 1680
rect 11020 1640 11026 1652
rect 20714 1640 20720 1652
rect 20772 1640 20778 1692
rect 1578 1572 1584 1624
rect 1636 1612 1642 1624
rect 11146 1612 11152 1624
rect 1636 1584 11152 1612
rect 1636 1572 1642 1584
rect 11146 1572 11152 1584
rect 11204 1572 11210 1624
rect 3326 1504 3332 1556
rect 3384 1544 3390 1556
rect 14366 1544 14372 1556
rect 3384 1516 14372 1544
rect 3384 1504 3390 1516
rect 14366 1504 14372 1516
rect 14424 1504 14430 1556
rect 10318 1436 10324 1488
rect 10376 1476 10382 1488
rect 19334 1476 19340 1488
rect 10376 1448 19340 1476
rect 10376 1436 10382 1448
rect 19334 1436 19340 1448
rect 19392 1436 19398 1488
rect 11054 1408 11060 1420
rect 9600 1380 11060 1408
rect 566 1300 572 1352
rect 624 1340 630 1352
rect 9600 1340 9628 1380
rect 11054 1368 11060 1380
rect 11112 1368 11118 1420
rect 16482 1368 16488 1420
rect 16540 1408 16546 1420
rect 16540 1380 18000 1408
rect 16540 1368 16546 1380
rect 624 1312 9628 1340
rect 624 1300 630 1312
rect 11330 1300 11336 1352
rect 11388 1340 11394 1352
rect 17972 1340 18000 1380
rect 22186 1340 22192 1352
rect 11388 1312 12434 1340
rect 17972 1312 22192 1340
rect 11388 1300 11394 1312
rect 5626 1232 5632 1284
rect 5684 1272 5690 1284
rect 11698 1272 11704 1284
rect 5684 1244 11704 1272
rect 5684 1232 5690 1244
rect 11698 1232 11704 1244
rect 11756 1232 11762 1284
rect 12406 1272 12434 1312
rect 22186 1300 22192 1312
rect 22244 1300 22250 1352
rect 25314 1272 25320 1284
rect 12406 1244 25320 1272
rect 25314 1232 25320 1244
rect 25372 1232 25378 1284
rect 13630 1164 13636 1216
rect 13688 1204 13694 1216
rect 21450 1204 21456 1216
rect 13688 1176 21456 1204
rect 13688 1164 13694 1176
rect 21450 1164 21456 1176
rect 21508 1164 21514 1216
rect 22094 1164 22100 1216
rect 22152 1204 22158 1216
rect 22462 1204 22468 1216
rect 22152 1176 22468 1204
rect 22152 1164 22158 1176
rect 22462 1164 22468 1176
rect 22520 1204 22526 1216
rect 35434 1204 35440 1216
rect 22520 1176 35440 1204
rect 22520 1164 22526 1176
rect 35434 1164 35440 1176
rect 35492 1164 35498 1216
rect 15746 1096 15752 1148
rect 15804 1136 15810 1148
rect 25958 1136 25964 1148
rect 15804 1108 25964 1136
rect 15804 1096 15810 1108
rect 25958 1096 25964 1108
rect 26016 1096 26022 1148
rect 3694 1028 3700 1080
rect 3752 1068 3758 1080
rect 18690 1068 18696 1080
rect 3752 1040 18696 1068
rect 3752 1028 3758 1040
rect 18690 1028 18696 1040
rect 18748 1028 18754 1080
rect 4798 960 4804 1012
rect 4856 1000 4862 1012
rect 20346 1000 20352 1012
rect 4856 972 20352 1000
rect 4856 960 4862 972
rect 20346 960 20352 972
rect 20404 960 20410 1012
rect 4706 892 4712 944
rect 4764 932 4770 944
rect 17862 932 17868 944
rect 4764 904 17868 932
rect 4764 892 4770 904
rect 17862 892 17868 904
rect 17920 892 17926 944
rect 3970 824 3976 876
rect 4028 864 4034 876
rect 21174 864 21180 876
rect 4028 836 21180 864
rect 4028 824 4034 836
rect 21174 824 21180 836
rect 21232 824 21238 876
rect 6638 756 6644 808
rect 6696 796 6702 808
rect 16482 796 16488 808
rect 6696 768 16488 796
rect 6696 756 6702 768
rect 16482 756 16488 768
rect 16540 756 16546 808
rect 6362 688 6368 740
rect 6420 728 6426 740
rect 34974 728 34980 740
rect 6420 700 34980 728
rect 6420 688 6426 700
rect 34974 688 34980 700
rect 35032 688 35038 740
rect 1486 552 1492 604
rect 1544 592 1550 604
rect 21266 592 21272 604
rect 1544 564 21272 592
rect 1544 552 1550 564
rect 21266 552 21272 564
rect 21324 552 21330 604
rect 3510 484 3516 536
rect 3568 524 3574 536
rect 18782 524 18788 536
rect 3568 496 18788 524
rect 3568 484 3574 496
rect 18782 484 18788 496
rect 18840 484 18846 536
rect 2222 416 2228 468
rect 2280 456 2286 468
rect 15470 456 15476 468
rect 2280 428 15476 456
rect 2280 416 2286 428
rect 15470 416 15476 428
rect 15528 416 15534 468
rect 3786 212 3792 264
rect 3844 252 3850 264
rect 18874 252 18880 264
rect 3844 224 18880 252
rect 3844 212 3850 224
rect 18874 212 18880 224
rect 18932 212 18938 264
rect 5902 144 5908 196
rect 5960 184 5966 196
rect 20806 184 20812 196
rect 5960 156 20812 184
rect 5960 144 5966 156
rect 20806 144 20812 156
rect 20864 144 20870 196
<< via1 >>
rect 7748 26936 7800 26988
rect 21732 26936 21784 26988
rect 10232 26868 10284 26920
rect 19708 26868 19760 26920
rect 9496 26596 9548 26648
rect 22928 26800 22980 26852
rect 23388 26800 23440 26852
rect 33692 26800 33744 26852
rect 16856 26528 16908 26580
rect 29828 26732 29880 26784
rect 20536 26596 20588 26648
rect 36544 26664 36596 26716
rect 25964 26596 26016 26648
rect 34612 26596 34664 26648
rect 17776 26528 17828 26580
rect 42892 26528 42944 26580
rect 17224 26460 17276 26512
rect 41604 26460 41656 26512
rect 1308 26324 1360 26376
rect 18880 26392 18932 26444
rect 19064 26392 19116 26444
rect 40960 26392 41012 26444
rect 14740 26324 14792 26376
rect 572 26256 624 26308
rect 22100 26256 22152 26308
rect 5264 26188 5316 26240
rect 20076 26188 20128 26240
rect 22376 26188 22428 26240
rect 23388 26188 23440 26240
rect 14188 26120 14240 26172
rect 19064 26120 19116 26172
rect 28264 26324 28316 26376
rect 45928 26324 45980 26376
rect 26976 26256 27028 26308
rect 36820 26256 36872 26308
rect 26884 26188 26936 26240
rect 37280 26188 37332 26240
rect 33876 26120 33928 26172
rect 17592 26052 17644 26104
rect 39120 26052 39172 26104
rect 12624 25984 12676 26036
rect 39764 25984 39816 26036
rect 8944 25916 8996 25968
rect 34704 25916 34756 25968
rect 7564 25848 7616 25900
rect 17868 25848 17920 25900
rect 21272 25848 21324 25900
rect 41880 25848 41932 25900
rect 6644 25780 6696 25832
rect 37004 25780 37056 25832
rect 3884 25712 3936 25764
rect 41144 25712 41196 25764
rect 8300 25644 8352 25696
rect 22100 25644 22152 25696
rect 22284 25644 22336 25696
rect 29552 25644 29604 25696
rect 2044 25576 2096 25628
rect 16212 25576 16264 25628
rect 17040 25576 17092 25628
rect 31944 25576 31996 25628
rect 2136 25508 2188 25560
rect 14556 25508 14608 25560
rect 14832 25508 14884 25560
rect 33784 25508 33836 25560
rect 9220 25440 9272 25492
rect 20812 25440 20864 25492
rect 21088 25440 21140 25492
rect 40316 25440 40368 25492
rect 17500 25372 17552 25424
rect 40408 25372 40460 25424
rect 15016 25304 15068 25356
rect 7104 25236 7156 25288
rect 16948 25236 17000 25288
rect 18696 25304 18748 25356
rect 43628 25304 43680 25356
rect 1860 25168 1912 25220
rect 6736 25100 6788 25152
rect 16396 25100 16448 25152
rect 20812 25168 20864 25220
rect 21916 25168 21968 25220
rect 22100 25236 22152 25288
rect 22560 25236 22612 25288
rect 22652 25236 22704 25288
rect 23940 25168 23992 25220
rect 30380 25236 30432 25288
rect 44364 25236 44416 25288
rect 36636 25168 36688 25220
rect 19892 25100 19944 25152
rect 19984 25100 20036 25152
rect 36176 25100 36228 25152
rect 4068 25032 4120 25084
rect 10048 25032 10100 25084
rect 12072 25032 12124 25084
rect 4528 24964 4580 25016
rect 15844 24964 15896 25016
rect 5724 24896 5776 24948
rect 13728 24896 13780 24948
rect 16948 25032 17000 25084
rect 23388 25032 23440 25084
rect 24584 25032 24636 25084
rect 26240 25032 26292 25084
rect 28724 25032 28776 25084
rect 39212 25032 39264 25084
rect 16488 24964 16540 25016
rect 18144 24896 18196 24948
rect 20260 24896 20312 24948
rect 20720 24896 20772 24948
rect 3332 24828 3384 24880
rect 4896 24828 4948 24880
rect 8392 24828 8444 24880
rect 11060 24828 11112 24880
rect 13636 24828 13688 24880
rect 17960 24828 18012 24880
rect 18512 24828 18564 24880
rect 20812 24828 20864 24880
rect 6552 24760 6604 24812
rect 21364 24760 21416 24812
rect 23480 24964 23532 25016
rect 35808 24964 35860 25016
rect 22836 24896 22888 24948
rect 26976 24896 27028 24948
rect 28816 24896 28868 24948
rect 31116 24896 31168 24948
rect 32680 24896 32732 24948
rect 42064 24896 42116 24948
rect 22560 24828 22612 24880
rect 24584 24828 24636 24880
rect 24676 24828 24728 24880
rect 29184 24828 29236 24880
rect 25964 24760 26016 24812
rect 26240 24760 26292 24812
rect 30656 24828 30708 24880
rect 13728 24692 13780 24744
rect 16304 24692 16356 24744
rect 17868 24692 17920 24744
rect 22560 24692 22612 24744
rect 22836 24692 22888 24744
rect 28356 24692 28408 24744
rect 12348 24624 12400 24676
rect 25780 24624 25832 24676
rect 26608 24624 26660 24676
rect 29920 24624 29972 24676
rect 14004 24556 14056 24608
rect 16856 24556 16908 24608
rect 16948 24556 17000 24608
rect 17132 24556 17184 24608
rect 17960 24556 18012 24608
rect 19800 24556 19852 24608
rect 20352 24556 20404 24608
rect 26056 24556 26108 24608
rect 29460 24556 29512 24608
rect 37464 24556 37516 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 848 24352 900 24404
rect 3516 24216 3568 24268
rect 3976 24352 4028 24404
rect 7472 24352 7524 24404
rect 11428 24352 11480 24404
rect 9312 24284 9364 24336
rect 7380 24216 7432 24268
rect 2228 24191 2280 24200
rect 2228 24157 2237 24191
rect 2237 24157 2271 24191
rect 2271 24157 2280 24191
rect 2228 24148 2280 24157
rect 4712 24148 4764 24200
rect 4804 24191 4856 24200
rect 4804 24157 4813 24191
rect 4813 24157 4847 24191
rect 4847 24157 4856 24191
rect 4804 24148 4856 24157
rect 6552 24191 6604 24200
rect 6552 24157 6561 24191
rect 6561 24157 6595 24191
rect 6595 24157 6604 24191
rect 6552 24148 6604 24157
rect 11520 24216 11572 24268
rect 9772 24191 9824 24200
rect 9772 24157 9781 24191
rect 9781 24157 9815 24191
rect 9815 24157 9824 24191
rect 9772 24148 9824 24157
rect 14464 24284 14516 24336
rect 16672 24352 16724 24404
rect 24768 24352 24820 24404
rect 25780 24395 25832 24404
rect 25780 24361 25789 24395
rect 25789 24361 25823 24395
rect 25823 24361 25832 24395
rect 25780 24352 25832 24361
rect 16856 24284 16908 24336
rect 18144 24284 18196 24336
rect 21456 24284 21508 24336
rect 24860 24284 24912 24336
rect 25964 24352 26016 24404
rect 14372 24216 14424 24268
rect 12532 24191 12584 24200
rect 12532 24157 12541 24191
rect 12541 24157 12575 24191
rect 12575 24157 12584 24191
rect 12532 24148 12584 24157
rect 14464 24191 14516 24200
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 18972 24216 19024 24268
rect 14464 24148 14516 24157
rect 1768 24055 1820 24064
rect 1768 24021 1777 24055
rect 1777 24021 1811 24055
rect 1811 24021 1820 24055
rect 1768 24012 1820 24021
rect 3516 24012 3568 24064
rect 10140 24080 10192 24132
rect 13820 24080 13872 24132
rect 7380 24012 7432 24064
rect 9128 24055 9180 24064
rect 9128 24021 9137 24055
rect 9137 24021 9171 24055
rect 9171 24021 9180 24055
rect 9128 24012 9180 24021
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 11796 24012 11848 24064
rect 12440 24012 12492 24064
rect 12532 24012 12584 24064
rect 14188 24012 14240 24064
rect 14280 24055 14332 24064
rect 14280 24021 14289 24055
rect 14289 24021 14323 24055
rect 14323 24021 14332 24055
rect 14280 24012 14332 24021
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 19616 24191 19668 24200
rect 19616 24157 19625 24191
rect 19625 24157 19659 24191
rect 19659 24157 19668 24191
rect 19616 24148 19668 24157
rect 16764 24080 16816 24132
rect 18420 24080 18472 24132
rect 19524 24080 19576 24132
rect 20628 24216 20680 24268
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 21548 24216 21600 24268
rect 22560 24216 22612 24268
rect 25136 24216 25188 24268
rect 26056 24216 26108 24268
rect 26424 24216 26476 24268
rect 27160 24327 27212 24336
rect 27160 24293 27169 24327
rect 27169 24293 27203 24327
rect 27203 24293 27212 24327
rect 27160 24284 27212 24293
rect 29092 24284 29144 24336
rect 27712 24259 27764 24268
rect 27712 24225 27721 24259
rect 27721 24225 27755 24259
rect 27755 24225 27764 24259
rect 27712 24216 27764 24225
rect 27804 24216 27856 24268
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20168 24148 20220 24200
rect 22284 24148 22336 24200
rect 24768 24148 24820 24200
rect 28356 24191 28408 24200
rect 28356 24157 28365 24191
rect 28365 24157 28399 24191
rect 28399 24157 28408 24191
rect 28356 24148 28408 24157
rect 29184 24216 29236 24268
rect 29276 24216 29328 24268
rect 29736 24259 29788 24268
rect 29736 24225 29745 24259
rect 29745 24225 29779 24259
rect 29779 24225 29788 24259
rect 29736 24216 29788 24225
rect 29920 24284 29972 24336
rect 32220 24216 32272 24268
rect 31024 24191 31076 24200
rect 31024 24157 31033 24191
rect 31033 24157 31067 24191
rect 31067 24157 31076 24191
rect 31024 24148 31076 24157
rect 27252 24080 27304 24132
rect 27436 24080 27488 24132
rect 34336 24191 34388 24200
rect 34336 24157 34345 24191
rect 34345 24157 34379 24191
rect 34379 24157 34388 24191
rect 34336 24148 34388 24157
rect 36636 24327 36688 24336
rect 36636 24293 36645 24327
rect 36645 24293 36679 24327
rect 36679 24293 36688 24327
rect 36636 24284 36688 24293
rect 37004 24327 37056 24336
rect 37004 24293 37013 24327
rect 37013 24293 37047 24327
rect 37047 24293 37056 24327
rect 37004 24284 37056 24293
rect 37372 24148 37424 24200
rect 37464 24191 37516 24200
rect 37464 24157 37473 24191
rect 37473 24157 37507 24191
rect 37507 24157 37516 24191
rect 37464 24148 37516 24157
rect 35624 24080 35676 24132
rect 45928 24352 45980 24404
rect 39396 24284 39448 24336
rect 44916 24284 44968 24336
rect 41420 24148 41472 24200
rect 41512 24191 41564 24200
rect 41512 24157 41521 24191
rect 41521 24157 41555 24191
rect 41555 24157 41564 24191
rect 41512 24148 41564 24157
rect 42800 24148 42852 24200
rect 43904 24191 43956 24200
rect 43904 24157 43913 24191
rect 43913 24157 43947 24191
rect 43947 24157 43956 24191
rect 43904 24148 43956 24157
rect 44456 24148 44508 24200
rect 42708 24080 42760 24132
rect 48412 24148 48464 24200
rect 49240 24148 49292 24200
rect 49332 24080 49384 24132
rect 17868 24012 17920 24064
rect 18788 24012 18840 24064
rect 19064 24055 19116 24064
rect 19064 24021 19073 24055
rect 19073 24021 19107 24055
rect 19107 24021 19116 24055
rect 19064 24012 19116 24021
rect 24492 24012 24544 24064
rect 24584 24055 24636 24064
rect 24584 24021 24593 24055
rect 24593 24021 24627 24055
rect 24627 24021 24636 24055
rect 24584 24012 24636 24021
rect 25872 24012 25924 24064
rect 26332 24012 26384 24064
rect 26516 24012 26568 24064
rect 29276 24055 29328 24064
rect 29276 24021 29285 24055
rect 29285 24021 29319 24055
rect 29319 24021 29328 24055
rect 29276 24012 29328 24021
rect 29368 24012 29420 24064
rect 32036 24012 32088 24064
rect 35440 24012 35492 24064
rect 37464 24012 37516 24064
rect 39488 24055 39540 24064
rect 39488 24021 39497 24055
rect 39497 24021 39531 24055
rect 39531 24021 39540 24055
rect 39488 24012 39540 24021
rect 39672 24012 39724 24064
rect 42892 24012 42944 24064
rect 43812 24012 43864 24064
rect 44548 24055 44600 24064
rect 44548 24021 44557 24055
rect 44557 24021 44591 24055
rect 44591 24021 44600 24055
rect 44548 24012 44600 24021
rect 48320 24012 48372 24064
rect 48504 24012 48556 24064
rect 48964 24012 49016 24064
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 1768 23808 1820 23860
rect 14464 23808 14516 23860
rect 16304 23808 16356 23860
rect 18972 23808 19024 23860
rect 19064 23808 19116 23860
rect 22284 23808 22336 23860
rect 24860 23808 24912 23860
rect 756 23740 808 23792
rect 2412 23604 2464 23656
rect 1952 23536 2004 23588
rect 2780 23604 2832 23656
rect 4160 23672 4212 23724
rect 9128 23740 9180 23792
rect 11796 23740 11848 23792
rect 12256 23783 12308 23792
rect 12256 23749 12265 23783
rect 12265 23749 12299 23783
rect 12299 23749 12308 23783
rect 12256 23740 12308 23749
rect 12348 23783 12400 23792
rect 12348 23749 12357 23783
rect 12357 23749 12391 23783
rect 12391 23749 12400 23783
rect 12348 23740 12400 23749
rect 5448 23647 5500 23656
rect 5448 23613 5457 23647
rect 5457 23613 5491 23647
rect 5491 23613 5500 23647
rect 5448 23604 5500 23613
rect 6736 23672 6788 23724
rect 7932 23604 7984 23656
rect 2596 23468 2648 23520
rect 4988 23536 5040 23588
rect 5356 23536 5408 23588
rect 9864 23715 9916 23724
rect 9864 23681 9873 23715
rect 9873 23681 9907 23715
rect 9907 23681 9916 23715
rect 9864 23672 9916 23681
rect 13912 23740 13964 23792
rect 15752 23740 15804 23792
rect 15936 23740 15988 23792
rect 17592 23740 17644 23792
rect 19156 23740 19208 23792
rect 19524 23740 19576 23792
rect 21364 23783 21416 23792
rect 21364 23749 21373 23783
rect 21373 23749 21407 23783
rect 21407 23749 21416 23783
rect 21364 23740 21416 23749
rect 22560 23740 22612 23792
rect 23296 23740 23348 23792
rect 25044 23740 25096 23792
rect 29368 23808 29420 23860
rect 31024 23808 31076 23860
rect 33692 23808 33744 23860
rect 27068 23740 27120 23792
rect 27712 23740 27764 23792
rect 9956 23604 10008 23656
rect 8116 23536 8168 23588
rect 12348 23604 12400 23656
rect 13360 23672 13412 23724
rect 14924 23715 14976 23724
rect 14924 23681 14933 23715
rect 14933 23681 14967 23715
rect 14967 23681 14976 23715
rect 14924 23672 14976 23681
rect 18512 23672 18564 23724
rect 20996 23715 21048 23724
rect 20996 23681 21005 23715
rect 21005 23681 21039 23715
rect 21039 23681 21048 23715
rect 20996 23672 21048 23681
rect 18328 23604 18380 23656
rect 18788 23647 18840 23656
rect 18788 23613 18797 23647
rect 18797 23613 18831 23647
rect 18831 23613 18840 23647
rect 18788 23604 18840 23613
rect 7656 23468 7708 23520
rect 7932 23468 7984 23520
rect 9680 23468 9732 23520
rect 12164 23468 12216 23520
rect 15200 23536 15252 23588
rect 15292 23536 15344 23588
rect 18236 23536 18288 23588
rect 18696 23536 18748 23588
rect 19156 23604 19208 23656
rect 20904 23604 20956 23656
rect 22376 23604 22428 23656
rect 22744 23604 22796 23656
rect 22928 23604 22980 23656
rect 24860 23647 24912 23656
rect 24860 23613 24869 23647
rect 24869 23613 24903 23647
rect 24903 23613 24912 23647
rect 24860 23604 24912 23613
rect 13912 23468 13964 23520
rect 18788 23468 18840 23520
rect 20076 23468 20128 23520
rect 20352 23536 20404 23588
rect 23388 23536 23440 23588
rect 26424 23604 26476 23656
rect 26608 23579 26660 23588
rect 26608 23545 26617 23579
rect 26617 23545 26651 23579
rect 26651 23545 26660 23579
rect 26608 23536 26660 23545
rect 24860 23468 24912 23520
rect 27436 23647 27488 23656
rect 27436 23613 27445 23647
rect 27445 23613 27479 23647
rect 27479 23613 27488 23647
rect 27436 23604 27488 23613
rect 27804 23604 27856 23656
rect 28816 23740 28868 23792
rect 28908 23740 28960 23792
rect 31392 23740 31444 23792
rect 29000 23672 29052 23724
rect 28816 23604 28868 23656
rect 29644 23647 29696 23656
rect 29644 23613 29653 23647
rect 29653 23613 29687 23647
rect 29687 23613 29696 23647
rect 29644 23604 29696 23613
rect 30748 23672 30800 23724
rect 32036 23740 32088 23792
rect 32220 23740 32272 23792
rect 32312 23715 32364 23724
rect 32312 23681 32321 23715
rect 32321 23681 32355 23715
rect 32355 23681 32364 23715
rect 32312 23672 32364 23681
rect 40316 23851 40368 23860
rect 40316 23817 40325 23851
rect 40325 23817 40359 23851
rect 40359 23817 40368 23851
rect 40316 23808 40368 23817
rect 41420 23808 41472 23860
rect 48412 23851 48464 23860
rect 48412 23817 48421 23851
rect 48421 23817 48455 23851
rect 48455 23817 48464 23851
rect 48412 23808 48464 23817
rect 35624 23672 35676 23724
rect 31116 23604 31168 23656
rect 31668 23604 31720 23656
rect 29460 23536 29512 23588
rect 29736 23536 29788 23588
rect 39672 23715 39724 23724
rect 39672 23681 39681 23715
rect 39681 23681 39715 23715
rect 39715 23681 39724 23715
rect 39672 23672 39724 23681
rect 40500 23604 40552 23656
rect 39948 23536 40000 23588
rect 42708 23783 42760 23792
rect 42708 23749 42717 23783
rect 42717 23749 42751 23783
rect 42751 23749 42760 23783
rect 42708 23740 42760 23749
rect 42892 23783 42944 23792
rect 42892 23749 42901 23783
rect 42901 23749 42935 23783
rect 42935 23749 42944 23783
rect 42892 23740 42944 23749
rect 41788 23672 41840 23724
rect 42800 23672 42852 23724
rect 43352 23672 43404 23724
rect 47308 23740 47360 23792
rect 44824 23715 44876 23724
rect 44824 23681 44833 23715
rect 44833 23681 44867 23715
rect 44867 23681 44876 23715
rect 44824 23672 44876 23681
rect 43444 23604 43496 23656
rect 27160 23468 27212 23520
rect 27252 23468 27304 23520
rect 29000 23468 29052 23520
rect 29276 23468 29328 23520
rect 31760 23468 31812 23520
rect 35992 23468 36044 23520
rect 37096 23511 37148 23520
rect 37096 23477 37105 23511
rect 37105 23477 37139 23511
rect 37139 23477 37148 23511
rect 37096 23468 37148 23477
rect 38568 23468 38620 23520
rect 41880 23579 41932 23588
rect 41880 23545 41889 23579
rect 41889 23545 41923 23579
rect 41923 23545 41932 23579
rect 41880 23536 41932 23545
rect 44916 23604 44968 23656
rect 47032 23672 47084 23724
rect 48872 23715 48924 23724
rect 48872 23681 48881 23715
rect 48881 23681 48915 23715
rect 48915 23681 48924 23715
rect 48872 23672 48924 23681
rect 45928 23647 45980 23656
rect 45928 23613 45937 23647
rect 45937 23613 45971 23647
rect 45971 23613 45980 23647
rect 45928 23604 45980 23613
rect 46940 23536 46992 23588
rect 44180 23468 44232 23520
rect 49056 23511 49108 23520
rect 49056 23477 49065 23511
rect 49065 23477 49099 23511
rect 49099 23477 49108 23511
rect 49056 23468 49108 23477
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 2872 23264 2924 23316
rect 4160 23264 4212 23316
rect 8024 23264 8076 23316
rect 12624 23264 12676 23316
rect 13544 23264 13596 23316
rect 14188 23264 14240 23316
rect 3608 23239 3660 23248
rect 3608 23205 3617 23239
rect 3617 23205 3651 23239
rect 3651 23205 3660 23239
rect 3608 23196 3660 23205
rect 7288 23196 7340 23248
rect 5264 23128 5316 23180
rect 6092 23171 6144 23180
rect 6092 23137 6101 23171
rect 6101 23137 6135 23171
rect 6135 23137 6144 23171
rect 6092 23128 6144 23137
rect 7840 23171 7892 23180
rect 7840 23137 7849 23171
rect 7849 23137 7883 23171
rect 7883 23137 7892 23171
rect 7840 23128 7892 23137
rect 10508 23171 10560 23180
rect 10508 23137 10517 23171
rect 10517 23137 10551 23171
rect 10551 23137 10560 23171
rect 10508 23128 10560 23137
rect 13912 23239 13964 23248
rect 13912 23205 13921 23239
rect 13921 23205 13955 23239
rect 13955 23205 13964 23239
rect 13912 23196 13964 23205
rect 14096 23196 14148 23248
rect 11796 23128 11848 23180
rect 11888 23128 11940 23180
rect 12808 23128 12860 23180
rect 13544 23128 13596 23180
rect 14740 23128 14792 23180
rect 16856 23128 16908 23180
rect 17776 23128 17828 23180
rect 20076 23171 20128 23180
rect 20076 23137 20085 23171
rect 20085 23137 20119 23171
rect 20119 23137 20128 23171
rect 20076 23128 20128 23137
rect 20904 23128 20956 23180
rect 22284 23171 22336 23180
rect 22284 23137 22293 23171
rect 22293 23137 22327 23171
rect 22327 23137 22336 23171
rect 22284 23128 22336 23137
rect 22652 23128 22704 23180
rect 23296 23128 23348 23180
rect 1860 23060 1912 23112
rect 2780 23035 2832 23044
rect 2780 23001 2789 23035
rect 2789 23001 2823 23035
rect 2823 23001 2832 23035
rect 2780 22992 2832 23001
rect 6184 23060 6236 23112
rect 8024 23060 8076 23112
rect 9496 23103 9548 23112
rect 9496 23069 9505 23103
rect 9505 23069 9539 23103
rect 9539 23069 9548 23103
rect 9496 23060 9548 23069
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 14648 23103 14700 23112
rect 14648 23069 14657 23103
rect 14657 23069 14691 23103
rect 14691 23069 14700 23103
rect 14648 23060 14700 23069
rect 15476 23103 15528 23112
rect 15476 23069 15485 23103
rect 15485 23069 15519 23103
rect 15519 23069 15528 23103
rect 15476 23060 15528 23069
rect 11060 22992 11112 23044
rect 11428 23035 11480 23044
rect 11428 23001 11437 23035
rect 11437 23001 11471 23035
rect 11471 23001 11480 23035
rect 11428 22992 11480 23001
rect 9036 22967 9088 22976
rect 9036 22933 9045 22967
rect 9045 22933 9079 22967
rect 9079 22933 9088 22967
rect 9036 22924 9088 22933
rect 9404 22924 9456 22976
rect 10784 22924 10836 22976
rect 12992 22992 13044 23044
rect 13360 22992 13412 23044
rect 23664 23060 23716 23112
rect 23848 23264 23900 23316
rect 24860 23264 24912 23316
rect 26056 23264 26108 23316
rect 29644 23264 29696 23316
rect 30196 23264 30248 23316
rect 32220 23264 32272 23316
rect 32312 23264 32364 23316
rect 24124 23196 24176 23248
rect 24768 23196 24820 23248
rect 25320 23196 25372 23248
rect 25780 23128 25832 23180
rect 25964 23128 26016 23180
rect 13728 22967 13780 22976
rect 13728 22933 13737 22967
rect 13737 22933 13771 22967
rect 13771 22933 13780 22967
rect 13728 22924 13780 22933
rect 14280 22967 14332 22976
rect 14280 22933 14289 22967
rect 14289 22933 14323 22967
rect 14323 22933 14332 22967
rect 14280 22924 14332 22933
rect 14740 22967 14792 22976
rect 14740 22933 14749 22967
rect 14749 22933 14783 22967
rect 14783 22933 14792 22967
rect 14740 22924 14792 22933
rect 17684 22992 17736 23044
rect 18420 22992 18472 23044
rect 20260 22992 20312 23044
rect 17224 22924 17276 22976
rect 18972 22924 19024 22976
rect 20628 22992 20680 23044
rect 21088 22924 21140 22976
rect 21180 22924 21232 22976
rect 21824 22967 21876 22976
rect 21824 22933 21833 22967
rect 21833 22933 21867 22967
rect 21867 22933 21876 22967
rect 21824 22924 21876 22933
rect 23296 22992 23348 23044
rect 24124 22924 24176 22976
rect 24952 23035 25004 23044
rect 24952 23001 24961 23035
rect 24961 23001 24995 23035
rect 24995 23001 25004 23035
rect 24952 22992 25004 23001
rect 26148 23060 26200 23112
rect 26700 23196 26752 23248
rect 27252 23196 27304 23248
rect 29092 23239 29144 23248
rect 29092 23205 29101 23239
rect 29101 23205 29135 23239
rect 29135 23205 29144 23239
rect 29092 23196 29144 23205
rect 31760 23196 31812 23248
rect 40500 23264 40552 23316
rect 41788 23307 41840 23316
rect 41788 23273 41797 23307
rect 41797 23273 41831 23307
rect 41831 23273 41840 23307
rect 41788 23264 41840 23273
rect 27160 23128 27212 23180
rect 28908 23128 28960 23180
rect 33416 23196 33468 23248
rect 36360 23196 36412 23248
rect 32496 23128 32548 23180
rect 37096 23128 37148 23180
rect 39580 23196 39632 23248
rect 41236 23196 41288 23248
rect 43168 23264 43220 23316
rect 43444 23264 43496 23316
rect 44364 23264 44416 23316
rect 46664 23264 46716 23316
rect 48872 23264 48924 23316
rect 49332 23307 49384 23316
rect 49332 23273 49341 23307
rect 49341 23273 49375 23307
rect 49375 23273 49384 23307
rect 49332 23264 49384 23273
rect 43628 23196 43680 23248
rect 46112 23239 46164 23248
rect 46112 23205 46121 23239
rect 46121 23205 46155 23239
rect 46155 23205 46164 23239
rect 46112 23196 46164 23205
rect 26700 22992 26752 23044
rect 25504 22924 25556 22976
rect 25596 22924 25648 22976
rect 25872 22924 25924 22976
rect 26056 22924 26108 22976
rect 26884 22967 26936 22976
rect 26884 22933 26893 22967
rect 26893 22933 26927 22967
rect 26927 22933 26936 22967
rect 26884 22924 26936 22933
rect 29276 23060 29328 23112
rect 31392 23060 31444 23112
rect 33140 23060 33192 23112
rect 27712 22992 27764 23044
rect 29000 22992 29052 23044
rect 29644 22992 29696 23044
rect 30104 22992 30156 23044
rect 35992 23103 36044 23112
rect 35992 23069 36001 23103
rect 36001 23069 36035 23103
rect 36035 23069 36044 23103
rect 35992 23060 36044 23069
rect 36820 23060 36872 23112
rect 40040 23103 40092 23112
rect 40040 23069 40049 23103
rect 40049 23069 40083 23103
rect 40083 23069 40092 23103
rect 40040 23060 40092 23069
rect 41144 23103 41196 23112
rect 41144 23069 41153 23103
rect 41153 23069 41187 23103
rect 41187 23069 41196 23103
rect 41144 23060 41196 23069
rect 44548 23128 44600 23180
rect 44180 23060 44232 23112
rect 44640 23103 44692 23112
rect 44640 23069 44649 23103
rect 44649 23069 44683 23103
rect 44683 23069 44692 23103
rect 44640 23060 44692 23069
rect 48504 23196 48556 23248
rect 48504 23060 48556 23112
rect 49332 23060 49384 23112
rect 29736 22924 29788 22976
rect 30196 22924 30248 22976
rect 33968 22992 34020 23044
rect 31576 22924 31628 22976
rect 31944 22924 31996 22976
rect 33048 22924 33100 22976
rect 33508 22924 33560 22976
rect 34796 22924 34848 22976
rect 37096 22967 37148 22976
rect 37096 22933 37105 22967
rect 37105 22933 37139 22967
rect 37139 22933 37148 22967
rect 37096 22924 37148 22933
rect 38292 22992 38344 23044
rect 40316 22992 40368 23044
rect 42800 22992 42852 23044
rect 39488 22967 39540 22976
rect 39488 22933 39497 22967
rect 39497 22933 39531 22967
rect 39531 22933 39540 22967
rect 39488 22924 39540 22933
rect 39764 22924 39816 22976
rect 41052 22924 41104 22976
rect 45836 22967 45888 22976
rect 45836 22933 45845 22967
rect 45845 22933 45879 22967
rect 45879 22933 45888 22967
rect 45836 22924 45888 22933
rect 47216 22924 47268 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 4528 22720 4580 22772
rect 2044 22584 2096 22636
rect 8576 22695 8628 22704
rect 8576 22661 8585 22695
rect 8585 22661 8619 22695
rect 8619 22661 8628 22695
rect 8576 22652 8628 22661
rect 388 22516 440 22568
rect 2228 22559 2280 22568
rect 2228 22525 2237 22559
rect 2237 22525 2271 22559
rect 2271 22525 2280 22559
rect 2228 22516 2280 22525
rect 4068 22559 4120 22568
rect 4068 22525 4077 22559
rect 4077 22525 4111 22559
rect 4111 22525 4120 22559
rect 4068 22516 4120 22525
rect 3424 22423 3476 22432
rect 3424 22389 3433 22423
rect 3433 22389 3467 22423
rect 3467 22389 3476 22423
rect 3424 22380 3476 22389
rect 7564 22627 7616 22636
rect 7564 22593 7573 22627
rect 7573 22593 7607 22627
rect 7607 22593 7616 22627
rect 7564 22584 7616 22593
rect 7748 22584 7800 22636
rect 10784 22652 10836 22704
rect 11980 22695 12032 22704
rect 11980 22661 11989 22695
rect 11989 22661 12023 22695
rect 12023 22661 12032 22695
rect 11980 22652 12032 22661
rect 12532 22695 12584 22704
rect 12532 22661 12541 22695
rect 12541 22661 12575 22695
rect 12575 22661 12584 22695
rect 12532 22652 12584 22661
rect 12992 22652 13044 22704
rect 11152 22584 11204 22636
rect 12256 22627 12308 22636
rect 12256 22593 12265 22627
rect 12265 22593 12299 22627
rect 12299 22593 12308 22627
rect 12256 22584 12308 22593
rect 14556 22584 14608 22636
rect 14832 22584 14884 22636
rect 14924 22627 14976 22636
rect 14924 22593 14933 22627
rect 14933 22593 14967 22627
rect 14967 22593 14976 22627
rect 14924 22584 14976 22593
rect 16120 22695 16172 22704
rect 16120 22661 16129 22695
rect 16129 22661 16163 22695
rect 16163 22661 16172 22695
rect 16120 22652 16172 22661
rect 17224 22652 17276 22704
rect 18420 22652 18472 22704
rect 16580 22584 16632 22636
rect 5080 22559 5132 22568
rect 5080 22525 5089 22559
rect 5089 22525 5123 22559
rect 5123 22525 5132 22559
rect 5080 22516 5132 22525
rect 6644 22516 6696 22568
rect 8668 22516 8720 22568
rect 6000 22448 6052 22500
rect 15476 22516 15528 22568
rect 16856 22559 16908 22568
rect 16856 22525 16865 22559
rect 16865 22525 16899 22559
rect 16899 22525 16908 22559
rect 16856 22516 16908 22525
rect 8392 22380 8444 22432
rect 9956 22380 10008 22432
rect 11336 22423 11388 22432
rect 11336 22389 11345 22423
rect 11345 22389 11379 22423
rect 11379 22389 11388 22423
rect 11336 22380 11388 22389
rect 11428 22380 11480 22432
rect 16120 22448 16172 22500
rect 18604 22720 18656 22772
rect 20076 22652 20128 22704
rect 20628 22652 20680 22704
rect 19616 22516 19668 22568
rect 19708 22559 19760 22568
rect 19708 22525 19717 22559
rect 19717 22525 19751 22559
rect 19751 22525 19760 22559
rect 19708 22516 19760 22525
rect 20996 22516 21048 22568
rect 22284 22584 22336 22636
rect 23388 22652 23440 22704
rect 23664 22652 23716 22704
rect 25228 22652 25280 22704
rect 29368 22720 29420 22772
rect 29460 22720 29512 22772
rect 30012 22720 30064 22772
rect 24768 22584 24820 22636
rect 25136 22584 25188 22636
rect 27160 22652 27212 22704
rect 28724 22695 28776 22704
rect 28724 22661 28733 22695
rect 28733 22661 28767 22695
rect 28767 22661 28776 22695
rect 28724 22652 28776 22661
rect 30104 22652 30156 22704
rect 14004 22423 14056 22432
rect 14004 22389 14013 22423
rect 14013 22389 14047 22423
rect 14047 22389 14056 22423
rect 14004 22380 14056 22389
rect 14832 22380 14884 22432
rect 20352 22380 20404 22432
rect 22652 22423 22704 22432
rect 22652 22389 22661 22423
rect 22661 22389 22695 22423
rect 22695 22389 22704 22423
rect 22652 22380 22704 22389
rect 23480 22516 23532 22568
rect 23940 22516 23992 22568
rect 24124 22516 24176 22568
rect 24676 22380 24728 22432
rect 25780 22559 25832 22568
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 25964 22559 26016 22568
rect 25964 22525 25973 22559
rect 25973 22525 26007 22559
rect 26007 22525 26016 22559
rect 25964 22516 26016 22525
rect 27160 22516 27212 22568
rect 25872 22380 25924 22432
rect 26332 22380 26384 22432
rect 26884 22380 26936 22432
rect 27620 22627 27672 22636
rect 27620 22593 27629 22627
rect 27629 22593 27663 22627
rect 27663 22593 27672 22627
rect 27620 22584 27672 22593
rect 28448 22627 28500 22636
rect 28448 22593 28457 22627
rect 28457 22593 28491 22627
rect 28491 22593 28500 22627
rect 28448 22584 28500 22593
rect 27712 22559 27764 22568
rect 27712 22525 27721 22559
rect 27721 22525 27755 22559
rect 27755 22525 27764 22559
rect 27712 22516 27764 22525
rect 31392 22720 31444 22772
rect 31760 22720 31812 22772
rect 32496 22720 32548 22772
rect 34336 22763 34388 22772
rect 34336 22729 34345 22763
rect 34345 22729 34379 22763
rect 34379 22729 34388 22763
rect 34336 22720 34388 22729
rect 35440 22720 35492 22772
rect 35900 22720 35952 22772
rect 36820 22720 36872 22772
rect 37372 22720 37424 22772
rect 38936 22720 38988 22772
rect 40500 22720 40552 22772
rect 43904 22720 43956 22772
rect 31208 22652 31260 22704
rect 31300 22652 31352 22704
rect 44640 22652 44692 22704
rect 45376 22652 45428 22704
rect 46940 22652 46992 22704
rect 47308 22652 47360 22704
rect 31484 22584 31536 22636
rect 33324 22584 33376 22636
rect 33968 22584 34020 22636
rect 37188 22584 37240 22636
rect 37464 22627 37516 22636
rect 37464 22593 37473 22627
rect 37473 22593 37507 22627
rect 37507 22593 37516 22627
rect 37464 22584 37516 22593
rect 38568 22627 38620 22636
rect 38568 22593 38577 22627
rect 38577 22593 38611 22627
rect 38611 22593 38620 22627
rect 38568 22584 38620 22593
rect 39212 22627 39264 22636
rect 39212 22593 39221 22627
rect 39221 22593 39255 22627
rect 39255 22593 39264 22627
rect 39212 22584 39264 22593
rect 39672 22627 39724 22636
rect 39672 22593 39681 22627
rect 39681 22593 39715 22627
rect 39715 22593 39724 22627
rect 39672 22584 39724 22593
rect 27528 22448 27580 22500
rect 31576 22516 31628 22568
rect 40040 22516 40092 22568
rect 29736 22448 29788 22500
rect 33048 22448 33100 22500
rect 28908 22380 28960 22432
rect 29920 22380 29972 22432
rect 30196 22423 30248 22432
rect 30196 22389 30205 22423
rect 30205 22389 30239 22423
rect 30239 22389 30248 22423
rect 30196 22380 30248 22389
rect 30288 22380 30340 22432
rect 31760 22423 31812 22432
rect 31760 22389 31769 22423
rect 31769 22389 31803 22423
rect 31803 22389 31812 22423
rect 31760 22380 31812 22389
rect 32496 22380 32548 22432
rect 34796 22448 34848 22500
rect 37004 22448 37056 22500
rect 41052 22584 41104 22636
rect 43720 22584 43772 22636
rect 44916 22584 44968 22636
rect 45008 22627 45060 22636
rect 45008 22593 45017 22627
rect 45017 22593 45051 22627
rect 45051 22593 45060 22627
rect 45008 22584 45060 22593
rect 45100 22584 45152 22636
rect 41880 22559 41932 22568
rect 41880 22525 41889 22559
rect 41889 22525 41923 22559
rect 41923 22525 41932 22559
rect 41880 22516 41932 22525
rect 43168 22516 43220 22568
rect 43996 22516 44048 22568
rect 45652 22516 45704 22568
rect 46480 22627 46532 22636
rect 46480 22593 46489 22627
rect 46489 22593 46523 22627
rect 46523 22593 46532 22627
rect 46480 22584 46532 22593
rect 48320 22584 48372 22636
rect 44364 22448 44416 22500
rect 44824 22448 44876 22500
rect 40132 22380 40184 22432
rect 40868 22380 40920 22432
rect 43444 22380 43496 22432
rect 44548 22423 44600 22432
rect 44548 22389 44557 22423
rect 44557 22389 44591 22423
rect 44591 22389 44600 22423
rect 44548 22380 44600 22389
rect 45192 22423 45244 22432
rect 45192 22389 45201 22423
rect 45201 22389 45235 22423
rect 45235 22389 45244 22423
rect 45192 22380 45244 22389
rect 46664 22423 46716 22432
rect 46664 22389 46673 22423
rect 46673 22389 46707 22423
rect 46707 22389 46716 22423
rect 46664 22380 46716 22389
rect 46940 22380 46992 22432
rect 48688 22380 48740 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 3332 22176 3384 22228
rect 4344 22176 4396 22228
rect 4620 22176 4672 22228
rect 14740 22176 14792 22228
rect 14832 22176 14884 22228
rect 16304 22176 16356 22228
rect 16580 22176 16632 22228
rect 17500 22176 17552 22228
rect 17960 22176 18012 22228
rect 19432 22176 19484 22228
rect 3976 22108 4028 22160
rect 4252 22108 4304 22160
rect 1492 22040 1544 22092
rect 3332 22040 3384 22092
rect 7012 22040 7064 22092
rect 11888 22108 11940 22160
rect 12716 22108 12768 22160
rect 16764 22108 16816 22160
rect 21272 22176 21324 22228
rect 22652 22176 22704 22228
rect 26148 22176 26200 22228
rect 10416 22040 10468 22092
rect 11244 22083 11296 22092
rect 11244 22049 11253 22083
rect 11253 22049 11287 22083
rect 11287 22049 11296 22083
rect 11244 22040 11296 22049
rect 13452 22083 13504 22092
rect 13452 22049 13461 22083
rect 13461 22049 13495 22083
rect 13495 22049 13504 22083
rect 13452 22040 13504 22049
rect 1584 22015 1636 22024
rect 1584 21981 1593 22015
rect 1593 21981 1627 22015
rect 1627 21981 1636 22015
rect 1584 21972 1636 21981
rect 3976 22015 4028 22024
rect 3976 21981 3985 22015
rect 3985 21981 4019 22015
rect 4019 21981 4028 22015
rect 3976 21972 4028 21981
rect 5540 21904 5592 21956
rect 6920 22015 6972 22024
rect 6920 21981 6929 22015
rect 6929 21981 6963 22015
rect 6963 21981 6972 22015
rect 6920 21972 6972 21981
rect 8392 21904 8444 21956
rect 3332 21836 3384 21888
rect 5816 21879 5868 21888
rect 5816 21845 5825 21879
rect 5825 21845 5859 21879
rect 5859 21845 5868 21879
rect 5816 21836 5868 21845
rect 6828 21836 6880 21888
rect 7380 21836 7432 21888
rect 8760 21879 8812 21888
rect 8760 21845 8769 21879
rect 8769 21845 8803 21879
rect 8803 21845 8812 21879
rect 8760 21836 8812 21845
rect 9036 21947 9088 21956
rect 9036 21913 9045 21947
rect 9045 21913 9079 21947
rect 9079 21913 9088 21947
rect 9036 21904 9088 21913
rect 10324 21904 10376 21956
rect 10692 22015 10744 22024
rect 10692 21981 10701 22015
rect 10701 21981 10735 22015
rect 10735 21981 10744 22015
rect 10692 21972 10744 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 13544 21904 13596 21956
rect 9312 21879 9364 21888
rect 9312 21845 9321 21879
rect 9321 21845 9355 21879
rect 9355 21845 9364 21879
rect 9312 21836 9364 21845
rect 9680 21879 9732 21888
rect 9680 21845 9689 21879
rect 9689 21845 9723 21879
rect 9723 21845 9732 21879
rect 9680 21836 9732 21845
rect 11152 21836 11204 21888
rect 14280 21972 14332 22024
rect 14648 21972 14700 22024
rect 15108 22040 15160 22092
rect 16856 22040 16908 22092
rect 17500 22040 17552 22092
rect 18052 22040 18104 22092
rect 19800 22108 19852 22160
rect 22100 22108 22152 22160
rect 23112 22108 23164 22160
rect 15200 22015 15252 22024
rect 15200 21981 15209 22015
rect 15209 21981 15243 22015
rect 15243 21981 15252 22015
rect 15200 21972 15252 21981
rect 19616 22040 19668 22092
rect 20076 22040 20128 22092
rect 20720 22040 20772 22092
rect 21456 22040 21508 22092
rect 22652 22040 22704 22092
rect 22744 22040 22796 22092
rect 23940 22083 23992 22092
rect 23940 22049 23949 22083
rect 23949 22049 23983 22083
rect 23983 22049 23992 22083
rect 23940 22040 23992 22049
rect 20260 21972 20312 22024
rect 20352 22015 20404 22024
rect 20352 21981 20361 22015
rect 20361 21981 20395 22015
rect 20395 21981 20404 22015
rect 20352 21972 20404 21981
rect 23572 21972 23624 22024
rect 25688 22108 25740 22160
rect 27252 22176 27304 22228
rect 27896 22176 27948 22228
rect 28448 22176 28500 22228
rect 29276 22219 29328 22228
rect 29276 22185 29285 22219
rect 29285 22185 29319 22219
rect 29319 22185 29328 22219
rect 29276 22176 29328 22185
rect 29644 22176 29696 22228
rect 30012 22176 30064 22228
rect 30288 22108 30340 22160
rect 25136 22083 25188 22092
rect 25136 22049 25145 22083
rect 25145 22049 25179 22083
rect 25179 22049 25188 22083
rect 25136 22040 25188 22049
rect 17684 21904 17736 21956
rect 16212 21836 16264 21888
rect 17592 21836 17644 21888
rect 19156 21836 19208 21888
rect 20628 21904 20680 21956
rect 19432 21836 19484 21888
rect 19616 21836 19668 21888
rect 22744 21836 22796 21888
rect 24400 21836 24452 21888
rect 26056 22040 26108 22092
rect 27528 22083 27580 22092
rect 27528 22049 27537 22083
rect 27537 22049 27571 22083
rect 27571 22049 27580 22083
rect 27528 22040 27580 22049
rect 30564 22176 30616 22228
rect 39672 22176 39724 22228
rect 40224 22176 40276 22228
rect 41696 22176 41748 22228
rect 43536 22176 43588 22228
rect 35072 22108 35124 22160
rect 45008 22108 45060 22160
rect 27344 21972 27396 22024
rect 28816 21972 28868 22024
rect 29828 21972 29880 22024
rect 33324 22040 33376 22092
rect 37004 22083 37056 22092
rect 37004 22049 37013 22083
rect 37013 22049 37047 22083
rect 37047 22049 37056 22083
rect 37004 22040 37056 22049
rect 37188 22040 37240 22092
rect 40408 22040 40460 22092
rect 41604 22083 41656 22092
rect 41604 22049 41613 22083
rect 41613 22049 41647 22083
rect 41647 22049 41656 22083
rect 41604 22040 41656 22049
rect 30932 22015 30984 22024
rect 30932 21981 30941 22015
rect 30941 21981 30975 22015
rect 30975 21981 30984 22015
rect 30932 21972 30984 21981
rect 33048 21972 33100 22024
rect 33416 22015 33468 22024
rect 33416 21981 33425 22015
rect 33425 21981 33459 22015
rect 33459 21981 33468 22015
rect 33416 21972 33468 21981
rect 34520 21972 34572 22024
rect 34980 21972 35032 22024
rect 25964 21904 26016 21956
rect 25320 21836 25372 21888
rect 25412 21836 25464 21888
rect 26332 21904 26384 21956
rect 27068 21904 27120 21956
rect 26240 21836 26292 21888
rect 34796 21904 34848 21956
rect 36084 21904 36136 21956
rect 37096 21947 37148 21956
rect 37096 21913 37105 21947
rect 37105 21913 37139 21947
rect 37139 21913 37148 21947
rect 37096 21904 37148 21913
rect 37832 21972 37884 22024
rect 38844 21972 38896 22024
rect 40684 21972 40736 22024
rect 45836 22040 45888 22092
rect 40132 21904 40184 21956
rect 40408 21904 40460 21956
rect 44364 22015 44416 22024
rect 44364 21981 44373 22015
rect 44373 21981 44407 22015
rect 44407 21981 44416 22015
rect 44364 21972 44416 21981
rect 46480 22176 46532 22228
rect 46020 22108 46072 22160
rect 48504 22040 48556 22092
rect 27620 21836 27672 21888
rect 28908 21879 28960 21888
rect 28908 21845 28917 21879
rect 28917 21845 28951 21879
rect 28951 21845 28960 21879
rect 28908 21836 28960 21845
rect 30012 21836 30064 21888
rect 30288 21836 30340 21888
rect 30748 21836 30800 21888
rect 33048 21836 33100 21888
rect 34336 21879 34388 21888
rect 34336 21845 34345 21879
rect 34345 21845 34379 21879
rect 34379 21845 34388 21879
rect 34336 21836 34388 21845
rect 34428 21836 34480 21888
rect 35624 21836 35676 21888
rect 37188 21836 37240 21888
rect 38752 21836 38804 21888
rect 43260 21879 43312 21888
rect 43260 21845 43269 21879
rect 43269 21845 43303 21879
rect 43303 21845 43312 21879
rect 43260 21836 43312 21845
rect 44180 21904 44232 21956
rect 47860 21972 47912 22024
rect 48688 22015 48740 22024
rect 48688 21981 48697 22015
rect 48697 21981 48731 22015
rect 48731 21981 48740 22015
rect 48688 21972 48740 21981
rect 45284 21904 45336 21956
rect 45468 21904 45520 21956
rect 45376 21879 45428 21888
rect 45376 21845 45385 21879
rect 45385 21845 45419 21879
rect 45419 21845 45428 21879
rect 45376 21836 45428 21845
rect 47400 21879 47452 21888
rect 47400 21845 47409 21879
rect 47409 21845 47443 21879
rect 47443 21845 47452 21879
rect 47400 21836 47452 21845
rect 47860 21836 47912 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 5724 21675 5776 21684
rect 5724 21641 5733 21675
rect 5733 21641 5767 21675
rect 5767 21641 5776 21675
rect 5724 21632 5776 21641
rect 7104 21632 7156 21684
rect 4436 21564 4488 21616
rect 6276 21564 6328 21616
rect 12072 21632 12124 21684
rect 23296 21632 23348 21684
rect 23940 21632 23992 21684
rect 9404 21564 9456 21616
rect 1676 21539 1728 21548
rect 1676 21505 1685 21539
rect 1685 21505 1719 21539
rect 1719 21505 1728 21539
rect 1676 21496 1728 21505
rect 3608 21539 3660 21548
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 5632 21539 5684 21548
rect 5632 21505 5641 21539
rect 5641 21505 5675 21539
rect 5675 21505 5684 21539
rect 5632 21496 5684 21505
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 4160 21471 4212 21480
rect 4160 21437 4169 21471
rect 4169 21437 4203 21471
rect 4203 21437 4212 21471
rect 4160 21428 4212 21437
rect 7104 21428 7156 21480
rect 7564 21428 7616 21480
rect 2504 21360 2556 21412
rect 7012 21360 7064 21412
rect 5448 21292 5500 21344
rect 6552 21335 6604 21344
rect 6552 21301 6561 21335
rect 6561 21301 6595 21335
rect 6595 21301 6604 21335
rect 6552 21292 6604 21301
rect 8024 21471 8076 21480
rect 8024 21437 8033 21471
rect 8033 21437 8067 21471
rect 8067 21437 8076 21471
rect 8024 21428 8076 21437
rect 8392 21428 8444 21480
rect 10324 21496 10376 21548
rect 12256 21564 12308 21616
rect 12716 21496 12768 21548
rect 10508 21428 10560 21480
rect 10968 21471 11020 21480
rect 10968 21437 10977 21471
rect 10977 21437 11011 21471
rect 11011 21437 11020 21471
rect 10968 21428 11020 21437
rect 12256 21471 12308 21480
rect 12256 21437 12265 21471
rect 12265 21437 12299 21471
rect 12299 21437 12308 21471
rect 12256 21428 12308 21437
rect 15108 21607 15160 21616
rect 15108 21573 15117 21607
rect 15117 21573 15151 21607
rect 15151 21573 15160 21607
rect 15108 21564 15160 21573
rect 14464 21496 14516 21548
rect 18420 21564 18472 21616
rect 18880 21564 18932 21616
rect 19064 21564 19116 21616
rect 20628 21564 20680 21616
rect 20996 21564 21048 21616
rect 21088 21607 21140 21616
rect 21088 21573 21097 21607
rect 21097 21573 21131 21607
rect 21131 21573 21140 21607
rect 21088 21564 21140 21573
rect 23664 21607 23716 21616
rect 23664 21573 23673 21607
rect 23673 21573 23707 21607
rect 23707 21573 23716 21607
rect 23664 21564 23716 21573
rect 25044 21632 25096 21684
rect 27528 21632 27580 21684
rect 28356 21632 28408 21684
rect 26056 21564 26108 21616
rect 26148 21607 26200 21616
rect 26148 21573 26157 21607
rect 26157 21573 26191 21607
rect 26191 21573 26200 21607
rect 26148 21564 26200 21573
rect 27896 21564 27948 21616
rect 27988 21564 28040 21616
rect 28724 21607 28776 21616
rect 28724 21573 28733 21607
rect 28733 21573 28767 21607
rect 28767 21573 28776 21607
rect 28724 21564 28776 21573
rect 30932 21632 30984 21684
rect 33048 21632 33100 21684
rect 36544 21632 36596 21684
rect 37096 21632 37148 21684
rect 37832 21632 37884 21684
rect 38292 21632 38344 21684
rect 43260 21632 43312 21684
rect 44088 21675 44140 21684
rect 44088 21641 44097 21675
rect 44097 21641 44131 21675
rect 44131 21641 44140 21675
rect 44088 21632 44140 21641
rect 44916 21632 44968 21684
rect 45284 21632 45336 21684
rect 45652 21632 45704 21684
rect 47032 21675 47084 21684
rect 47032 21641 47041 21675
rect 47041 21641 47075 21675
rect 47075 21641 47084 21675
rect 47032 21632 47084 21641
rect 47768 21632 47820 21684
rect 15936 21539 15988 21548
rect 15936 21505 15945 21539
rect 15945 21505 15979 21539
rect 15979 21505 15988 21539
rect 15936 21496 15988 21505
rect 16488 21496 16540 21548
rect 17132 21496 17184 21548
rect 9588 21360 9640 21412
rect 8668 21292 8720 21344
rect 13544 21428 13596 21480
rect 13728 21428 13780 21480
rect 14832 21428 14884 21480
rect 15108 21428 15160 21480
rect 15752 21428 15804 21480
rect 16120 21428 16172 21480
rect 14372 21360 14424 21412
rect 16764 21428 16816 21480
rect 17776 21496 17828 21548
rect 20260 21496 20312 21548
rect 17316 21471 17368 21480
rect 17316 21437 17325 21471
rect 17325 21437 17359 21471
rect 17359 21437 17368 21471
rect 17316 21428 17368 21437
rect 17500 21428 17552 21480
rect 13544 21292 13596 21344
rect 14924 21292 14976 21344
rect 15384 21292 15436 21344
rect 17960 21360 18012 21412
rect 16304 21292 16356 21344
rect 19064 21428 19116 21480
rect 21640 21428 21692 21480
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 25320 21496 25372 21548
rect 27436 21496 27488 21548
rect 27528 21496 27580 21548
rect 28080 21496 28132 21548
rect 28448 21539 28500 21548
rect 28448 21505 28457 21539
rect 28457 21505 28491 21539
rect 28491 21505 28500 21539
rect 28448 21496 28500 21505
rect 29736 21496 29788 21548
rect 30656 21496 30708 21548
rect 30748 21496 30800 21548
rect 31116 21539 31168 21548
rect 31116 21505 31125 21539
rect 31125 21505 31159 21539
rect 31159 21505 31168 21539
rect 31116 21496 31168 21505
rect 31760 21607 31812 21616
rect 31760 21573 31769 21607
rect 31769 21573 31803 21607
rect 31803 21573 31812 21607
rect 31760 21564 31812 21573
rect 32588 21564 32640 21616
rect 32772 21564 32824 21616
rect 32864 21564 32916 21616
rect 33324 21496 33376 21548
rect 34428 21496 34480 21548
rect 35624 21496 35676 21548
rect 35900 21496 35952 21548
rect 37740 21539 37792 21548
rect 37740 21505 37749 21539
rect 37749 21505 37783 21539
rect 37783 21505 37792 21539
rect 37740 21496 37792 21505
rect 38752 21539 38804 21548
rect 38752 21505 38761 21539
rect 38761 21505 38795 21539
rect 38795 21505 38804 21539
rect 38752 21496 38804 21505
rect 39488 21496 39540 21548
rect 39856 21539 39908 21548
rect 39856 21505 39865 21539
rect 39865 21505 39899 21539
rect 39899 21505 39908 21539
rect 39856 21496 39908 21505
rect 22376 21428 22428 21480
rect 23388 21471 23440 21480
rect 23388 21437 23397 21471
rect 23397 21437 23431 21471
rect 23431 21437 23440 21471
rect 23388 21428 23440 21437
rect 23664 21428 23716 21480
rect 27712 21428 27764 21480
rect 22284 21360 22336 21412
rect 23112 21360 23164 21412
rect 23296 21360 23348 21412
rect 19708 21292 19760 21344
rect 20260 21292 20312 21344
rect 21272 21292 21324 21344
rect 21640 21292 21692 21344
rect 22008 21292 22060 21344
rect 24676 21360 24728 21412
rect 25136 21403 25188 21412
rect 25136 21369 25145 21403
rect 25145 21369 25179 21403
rect 25179 21369 25188 21403
rect 25136 21360 25188 21369
rect 24124 21292 24176 21344
rect 24400 21292 24452 21344
rect 26516 21360 26568 21412
rect 26608 21360 26660 21412
rect 27068 21360 27120 21412
rect 27344 21360 27396 21412
rect 27896 21428 27948 21480
rect 29920 21428 29972 21480
rect 34980 21428 35032 21480
rect 37004 21428 37056 21480
rect 27988 21360 28040 21412
rect 30104 21360 30156 21412
rect 25688 21335 25740 21344
rect 25688 21301 25697 21335
rect 25697 21301 25731 21335
rect 25731 21301 25740 21335
rect 25688 21292 25740 21301
rect 27252 21335 27304 21344
rect 27252 21301 27261 21335
rect 27261 21301 27295 21335
rect 27295 21301 27304 21335
rect 27252 21292 27304 21301
rect 27528 21292 27580 21344
rect 31944 21360 31996 21412
rect 41788 21496 41840 21548
rect 42524 21496 42576 21548
rect 43628 21496 43680 21548
rect 43996 21496 44048 21548
rect 47216 21539 47268 21548
rect 47216 21505 47225 21539
rect 47225 21505 47259 21539
rect 47259 21505 47268 21539
rect 47216 21496 47268 21505
rect 47768 21496 47820 21548
rect 44456 21428 44508 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 31852 21335 31904 21344
rect 31852 21301 31861 21335
rect 31861 21301 31895 21335
rect 31895 21301 31904 21335
rect 31852 21292 31904 21301
rect 32128 21292 32180 21344
rect 32588 21292 32640 21344
rect 33508 21292 33560 21344
rect 35256 21292 35308 21344
rect 35992 21292 36044 21344
rect 36544 21292 36596 21344
rect 37004 21335 37056 21344
rect 37004 21301 37013 21335
rect 37013 21301 37047 21335
rect 37047 21301 37056 21335
rect 37004 21292 37056 21301
rect 38200 21292 38252 21344
rect 39488 21292 39540 21344
rect 40224 21292 40276 21344
rect 41328 21360 41380 21412
rect 42800 21335 42852 21344
rect 42800 21301 42809 21335
rect 42809 21301 42843 21335
rect 42843 21301 42852 21335
rect 42800 21292 42852 21301
rect 43536 21335 43588 21344
rect 43536 21301 43545 21335
rect 43545 21301 43579 21335
rect 43579 21301 43588 21335
rect 43536 21292 43588 21301
rect 44732 21335 44784 21344
rect 44732 21301 44741 21335
rect 44741 21301 44775 21335
rect 44775 21301 44784 21335
rect 44732 21292 44784 21301
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 3608 21088 3660 21140
rect 3792 21088 3844 21140
rect 7564 21020 7616 21072
rect 9956 21020 10008 21072
rect 2044 20995 2096 21004
rect 2044 20961 2053 20995
rect 2053 20961 2087 20995
rect 2087 20961 2096 20995
rect 2044 20952 2096 20961
rect 3792 20952 3844 21004
rect 6828 20952 6880 21004
rect 2228 20884 2280 20936
rect 4068 20927 4120 20936
rect 4068 20893 4077 20927
rect 4077 20893 4111 20927
rect 4111 20893 4120 20927
rect 4068 20884 4120 20893
rect 6184 20927 6236 20936
rect 6184 20893 6193 20927
rect 6193 20893 6227 20927
rect 6227 20893 6236 20927
rect 6184 20884 6236 20893
rect 7564 20884 7616 20936
rect 7840 20952 7892 21004
rect 9404 20952 9456 21004
rect 10048 20995 10100 21004
rect 10048 20961 10057 20995
rect 10057 20961 10091 20995
rect 10091 20961 10100 20995
rect 10048 20952 10100 20961
rect 14372 21088 14424 21140
rect 15108 21088 15160 21140
rect 15752 21131 15804 21140
rect 15752 21097 15761 21131
rect 15761 21097 15795 21131
rect 15795 21097 15804 21131
rect 15752 21088 15804 21097
rect 10508 21020 10560 21072
rect 11980 20927 12032 20936
rect 2596 20816 2648 20868
rect 5816 20816 5868 20868
rect 6460 20859 6512 20868
rect 6460 20825 6469 20859
rect 6469 20825 6503 20859
rect 6503 20825 6512 20859
rect 6460 20816 6512 20825
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 12808 20995 12860 21004
rect 12808 20961 12817 20995
rect 12817 20961 12851 20995
rect 12851 20961 12860 20995
rect 12808 20952 12860 20961
rect 16580 21088 16632 21140
rect 14648 20952 14700 21004
rect 14372 20884 14424 20936
rect 10508 20816 10560 20868
rect 5540 20748 5592 20800
rect 5724 20791 5776 20800
rect 5724 20757 5733 20791
rect 5733 20757 5767 20791
rect 5767 20757 5776 20791
rect 5724 20748 5776 20757
rect 5908 20791 5960 20800
rect 5908 20757 5917 20791
rect 5917 20757 5951 20791
rect 5951 20757 5960 20791
rect 5908 20748 5960 20757
rect 7840 20748 7892 20800
rect 10140 20748 10192 20800
rect 11244 20748 11296 20800
rect 11336 20791 11388 20800
rect 11336 20757 11345 20791
rect 11345 20757 11379 20791
rect 11379 20757 11388 20791
rect 11336 20748 11388 20757
rect 11520 20748 11572 20800
rect 11704 20791 11756 20800
rect 11704 20757 11713 20791
rect 11713 20757 11747 20791
rect 11747 20757 11756 20791
rect 11704 20748 11756 20757
rect 14648 20816 14700 20868
rect 15200 20952 15252 21004
rect 16396 21020 16448 21072
rect 16304 20995 16356 21004
rect 16304 20961 16313 20995
rect 16313 20961 16347 20995
rect 16347 20961 16356 20995
rect 16304 20952 16356 20961
rect 20168 21088 20220 21140
rect 17316 21020 17368 21072
rect 17868 21020 17920 21072
rect 16120 20884 16172 20936
rect 16580 20884 16632 20936
rect 17500 20995 17552 21004
rect 17500 20961 17509 20995
rect 17509 20961 17543 20995
rect 17543 20961 17552 20995
rect 17500 20952 17552 20961
rect 18604 20995 18656 21004
rect 18604 20961 18613 20995
rect 18613 20961 18647 20995
rect 18647 20961 18656 20995
rect 18604 20952 18656 20961
rect 21088 21020 21140 21072
rect 23480 21088 23532 21140
rect 23572 21088 23624 21140
rect 27252 21088 27304 21140
rect 27712 21131 27764 21140
rect 27712 21097 27721 21131
rect 27721 21097 27755 21131
rect 27755 21097 27764 21131
rect 27712 21088 27764 21097
rect 28448 21088 28500 21140
rect 29276 21088 29328 21140
rect 30748 21088 30800 21140
rect 31484 21088 31536 21140
rect 25412 21020 25464 21072
rect 27436 21020 27488 21072
rect 28724 21020 28776 21072
rect 28816 21063 28868 21072
rect 28816 21029 28825 21063
rect 28825 21029 28859 21063
rect 28859 21029 28868 21063
rect 28816 21020 28868 21029
rect 14832 20816 14884 20868
rect 15660 20816 15712 20868
rect 15844 20816 15896 20868
rect 16856 20816 16908 20868
rect 17408 20884 17460 20936
rect 18420 20884 18472 20936
rect 18972 20884 19024 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 19064 20816 19116 20868
rect 19984 20816 20036 20868
rect 20996 20816 21048 20868
rect 21364 20816 21416 20868
rect 23572 20952 23624 21004
rect 22560 20884 22612 20936
rect 23204 20884 23256 20936
rect 16120 20791 16172 20800
rect 16120 20757 16129 20791
rect 16129 20757 16163 20791
rect 16163 20757 16172 20791
rect 16120 20748 16172 20757
rect 16948 20791 17000 20800
rect 16948 20757 16957 20791
rect 16957 20757 16991 20791
rect 16991 20757 17000 20791
rect 16948 20748 17000 20757
rect 17408 20791 17460 20800
rect 17408 20757 17417 20791
rect 17417 20757 17451 20791
rect 17451 20757 17460 20791
rect 17408 20748 17460 20757
rect 18880 20748 18932 20800
rect 20720 20748 20772 20800
rect 21272 20748 21324 20800
rect 21824 20791 21876 20800
rect 21824 20757 21833 20791
rect 21833 20757 21867 20791
rect 21867 20757 21876 20791
rect 21824 20748 21876 20757
rect 23572 20816 23624 20868
rect 22560 20748 22612 20800
rect 22744 20748 22796 20800
rect 23204 20748 23256 20800
rect 23480 20748 23532 20800
rect 23940 20952 23992 21004
rect 25136 20952 25188 21004
rect 25228 20995 25280 21004
rect 25228 20961 25237 20995
rect 25237 20961 25271 20995
rect 25271 20961 25280 20995
rect 25228 20952 25280 20961
rect 25320 20952 25372 21004
rect 24124 20884 24176 20936
rect 25964 20927 26016 20936
rect 25964 20893 25973 20927
rect 25973 20893 26007 20927
rect 26007 20893 26016 20927
rect 25964 20884 26016 20893
rect 27344 20884 27396 20936
rect 27712 20884 27764 20936
rect 27988 20884 28040 20936
rect 31852 21088 31904 21140
rect 32864 21088 32916 21140
rect 34704 21088 34756 21140
rect 32496 21020 32548 21072
rect 32128 20952 32180 21004
rect 32588 20952 32640 21004
rect 37188 21020 37240 21072
rect 38844 21131 38896 21140
rect 38844 21097 38853 21131
rect 38853 21097 38887 21131
rect 38887 21097 38896 21131
rect 38844 21088 38896 21097
rect 40684 21131 40736 21140
rect 40684 21097 40693 21131
rect 40693 21097 40727 21131
rect 40727 21097 40736 21131
rect 40684 21088 40736 21097
rect 41972 21088 42024 21140
rect 44088 21088 44140 21140
rect 48596 21088 48648 21140
rect 49332 21131 49384 21140
rect 49332 21097 49341 21131
rect 49341 21097 49375 21131
rect 49375 21097 49384 21131
rect 49332 21088 49384 21097
rect 26148 20816 26200 20868
rect 26240 20859 26292 20868
rect 26240 20825 26249 20859
rect 26249 20825 26283 20859
rect 26283 20825 26292 20859
rect 26240 20816 26292 20825
rect 27804 20816 27856 20868
rect 24676 20791 24728 20800
rect 24676 20757 24685 20791
rect 24685 20757 24719 20791
rect 24719 20757 24728 20791
rect 24676 20748 24728 20757
rect 27528 20748 27580 20800
rect 28080 20748 28132 20800
rect 28816 20748 28868 20800
rect 29276 20791 29328 20800
rect 29276 20757 29285 20791
rect 29285 20757 29319 20791
rect 29319 20757 29328 20791
rect 29276 20748 29328 20757
rect 30104 20816 30156 20868
rect 30656 20859 30708 20868
rect 30656 20825 30665 20859
rect 30665 20825 30699 20859
rect 30699 20825 30708 20859
rect 31668 20927 31720 20936
rect 31668 20893 31677 20927
rect 31677 20893 31711 20927
rect 31711 20893 31720 20927
rect 31668 20884 31720 20893
rect 31944 20884 31996 20936
rect 33508 20927 33560 20936
rect 33508 20893 33517 20927
rect 33517 20893 33551 20927
rect 33551 20893 33560 20927
rect 33508 20884 33560 20893
rect 35440 20884 35492 20936
rect 30656 20816 30708 20825
rect 31116 20748 31168 20800
rect 31760 20748 31812 20800
rect 32220 20748 32272 20800
rect 36176 20952 36228 21004
rect 36268 20884 36320 20936
rect 38200 20927 38252 20936
rect 38200 20893 38209 20927
rect 38209 20893 38243 20927
rect 38243 20893 38252 20927
rect 38200 20884 38252 20893
rect 39212 20884 39264 20936
rect 39488 20927 39540 20936
rect 39488 20893 39497 20927
rect 39497 20893 39531 20927
rect 39531 20893 39540 20927
rect 39488 20884 39540 20893
rect 40040 20927 40092 20936
rect 40040 20893 40049 20927
rect 40049 20893 40083 20927
rect 40083 20893 40092 20927
rect 40040 20884 40092 20893
rect 42064 20884 42116 20936
rect 43444 20884 43496 20936
rect 48596 20884 48648 20936
rect 41328 20816 41380 20868
rect 42708 20859 42760 20868
rect 42708 20825 42717 20859
rect 42717 20825 42751 20859
rect 42751 20825 42760 20859
rect 42708 20816 42760 20825
rect 43904 20816 43956 20868
rect 34152 20791 34204 20800
rect 34152 20757 34161 20791
rect 34161 20757 34195 20791
rect 34195 20757 34204 20791
rect 34152 20748 34204 20757
rect 37740 20791 37792 20800
rect 37740 20757 37749 20791
rect 37749 20757 37783 20791
rect 37783 20757 37792 20791
rect 37740 20748 37792 20757
rect 39304 20791 39356 20800
rect 39304 20757 39313 20791
rect 39313 20757 39347 20791
rect 39347 20757 39356 20791
rect 39304 20748 39356 20757
rect 42064 20791 42116 20800
rect 42064 20757 42073 20791
rect 42073 20757 42107 20791
rect 42107 20757 42116 20791
rect 42064 20748 42116 20757
rect 43352 20791 43404 20800
rect 43352 20757 43361 20791
rect 43361 20757 43395 20791
rect 43395 20757 43404 20791
rect 43352 20748 43404 20757
rect 47768 20791 47820 20800
rect 47768 20757 47777 20791
rect 47777 20757 47811 20791
rect 47811 20757 47820 20791
rect 47768 20748 47820 20757
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 3792 20544 3844 20596
rect 10692 20544 10744 20596
rect 11060 20544 11112 20596
rect 12348 20587 12400 20596
rect 12348 20553 12357 20587
rect 12357 20553 12391 20587
rect 12391 20553 12400 20587
rect 12348 20544 12400 20553
rect 4252 20476 4304 20528
rect 1124 20408 1176 20460
rect 3976 20408 4028 20460
rect 5632 20408 5684 20460
rect 1400 20340 1452 20392
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 5264 20340 5316 20392
rect 10876 20476 10928 20528
rect 6920 20408 6972 20460
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 8668 20383 8720 20392
rect 8668 20349 8677 20383
rect 8677 20349 8711 20383
rect 8711 20349 8720 20383
rect 8668 20340 8720 20349
rect 10508 20408 10560 20460
rect 11796 20408 11848 20460
rect 12900 20476 12952 20528
rect 14096 20476 14148 20528
rect 14464 20476 14516 20528
rect 16856 20587 16908 20596
rect 16856 20553 16865 20587
rect 16865 20553 16899 20587
rect 16899 20553 16908 20587
rect 16856 20544 16908 20553
rect 17316 20544 17368 20596
rect 17592 20587 17644 20596
rect 17592 20553 17601 20587
rect 17601 20553 17635 20587
rect 17635 20553 17644 20587
rect 17592 20544 17644 20553
rect 16396 20476 16448 20528
rect 18144 20476 18196 20528
rect 18328 20476 18380 20528
rect 19432 20544 19484 20596
rect 6552 20272 6604 20324
rect 6736 20272 6788 20324
rect 10784 20340 10836 20392
rect 11060 20340 11112 20392
rect 11428 20340 11480 20392
rect 15476 20408 15528 20460
rect 16304 20408 16356 20460
rect 17224 20408 17276 20460
rect 17592 20408 17644 20460
rect 18604 20408 18656 20460
rect 18972 20451 19024 20460
rect 18972 20417 18981 20451
rect 18981 20417 19015 20451
rect 19015 20417 19024 20451
rect 18972 20408 19024 20417
rect 19432 20408 19484 20460
rect 20904 20544 20956 20596
rect 22192 20544 22244 20596
rect 23572 20587 23624 20596
rect 23572 20553 23581 20587
rect 23581 20553 23615 20587
rect 23615 20553 23624 20587
rect 23572 20544 23624 20553
rect 24124 20587 24176 20596
rect 24124 20553 24133 20587
rect 24133 20553 24167 20587
rect 24167 20553 24176 20587
rect 24124 20544 24176 20553
rect 21640 20476 21692 20528
rect 21824 20476 21876 20528
rect 21272 20408 21324 20460
rect 23940 20476 23992 20528
rect 25136 20476 25188 20528
rect 26608 20476 26660 20528
rect 26792 20587 26844 20596
rect 26792 20553 26801 20587
rect 26801 20553 26835 20587
rect 26835 20553 26844 20587
rect 26792 20544 26844 20553
rect 26976 20476 27028 20528
rect 27160 20476 27212 20528
rect 27436 20544 27488 20596
rect 34152 20544 34204 20596
rect 34612 20587 34664 20596
rect 34612 20553 34621 20587
rect 34621 20553 34655 20587
rect 34655 20553 34664 20587
rect 34612 20544 34664 20553
rect 35900 20544 35952 20596
rect 36728 20544 36780 20596
rect 27804 20476 27856 20528
rect 29736 20476 29788 20528
rect 31760 20519 31812 20528
rect 31760 20485 31769 20519
rect 31769 20485 31803 20519
rect 31803 20485 31812 20519
rect 31760 20476 31812 20485
rect 22008 20451 22060 20460
rect 22008 20417 22017 20451
rect 22017 20417 22051 20451
rect 22051 20417 22060 20451
rect 22008 20408 22060 20417
rect 22192 20408 22244 20460
rect 9956 20272 10008 20324
rect 5724 20204 5776 20256
rect 5908 20204 5960 20256
rect 8116 20204 8168 20256
rect 8392 20247 8444 20256
rect 8392 20213 8401 20247
rect 8401 20213 8435 20247
rect 8435 20213 8444 20247
rect 8392 20204 8444 20213
rect 8576 20204 8628 20256
rect 9312 20204 9364 20256
rect 9680 20204 9732 20256
rect 10416 20247 10468 20256
rect 10416 20213 10425 20247
rect 10425 20213 10459 20247
rect 10459 20213 10468 20247
rect 10416 20204 10468 20213
rect 12992 20383 13044 20392
rect 12992 20349 13001 20383
rect 13001 20349 13035 20383
rect 13035 20349 13044 20383
rect 12992 20340 13044 20349
rect 13544 20383 13596 20392
rect 13544 20349 13553 20383
rect 13553 20349 13587 20383
rect 13587 20349 13596 20383
rect 13544 20340 13596 20349
rect 16488 20340 16540 20392
rect 16396 20272 16448 20324
rect 16948 20272 17000 20324
rect 17408 20272 17460 20324
rect 17960 20340 18012 20392
rect 18788 20340 18840 20392
rect 19064 20383 19116 20392
rect 19064 20349 19073 20383
rect 19073 20349 19107 20383
rect 19107 20349 19116 20383
rect 19064 20340 19116 20349
rect 20536 20340 20588 20392
rect 21456 20383 21508 20392
rect 21456 20349 21465 20383
rect 21465 20349 21499 20383
rect 21499 20349 21508 20383
rect 21456 20340 21508 20349
rect 22468 20340 22520 20392
rect 22744 20340 22796 20392
rect 23572 20408 23624 20460
rect 26516 20451 26568 20460
rect 26516 20417 26525 20451
rect 26525 20417 26559 20451
rect 26559 20417 26568 20451
rect 26516 20408 26568 20417
rect 27436 20340 27488 20392
rect 17868 20272 17920 20324
rect 18144 20272 18196 20324
rect 18972 20272 19024 20324
rect 15660 20247 15712 20256
rect 15660 20213 15669 20247
rect 15669 20213 15703 20247
rect 15703 20213 15712 20247
rect 15660 20204 15712 20213
rect 16488 20204 16540 20256
rect 17684 20204 17736 20256
rect 18512 20247 18564 20256
rect 18512 20213 18521 20247
rect 18521 20213 18555 20247
rect 18555 20213 18564 20247
rect 18512 20204 18564 20213
rect 19156 20204 19208 20256
rect 21640 20272 21692 20324
rect 23388 20272 23440 20324
rect 27252 20272 27304 20324
rect 22836 20204 22888 20256
rect 22928 20204 22980 20256
rect 23664 20204 23716 20256
rect 24860 20204 24912 20256
rect 25412 20204 25464 20256
rect 27160 20247 27212 20256
rect 27160 20213 27169 20247
rect 27169 20213 27203 20247
rect 27203 20213 27212 20247
rect 27160 20204 27212 20213
rect 28448 20451 28500 20460
rect 28448 20417 28457 20451
rect 28457 20417 28491 20451
rect 28491 20417 28500 20451
rect 28448 20408 28500 20417
rect 31024 20451 31076 20460
rect 31024 20417 31033 20451
rect 31033 20417 31067 20451
rect 31067 20417 31076 20451
rect 31024 20408 31076 20417
rect 27804 20383 27856 20392
rect 27804 20349 27813 20383
rect 27813 20349 27847 20383
rect 27847 20349 27856 20383
rect 27804 20340 27856 20349
rect 30656 20315 30708 20324
rect 30656 20281 30665 20315
rect 30665 20281 30699 20315
rect 30699 20281 30708 20315
rect 30656 20272 30708 20281
rect 31116 20383 31168 20392
rect 31116 20349 31125 20383
rect 31125 20349 31159 20383
rect 31159 20349 31168 20383
rect 31116 20340 31168 20349
rect 32312 20451 32364 20460
rect 32312 20417 32321 20451
rect 32321 20417 32355 20451
rect 32355 20417 32364 20451
rect 32312 20408 32364 20417
rect 33416 20451 33468 20460
rect 33416 20417 33425 20451
rect 33425 20417 33459 20451
rect 33459 20417 33468 20451
rect 33416 20408 33468 20417
rect 35532 20408 35584 20460
rect 35992 20451 36044 20460
rect 35992 20417 36001 20451
rect 36001 20417 36035 20451
rect 36035 20417 36044 20451
rect 35992 20408 36044 20417
rect 37372 20408 37424 20460
rect 31300 20383 31352 20392
rect 31300 20349 31309 20383
rect 31309 20349 31343 20383
rect 31343 20349 31352 20383
rect 31300 20340 31352 20349
rect 34060 20383 34112 20392
rect 34060 20349 34069 20383
rect 34069 20349 34103 20383
rect 34103 20349 34112 20383
rect 34060 20340 34112 20349
rect 34336 20383 34388 20392
rect 34336 20349 34345 20383
rect 34345 20349 34379 20383
rect 34379 20349 34388 20383
rect 34336 20340 34388 20349
rect 36636 20340 36688 20392
rect 39028 20451 39080 20460
rect 39028 20417 39037 20451
rect 39037 20417 39071 20451
rect 39071 20417 39080 20451
rect 39028 20408 39080 20417
rect 41512 20476 41564 20528
rect 43444 20587 43496 20596
rect 43444 20553 43453 20587
rect 43453 20553 43487 20587
rect 43487 20553 43496 20587
rect 43444 20544 43496 20553
rect 48872 20544 48924 20596
rect 44548 20476 44600 20528
rect 49240 20519 49292 20528
rect 49240 20485 49249 20519
rect 49249 20485 49283 20519
rect 49283 20485 49292 20519
rect 49240 20476 49292 20485
rect 40316 20451 40368 20460
rect 40316 20417 40325 20451
rect 40325 20417 40359 20451
rect 40359 20417 40368 20451
rect 40316 20408 40368 20417
rect 41236 20451 41288 20460
rect 41236 20417 41245 20451
rect 41245 20417 41279 20451
rect 41279 20417 41288 20451
rect 41236 20408 41288 20417
rect 39488 20340 39540 20392
rect 41420 20340 41472 20392
rect 29276 20204 29328 20256
rect 29368 20204 29420 20256
rect 31392 20204 31444 20256
rect 31944 20247 31996 20256
rect 31944 20213 31953 20247
rect 31953 20213 31987 20247
rect 31987 20213 31996 20247
rect 31944 20204 31996 20213
rect 32220 20204 32272 20256
rect 33048 20204 33100 20256
rect 42708 20272 42760 20324
rect 37004 20247 37056 20256
rect 37004 20213 37013 20247
rect 37013 20213 37047 20247
rect 37047 20213 37056 20247
rect 37004 20204 37056 20213
rect 40592 20204 40644 20256
rect 40868 20204 40920 20256
rect 43628 20247 43680 20256
rect 43628 20213 43637 20247
rect 43637 20213 43671 20247
rect 43671 20213 43680 20247
rect 43628 20204 43680 20213
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 3792 20000 3844 20052
rect 1492 19864 1544 19916
rect 8576 20000 8628 20052
rect 9036 20043 9088 20052
rect 9036 20009 9045 20043
rect 9045 20009 9079 20043
rect 9079 20009 9088 20043
rect 9036 20000 9088 20009
rect 9404 20000 9456 20052
rect 8116 19932 8168 19984
rect 1032 19796 1084 19848
rect 3424 19796 3476 19848
rect 4436 19796 4488 19848
rect 6184 19864 6236 19916
rect 6552 19864 6604 19916
rect 8668 19864 8720 19916
rect 13176 19907 13228 19916
rect 13176 19873 13185 19907
rect 13185 19873 13219 19907
rect 13219 19873 13228 19907
rect 13176 19864 13228 19873
rect 14096 19932 14148 19984
rect 14280 19932 14332 19984
rect 16856 20000 16908 20052
rect 17592 20000 17644 20052
rect 17776 20000 17828 20052
rect 19156 20000 19208 20052
rect 19248 20000 19300 20052
rect 13452 19864 13504 19916
rect 15292 19864 15344 19916
rect 15660 19864 15712 19916
rect 16764 19864 16816 19916
rect 17684 19932 17736 19984
rect 20628 20000 20680 20052
rect 20720 20000 20772 20052
rect 22008 20000 22060 20052
rect 24952 20000 25004 20052
rect 22284 19975 22336 19984
rect 22284 19941 22293 19975
rect 22293 19941 22327 19975
rect 22327 19941 22336 19975
rect 22284 19932 22336 19941
rect 23112 19932 23164 19984
rect 27160 20000 27212 20052
rect 27712 20000 27764 20052
rect 28448 20000 28500 20052
rect 29552 20000 29604 20052
rect 31392 20000 31444 20052
rect 31944 20000 31996 20052
rect 32588 20000 32640 20052
rect 35532 20043 35584 20052
rect 35532 20009 35541 20043
rect 35541 20009 35575 20043
rect 35575 20009 35584 20043
rect 35532 20000 35584 20009
rect 40040 20000 40092 20052
rect 3700 19728 3752 19780
rect 4160 19728 4212 19780
rect 9220 19796 9272 19848
rect 9588 19796 9640 19848
rect 11704 19796 11756 19848
rect 4804 19728 4856 19780
rect 3424 19703 3476 19712
rect 3424 19669 3433 19703
rect 3433 19669 3467 19703
rect 3467 19669 3476 19703
rect 3424 19660 3476 19669
rect 4252 19660 4304 19712
rect 6828 19728 6880 19780
rect 7104 19771 7156 19780
rect 7104 19737 7113 19771
rect 7113 19737 7147 19771
rect 7147 19737 7156 19771
rect 7104 19728 7156 19737
rect 5632 19660 5684 19712
rect 6184 19660 6236 19712
rect 6460 19660 6512 19712
rect 6736 19660 6788 19712
rect 8668 19728 8720 19780
rect 10324 19771 10376 19780
rect 10324 19737 10333 19771
rect 10333 19737 10367 19771
rect 10367 19737 10376 19771
rect 10324 19728 10376 19737
rect 7748 19660 7800 19712
rect 9128 19660 9180 19712
rect 10784 19728 10836 19780
rect 11888 19728 11940 19780
rect 12808 19728 12860 19780
rect 13820 19839 13872 19848
rect 13820 19805 13829 19839
rect 13829 19805 13863 19839
rect 13863 19805 13872 19839
rect 13820 19796 13872 19805
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 16948 19796 17000 19848
rect 14648 19771 14700 19780
rect 11336 19660 11388 19712
rect 12072 19660 12124 19712
rect 13452 19660 13504 19712
rect 14648 19737 14657 19771
rect 14657 19737 14691 19771
rect 14691 19737 14700 19771
rect 14648 19728 14700 19737
rect 13728 19660 13780 19712
rect 14464 19660 14516 19712
rect 15476 19660 15528 19712
rect 15660 19660 15712 19712
rect 17868 19864 17920 19916
rect 19064 19864 19116 19916
rect 19524 19864 19576 19916
rect 20076 19864 20128 19916
rect 17316 19839 17368 19848
rect 17316 19805 17325 19839
rect 17325 19805 17359 19839
rect 17359 19805 17368 19839
rect 17316 19796 17368 19805
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 20260 19839 20312 19848
rect 20260 19805 20269 19839
rect 20269 19805 20303 19839
rect 20303 19805 20312 19839
rect 20260 19796 20312 19805
rect 17776 19728 17828 19780
rect 19800 19728 19852 19780
rect 20536 19771 20588 19780
rect 20536 19737 20545 19771
rect 20545 19737 20579 19771
rect 20579 19737 20588 19771
rect 20536 19728 20588 19737
rect 20996 19728 21048 19780
rect 17408 19660 17460 19712
rect 18512 19703 18564 19712
rect 18512 19669 18521 19703
rect 18521 19669 18555 19703
rect 18555 19669 18564 19703
rect 18512 19660 18564 19669
rect 21180 19660 21232 19712
rect 22376 19660 22428 19712
rect 25228 19907 25280 19916
rect 25228 19873 25237 19907
rect 25237 19873 25271 19907
rect 25271 19873 25280 19907
rect 25228 19864 25280 19873
rect 33140 19932 33192 19984
rect 40960 19932 41012 19984
rect 41236 20000 41288 20052
rect 42156 20000 42208 20052
rect 46756 19932 46808 19984
rect 29828 19864 29880 19916
rect 30288 19907 30340 19916
rect 30288 19873 30297 19907
rect 30297 19873 30331 19907
rect 30331 19873 30340 19907
rect 30288 19864 30340 19873
rect 31024 19864 31076 19916
rect 25320 19796 25372 19848
rect 25780 19796 25832 19848
rect 30104 19796 30156 19848
rect 32220 19796 32272 19848
rect 34060 19864 34112 19916
rect 23848 19660 23900 19712
rect 24308 19660 24360 19712
rect 24676 19703 24728 19712
rect 24676 19669 24685 19703
rect 24685 19669 24719 19703
rect 24719 19669 24728 19703
rect 24676 19660 24728 19669
rect 25044 19703 25096 19712
rect 25044 19669 25053 19703
rect 25053 19669 25087 19703
rect 25087 19669 25096 19703
rect 25044 19660 25096 19669
rect 26608 19728 26660 19780
rect 27436 19728 27488 19780
rect 27160 19660 27212 19712
rect 30472 19728 30524 19780
rect 30564 19728 30616 19780
rect 33048 19728 33100 19780
rect 46664 19864 46716 19916
rect 34428 19796 34480 19848
rect 29368 19660 29420 19712
rect 29828 19660 29880 19712
rect 30196 19703 30248 19712
rect 30196 19669 30205 19703
rect 30205 19669 30239 19703
rect 30239 19669 30248 19703
rect 30196 19660 30248 19669
rect 30932 19660 30984 19712
rect 32128 19660 32180 19712
rect 32220 19660 32272 19712
rect 37096 19839 37148 19848
rect 37096 19805 37105 19839
rect 37105 19805 37139 19839
rect 37139 19805 37148 19839
rect 37096 19796 37148 19805
rect 37004 19728 37056 19780
rect 39396 19796 39448 19848
rect 40868 19839 40920 19848
rect 40868 19805 40877 19839
rect 40877 19805 40911 19839
rect 40911 19805 40920 19839
rect 40868 19796 40920 19805
rect 41696 19839 41748 19848
rect 41696 19805 41705 19839
rect 41705 19805 41739 19839
rect 41739 19805 41748 19839
rect 41696 19796 41748 19805
rect 37648 19728 37700 19780
rect 38568 19728 38620 19780
rect 40592 19728 40644 19780
rect 34060 19703 34112 19712
rect 34060 19669 34069 19703
rect 34069 19669 34103 19703
rect 34103 19669 34112 19703
rect 34060 19660 34112 19669
rect 35164 19660 35216 19712
rect 35992 19660 36044 19712
rect 37556 19660 37608 19712
rect 38660 19660 38712 19712
rect 40960 19703 41012 19712
rect 40960 19669 40969 19703
rect 40969 19669 41003 19703
rect 41003 19669 41012 19703
rect 40960 19660 41012 19669
rect 41604 19660 41656 19712
rect 42524 19703 42576 19712
rect 42524 19669 42533 19703
rect 42533 19669 42567 19703
rect 42567 19669 42576 19703
rect 42524 19660 42576 19669
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 664 19388 716 19440
rect 5724 19499 5776 19508
rect 5724 19465 5733 19499
rect 5733 19465 5767 19499
rect 5767 19465 5776 19499
rect 5724 19456 5776 19465
rect 6184 19456 6236 19508
rect 6736 19456 6788 19508
rect 7196 19456 7248 19508
rect 7656 19456 7708 19508
rect 9128 19456 9180 19508
rect 3700 19388 3752 19440
rect 3976 19388 4028 19440
rect 4344 19431 4396 19440
rect 4344 19397 4353 19431
rect 4353 19397 4387 19431
rect 4387 19397 4396 19431
rect 4344 19388 4396 19397
rect 2136 19320 2188 19372
rect 4620 19320 4672 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 2872 19252 2924 19304
rect 6368 19388 6420 19440
rect 7564 19388 7616 19440
rect 9496 19456 9548 19508
rect 10600 19456 10652 19508
rect 10692 19456 10744 19508
rect 2136 19116 2188 19168
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 10324 19320 10376 19372
rect 11520 19320 11572 19372
rect 7840 19252 7892 19304
rect 9128 19252 9180 19304
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 10784 19252 10836 19304
rect 11980 19388 12032 19440
rect 11888 19320 11940 19372
rect 12440 19320 12492 19372
rect 13544 19431 13596 19440
rect 13544 19397 13553 19431
rect 13553 19397 13587 19431
rect 13587 19397 13596 19431
rect 13544 19388 13596 19397
rect 16212 19388 16264 19440
rect 16304 19388 16356 19440
rect 18788 19456 18840 19508
rect 20352 19456 20404 19508
rect 21456 19499 21508 19508
rect 21456 19465 21465 19499
rect 21465 19465 21499 19499
rect 21499 19465 21508 19499
rect 21456 19456 21508 19465
rect 21916 19456 21968 19508
rect 23296 19456 23348 19508
rect 23480 19456 23532 19508
rect 24124 19456 24176 19508
rect 17776 19388 17828 19440
rect 19156 19388 19208 19440
rect 20996 19388 21048 19440
rect 21272 19388 21324 19440
rect 24676 19388 24728 19440
rect 24860 19456 24912 19508
rect 29644 19456 29696 19508
rect 11980 19252 12032 19304
rect 12256 19252 12308 19304
rect 14924 19320 14976 19372
rect 15292 19320 15344 19372
rect 17592 19320 17644 19372
rect 14832 19295 14884 19304
rect 14832 19261 14841 19295
rect 14841 19261 14875 19295
rect 14875 19261 14884 19295
rect 14832 19252 14884 19261
rect 15936 19295 15988 19304
rect 15936 19261 15945 19295
rect 15945 19261 15979 19295
rect 15979 19261 15988 19295
rect 15936 19252 15988 19261
rect 16028 19295 16080 19304
rect 16028 19261 16037 19295
rect 16037 19261 16071 19295
rect 16071 19261 16080 19295
rect 16028 19252 16080 19261
rect 16120 19252 16172 19304
rect 17500 19252 17552 19304
rect 17684 19252 17736 19304
rect 17960 19252 18012 19304
rect 6092 19184 6144 19236
rect 11612 19184 11664 19236
rect 8944 19159 8996 19168
rect 8944 19125 8953 19159
rect 8953 19125 8987 19159
rect 8987 19125 8996 19159
rect 8944 19116 8996 19125
rect 9496 19116 9548 19168
rect 13820 19184 13872 19236
rect 14280 19227 14332 19236
rect 14280 19193 14289 19227
rect 14289 19193 14323 19227
rect 14323 19193 14332 19227
rect 14280 19184 14332 19193
rect 12532 19116 12584 19168
rect 16672 19116 16724 19168
rect 16764 19116 16816 19168
rect 17868 19116 17920 19168
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19616 19320 19668 19372
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 22376 19363 22428 19372
rect 22376 19329 22385 19363
rect 22385 19329 22419 19363
rect 22419 19329 22428 19363
rect 22376 19320 22428 19329
rect 18236 19252 18288 19304
rect 18788 19252 18840 19304
rect 18696 19184 18748 19236
rect 21364 19252 21416 19304
rect 22744 19252 22796 19304
rect 22928 19320 22980 19372
rect 24124 19363 24176 19372
rect 24124 19329 24133 19363
rect 24133 19329 24167 19363
rect 24167 19329 24176 19363
rect 24124 19320 24176 19329
rect 24952 19431 25004 19440
rect 24952 19397 24961 19431
rect 24961 19397 24995 19431
rect 24995 19397 25004 19431
rect 24952 19388 25004 19397
rect 25504 19388 25556 19440
rect 24400 19295 24452 19304
rect 24400 19261 24409 19295
rect 24409 19261 24443 19295
rect 24443 19261 24452 19295
rect 24400 19252 24452 19261
rect 25596 19320 25648 19372
rect 26792 19388 26844 19440
rect 27712 19388 27764 19440
rect 28908 19388 28960 19440
rect 32312 19456 32364 19508
rect 36636 19499 36688 19508
rect 36636 19465 36645 19499
rect 36645 19465 36679 19499
rect 36679 19465 36688 19499
rect 36636 19456 36688 19465
rect 31300 19388 31352 19440
rect 40224 19456 40276 19508
rect 41236 19456 41288 19508
rect 41512 19456 41564 19508
rect 25780 19295 25832 19304
rect 25780 19261 25789 19295
rect 25789 19261 25823 19295
rect 25823 19261 25832 19295
rect 25780 19252 25832 19261
rect 29736 19320 29788 19372
rect 19524 19116 19576 19168
rect 19984 19116 20036 19168
rect 26792 19184 26844 19236
rect 22652 19116 22704 19168
rect 22836 19116 22888 19168
rect 23572 19116 23624 19168
rect 24492 19116 24544 19168
rect 26516 19159 26568 19168
rect 26516 19125 26525 19159
rect 26525 19125 26559 19159
rect 26559 19125 26568 19159
rect 26516 19116 26568 19125
rect 27620 19295 27672 19304
rect 27620 19261 27629 19295
rect 27629 19261 27663 19295
rect 27663 19261 27672 19295
rect 27620 19252 27672 19261
rect 27344 19184 27396 19236
rect 28356 19295 28408 19304
rect 28356 19261 28365 19295
rect 28365 19261 28399 19295
rect 28399 19261 28408 19295
rect 28356 19252 28408 19261
rect 29276 19252 29328 19304
rect 30472 19320 30524 19372
rect 31760 19320 31812 19372
rect 32128 19320 32180 19372
rect 38384 19388 38436 19440
rect 40500 19388 40552 19440
rect 31944 19252 31996 19304
rect 33140 19252 33192 19304
rect 35532 19363 35584 19372
rect 35532 19329 35541 19363
rect 35541 19329 35575 19363
rect 35575 19329 35584 19363
rect 35532 19320 35584 19329
rect 35992 19363 36044 19372
rect 35992 19329 36001 19363
rect 36001 19329 36035 19363
rect 36035 19329 36044 19363
rect 35992 19320 36044 19329
rect 38476 19320 38528 19372
rect 38568 19320 38620 19372
rect 40224 19320 40276 19372
rect 36636 19252 36688 19304
rect 39120 19252 39172 19304
rect 30932 19184 30984 19236
rect 31300 19184 31352 19236
rect 31484 19184 31536 19236
rect 33048 19184 33100 19236
rect 28816 19116 28868 19168
rect 31760 19159 31812 19168
rect 31760 19125 31769 19159
rect 31769 19125 31803 19159
rect 31803 19125 31812 19159
rect 31760 19116 31812 19125
rect 32312 19116 32364 19168
rect 34612 19184 34664 19236
rect 39396 19184 39448 19236
rect 41788 19252 41840 19304
rect 45468 19184 45520 19236
rect 34336 19159 34388 19168
rect 34336 19125 34345 19159
rect 34345 19125 34379 19159
rect 34379 19125 34388 19159
rect 34336 19116 34388 19125
rect 36636 19116 36688 19168
rect 39488 19159 39540 19168
rect 39488 19125 39497 19159
rect 39497 19125 39531 19159
rect 39531 19125 39540 19159
rect 39488 19116 39540 19125
rect 40776 19159 40828 19168
rect 40776 19125 40785 19159
rect 40785 19125 40819 19159
rect 40819 19125 40828 19159
rect 40776 19116 40828 19125
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 2412 18912 2464 18964
rect 6736 18912 6788 18964
rect 480 18844 532 18896
rect 6368 18844 6420 18896
rect 1400 18776 1452 18828
rect 3424 18819 3476 18828
rect 3424 18785 3433 18819
rect 3433 18785 3467 18819
rect 3467 18785 3476 18819
rect 3424 18776 3476 18785
rect 3608 18776 3660 18828
rect 6276 18819 6328 18828
rect 6276 18785 6285 18819
rect 6285 18785 6319 18819
rect 6319 18785 6328 18819
rect 6276 18776 6328 18785
rect 7380 18912 7432 18964
rect 7840 18912 7892 18964
rect 8944 18912 8996 18964
rect 12440 18912 12492 18964
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 13636 18912 13688 18964
rect 13912 18912 13964 18964
rect 14832 18912 14884 18964
rect 16580 18912 16632 18964
rect 17224 18912 17276 18964
rect 7932 18844 7984 18896
rect 9956 18844 10008 18896
rect 12348 18844 12400 18896
rect 14004 18844 14056 18896
rect 16212 18844 16264 18896
rect 8300 18776 8352 18828
rect 8392 18776 8444 18828
rect 3516 18708 3568 18760
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 9128 18708 9180 18760
rect 9220 18708 9272 18760
rect 11704 18776 11756 18828
rect 14372 18776 14424 18828
rect 14464 18819 14516 18828
rect 14464 18785 14473 18819
rect 14473 18785 14507 18819
rect 14507 18785 14516 18819
rect 14464 18776 14516 18785
rect 15752 18776 15804 18828
rect 16580 18776 16632 18828
rect 17684 18912 17736 18964
rect 19892 18912 19944 18964
rect 22376 18912 22428 18964
rect 23388 18912 23440 18964
rect 24768 18912 24820 18964
rect 17500 18844 17552 18896
rect 12716 18708 12768 18760
rect 17776 18776 17828 18828
rect 18144 18819 18196 18828
rect 18144 18785 18153 18819
rect 18153 18785 18187 18819
rect 18187 18785 18196 18819
rect 18144 18776 18196 18785
rect 17040 18708 17092 18760
rect 19984 18776 20036 18828
rect 20260 18776 20312 18828
rect 20904 18776 20956 18828
rect 23572 18844 23624 18896
rect 25320 18912 25372 18964
rect 25504 18912 25556 18964
rect 27528 18912 27580 18964
rect 27620 18912 27672 18964
rect 29828 18912 29880 18964
rect 33324 18912 33376 18964
rect 33692 18912 33744 18964
rect 34244 18912 34296 18964
rect 35624 18912 35676 18964
rect 35716 18912 35768 18964
rect 19064 18708 19116 18760
rect 19432 18708 19484 18760
rect 20720 18708 20772 18760
rect 23572 18708 23624 18760
rect 23848 18776 23900 18828
rect 24676 18776 24728 18828
rect 26792 18844 26844 18896
rect 37096 18912 37148 18964
rect 7932 18640 7984 18692
rect 8024 18683 8076 18692
rect 8024 18649 8033 18683
rect 8033 18649 8067 18683
rect 8067 18649 8076 18683
rect 8024 18640 8076 18649
rect 9404 18640 9456 18692
rect 10600 18683 10652 18692
rect 10600 18649 10609 18683
rect 10609 18649 10643 18683
rect 10643 18649 10652 18683
rect 10600 18640 10652 18649
rect 11152 18683 11204 18692
rect 11152 18649 11161 18683
rect 11161 18649 11195 18683
rect 11195 18649 11204 18683
rect 11152 18640 11204 18649
rect 15016 18683 15068 18692
rect 15016 18649 15025 18683
rect 15025 18649 15059 18683
rect 15059 18649 15068 18683
rect 15016 18640 15068 18649
rect 15476 18640 15528 18692
rect 16304 18640 16356 18692
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 5724 18572 5776 18624
rect 7564 18572 7616 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 7840 18572 7892 18624
rect 8760 18615 8812 18624
rect 8760 18581 8769 18615
rect 8769 18581 8803 18615
rect 8803 18581 8812 18615
rect 8760 18572 8812 18581
rect 8852 18572 8904 18624
rect 10324 18572 10376 18624
rect 11060 18572 11112 18624
rect 11336 18572 11388 18624
rect 11980 18572 12032 18624
rect 15292 18572 15344 18624
rect 15752 18572 15804 18624
rect 16764 18640 16816 18692
rect 17868 18640 17920 18692
rect 22652 18640 22704 18692
rect 24308 18640 24360 18692
rect 24952 18640 25004 18692
rect 18236 18572 18288 18624
rect 18420 18572 18472 18624
rect 18788 18615 18840 18624
rect 18788 18581 18797 18615
rect 18797 18581 18831 18615
rect 18831 18581 18840 18615
rect 18788 18572 18840 18581
rect 19156 18572 19208 18624
rect 19432 18572 19484 18624
rect 20628 18572 20680 18624
rect 22744 18572 22796 18624
rect 23664 18572 23716 18624
rect 23848 18572 23900 18624
rect 25228 18615 25280 18624
rect 25228 18581 25237 18615
rect 25237 18581 25271 18615
rect 25271 18581 25280 18615
rect 25228 18572 25280 18581
rect 25780 18776 25832 18828
rect 25872 18776 25924 18828
rect 26148 18776 26200 18828
rect 26240 18776 26292 18828
rect 28264 18776 28316 18828
rect 28816 18708 28868 18760
rect 29092 18819 29144 18828
rect 29092 18785 29101 18819
rect 29101 18785 29135 18819
rect 29135 18785 29144 18819
rect 29092 18776 29144 18785
rect 29460 18776 29512 18828
rect 26240 18640 26292 18692
rect 30840 18751 30892 18760
rect 30840 18717 30849 18751
rect 30849 18717 30883 18751
rect 30883 18717 30892 18751
rect 30840 18708 30892 18717
rect 31208 18776 31260 18828
rect 32220 18708 32272 18760
rect 32312 18751 32364 18760
rect 32312 18717 32321 18751
rect 32321 18717 32355 18751
rect 32355 18717 32364 18751
rect 32312 18708 32364 18717
rect 32496 18708 32548 18760
rect 33784 18708 33836 18760
rect 27160 18572 27212 18624
rect 27804 18572 27856 18624
rect 28264 18572 28316 18624
rect 29368 18572 29420 18624
rect 30196 18572 30248 18624
rect 30380 18615 30432 18624
rect 30380 18581 30389 18615
rect 30389 18581 30423 18615
rect 30423 18581 30432 18615
rect 30380 18572 30432 18581
rect 30564 18572 30616 18624
rect 31760 18683 31812 18692
rect 31760 18649 31769 18683
rect 31769 18649 31803 18683
rect 31803 18649 31812 18683
rect 31760 18640 31812 18649
rect 33692 18640 33744 18692
rect 34336 18640 34388 18692
rect 34888 18751 34940 18760
rect 34888 18717 34897 18751
rect 34897 18717 34931 18751
rect 34931 18717 34940 18751
rect 34888 18708 34940 18717
rect 39580 18912 39632 18964
rect 43536 18912 43588 18964
rect 37464 18751 37516 18760
rect 37464 18717 37473 18751
rect 37473 18717 37507 18751
rect 37507 18717 37516 18751
rect 37464 18708 37516 18717
rect 40224 18887 40276 18896
rect 40224 18853 40233 18887
rect 40233 18853 40267 18887
rect 40267 18853 40276 18887
rect 40224 18844 40276 18853
rect 32956 18615 33008 18624
rect 32956 18581 32965 18615
rect 32965 18581 32999 18615
rect 32999 18581 33008 18615
rect 32956 18572 33008 18581
rect 33508 18572 33560 18624
rect 34888 18572 34940 18624
rect 35624 18572 35676 18624
rect 37832 18572 37884 18624
rect 38752 18615 38804 18624
rect 38752 18581 38761 18615
rect 38761 18581 38795 18615
rect 38795 18581 38804 18615
rect 38752 18572 38804 18581
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 3424 18368 3476 18420
rect 5816 18300 5868 18352
rect 3332 18232 3384 18284
rect 7380 18300 7432 18352
rect 7472 18343 7524 18352
rect 7472 18309 7481 18343
rect 7481 18309 7515 18343
rect 7515 18309 7524 18343
rect 7472 18300 7524 18309
rect 7932 18300 7984 18352
rect 2044 18207 2096 18216
rect 2044 18173 2053 18207
rect 2053 18173 2087 18207
rect 2087 18173 2096 18207
rect 2044 18164 2096 18173
rect 3884 18207 3936 18216
rect 3884 18173 3893 18207
rect 3893 18173 3927 18207
rect 3927 18173 3936 18207
rect 3884 18164 3936 18173
rect 5724 18207 5776 18216
rect 5724 18173 5733 18207
rect 5733 18173 5767 18207
rect 5767 18173 5776 18207
rect 5724 18164 5776 18173
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 6092 18164 6144 18216
rect 7288 18164 7340 18216
rect 7932 18096 7984 18148
rect 8208 18164 8260 18216
rect 10876 18368 10928 18420
rect 11520 18368 11572 18420
rect 12900 18368 12952 18420
rect 9588 18300 9640 18352
rect 8944 18275 8996 18284
rect 8944 18241 8953 18275
rect 8953 18241 8987 18275
rect 8987 18241 8996 18275
rect 8944 18232 8996 18241
rect 9404 18232 9456 18284
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 11612 18300 11664 18352
rect 12440 18300 12492 18352
rect 14648 18368 14700 18420
rect 15108 18368 15160 18420
rect 14372 18300 14424 18352
rect 13912 18232 13964 18284
rect 15200 18275 15252 18284
rect 15200 18241 15209 18275
rect 15209 18241 15243 18275
rect 15243 18241 15252 18275
rect 15200 18232 15252 18241
rect 15292 18232 15344 18284
rect 10600 18164 10652 18216
rect 10876 18164 10928 18216
rect 10968 18207 11020 18216
rect 10968 18173 10977 18207
rect 10977 18173 11011 18207
rect 11011 18173 11020 18207
rect 10968 18164 11020 18173
rect 12256 18164 12308 18216
rect 13452 18164 13504 18216
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 15752 18164 15804 18216
rect 16120 18275 16172 18284
rect 16120 18241 16129 18275
rect 16129 18241 16163 18275
rect 16163 18241 16172 18275
rect 16120 18232 16172 18241
rect 16212 18232 16264 18284
rect 17132 18232 17184 18284
rect 17868 18232 17920 18284
rect 19800 18300 19852 18352
rect 22652 18343 22704 18352
rect 22652 18309 22661 18343
rect 22661 18309 22695 18343
rect 22695 18309 22704 18343
rect 22652 18300 22704 18309
rect 23296 18300 23348 18352
rect 23848 18300 23900 18352
rect 24676 18300 24728 18352
rect 29368 18368 29420 18420
rect 25964 18300 26016 18352
rect 26148 18300 26200 18352
rect 27620 18300 27672 18352
rect 18144 18232 18196 18284
rect 18972 18232 19024 18284
rect 19524 18275 19576 18284
rect 19524 18241 19533 18275
rect 19533 18241 19567 18275
rect 19567 18241 19576 18275
rect 19524 18232 19576 18241
rect 16580 18164 16632 18216
rect 19156 18164 19208 18216
rect 19248 18164 19300 18216
rect 19984 18164 20036 18216
rect 16764 18096 16816 18148
rect 17132 18096 17184 18148
rect 19524 18096 19576 18148
rect 22008 18275 22060 18284
rect 22008 18241 22017 18275
rect 22017 18241 22051 18275
rect 22051 18241 22060 18275
rect 22008 18232 22060 18241
rect 23112 18275 23164 18284
rect 23112 18241 23121 18275
rect 23121 18241 23155 18275
rect 23155 18241 23164 18275
rect 23112 18232 23164 18241
rect 25228 18232 25280 18284
rect 27528 18232 27580 18284
rect 27988 18232 28040 18284
rect 28356 18300 28408 18352
rect 29736 18368 29788 18420
rect 32128 18411 32180 18420
rect 32128 18377 32137 18411
rect 32137 18377 32171 18411
rect 32171 18377 32180 18411
rect 32128 18368 32180 18377
rect 30104 18300 30156 18352
rect 32036 18300 32088 18352
rect 29460 18232 29512 18284
rect 30564 18232 30616 18284
rect 33600 18368 33652 18420
rect 36912 18368 36964 18420
rect 37740 18300 37792 18352
rect 34244 18232 34296 18284
rect 35808 18275 35860 18284
rect 35808 18241 35817 18275
rect 35817 18241 35851 18275
rect 35851 18241 35860 18275
rect 35808 18232 35860 18241
rect 37188 18232 37240 18284
rect 38660 18232 38712 18284
rect 25136 18164 25188 18216
rect 26148 18164 26200 18216
rect 27160 18207 27212 18216
rect 27160 18173 27169 18207
rect 27169 18173 27203 18207
rect 27203 18173 27212 18207
rect 27160 18164 27212 18173
rect 32956 18164 33008 18216
rect 33416 18164 33468 18216
rect 34520 18207 34572 18216
rect 34520 18173 34529 18207
rect 34529 18173 34563 18207
rect 34563 18173 34572 18207
rect 34520 18164 34572 18173
rect 22468 18096 22520 18148
rect 26516 18096 26568 18148
rect 6000 18028 6052 18080
rect 7104 18028 7156 18080
rect 8116 18028 8168 18080
rect 8576 18028 8628 18080
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 8760 18028 8812 18080
rect 12900 18028 12952 18080
rect 14372 18028 14424 18080
rect 14924 18028 14976 18080
rect 18420 18028 18472 18080
rect 20076 18028 20128 18080
rect 20168 18071 20220 18080
rect 20168 18037 20177 18071
rect 20177 18037 20211 18071
rect 20211 18037 20220 18071
rect 20168 18028 20220 18037
rect 20352 18028 20404 18080
rect 23112 18028 23164 18080
rect 23388 18028 23440 18080
rect 23480 18028 23532 18080
rect 25504 18028 25556 18080
rect 27068 18028 27120 18080
rect 27804 18028 27856 18080
rect 30564 18096 30616 18148
rect 36820 18164 36872 18216
rect 39856 18164 39908 18216
rect 46848 18096 46900 18148
rect 30840 18028 30892 18080
rect 31668 18028 31720 18080
rect 36452 18071 36504 18080
rect 36452 18037 36461 18071
rect 36461 18037 36495 18071
rect 36495 18037 36504 18071
rect 36452 18028 36504 18037
rect 36728 18028 36780 18080
rect 37188 18028 37240 18080
rect 37648 18071 37700 18080
rect 37648 18037 37657 18071
rect 37657 18037 37691 18071
rect 37691 18037 37700 18071
rect 37648 18028 37700 18037
rect 38384 18071 38436 18080
rect 38384 18037 38393 18071
rect 38393 18037 38427 18071
rect 38427 18037 38436 18071
rect 38384 18028 38436 18037
rect 38936 18071 38988 18080
rect 38936 18037 38945 18071
rect 38945 18037 38979 18071
rect 38979 18037 38988 18071
rect 38936 18028 38988 18037
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 1308 17824 1360 17876
rect 1584 17824 1636 17876
rect 2780 17824 2832 17876
rect 7472 17824 7524 17876
rect 10968 17824 11020 17876
rect 1216 17688 1268 17740
rect 6552 17756 6604 17808
rect 11888 17756 11940 17808
rect 12072 17756 12124 17808
rect 12808 17824 12860 17876
rect 14556 17824 14608 17876
rect 14832 17824 14884 17876
rect 15292 17824 15344 17876
rect 16304 17824 16356 17876
rect 16580 17824 16632 17876
rect 17224 17824 17276 17876
rect 18420 17824 18472 17876
rect 3608 17731 3660 17740
rect 3608 17697 3617 17731
rect 3617 17697 3651 17731
rect 3651 17697 3660 17731
rect 3608 17688 3660 17697
rect 4804 17731 4856 17740
rect 4804 17697 4813 17731
rect 4813 17697 4847 17731
rect 4847 17697 4856 17731
rect 4804 17688 4856 17697
rect 3884 17663 3936 17672
rect 3884 17629 3893 17663
rect 3893 17629 3927 17663
rect 3927 17629 3936 17663
rect 3884 17620 3936 17629
rect 4344 17663 4396 17672
rect 4344 17629 4353 17663
rect 4353 17629 4387 17663
rect 4387 17629 4396 17663
rect 4344 17620 4396 17629
rect 6184 17620 6236 17672
rect 6920 17688 6972 17740
rect 9128 17688 9180 17740
rect 9496 17688 9548 17740
rect 10600 17688 10652 17740
rect 11520 17688 11572 17740
rect 11612 17688 11664 17740
rect 11796 17688 11848 17740
rect 12348 17731 12400 17740
rect 12348 17697 12357 17731
rect 12357 17697 12391 17731
rect 12391 17697 12400 17731
rect 12348 17688 12400 17697
rect 13728 17688 13780 17740
rect 14924 17688 14976 17740
rect 15844 17731 15896 17740
rect 15844 17697 15853 17731
rect 15853 17697 15887 17731
rect 15887 17697 15896 17731
rect 15844 17688 15896 17697
rect 17684 17756 17736 17808
rect 18144 17756 18196 17808
rect 21180 17824 21232 17876
rect 22192 17824 22244 17876
rect 22468 17824 22520 17876
rect 24308 17824 24360 17876
rect 30380 17824 30432 17876
rect 37464 17824 37516 17876
rect 38660 17824 38712 17876
rect 45376 17824 45428 17876
rect 17776 17688 17828 17740
rect 9956 17620 10008 17672
rect 2504 17552 2556 17604
rect 4252 17552 4304 17604
rect 5172 17552 5224 17604
rect 1400 17484 1452 17536
rect 6828 17484 6880 17536
rect 6920 17484 6972 17536
rect 8852 17552 8904 17604
rect 8944 17552 8996 17604
rect 9128 17595 9180 17604
rect 9128 17561 9137 17595
rect 9137 17561 9171 17595
rect 9171 17561 9180 17595
rect 9128 17552 9180 17561
rect 9220 17552 9272 17604
rect 11520 17552 11572 17604
rect 7840 17527 7892 17536
rect 7840 17493 7849 17527
rect 7849 17493 7883 17527
rect 7883 17493 7892 17527
rect 7840 17484 7892 17493
rect 10600 17484 10652 17536
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 12532 17552 12584 17604
rect 14556 17620 14608 17672
rect 17408 17620 17460 17672
rect 18144 17620 18196 17672
rect 15844 17552 15896 17604
rect 16120 17595 16172 17604
rect 16120 17561 16129 17595
rect 16129 17561 16163 17595
rect 16163 17561 16172 17595
rect 16120 17552 16172 17561
rect 17500 17552 17552 17604
rect 17868 17552 17920 17604
rect 22008 17756 22060 17808
rect 20628 17688 20680 17740
rect 26148 17756 26200 17808
rect 28448 17756 28500 17808
rect 18972 17620 19024 17672
rect 21640 17620 21692 17672
rect 18880 17552 18932 17604
rect 19248 17552 19300 17604
rect 21272 17552 21324 17604
rect 24676 17688 24728 17740
rect 25780 17688 25832 17740
rect 27988 17688 28040 17740
rect 30196 17756 30248 17808
rect 31576 17756 31628 17808
rect 29460 17688 29512 17740
rect 31024 17688 31076 17740
rect 22008 17620 22060 17672
rect 23388 17620 23440 17672
rect 23664 17620 23716 17672
rect 23756 17620 23808 17672
rect 26792 17620 26844 17672
rect 26976 17620 27028 17672
rect 28448 17620 28500 17672
rect 30840 17620 30892 17672
rect 32036 17663 32088 17672
rect 32036 17629 32045 17663
rect 32045 17629 32079 17663
rect 32079 17629 32088 17663
rect 32036 17620 32088 17629
rect 12624 17527 12676 17536
rect 12624 17493 12633 17527
rect 12633 17493 12667 17527
rect 12667 17493 12676 17527
rect 12624 17484 12676 17493
rect 13268 17527 13320 17536
rect 13268 17493 13277 17527
rect 13277 17493 13311 17527
rect 13311 17493 13320 17527
rect 13268 17484 13320 17493
rect 14372 17484 14424 17536
rect 14464 17484 14516 17536
rect 16856 17484 16908 17536
rect 17592 17527 17644 17536
rect 17592 17493 17601 17527
rect 17601 17493 17635 17527
rect 17635 17493 17644 17527
rect 17592 17484 17644 17493
rect 19432 17484 19484 17536
rect 19616 17527 19668 17536
rect 19616 17493 19625 17527
rect 19625 17493 19659 17527
rect 19659 17493 19668 17527
rect 19616 17484 19668 17493
rect 20260 17484 20312 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 20904 17484 20956 17536
rect 22468 17484 22520 17536
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 24308 17484 24360 17536
rect 27068 17552 27120 17604
rect 27436 17552 27488 17604
rect 29276 17595 29328 17604
rect 29276 17561 29285 17595
rect 29285 17561 29319 17595
rect 29319 17561 29328 17595
rect 29276 17552 29328 17561
rect 32864 17756 32916 17808
rect 36636 17756 36688 17808
rect 36912 17799 36964 17808
rect 36912 17765 36921 17799
rect 36921 17765 36955 17799
rect 36955 17765 36964 17799
rect 36912 17756 36964 17765
rect 36268 17688 36320 17740
rect 33324 17620 33376 17672
rect 34612 17620 34664 17672
rect 35900 17620 35952 17672
rect 37004 17620 37056 17672
rect 37464 17620 37516 17672
rect 39304 17552 39356 17604
rect 28264 17484 28316 17536
rect 29644 17484 29696 17536
rect 30104 17527 30156 17536
rect 30104 17493 30113 17527
rect 30113 17493 30147 17527
rect 30147 17493 30156 17527
rect 30104 17484 30156 17493
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 30564 17484 30616 17536
rect 31208 17484 31260 17536
rect 32680 17527 32732 17536
rect 32680 17493 32689 17527
rect 32689 17493 32723 17527
rect 32723 17493 32732 17527
rect 32680 17484 32732 17493
rect 34060 17527 34112 17536
rect 34060 17493 34069 17527
rect 34069 17493 34103 17527
rect 34103 17493 34112 17527
rect 34060 17484 34112 17493
rect 34612 17484 34664 17536
rect 36084 17484 36136 17536
rect 37372 17527 37424 17536
rect 37372 17493 37381 17527
rect 37381 17493 37415 17527
rect 37415 17493 37424 17527
rect 37372 17484 37424 17493
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 7656 17280 7708 17332
rect 8024 17323 8076 17332
rect 8024 17289 8033 17323
rect 8033 17289 8067 17323
rect 8067 17289 8076 17323
rect 8024 17280 8076 17289
rect 8576 17280 8628 17332
rect 9864 17280 9916 17332
rect 10232 17280 10284 17332
rect 10968 17280 11020 17332
rect 14096 17280 14148 17332
rect 14188 17323 14240 17332
rect 14188 17289 14197 17323
rect 14197 17289 14231 17323
rect 14231 17289 14240 17323
rect 14188 17280 14240 17289
rect 14832 17280 14884 17332
rect 17500 17280 17552 17332
rect 10600 17212 10652 17264
rect 1768 17187 1820 17196
rect 1768 17153 1777 17187
rect 1777 17153 1811 17187
rect 1811 17153 1820 17187
rect 1768 17144 1820 17153
rect 4252 17144 4304 17196
rect 6368 17144 6420 17196
rect 6552 17187 6604 17196
rect 6552 17153 6561 17187
rect 6561 17153 6595 17187
rect 6595 17153 6604 17187
rect 6552 17144 6604 17153
rect 7196 17187 7248 17196
rect 7196 17153 7205 17187
rect 7205 17153 7239 17187
rect 7239 17153 7248 17187
rect 7196 17144 7248 17153
rect 1308 17076 1360 17128
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 5908 17119 5960 17128
rect 5908 17085 5917 17119
rect 5917 17085 5951 17119
rect 5951 17085 5960 17119
rect 5908 17076 5960 17085
rect 6828 17076 6880 17128
rect 6920 17076 6972 17128
rect 8576 17144 8628 17196
rect 11980 17212 12032 17264
rect 15108 17212 15160 17264
rect 17132 17212 17184 17264
rect 17224 17212 17276 17264
rect 11060 17144 11112 17196
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 14280 17144 14332 17196
rect 15660 17144 15712 17196
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 7472 17076 7524 17128
rect 8208 17119 8260 17128
rect 8208 17085 8217 17119
rect 8217 17085 8251 17119
rect 8251 17085 8260 17119
rect 8208 17076 8260 17085
rect 9312 17119 9364 17128
rect 9312 17085 9321 17119
rect 9321 17085 9355 17119
rect 9355 17085 9364 17119
rect 9312 17076 9364 17085
rect 9496 17119 9548 17128
rect 9496 17085 9505 17119
rect 9505 17085 9539 17119
rect 9539 17085 9548 17119
rect 9496 17076 9548 17085
rect 10324 17076 10376 17128
rect 10600 17076 10652 17128
rect 5724 17008 5776 17060
rect 10784 17008 10836 17060
rect 12624 17076 12676 17128
rect 14648 17076 14700 17128
rect 14832 17119 14884 17128
rect 14832 17085 14841 17119
rect 14841 17085 14875 17119
rect 14875 17085 14884 17119
rect 14832 17076 14884 17085
rect 15752 17076 15804 17128
rect 16028 17119 16080 17128
rect 16028 17085 16037 17119
rect 16037 17085 16071 17119
rect 16071 17085 16080 17119
rect 16028 17076 16080 17085
rect 16212 17119 16264 17128
rect 16212 17085 16221 17119
rect 16221 17085 16255 17119
rect 16255 17085 16264 17119
rect 16212 17076 16264 17085
rect 17868 17212 17920 17264
rect 18328 17280 18380 17332
rect 19800 17212 19852 17264
rect 20352 17212 20404 17264
rect 19616 17144 19668 17196
rect 20720 17280 20772 17332
rect 21180 17212 21232 17264
rect 22192 17280 22244 17332
rect 22468 17323 22520 17332
rect 22468 17289 22477 17323
rect 22477 17289 22511 17323
rect 22511 17289 22520 17323
rect 22468 17280 22520 17289
rect 23204 17280 23256 17332
rect 23756 17280 23808 17332
rect 9956 16940 10008 16992
rect 10324 16940 10376 16992
rect 10416 16983 10468 16992
rect 10416 16949 10425 16983
rect 10425 16949 10459 16983
rect 10459 16949 10468 16983
rect 10416 16940 10468 16949
rect 11980 16940 12032 16992
rect 12624 16940 12676 16992
rect 13452 16983 13504 16992
rect 13452 16949 13461 16983
rect 13461 16949 13495 16983
rect 13495 16949 13504 16983
rect 13452 16940 13504 16949
rect 13636 16940 13688 16992
rect 14096 16983 14148 16992
rect 14096 16949 14105 16983
rect 14105 16949 14139 16983
rect 14139 16949 14148 16983
rect 14096 16940 14148 16949
rect 15384 17008 15436 17060
rect 17592 17008 17644 17060
rect 19156 17008 19208 17060
rect 16764 16940 16816 16992
rect 16856 16940 16908 16992
rect 20168 17076 20220 17128
rect 21640 17144 21692 17196
rect 23756 17144 23808 17196
rect 24308 17212 24360 17264
rect 27344 17280 27396 17332
rect 27068 17212 27120 17264
rect 28448 17212 28500 17264
rect 29460 17212 29512 17264
rect 32036 17280 32088 17332
rect 34520 17280 34572 17332
rect 35900 17323 35952 17332
rect 35900 17289 35909 17323
rect 35909 17289 35943 17323
rect 35943 17289 35952 17323
rect 35900 17280 35952 17289
rect 30840 17212 30892 17264
rect 31668 17212 31720 17264
rect 24676 17187 24728 17196
rect 24676 17153 24685 17187
rect 24685 17153 24719 17187
rect 24719 17153 24728 17187
rect 24676 17144 24728 17153
rect 26792 17187 26844 17196
rect 26792 17153 26801 17187
rect 26801 17153 26835 17187
rect 26835 17153 26844 17187
rect 26792 17144 26844 17153
rect 27528 17144 27580 17196
rect 30288 17144 30340 17196
rect 31116 17144 31168 17196
rect 20260 16940 20312 16992
rect 20904 16940 20956 16992
rect 21456 17008 21508 17060
rect 22468 17076 22520 17128
rect 22100 17051 22152 17060
rect 22100 17017 22109 17051
rect 22109 17017 22143 17051
rect 22143 17017 22152 17051
rect 22100 17008 22152 17017
rect 23664 17008 23716 17060
rect 22744 16940 22796 16992
rect 23480 16983 23532 16992
rect 23480 16949 23489 16983
rect 23489 16949 23523 16983
rect 23523 16949 23532 16983
rect 23480 16940 23532 16949
rect 24124 17119 24176 17128
rect 24124 17085 24133 17119
rect 24133 17085 24167 17119
rect 24167 17085 24176 17119
rect 24124 17076 24176 17085
rect 24400 17076 24452 17128
rect 26148 17076 26200 17128
rect 27252 17119 27304 17128
rect 27252 17085 27261 17119
rect 27261 17085 27295 17119
rect 27295 17085 27304 17119
rect 27252 17076 27304 17085
rect 28908 17076 28960 17128
rect 29184 17076 29236 17128
rect 31300 17076 31352 17128
rect 31944 17008 31996 17060
rect 34060 17144 34112 17196
rect 34520 17144 34572 17196
rect 41604 17280 41656 17332
rect 32772 17076 32824 17128
rect 37280 17144 37332 17196
rect 47400 17212 47452 17264
rect 34796 17076 34848 17128
rect 35992 17076 36044 17128
rect 39212 17076 39264 17128
rect 38936 17008 38988 17060
rect 30564 16940 30616 16992
rect 32404 16940 32456 16992
rect 34704 16983 34756 16992
rect 34704 16949 34713 16983
rect 34713 16949 34747 16983
rect 34747 16949 34756 16983
rect 34704 16940 34756 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 3424 16711 3476 16720
rect 3424 16677 3433 16711
rect 3433 16677 3467 16711
rect 3467 16677 3476 16711
rect 3424 16668 3476 16677
rect 3608 16668 3660 16720
rect 8116 16668 8168 16720
rect 8576 16668 8628 16720
rect 2412 16600 2464 16652
rect 3792 16600 3844 16652
rect 1308 16464 1360 16516
rect 4988 16575 5040 16584
rect 4988 16541 4997 16575
rect 4997 16541 5031 16575
rect 5031 16541 5040 16575
rect 4988 16532 5040 16541
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 9404 16736 9456 16788
rect 11060 16736 11112 16788
rect 13360 16736 13412 16788
rect 14740 16736 14792 16788
rect 15568 16736 15620 16788
rect 15844 16736 15896 16788
rect 20076 16736 20128 16788
rect 9312 16668 9364 16720
rect 8760 16600 8812 16652
rect 9956 16600 10008 16652
rect 10324 16600 10376 16652
rect 10876 16643 10928 16652
rect 10876 16609 10885 16643
rect 10885 16609 10919 16643
rect 10919 16609 10928 16643
rect 10876 16600 10928 16609
rect 11060 16643 11112 16652
rect 11060 16609 11069 16643
rect 11069 16609 11103 16643
rect 11103 16609 11112 16643
rect 11060 16600 11112 16609
rect 16856 16668 16908 16720
rect 17132 16711 17184 16720
rect 17132 16677 17141 16711
rect 17141 16677 17175 16711
rect 17175 16677 17184 16711
rect 17132 16668 17184 16677
rect 12992 16600 13044 16652
rect 5816 16464 5868 16516
rect 6460 16464 6512 16516
rect 4620 16396 4672 16448
rect 5264 16396 5316 16448
rect 6092 16396 6144 16448
rect 6920 16396 6972 16448
rect 7288 16396 7340 16448
rect 9496 16532 9548 16584
rect 9588 16532 9640 16584
rect 13268 16532 13320 16584
rect 13360 16575 13412 16584
rect 13360 16541 13369 16575
rect 13369 16541 13403 16575
rect 13403 16541 13412 16575
rect 13360 16532 13412 16541
rect 13636 16643 13688 16652
rect 13636 16609 13645 16643
rect 13645 16609 13679 16643
rect 13679 16609 13688 16643
rect 13636 16600 13688 16609
rect 13820 16600 13872 16652
rect 15016 16600 15068 16652
rect 16396 16600 16448 16652
rect 19248 16668 19300 16720
rect 20720 16668 20772 16720
rect 21456 16668 21508 16720
rect 18880 16600 18932 16652
rect 18972 16643 19024 16652
rect 18972 16609 18981 16643
rect 18981 16609 19015 16643
rect 19015 16609 19024 16643
rect 18972 16600 19024 16609
rect 19708 16600 19760 16652
rect 14280 16532 14332 16584
rect 15936 16532 15988 16584
rect 16120 16532 16172 16584
rect 16304 16532 16356 16584
rect 17868 16532 17920 16584
rect 9036 16464 9088 16516
rect 10876 16464 10928 16516
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 8300 16439 8352 16448
rect 8300 16405 8309 16439
rect 8309 16405 8343 16439
rect 8343 16405 8352 16439
rect 8300 16396 8352 16405
rect 8760 16396 8812 16448
rect 9680 16396 9732 16448
rect 10508 16396 10560 16448
rect 11796 16439 11848 16448
rect 11796 16405 11805 16439
rect 11805 16405 11839 16439
rect 11839 16405 11848 16439
rect 11796 16396 11848 16405
rect 11980 16396 12032 16448
rect 13912 16464 13964 16516
rect 14740 16507 14792 16516
rect 14740 16473 14749 16507
rect 14749 16473 14783 16507
rect 14783 16473 14792 16507
rect 14740 16464 14792 16473
rect 14924 16464 14976 16516
rect 17684 16464 17736 16516
rect 14004 16396 14056 16448
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 14280 16439 14332 16448
rect 14280 16405 14289 16439
rect 14289 16405 14323 16439
rect 14323 16405 14332 16439
rect 14280 16396 14332 16405
rect 15292 16396 15344 16448
rect 18328 16396 18380 16448
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 18972 16396 19024 16448
rect 19984 16396 20036 16448
rect 20996 16600 21048 16652
rect 21548 16532 21600 16584
rect 21732 16600 21784 16652
rect 22100 16600 22152 16652
rect 22560 16736 22612 16788
rect 23572 16736 23624 16788
rect 23664 16736 23716 16788
rect 24124 16736 24176 16788
rect 25044 16736 25096 16788
rect 27620 16736 27672 16788
rect 28908 16736 28960 16788
rect 29460 16736 29512 16788
rect 29644 16779 29696 16788
rect 29644 16745 29653 16779
rect 29653 16745 29687 16779
rect 29687 16745 29696 16779
rect 29644 16736 29696 16745
rect 31300 16736 31352 16788
rect 35164 16736 35216 16788
rect 22468 16600 22520 16652
rect 24860 16668 24912 16720
rect 26608 16668 26660 16720
rect 30472 16668 30524 16720
rect 23296 16532 23348 16584
rect 23940 16643 23992 16652
rect 23940 16609 23949 16643
rect 23949 16609 23983 16643
rect 23983 16609 23992 16643
rect 23940 16600 23992 16609
rect 21916 16464 21968 16516
rect 22284 16464 22336 16516
rect 22744 16464 22796 16516
rect 23848 16532 23900 16584
rect 25320 16643 25372 16652
rect 25320 16609 25329 16643
rect 25329 16609 25363 16643
rect 25363 16609 25372 16643
rect 25320 16600 25372 16609
rect 26516 16643 26568 16652
rect 26516 16609 26525 16643
rect 26525 16609 26559 16643
rect 26559 16609 26568 16643
rect 26516 16600 26568 16609
rect 26792 16600 26844 16652
rect 27436 16600 27488 16652
rect 27988 16600 28040 16652
rect 29184 16600 29236 16652
rect 29644 16600 29696 16652
rect 25136 16532 25188 16584
rect 27160 16532 27212 16584
rect 27252 16532 27304 16584
rect 28356 16532 28408 16584
rect 28908 16532 28960 16584
rect 29736 16532 29788 16584
rect 30656 16643 30708 16652
rect 30656 16609 30665 16643
rect 30665 16609 30699 16643
rect 30699 16609 30708 16643
rect 30656 16600 30708 16609
rect 31392 16600 31444 16652
rect 32312 16600 32364 16652
rect 37832 16668 37884 16720
rect 33876 16600 33928 16652
rect 32588 16532 32640 16584
rect 33324 16532 33376 16584
rect 34612 16532 34664 16584
rect 22468 16396 22520 16448
rect 22836 16396 22888 16448
rect 24768 16439 24820 16448
rect 24768 16405 24777 16439
rect 24777 16405 24811 16439
rect 24811 16405 24820 16439
rect 24768 16396 24820 16405
rect 25136 16439 25188 16448
rect 25136 16405 25145 16439
rect 25145 16405 25179 16439
rect 25179 16405 25188 16439
rect 25136 16396 25188 16405
rect 25412 16396 25464 16448
rect 25504 16396 25556 16448
rect 25688 16396 25740 16448
rect 25780 16396 25832 16448
rect 26608 16396 26660 16448
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 28724 16464 28776 16516
rect 28448 16396 28500 16448
rect 28816 16396 28868 16448
rect 29092 16439 29144 16448
rect 29092 16405 29101 16439
rect 29101 16405 29135 16439
rect 29135 16405 29144 16439
rect 29092 16396 29144 16405
rect 34980 16507 35032 16516
rect 34980 16473 34989 16507
rect 34989 16473 35023 16507
rect 35023 16473 35032 16507
rect 34980 16464 35032 16473
rect 30104 16396 30156 16448
rect 33232 16396 33284 16448
rect 35072 16439 35124 16448
rect 35072 16405 35081 16439
rect 35081 16405 35115 16439
rect 35115 16405 35124 16439
rect 35072 16396 35124 16405
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 8668 16192 8720 16244
rect 9036 16192 9088 16244
rect 9220 16235 9272 16244
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 4712 16124 4764 16176
rect 9496 16192 9548 16244
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 6552 16056 6604 16108
rect 6644 16056 6696 16108
rect 7932 16099 7984 16108
rect 7932 16065 7941 16099
rect 7941 16065 7975 16099
rect 7975 16065 7984 16099
rect 7932 16056 7984 16065
rect 1308 15988 1360 16040
rect 4712 15988 4764 16040
rect 7656 15988 7708 16040
rect 1860 15920 1912 15972
rect 7564 15963 7616 15972
rect 7564 15929 7573 15963
rect 7573 15929 7607 15963
rect 7607 15929 7616 15963
rect 7564 15920 7616 15929
rect 7748 15920 7800 15972
rect 10968 16192 11020 16244
rect 11428 16192 11480 16244
rect 12992 16192 13044 16244
rect 14372 16192 14424 16244
rect 14648 16192 14700 16244
rect 10600 16124 10652 16176
rect 11060 16167 11112 16176
rect 11060 16133 11069 16167
rect 11069 16133 11103 16167
rect 11103 16133 11112 16167
rect 11060 16124 11112 16133
rect 11980 16124 12032 16176
rect 12900 16124 12952 16176
rect 14280 16124 14332 16176
rect 12072 16056 12124 16108
rect 9588 15988 9640 16040
rect 10600 16031 10652 16040
rect 10600 15997 10609 16031
rect 10609 15997 10643 16031
rect 10643 15997 10652 16031
rect 10600 15988 10652 15997
rect 11428 15988 11480 16040
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13912 15988 13964 16040
rect 4988 15852 5040 15904
rect 8760 15895 8812 15904
rect 8760 15861 8769 15895
rect 8769 15861 8803 15895
rect 8803 15861 8812 15895
rect 8760 15852 8812 15861
rect 9680 15920 9732 15972
rect 15200 16056 15252 16108
rect 18972 16192 19024 16244
rect 19432 16192 19484 16244
rect 23480 16192 23532 16244
rect 17224 16124 17276 16176
rect 17684 16124 17736 16176
rect 22284 16124 22336 16176
rect 23388 16124 23440 16176
rect 15936 15988 15988 16040
rect 16856 16031 16908 16040
rect 16856 15997 16865 16031
rect 16865 15997 16899 16031
rect 16899 15997 16908 16031
rect 16856 15988 16908 15997
rect 17132 16031 17184 16040
rect 17132 15997 17141 16031
rect 17141 15997 17175 16031
rect 17175 15997 17184 16031
rect 17132 15988 17184 15997
rect 17500 15988 17552 16040
rect 19432 16056 19484 16108
rect 21456 16056 21508 16108
rect 22100 16056 22152 16108
rect 23112 16056 23164 16108
rect 23204 16099 23256 16108
rect 23204 16065 23213 16099
rect 23213 16065 23247 16099
rect 23247 16065 23256 16099
rect 23204 16056 23256 16065
rect 23572 16056 23624 16108
rect 23940 16192 23992 16244
rect 27160 16192 27212 16244
rect 31208 16192 31260 16244
rect 31852 16192 31904 16244
rect 32680 16192 32732 16244
rect 26700 16124 26752 16176
rect 24676 16056 24728 16108
rect 27068 16056 27120 16108
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27528 16124 27580 16176
rect 18972 15988 19024 16040
rect 20628 15988 20680 16040
rect 21180 16031 21232 16040
rect 21180 15997 21189 16031
rect 21189 15997 21223 16031
rect 21223 15997 21232 16031
rect 21180 15988 21232 15997
rect 22744 15988 22796 16040
rect 24768 15988 24820 16040
rect 28264 16099 28316 16108
rect 28264 16065 28273 16099
rect 28273 16065 28307 16099
rect 28307 16065 28316 16099
rect 28264 16056 28316 16065
rect 30104 16056 30156 16108
rect 30564 16056 30616 16108
rect 30932 16056 30984 16108
rect 31668 16056 31720 16108
rect 31760 16099 31812 16108
rect 31760 16065 31769 16099
rect 31769 16065 31803 16099
rect 31803 16065 31812 16099
rect 31760 16056 31812 16065
rect 14464 15963 14516 15972
rect 14464 15929 14473 15963
rect 14473 15929 14507 15963
rect 14507 15929 14516 15963
rect 14464 15920 14516 15929
rect 15016 15920 15068 15972
rect 9220 15852 9272 15904
rect 10048 15895 10100 15904
rect 10048 15861 10057 15895
rect 10057 15861 10091 15895
rect 10091 15861 10100 15895
rect 10048 15852 10100 15861
rect 11796 15852 11848 15904
rect 12440 15852 12492 15904
rect 13820 15852 13872 15904
rect 14188 15852 14240 15904
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 16304 15895 16356 15904
rect 16304 15861 16313 15895
rect 16313 15861 16347 15895
rect 16347 15861 16356 15895
rect 16304 15852 16356 15861
rect 19064 15963 19116 15972
rect 19064 15929 19073 15963
rect 19073 15929 19107 15963
rect 19107 15929 19116 15963
rect 19064 15920 19116 15929
rect 19248 15920 19300 15972
rect 21640 15963 21692 15972
rect 21640 15929 21649 15963
rect 21649 15929 21683 15963
rect 21683 15929 21692 15963
rect 21640 15920 21692 15929
rect 22284 15920 22336 15972
rect 19984 15852 20036 15904
rect 20076 15852 20128 15904
rect 22560 15852 22612 15904
rect 23020 15895 23072 15904
rect 23020 15861 23029 15895
rect 23029 15861 23063 15895
rect 23063 15861 23072 15895
rect 23020 15852 23072 15861
rect 23112 15852 23164 15904
rect 24400 15895 24452 15904
rect 24400 15861 24409 15895
rect 24409 15861 24443 15895
rect 24443 15861 24452 15895
rect 24400 15852 24452 15861
rect 24492 15852 24544 15904
rect 24768 15852 24820 15904
rect 26148 15920 26200 15972
rect 31484 15988 31536 16040
rect 36452 15988 36504 16040
rect 32404 15920 32456 15972
rect 29000 15852 29052 15904
rect 29552 15852 29604 15904
rect 31576 15895 31628 15904
rect 31576 15861 31585 15895
rect 31585 15861 31619 15895
rect 31619 15861 31628 15895
rect 31576 15852 31628 15861
rect 31668 15852 31720 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 1124 15648 1176 15700
rect 2872 15648 2924 15700
rect 6368 15648 6420 15700
rect 3608 15623 3660 15632
rect 3608 15589 3617 15623
rect 3617 15589 3651 15623
rect 3651 15589 3660 15623
rect 3608 15580 3660 15589
rect 1308 15512 1360 15564
rect 2320 15512 2372 15564
rect 4804 15512 4856 15564
rect 6276 15580 6328 15632
rect 14280 15648 14332 15700
rect 15016 15648 15068 15700
rect 15752 15648 15804 15700
rect 16672 15648 16724 15700
rect 18972 15648 19024 15700
rect 19340 15648 19392 15700
rect 19892 15648 19944 15700
rect 7656 15512 7708 15564
rect 1860 15444 1912 15496
rect 940 15376 992 15428
rect 4896 15444 4948 15496
rect 6736 15444 6788 15496
rect 9496 15580 9548 15632
rect 9404 15512 9456 15564
rect 9864 15580 9916 15632
rect 16396 15580 16448 15632
rect 14004 15512 14056 15564
rect 18328 15580 18380 15632
rect 3424 15419 3476 15428
rect 3424 15385 3433 15419
rect 3433 15385 3467 15419
rect 3467 15385 3476 15419
rect 3424 15376 3476 15385
rect 3608 15376 3660 15428
rect 2412 15308 2464 15360
rect 4068 15308 4120 15360
rect 6552 15376 6604 15428
rect 6828 15376 6880 15428
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 7932 15419 7984 15428
rect 7932 15385 7941 15419
rect 7941 15385 7975 15419
rect 7975 15385 7984 15419
rect 7932 15376 7984 15385
rect 6184 15308 6236 15360
rect 7196 15308 7248 15360
rect 9312 15444 9364 15496
rect 11336 15444 11388 15496
rect 9036 15376 9088 15428
rect 13268 15444 13320 15496
rect 14648 15444 14700 15496
rect 16948 15487 17000 15496
rect 16948 15453 16957 15487
rect 16957 15453 16991 15487
rect 16991 15453 17000 15487
rect 16948 15444 17000 15453
rect 18788 15512 18840 15564
rect 20076 15512 20128 15564
rect 20168 15555 20220 15564
rect 20168 15521 20177 15555
rect 20177 15521 20211 15555
rect 20211 15521 20220 15555
rect 20168 15512 20220 15521
rect 20536 15623 20588 15632
rect 20536 15589 20545 15623
rect 20545 15589 20579 15623
rect 20579 15589 20588 15623
rect 20536 15580 20588 15589
rect 20904 15512 20956 15564
rect 19248 15444 19300 15496
rect 19708 15444 19760 15496
rect 22008 15512 22060 15564
rect 22284 15512 22336 15564
rect 23940 15555 23992 15564
rect 23940 15521 23949 15555
rect 23949 15521 23983 15555
rect 23983 15521 23992 15555
rect 23940 15512 23992 15521
rect 25136 15648 25188 15700
rect 24860 15555 24912 15564
rect 24860 15521 24869 15555
rect 24869 15521 24903 15555
rect 24903 15521 24912 15555
rect 24860 15512 24912 15521
rect 25688 15512 25740 15564
rect 26608 15512 26660 15564
rect 27804 15691 27856 15700
rect 27804 15657 27813 15691
rect 27813 15657 27847 15691
rect 27847 15657 27856 15691
rect 27804 15648 27856 15657
rect 27988 15691 28040 15700
rect 27988 15657 27997 15691
rect 27997 15657 28031 15691
rect 28031 15657 28040 15691
rect 27988 15648 28040 15657
rect 27344 15580 27396 15632
rect 31668 15648 31720 15700
rect 31760 15648 31812 15700
rect 28264 15580 28316 15632
rect 31852 15580 31904 15632
rect 32220 15580 32272 15632
rect 23204 15444 23256 15496
rect 8944 15308 8996 15360
rect 9588 15351 9640 15360
rect 9588 15317 9597 15351
rect 9597 15317 9631 15351
rect 9631 15317 9640 15351
rect 9588 15308 9640 15317
rect 9680 15308 9732 15360
rect 10692 15308 10744 15360
rect 11888 15419 11940 15428
rect 11888 15385 11897 15419
rect 11897 15385 11931 15419
rect 11931 15385 11940 15419
rect 11888 15376 11940 15385
rect 12624 15376 12676 15428
rect 13176 15376 13228 15428
rect 14556 15376 14608 15428
rect 15108 15376 15160 15428
rect 15660 15376 15712 15428
rect 16856 15376 16908 15428
rect 17684 15376 17736 15428
rect 20812 15376 20864 15428
rect 21916 15376 21968 15428
rect 22560 15376 22612 15428
rect 24216 15376 24268 15428
rect 25412 15444 25464 15496
rect 27712 15487 27764 15496
rect 27712 15453 27721 15487
rect 27721 15453 27755 15487
rect 27755 15453 27764 15487
rect 27712 15444 27764 15453
rect 11152 15308 11204 15360
rect 11704 15308 11756 15360
rect 12532 15308 12584 15360
rect 14096 15351 14148 15360
rect 14096 15317 14105 15351
rect 14105 15317 14139 15351
rect 14139 15317 14148 15351
rect 14096 15308 14148 15317
rect 16764 15308 16816 15360
rect 18512 15308 18564 15360
rect 18696 15351 18748 15360
rect 18696 15317 18705 15351
rect 18705 15317 18739 15351
rect 18739 15317 18748 15351
rect 18696 15308 18748 15317
rect 20444 15308 20496 15360
rect 21088 15308 21140 15360
rect 21640 15308 21692 15360
rect 23388 15308 23440 15360
rect 23756 15351 23808 15360
rect 23756 15317 23765 15351
rect 23765 15317 23799 15351
rect 23799 15317 23808 15351
rect 23756 15308 23808 15317
rect 24768 15308 24820 15360
rect 27252 15376 27304 15428
rect 26332 15308 26384 15360
rect 37280 15512 37332 15564
rect 27988 15444 28040 15496
rect 28632 15487 28684 15496
rect 28632 15453 28641 15487
rect 28641 15453 28675 15487
rect 28675 15453 28684 15487
rect 28632 15444 28684 15453
rect 29644 15444 29696 15496
rect 30012 15487 30064 15496
rect 30012 15453 30021 15487
rect 30021 15453 30055 15487
rect 30055 15453 30064 15487
rect 30012 15444 30064 15453
rect 30104 15444 30156 15496
rect 28724 15308 28776 15360
rect 31116 15376 31168 15428
rect 31668 15444 31720 15496
rect 32036 15444 32088 15496
rect 33876 15444 33928 15496
rect 38752 15444 38804 15496
rect 41236 15376 41288 15428
rect 31024 15308 31076 15360
rect 32220 15308 32272 15360
rect 32496 15308 32548 15360
rect 32588 15351 32640 15360
rect 32588 15317 32597 15351
rect 32597 15317 32631 15351
rect 32631 15317 32640 15351
rect 32588 15308 32640 15317
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 4436 15104 4488 15156
rect 5724 15147 5776 15156
rect 5724 15113 5733 15147
rect 5733 15113 5767 15147
rect 5767 15113 5776 15147
rect 5724 15104 5776 15113
rect 7656 15104 7708 15156
rect 7932 15104 7984 15156
rect 8024 15147 8076 15156
rect 8024 15113 8033 15147
rect 8033 15113 8067 15147
rect 8067 15113 8076 15147
rect 8024 15104 8076 15113
rect 8760 15104 8812 15156
rect 10600 15104 10652 15156
rect 11704 15104 11756 15156
rect 12256 15147 12308 15156
rect 12256 15113 12265 15147
rect 12265 15113 12299 15147
rect 12299 15113 12308 15147
rect 12256 15104 12308 15113
rect 14096 15104 14148 15156
rect 14188 15104 14240 15156
rect 14832 15104 14884 15156
rect 16028 15104 16080 15156
rect 16488 15104 16540 15156
rect 16764 15104 16816 15156
rect 17316 15104 17368 15156
rect 18236 15104 18288 15156
rect 664 15036 716 15088
rect 5540 15036 5592 15088
rect 8944 15036 8996 15088
rect 10416 15036 10468 15088
rect 2688 14968 2740 15020
rect 1308 14900 1360 14952
rect 3700 14968 3752 15020
rect 3976 14900 4028 14952
rect 4068 14900 4120 14952
rect 4712 14943 4764 14952
rect 4712 14909 4721 14943
rect 4721 14909 4755 14943
rect 4755 14909 4764 14943
rect 4712 14900 4764 14909
rect 5356 14900 5408 14952
rect 6828 14968 6880 15020
rect 7656 14968 7708 15020
rect 9220 14968 9272 15020
rect 7104 14900 7156 14952
rect 8576 14900 8628 14952
rect 9588 14900 9640 14952
rect 9864 14968 9916 15020
rect 10968 14968 11020 15020
rect 10416 14900 10468 14952
rect 10600 14900 10652 14952
rect 1768 14832 1820 14884
rect 8024 14832 8076 14884
rect 13176 15036 13228 15088
rect 13636 15036 13688 15088
rect 20628 15104 20680 15156
rect 21548 15104 21600 15156
rect 28632 15104 28684 15156
rect 29184 15104 29236 15156
rect 33508 15104 33560 15156
rect 20996 15036 21048 15088
rect 23848 15036 23900 15088
rect 24308 15036 24360 15088
rect 12440 14968 12492 15020
rect 13912 14968 13964 15020
rect 14188 14968 14240 15020
rect 12532 14900 12584 14952
rect 14464 14900 14516 14952
rect 15016 14943 15068 14952
rect 15016 14909 15025 14943
rect 15025 14909 15059 14943
rect 15059 14909 15068 14943
rect 15016 14900 15068 14909
rect 16580 14968 16632 15020
rect 18788 14900 18840 14952
rect 19064 14900 19116 14952
rect 2688 14764 2740 14816
rect 2780 14764 2832 14816
rect 3424 14807 3476 14816
rect 3424 14773 3433 14807
rect 3433 14773 3467 14807
rect 3467 14773 3476 14807
rect 3424 14764 3476 14773
rect 5080 14764 5132 14816
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 5540 14764 5592 14816
rect 6000 14764 6052 14816
rect 6736 14764 6788 14816
rect 7196 14807 7248 14816
rect 7196 14773 7205 14807
rect 7205 14773 7239 14807
rect 7239 14773 7248 14807
rect 7196 14764 7248 14773
rect 7288 14764 7340 14816
rect 8760 14807 8812 14816
rect 8760 14773 8769 14807
rect 8769 14773 8803 14807
rect 8803 14773 8812 14807
rect 8760 14764 8812 14773
rect 9036 14764 9088 14816
rect 9772 14764 9824 14816
rect 9864 14764 9916 14816
rect 10600 14764 10652 14816
rect 17132 14832 17184 14884
rect 18052 14832 18104 14884
rect 18236 14832 18288 14884
rect 18512 14832 18564 14884
rect 11796 14807 11848 14816
rect 11796 14773 11805 14807
rect 11805 14773 11839 14807
rect 11839 14773 11848 14807
rect 11796 14764 11848 14773
rect 13268 14764 13320 14816
rect 13636 14764 13688 14816
rect 14372 14764 14424 14816
rect 14648 14764 14700 14816
rect 18696 14764 18748 14816
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 24216 14968 24268 15020
rect 24768 15036 24820 15088
rect 27712 15036 27764 15088
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 27620 14968 27672 14977
rect 28724 15011 28776 15020
rect 28724 14977 28733 15011
rect 28733 14977 28767 15011
rect 28767 14977 28776 15011
rect 28724 14968 28776 14977
rect 29460 14968 29512 15020
rect 30932 15011 30984 15020
rect 30932 14977 30941 15011
rect 30941 14977 30975 15011
rect 30975 14977 30984 15011
rect 30932 14968 30984 14977
rect 31116 15036 31168 15088
rect 41420 15036 41472 15088
rect 33600 14968 33652 15020
rect 19708 14943 19760 14952
rect 19708 14909 19717 14943
rect 19717 14909 19751 14943
rect 19751 14909 19760 14943
rect 19708 14900 19760 14909
rect 19984 14900 20036 14952
rect 21088 14832 21140 14884
rect 21916 14832 21968 14884
rect 20628 14764 20680 14816
rect 21732 14764 21784 14816
rect 22560 14943 22612 14952
rect 22560 14909 22569 14943
rect 22569 14909 22603 14943
rect 22603 14909 22612 14943
rect 22560 14900 22612 14909
rect 23296 14900 23348 14952
rect 28448 14900 28500 14952
rect 31300 14900 31352 14952
rect 24860 14764 24912 14816
rect 26884 14832 26936 14884
rect 27252 14832 27304 14884
rect 44824 14832 44876 14884
rect 25320 14764 25372 14816
rect 25872 14764 25924 14816
rect 26608 14807 26660 14816
rect 26608 14773 26617 14807
rect 26617 14773 26651 14807
rect 26651 14773 26660 14807
rect 26608 14764 26660 14773
rect 27068 14807 27120 14816
rect 27068 14773 27077 14807
rect 27077 14773 27111 14807
rect 27111 14773 27120 14807
rect 27068 14764 27120 14773
rect 29368 14807 29420 14816
rect 29368 14773 29377 14807
rect 29377 14773 29411 14807
rect 29411 14773 29420 14807
rect 29368 14764 29420 14773
rect 30380 14764 30432 14816
rect 31576 14807 31628 14816
rect 31576 14773 31585 14807
rect 31585 14773 31619 14807
rect 31619 14773 31628 14807
rect 31576 14764 31628 14773
rect 31668 14764 31720 14816
rect 33600 14764 33652 14816
rect 40408 14764 40460 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 1768 14560 1820 14612
rect 2136 14560 2188 14612
rect 3516 14560 3568 14612
rect 1308 14424 1360 14476
rect 6276 14560 6328 14612
rect 6644 14560 6696 14612
rect 7196 14492 7248 14544
rect 7840 14560 7892 14612
rect 9404 14560 9456 14612
rect 10232 14560 10284 14612
rect 12440 14560 12492 14612
rect 12532 14560 12584 14612
rect 13912 14603 13964 14612
rect 13912 14569 13921 14603
rect 13921 14569 13955 14603
rect 13955 14569 13964 14603
rect 13912 14560 13964 14569
rect 8668 14492 8720 14544
rect 18788 14560 18840 14612
rect 22560 14560 22612 14612
rect 29000 14560 29052 14612
rect 29736 14560 29788 14612
rect 30932 14560 30984 14612
rect 21548 14492 21600 14544
rect 5080 14467 5132 14476
rect 5080 14433 5089 14467
rect 5089 14433 5123 14467
rect 5123 14433 5132 14467
rect 5080 14424 5132 14433
rect 5724 14424 5776 14476
rect 3608 14356 3660 14408
rect 4804 14356 4856 14408
rect 4988 14331 5040 14340
rect 4988 14297 4997 14331
rect 4997 14297 5031 14331
rect 5031 14297 5040 14331
rect 4988 14288 5040 14297
rect 5632 14288 5684 14340
rect 3608 14263 3660 14272
rect 3608 14229 3617 14263
rect 3617 14229 3651 14263
rect 3651 14229 3660 14263
rect 3608 14220 3660 14229
rect 5448 14220 5500 14272
rect 5540 14220 5592 14272
rect 6552 14288 6604 14340
rect 6368 14220 6420 14272
rect 7932 14288 7984 14340
rect 8484 14356 8536 14408
rect 8944 14399 8996 14408
rect 8944 14365 8953 14399
rect 8953 14365 8987 14399
rect 8987 14365 8996 14399
rect 8944 14356 8996 14365
rect 9588 14356 9640 14408
rect 10692 14356 10744 14408
rect 10968 14467 11020 14476
rect 10968 14433 10977 14467
rect 10977 14433 11011 14467
rect 11011 14433 11020 14467
rect 10968 14424 11020 14433
rect 14188 14467 14240 14476
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 14556 14424 14608 14476
rect 15384 14424 15436 14476
rect 16948 14424 17000 14476
rect 19708 14424 19760 14476
rect 20260 14424 20312 14476
rect 21364 14424 21416 14476
rect 21456 14424 21508 14476
rect 24216 14492 24268 14544
rect 24584 14492 24636 14544
rect 10600 14288 10652 14340
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 13360 14356 13412 14408
rect 13912 14356 13964 14408
rect 14648 14399 14700 14408
rect 14648 14365 14657 14399
rect 14657 14365 14691 14399
rect 14691 14365 14700 14399
rect 14648 14356 14700 14365
rect 18696 14356 18748 14408
rect 19524 14356 19576 14408
rect 19800 14356 19852 14408
rect 11428 14331 11480 14340
rect 11428 14297 11437 14331
rect 11437 14297 11471 14331
rect 11471 14297 11480 14331
rect 11428 14288 11480 14297
rect 7564 14220 7616 14272
rect 10692 14220 10744 14272
rect 12624 14288 12676 14340
rect 13820 14288 13872 14340
rect 15660 14288 15712 14340
rect 16948 14288 17000 14340
rect 17316 14288 17368 14340
rect 17408 14331 17460 14340
rect 17408 14297 17417 14331
rect 17417 14297 17451 14331
rect 17451 14297 17460 14331
rect 17408 14288 17460 14297
rect 17684 14288 17736 14340
rect 19064 14288 19116 14340
rect 19432 14331 19484 14340
rect 19432 14297 19441 14331
rect 19441 14297 19475 14331
rect 19475 14297 19484 14331
rect 19432 14288 19484 14297
rect 21916 14467 21968 14476
rect 21916 14433 21925 14467
rect 21925 14433 21959 14467
rect 21959 14433 21968 14467
rect 21916 14424 21968 14433
rect 22284 14424 22336 14476
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 23480 14424 23532 14476
rect 24492 14424 24544 14476
rect 22100 14356 22152 14408
rect 24584 14356 24636 14408
rect 25504 14356 25556 14408
rect 26792 14492 26844 14544
rect 28448 14492 28500 14544
rect 28816 14492 28868 14544
rect 42524 14560 42576 14612
rect 31852 14492 31904 14544
rect 37648 14492 37700 14544
rect 25872 14467 25924 14476
rect 25872 14433 25881 14467
rect 25881 14433 25915 14467
rect 25915 14433 25924 14467
rect 25872 14424 25924 14433
rect 26700 14424 26752 14476
rect 30288 14424 30340 14476
rect 30748 14424 30800 14476
rect 29368 14356 29420 14408
rect 12808 14220 12860 14272
rect 13084 14220 13136 14272
rect 15844 14220 15896 14272
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 17500 14220 17552 14272
rect 18052 14220 18104 14272
rect 19892 14220 19944 14272
rect 21364 14263 21416 14272
rect 21364 14229 21373 14263
rect 21373 14229 21407 14263
rect 21407 14229 21416 14263
rect 21364 14220 21416 14229
rect 21732 14220 21784 14272
rect 22284 14288 22336 14340
rect 23296 14288 23348 14340
rect 24216 14288 24268 14340
rect 29736 14399 29788 14408
rect 29736 14365 29745 14399
rect 29745 14365 29779 14399
rect 29779 14365 29788 14399
rect 29736 14356 29788 14365
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 46204 14288 46256 14340
rect 21916 14220 21968 14272
rect 22468 14220 22520 14272
rect 22928 14220 22980 14272
rect 23112 14220 23164 14272
rect 23756 14220 23808 14272
rect 24308 14220 24360 14272
rect 24768 14263 24820 14272
rect 24768 14229 24777 14263
rect 24777 14229 24811 14263
rect 24811 14229 24820 14263
rect 24768 14220 24820 14229
rect 24952 14220 25004 14272
rect 25688 14263 25740 14272
rect 25688 14229 25697 14263
rect 25697 14229 25731 14263
rect 25731 14229 25740 14263
rect 25688 14220 25740 14229
rect 26516 14220 26568 14272
rect 26700 14220 26752 14272
rect 27712 14220 27764 14272
rect 28816 14220 28868 14272
rect 29276 14220 29328 14272
rect 29368 14263 29420 14272
rect 29368 14229 29377 14263
rect 29377 14229 29411 14263
rect 29411 14229 29420 14263
rect 29368 14220 29420 14229
rect 30288 14220 30340 14272
rect 47860 14220 47912 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 3608 14016 3660 14068
rect 4528 14016 4580 14068
rect 4988 14016 5040 14068
rect 3884 13948 3936 14000
rect 296 13880 348 13932
rect 1492 13880 1544 13932
rect 1584 13923 1636 13932
rect 1584 13889 1593 13923
rect 1593 13889 1627 13923
rect 1627 13889 1636 13923
rect 1584 13880 1636 13889
rect 2136 13880 2188 13932
rect 4160 13948 4212 14000
rect 5540 13948 5592 14000
rect 6920 14016 6972 14068
rect 7748 14016 7800 14068
rect 8024 14016 8076 14068
rect 8392 14016 8444 14068
rect 9680 14016 9732 14068
rect 6368 13948 6420 14000
rect 6644 13948 6696 14000
rect 13268 14016 13320 14068
rect 16672 14059 16724 14068
rect 16672 14025 16681 14059
rect 16681 14025 16715 14059
rect 16715 14025 16724 14059
rect 16672 14016 16724 14025
rect 17132 14016 17184 14068
rect 18052 14016 18104 14068
rect 19800 14016 19852 14068
rect 20260 14016 20312 14068
rect 20812 14016 20864 14068
rect 20904 14016 20956 14068
rect 21548 14016 21600 14068
rect 21732 14016 21784 14068
rect 22284 14016 22336 14068
rect 22468 14016 22520 14068
rect 22744 14016 22796 14068
rect 23480 14016 23532 14068
rect 23572 14016 23624 14068
rect 24216 14059 24268 14068
rect 24216 14025 24225 14059
rect 24225 14025 24259 14059
rect 24259 14025 24268 14059
rect 24216 14016 24268 14025
rect 25504 14059 25556 14068
rect 25504 14025 25513 14059
rect 25513 14025 25547 14059
rect 25547 14025 25556 14059
rect 25504 14016 25556 14025
rect 25688 14016 25740 14068
rect 26424 14016 26476 14068
rect 29276 14016 29328 14068
rect 1308 13812 1360 13864
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 3516 13812 3568 13821
rect 6276 13880 6328 13932
rect 7196 13812 7248 13864
rect 7564 13880 7616 13932
rect 8392 13880 8444 13932
rect 7656 13812 7708 13864
rect 8576 13880 8628 13932
rect 11152 13948 11204 14000
rect 14648 13948 14700 14000
rect 3792 13744 3844 13796
rect 6552 13744 6604 13796
rect 3976 13676 4028 13728
rect 4712 13676 4764 13728
rect 5356 13676 5408 13728
rect 6276 13676 6328 13728
rect 6644 13676 6696 13728
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 10140 13812 10192 13864
rect 11244 13880 11296 13932
rect 13636 13880 13688 13932
rect 10968 13744 11020 13796
rect 11336 13744 11388 13796
rect 12532 13744 12584 13796
rect 12900 13812 12952 13864
rect 13268 13744 13320 13796
rect 14924 13880 14976 13932
rect 15200 13880 15252 13932
rect 17040 13880 17092 13932
rect 17316 13948 17368 14000
rect 17684 13948 17736 14000
rect 15016 13812 15068 13864
rect 15752 13855 15804 13864
rect 15752 13821 15761 13855
rect 15761 13821 15795 13855
rect 15795 13821 15804 13855
rect 15752 13812 15804 13821
rect 16396 13812 16448 13864
rect 20628 13948 20680 14000
rect 22560 13948 22612 14000
rect 24952 13948 25004 14000
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 21456 13880 21508 13932
rect 21916 13923 21968 13932
rect 21916 13889 21925 13923
rect 21925 13889 21959 13923
rect 21959 13889 21968 13923
rect 21916 13880 21968 13889
rect 10140 13676 10192 13728
rect 10600 13676 10652 13728
rect 11060 13719 11112 13728
rect 11060 13685 11069 13719
rect 11069 13685 11103 13719
rect 11103 13685 11112 13719
rect 11060 13676 11112 13685
rect 11612 13676 11664 13728
rect 11888 13676 11940 13728
rect 12072 13676 12124 13728
rect 13084 13676 13136 13728
rect 13636 13676 13688 13728
rect 15568 13744 15620 13796
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 18880 13812 18932 13821
rect 19524 13812 19576 13864
rect 19984 13812 20036 13864
rect 20076 13855 20128 13864
rect 20076 13821 20085 13855
rect 20085 13821 20119 13855
rect 20119 13821 20128 13855
rect 20076 13812 20128 13821
rect 18604 13744 18656 13796
rect 20260 13744 20312 13796
rect 20812 13744 20864 13796
rect 14096 13676 14148 13728
rect 18144 13676 18196 13728
rect 18696 13676 18748 13728
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23112 13812 23164 13821
rect 22008 13744 22060 13796
rect 22744 13744 22796 13796
rect 23940 13812 23992 13864
rect 24584 13880 24636 13932
rect 24768 13812 24820 13864
rect 24860 13812 24912 13864
rect 25596 13812 25648 13864
rect 26608 13880 26660 13932
rect 28540 13923 28592 13932
rect 28540 13889 28549 13923
rect 28549 13889 28583 13923
rect 28583 13889 28592 13923
rect 28540 13880 28592 13889
rect 29828 13923 29880 13932
rect 29828 13889 29837 13923
rect 29837 13889 29871 13923
rect 29871 13889 29880 13923
rect 29828 13880 29880 13889
rect 40040 13948 40092 14000
rect 42800 13948 42852 14000
rect 30472 13923 30524 13932
rect 30472 13889 30481 13923
rect 30481 13889 30515 13923
rect 30515 13889 30524 13923
rect 30472 13880 30524 13889
rect 23296 13744 23348 13796
rect 25228 13744 25280 13796
rect 25964 13744 26016 13796
rect 28908 13744 28960 13796
rect 36544 13744 36596 13796
rect 22652 13719 22704 13728
rect 22652 13685 22661 13719
rect 22661 13685 22695 13719
rect 22695 13685 22704 13719
rect 22652 13676 22704 13685
rect 22928 13676 22980 13728
rect 23480 13676 23532 13728
rect 23756 13676 23808 13728
rect 24032 13676 24084 13728
rect 24952 13676 25004 13728
rect 27804 13719 27856 13728
rect 27804 13685 27813 13719
rect 27813 13685 27847 13719
rect 27847 13685 27856 13719
rect 27804 13676 27856 13685
rect 29920 13676 29972 13728
rect 39672 13676 39724 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 3792 13472 3844 13524
rect 4252 13472 4304 13524
rect 4344 13472 4396 13524
rect 6092 13472 6144 13524
rect 5172 13404 5224 13456
rect 9956 13404 10008 13456
rect 2044 13379 2096 13388
rect 2044 13345 2053 13379
rect 2053 13345 2087 13379
rect 2087 13345 2096 13379
rect 2044 13336 2096 13345
rect 3424 13336 3476 13388
rect 3884 13336 3936 13388
rect 4988 13379 5040 13388
rect 4988 13345 4997 13379
rect 4997 13345 5031 13379
rect 5031 13345 5040 13379
rect 4988 13336 5040 13345
rect 5264 13336 5316 13388
rect 6276 13379 6328 13388
rect 6276 13345 6285 13379
rect 6285 13345 6319 13379
rect 6319 13345 6328 13379
rect 6276 13336 6328 13345
rect 9220 13336 9272 13388
rect 10600 13336 10652 13388
rect 11612 13472 11664 13524
rect 12716 13472 12768 13524
rect 13268 13404 13320 13456
rect 16304 13515 16356 13524
rect 16304 13481 16313 13515
rect 16313 13481 16347 13515
rect 16347 13481 16356 13515
rect 16304 13472 16356 13481
rect 16488 13515 16540 13524
rect 16488 13481 16497 13515
rect 16497 13481 16531 13515
rect 16531 13481 16540 13515
rect 16488 13472 16540 13481
rect 16672 13472 16724 13524
rect 17040 13472 17092 13524
rect 17316 13472 17368 13524
rect 16764 13404 16816 13456
rect 11796 13336 11848 13388
rect 12256 13336 12308 13388
rect 14648 13336 14700 13388
rect 14924 13336 14976 13388
rect 15016 13336 15068 13388
rect 16672 13336 16724 13388
rect 16856 13336 16908 13388
rect 17592 13379 17644 13388
rect 17592 13345 17601 13379
rect 17601 13345 17635 13379
rect 17635 13345 17644 13379
rect 17592 13336 17644 13345
rect 572 13268 624 13320
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 3240 13268 3292 13320
rect 4160 13268 4212 13320
rect 9496 13268 9548 13320
rect 10048 13268 10100 13320
rect 11520 13268 11572 13320
rect 15660 13268 15712 13320
rect 388 13200 440 13252
rect 1768 13132 1820 13184
rect 1952 13132 2004 13184
rect 3516 13132 3568 13184
rect 5080 13200 5132 13252
rect 6644 13200 6696 13252
rect 7012 13200 7064 13252
rect 7656 13200 7708 13252
rect 10876 13200 10928 13252
rect 11888 13200 11940 13252
rect 12072 13200 12124 13252
rect 5448 13132 5500 13184
rect 7748 13132 7800 13184
rect 9404 13132 9456 13184
rect 10048 13132 10100 13184
rect 10416 13132 10468 13184
rect 12624 13200 12676 13252
rect 14648 13200 14700 13252
rect 12532 13132 12584 13184
rect 13084 13132 13136 13184
rect 14004 13132 14056 13184
rect 14464 13132 14516 13184
rect 17316 13268 17368 13320
rect 17776 13268 17828 13320
rect 18512 13404 18564 13456
rect 18236 13336 18288 13388
rect 18696 13336 18748 13388
rect 19156 13472 19208 13524
rect 21916 13472 21968 13524
rect 30840 13472 30892 13524
rect 19156 13336 19208 13388
rect 19616 13379 19668 13388
rect 19616 13345 19625 13379
rect 19625 13345 19659 13379
rect 19659 13345 19668 13379
rect 19616 13336 19668 13345
rect 21548 13404 21600 13456
rect 22560 13404 22612 13456
rect 20536 13336 20588 13388
rect 22100 13336 22152 13388
rect 19708 13268 19760 13320
rect 22192 13268 22244 13320
rect 16488 13200 16540 13252
rect 16580 13200 16632 13252
rect 18696 13200 18748 13252
rect 19340 13200 19392 13252
rect 20536 13243 20588 13252
rect 20536 13209 20545 13243
rect 20545 13209 20579 13243
rect 20579 13209 20588 13243
rect 20536 13200 20588 13209
rect 20996 13200 21048 13252
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 17868 13132 17920 13184
rect 19524 13132 19576 13184
rect 26056 13404 26108 13456
rect 29736 13404 29788 13456
rect 23480 13336 23532 13388
rect 24124 13336 24176 13388
rect 24216 13336 24268 13388
rect 24584 13336 24636 13388
rect 25136 13379 25188 13388
rect 25136 13345 25145 13379
rect 25145 13345 25179 13379
rect 25179 13345 25188 13379
rect 25136 13336 25188 13345
rect 23112 13268 23164 13320
rect 24952 13311 25004 13320
rect 24952 13277 24961 13311
rect 24961 13277 24995 13311
rect 24995 13277 25004 13311
rect 24952 13268 25004 13277
rect 27804 13336 27856 13388
rect 28632 13336 28684 13388
rect 42708 13472 42760 13524
rect 26700 13268 26752 13320
rect 37556 13268 37608 13320
rect 22836 13200 22888 13252
rect 23296 13200 23348 13252
rect 28908 13243 28960 13252
rect 28908 13209 28917 13243
rect 28917 13209 28951 13243
rect 28951 13209 28960 13243
rect 28908 13200 28960 13209
rect 23480 13132 23532 13184
rect 23664 13132 23716 13184
rect 24032 13132 24084 13184
rect 26148 13132 26200 13184
rect 26240 13132 26292 13184
rect 26516 13132 26568 13184
rect 27712 13132 27764 13184
rect 27896 13132 27948 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 3700 12928 3752 12980
rect 4160 12928 4212 12980
rect 4804 12928 4856 12980
rect 5264 12928 5316 12980
rect 5724 12928 5776 12980
rect 6828 12928 6880 12980
rect 11796 12928 11848 12980
rect 11980 12971 12032 12980
rect 11980 12937 11989 12971
rect 11989 12937 12023 12971
rect 12023 12937 12032 12971
rect 11980 12928 12032 12937
rect 12072 12928 12124 12980
rect 3240 12860 3292 12912
rect 4436 12903 4488 12912
rect 4436 12869 4445 12903
rect 4445 12869 4479 12903
rect 4479 12869 4488 12903
rect 4436 12860 4488 12869
rect 6184 12860 6236 12912
rect 7656 12860 7708 12912
rect 8024 12860 8076 12912
rect 9404 12860 9456 12912
rect 9680 12860 9732 12912
rect 10232 12860 10284 12912
rect 10784 12903 10836 12912
rect 10784 12869 10793 12903
rect 10793 12869 10827 12903
rect 10827 12869 10836 12903
rect 10784 12860 10836 12869
rect 11704 12860 11756 12912
rect 13360 12860 13412 12912
rect 16488 12928 16540 12980
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 17776 12928 17828 12980
rect 14464 12860 14516 12912
rect 14832 12903 14884 12912
rect 14832 12869 14841 12903
rect 14841 12869 14875 12903
rect 14875 12869 14884 12903
rect 14832 12860 14884 12869
rect 16764 12860 16816 12912
rect 18880 12928 18932 12980
rect 22192 12928 22244 12980
rect 1124 12724 1176 12776
rect 1676 12724 1728 12776
rect 3700 12792 3752 12844
rect 4160 12835 4212 12844
rect 4160 12801 4169 12835
rect 4169 12801 4203 12835
rect 4203 12801 4212 12835
rect 4160 12792 4212 12801
rect 5724 12792 5776 12844
rect 6276 12792 6328 12844
rect 6552 12835 6604 12844
rect 3332 12656 3384 12708
rect 3516 12588 3568 12640
rect 4068 12656 4120 12708
rect 6092 12724 6144 12776
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7196 12835 7248 12844
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 10140 12792 10192 12844
rect 11336 12792 11388 12844
rect 11520 12792 11572 12844
rect 7656 12767 7708 12776
rect 7656 12733 7665 12767
rect 7665 12733 7699 12767
rect 7699 12733 7708 12767
rect 7656 12724 7708 12733
rect 8944 12724 8996 12776
rect 9864 12724 9916 12776
rect 10600 12724 10652 12776
rect 11060 12767 11112 12776
rect 11060 12733 11069 12767
rect 11069 12733 11103 12767
rect 11103 12733 11112 12767
rect 11060 12724 11112 12733
rect 11704 12724 11756 12776
rect 12716 12792 12768 12844
rect 15200 12792 15252 12844
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 13268 12724 13320 12776
rect 14556 12724 14608 12776
rect 3884 12588 3936 12640
rect 4160 12588 4212 12640
rect 9588 12656 9640 12708
rect 4620 12588 4672 12640
rect 5172 12588 5224 12640
rect 5632 12588 5684 12640
rect 6552 12588 6604 12640
rect 9220 12588 9272 12640
rect 9956 12588 10008 12640
rect 10140 12588 10192 12640
rect 10324 12588 10376 12640
rect 10692 12588 10744 12640
rect 11520 12588 11572 12640
rect 12624 12656 12676 12708
rect 13084 12656 13136 12708
rect 13176 12699 13228 12708
rect 13176 12665 13185 12699
rect 13185 12665 13219 12699
rect 13219 12665 13228 12699
rect 13176 12656 13228 12665
rect 13360 12656 13412 12708
rect 15844 12656 15896 12708
rect 13820 12588 13872 12640
rect 14372 12631 14424 12640
rect 14372 12597 14381 12631
rect 14381 12597 14415 12631
rect 14415 12597 14424 12631
rect 14372 12588 14424 12597
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 16212 12767 16264 12776
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 17316 12792 17368 12844
rect 16488 12724 16540 12776
rect 17592 12656 17644 12708
rect 16488 12588 16540 12640
rect 16948 12588 17000 12640
rect 17868 12767 17920 12776
rect 17868 12733 17877 12767
rect 17877 12733 17911 12767
rect 17911 12733 17920 12767
rect 17868 12724 17920 12733
rect 19616 12860 19668 12912
rect 21548 12860 21600 12912
rect 18604 12792 18656 12844
rect 19524 12792 19576 12844
rect 19708 12835 19760 12844
rect 19708 12801 19717 12835
rect 19717 12801 19751 12835
rect 19751 12801 19760 12835
rect 19708 12792 19760 12801
rect 22008 12792 22060 12844
rect 19156 12724 19208 12776
rect 22376 12724 22428 12776
rect 23296 12860 23348 12912
rect 25228 12860 25280 12912
rect 26056 12928 26108 12980
rect 36728 12928 36780 12980
rect 25964 12860 26016 12912
rect 24308 12792 24360 12844
rect 18880 12656 18932 12708
rect 22284 12699 22336 12708
rect 22284 12665 22293 12699
rect 22293 12665 22327 12699
rect 22327 12665 22336 12699
rect 22284 12656 22336 12665
rect 22468 12656 22520 12708
rect 23296 12724 23348 12776
rect 31576 12792 31628 12844
rect 28908 12767 28960 12776
rect 28908 12733 28917 12767
rect 28917 12733 28951 12767
rect 28951 12733 28960 12767
rect 28908 12724 28960 12733
rect 20076 12588 20128 12640
rect 20168 12588 20220 12640
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 22560 12588 22612 12640
rect 24860 12656 24912 12708
rect 24308 12588 24360 12640
rect 27068 12588 27120 12640
rect 28356 12588 28408 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 2228 12427 2280 12436
rect 2228 12393 2237 12427
rect 2237 12393 2271 12427
rect 2271 12393 2280 12427
rect 2228 12384 2280 12393
rect 4252 12384 4304 12436
rect 2412 12316 2464 12368
rect 6276 12384 6328 12436
rect 8576 12384 8628 12436
rect 9036 12427 9088 12436
rect 9036 12393 9045 12427
rect 9045 12393 9079 12427
rect 9079 12393 9088 12427
rect 9036 12384 9088 12393
rect 9496 12384 9548 12436
rect 5172 12316 5224 12368
rect 5448 12316 5500 12368
rect 6736 12316 6788 12368
rect 7288 12316 7340 12368
rect 7840 12316 7892 12368
rect 1860 12180 1912 12232
rect 2412 12180 2464 12232
rect 2228 12112 2280 12164
rect 4344 12223 4396 12232
rect 4344 12189 4353 12223
rect 4353 12189 4387 12223
rect 4387 12189 4396 12223
rect 4344 12180 4396 12189
rect 4804 12180 4856 12232
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 7840 12180 7892 12232
rect 11612 12384 11664 12436
rect 10876 12316 10928 12368
rect 13544 12384 13596 12436
rect 14740 12384 14792 12436
rect 9956 12291 10008 12300
rect 9956 12257 9965 12291
rect 9965 12257 9999 12291
rect 9999 12257 10008 12291
rect 9956 12248 10008 12257
rect 10416 12248 10468 12300
rect 9404 12180 9456 12232
rect 4528 12112 4580 12164
rect 1584 12087 1636 12096
rect 1584 12053 1593 12087
rect 1593 12053 1627 12087
rect 1627 12053 1636 12087
rect 1584 12044 1636 12053
rect 1860 12044 1912 12096
rect 4620 12044 4672 12096
rect 4988 12044 5040 12096
rect 6184 12112 6236 12164
rect 6368 12044 6420 12096
rect 8024 12044 8076 12096
rect 8484 12044 8536 12096
rect 9036 12044 9088 12096
rect 9404 12044 9456 12096
rect 10048 12112 10100 12164
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 10600 12180 10652 12232
rect 11520 12180 11572 12232
rect 12348 12291 12400 12300
rect 12348 12257 12357 12291
rect 12357 12257 12391 12291
rect 12391 12257 12400 12291
rect 12348 12248 12400 12257
rect 11980 12180 12032 12232
rect 12624 12248 12676 12300
rect 12900 12248 12952 12300
rect 13544 12291 13596 12300
rect 13544 12257 13553 12291
rect 13553 12257 13587 12291
rect 13587 12257 13596 12291
rect 13544 12248 13596 12257
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10692 12044 10744 12096
rect 11888 12112 11940 12164
rect 16948 12384 17000 12436
rect 17040 12384 17092 12436
rect 15200 12316 15252 12368
rect 15660 12316 15712 12368
rect 14924 12248 14976 12300
rect 16856 12248 16908 12300
rect 18052 12316 18104 12368
rect 18880 12427 18932 12436
rect 18880 12393 18889 12427
rect 18889 12393 18923 12427
rect 18923 12393 18932 12427
rect 18880 12384 18932 12393
rect 18604 12248 18656 12300
rect 20352 12384 20404 12436
rect 20720 12384 20772 12436
rect 21640 12384 21692 12436
rect 21732 12384 21784 12436
rect 25228 12384 25280 12436
rect 27620 12384 27672 12436
rect 28448 12427 28500 12436
rect 28448 12393 28457 12427
rect 28457 12393 28491 12427
rect 28491 12393 28500 12427
rect 28448 12384 28500 12393
rect 29276 12384 29328 12436
rect 29736 12384 29788 12436
rect 24124 12316 24176 12368
rect 22560 12248 22612 12300
rect 24308 12248 24360 12300
rect 24584 12248 24636 12300
rect 18512 12180 18564 12232
rect 19984 12180 20036 12232
rect 24400 12180 24452 12232
rect 26792 12180 26844 12232
rect 27712 12316 27764 12368
rect 35992 12316 36044 12368
rect 27344 12248 27396 12300
rect 29644 12248 29696 12300
rect 31668 12180 31720 12232
rect 12624 12044 12676 12096
rect 12808 12044 12860 12096
rect 13636 12044 13688 12096
rect 15200 12112 15252 12164
rect 16403 12155 16455 12164
rect 16403 12121 16405 12155
rect 16405 12121 16439 12155
rect 16439 12121 16455 12155
rect 16403 12112 16455 12121
rect 16856 12112 16908 12164
rect 15016 12044 15068 12096
rect 15844 12044 15896 12096
rect 16580 12044 16632 12096
rect 16672 12044 16724 12096
rect 18236 12044 18288 12096
rect 19524 12044 19576 12096
rect 19616 12044 19668 12096
rect 19800 12044 19852 12096
rect 20260 12044 20312 12096
rect 21732 12112 21784 12164
rect 21640 12044 21692 12096
rect 21824 12087 21876 12096
rect 21824 12053 21833 12087
rect 21833 12053 21867 12087
rect 21867 12053 21876 12087
rect 21824 12044 21876 12053
rect 22560 12155 22612 12164
rect 22560 12121 22569 12155
rect 22569 12121 22603 12155
rect 22603 12121 22612 12155
rect 22560 12112 22612 12121
rect 22836 12044 22888 12096
rect 24032 12087 24084 12096
rect 24032 12053 24041 12087
rect 24041 12053 24075 12087
rect 24075 12053 24084 12087
rect 24032 12044 24084 12053
rect 24676 12112 24728 12164
rect 24584 12044 24636 12096
rect 27620 12044 27672 12096
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 940 11840 992 11892
rect 2596 11883 2648 11892
rect 2596 11849 2605 11883
rect 2605 11849 2639 11883
rect 2639 11849 2648 11883
rect 2596 11840 2648 11849
rect 5448 11840 5500 11892
rect 1308 11772 1360 11824
rect 5264 11772 5316 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2780 11704 2832 11756
rect 3332 11704 3384 11756
rect 3608 11704 3660 11756
rect 5172 11704 5224 11756
rect 5632 11815 5684 11824
rect 5632 11781 5641 11815
rect 5641 11781 5675 11815
rect 5675 11781 5684 11815
rect 5632 11772 5684 11781
rect 5724 11772 5776 11824
rect 6000 11772 6052 11824
rect 6828 11772 6880 11824
rect 9588 11840 9640 11892
rect 11428 11840 11480 11892
rect 11520 11840 11572 11892
rect 11888 11840 11940 11892
rect 11980 11883 12032 11892
rect 11980 11849 11989 11883
rect 11989 11849 12023 11883
rect 12023 11849 12032 11883
rect 11980 11840 12032 11849
rect 7472 11815 7524 11824
rect 7472 11781 7481 11815
rect 7481 11781 7515 11815
rect 7515 11781 7524 11815
rect 7472 11772 7524 11781
rect 8484 11772 8536 11824
rect 9312 11772 9364 11824
rect 10968 11815 11020 11824
rect 10968 11781 10977 11815
rect 10977 11781 11011 11815
rect 11011 11781 11020 11815
rect 10968 11772 11020 11781
rect 12072 11772 12124 11824
rect 3240 11636 3292 11688
rect 4620 11636 4672 11688
rect 4988 11636 5040 11688
rect 5264 11636 5316 11688
rect 5724 11679 5776 11688
rect 5724 11645 5733 11679
rect 5733 11645 5767 11679
rect 5767 11645 5776 11679
rect 5724 11636 5776 11645
rect 9128 11704 9180 11756
rect 9680 11704 9732 11756
rect 11244 11704 11296 11756
rect 11888 11704 11940 11756
rect 12348 11840 12400 11892
rect 12440 11840 12492 11892
rect 14188 11840 14240 11892
rect 14372 11840 14424 11892
rect 12256 11772 12308 11824
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12808 11704 12860 11756
rect 13452 11815 13504 11824
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 15292 11772 15344 11824
rect 15476 11883 15528 11892
rect 15476 11849 15485 11883
rect 15485 11849 15519 11883
rect 15519 11849 15528 11883
rect 15476 11840 15528 11849
rect 16028 11840 16080 11892
rect 16212 11840 16264 11892
rect 16304 11840 16356 11892
rect 16580 11840 16632 11892
rect 17684 11840 17736 11892
rect 17500 11772 17552 11824
rect 18328 11840 18380 11892
rect 18880 11840 18932 11892
rect 6828 11636 6880 11688
rect 388 11568 440 11620
rect 572 11500 624 11552
rect 2596 11500 2648 11552
rect 3700 11543 3752 11552
rect 3700 11509 3709 11543
rect 3709 11509 3743 11543
rect 3743 11509 3752 11543
rect 3700 11500 3752 11509
rect 4252 11500 4304 11552
rect 6736 11568 6788 11620
rect 8576 11568 8628 11620
rect 9128 11568 9180 11620
rect 11704 11636 11756 11688
rect 12256 11636 12308 11688
rect 13912 11636 13964 11688
rect 14924 11704 14976 11756
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 16396 11704 16448 11756
rect 15936 11679 15988 11688
rect 12900 11568 12952 11620
rect 6920 11500 6972 11552
rect 7840 11500 7892 11552
rect 12440 11500 12492 11552
rect 15936 11645 15945 11679
rect 15945 11645 15979 11679
rect 15979 11645 15988 11679
rect 15936 11636 15988 11645
rect 16764 11636 16816 11688
rect 19616 11704 19668 11756
rect 20260 11840 20312 11892
rect 20996 11840 21048 11892
rect 21548 11840 21600 11892
rect 20352 11772 20404 11824
rect 22008 11772 22060 11824
rect 22100 11772 22152 11824
rect 23020 11772 23072 11824
rect 24584 11883 24636 11892
rect 24584 11849 24593 11883
rect 24593 11849 24627 11883
rect 24627 11849 24636 11883
rect 24584 11840 24636 11849
rect 25872 11840 25924 11892
rect 27804 11840 27856 11892
rect 30380 11840 30432 11892
rect 34520 11840 34572 11892
rect 24216 11772 24268 11824
rect 24952 11772 25004 11824
rect 25136 11772 25188 11824
rect 25228 11772 25280 11824
rect 33416 11772 33468 11824
rect 20628 11704 20680 11756
rect 21180 11704 21232 11756
rect 22468 11747 22520 11756
rect 22468 11713 22477 11747
rect 22477 11713 22511 11747
rect 22511 11713 22520 11747
rect 22468 11704 22520 11713
rect 26240 11704 26292 11756
rect 27160 11747 27212 11756
rect 27160 11713 27169 11747
rect 27169 11713 27203 11747
rect 27203 11713 27212 11747
rect 27160 11704 27212 11713
rect 32404 11704 32456 11756
rect 40040 11704 40092 11756
rect 14924 11611 14976 11620
rect 14924 11577 14933 11611
rect 14933 11577 14967 11611
rect 14967 11577 14976 11611
rect 14924 11568 14976 11577
rect 15660 11568 15712 11620
rect 17040 11568 17092 11620
rect 17592 11679 17644 11688
rect 17592 11645 17601 11679
rect 17601 11645 17635 11679
rect 17635 11645 17644 11679
rect 17592 11636 17644 11645
rect 17868 11568 17920 11620
rect 16672 11500 16724 11552
rect 17408 11500 17460 11552
rect 19248 11636 19300 11688
rect 19524 11636 19576 11688
rect 21088 11636 21140 11688
rect 21824 11636 21876 11688
rect 22284 11636 22336 11688
rect 19616 11568 19668 11620
rect 21732 11568 21784 11620
rect 22100 11611 22152 11620
rect 22100 11577 22109 11611
rect 22109 11577 22143 11611
rect 22143 11577 22152 11611
rect 22100 11568 22152 11577
rect 19708 11500 19760 11552
rect 19800 11500 19852 11552
rect 20720 11500 20772 11552
rect 23848 11500 23900 11552
rect 23940 11500 23992 11552
rect 24952 11568 25004 11620
rect 25872 11568 25924 11620
rect 32220 11568 32272 11620
rect 24584 11500 24636 11552
rect 27712 11500 27764 11552
rect 27804 11543 27856 11552
rect 27804 11509 27813 11543
rect 27813 11509 27847 11543
rect 27847 11509 27856 11543
rect 27804 11500 27856 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 3516 11296 3568 11348
rect 5816 11296 5868 11348
rect 7380 11296 7432 11348
rect 7564 11296 7616 11348
rect 12440 11296 12492 11348
rect 13268 11296 13320 11348
rect 13544 11296 13596 11348
rect 13820 11339 13872 11348
rect 13820 11305 13829 11339
rect 13829 11305 13863 11339
rect 13863 11305 13872 11339
rect 13820 11296 13872 11305
rect 14464 11296 14516 11348
rect 2412 11228 2464 11280
rect 1400 11160 1452 11212
rect 2596 11160 2648 11212
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 7104 11228 7156 11280
rect 2136 11092 2188 11144
rect 2412 11092 2464 11144
rect 3516 11092 3568 11144
rect 4068 11135 4120 11144
rect 4068 11101 4077 11135
rect 4077 11101 4111 11135
rect 4111 11101 4120 11135
rect 4068 11092 4120 11101
rect 6184 11092 6236 11144
rect 7196 11160 7248 11212
rect 7748 11160 7800 11212
rect 7380 11092 7432 11144
rect 7840 11092 7892 11144
rect 8576 11160 8628 11212
rect 9312 11228 9364 11280
rect 10784 11228 10836 11280
rect 11152 11228 11204 11280
rect 12808 11228 12860 11280
rect 9956 11203 10008 11212
rect 9956 11169 9965 11203
rect 9965 11169 9999 11203
rect 9999 11169 10008 11203
rect 9956 11160 10008 11169
rect 8484 11092 8536 11144
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 9220 11092 9272 11144
rect 10048 11092 10100 11144
rect 11428 11160 11480 11212
rect 12164 11160 12216 11212
rect 12256 11160 12308 11212
rect 14188 11228 14240 11280
rect 14556 11228 14608 11280
rect 16948 11296 17000 11348
rect 17776 11296 17828 11348
rect 25136 11296 25188 11348
rect 25504 11296 25556 11348
rect 27160 11296 27212 11348
rect 13820 11160 13872 11212
rect 16120 11160 16172 11212
rect 17408 11160 17460 11212
rect 17868 11160 17920 11212
rect 18604 11228 18656 11280
rect 20628 11271 20680 11280
rect 20628 11237 20637 11271
rect 20637 11237 20671 11271
rect 20671 11237 20680 11271
rect 20628 11228 20680 11237
rect 22284 11228 22336 11280
rect 10784 11092 10836 11144
rect 10968 11092 11020 11144
rect 14464 11092 14516 11144
rect 18880 11092 18932 11144
rect 19616 11160 19668 11212
rect 19708 11160 19760 11212
rect 20260 11160 20312 11212
rect 21916 11160 21968 11212
rect 22468 11160 22520 11212
rect 22744 11203 22796 11212
rect 22744 11169 22753 11203
rect 22753 11169 22787 11203
rect 22787 11169 22796 11203
rect 22744 11160 22796 11169
rect 23388 11160 23440 11212
rect 26700 11228 26752 11280
rect 27436 11271 27488 11280
rect 27436 11237 27445 11271
rect 27445 11237 27479 11271
rect 27479 11237 27488 11271
rect 27436 11228 27488 11237
rect 28724 11228 28776 11280
rect 29644 11228 29696 11280
rect 19432 11135 19484 11144
rect 19432 11101 19441 11135
rect 19441 11101 19475 11135
rect 19475 11101 19484 11135
rect 19432 11092 19484 11101
rect 23572 11135 23624 11144
rect 23572 11101 23581 11135
rect 23581 11101 23615 11135
rect 23615 11101 23624 11135
rect 23572 11092 23624 11101
rect 24584 11135 24636 11144
rect 24584 11101 24593 11135
rect 24593 11101 24627 11135
rect 24627 11101 24636 11135
rect 24584 11092 24636 11101
rect 25964 11160 26016 11212
rect 27068 11092 27120 11144
rect 27160 11092 27212 11144
rect 32220 11296 32272 11348
rect 4160 11024 4212 11076
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 9404 11024 9456 11076
rect 2780 10956 2832 11008
rect 6552 10956 6604 11008
rect 7564 10956 7616 11008
rect 7748 10956 7800 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 11796 11067 11848 11076
rect 11796 11033 11805 11067
rect 11805 11033 11839 11067
rect 11839 11033 11848 11067
rect 11796 11024 11848 11033
rect 12808 11024 12860 11076
rect 14372 11024 14424 11076
rect 14924 11067 14976 11076
rect 14924 11033 14933 11067
rect 14933 11033 14967 11067
rect 14967 11033 14976 11067
rect 14924 11024 14976 11033
rect 11980 10956 12032 11008
rect 12440 10956 12492 11008
rect 12716 10956 12768 11008
rect 13820 10956 13872 11008
rect 14832 10956 14884 11008
rect 15384 11024 15436 11076
rect 16764 11067 16816 11076
rect 16764 11033 16773 11067
rect 16773 11033 16807 11067
rect 16807 11033 16816 11067
rect 16764 11024 16816 11033
rect 16856 10956 16908 11008
rect 18696 11024 18748 11076
rect 19524 11024 19576 11076
rect 19616 11024 19668 11076
rect 21180 11024 21232 11076
rect 21364 11024 21416 11076
rect 23112 11024 23164 11076
rect 24216 11024 24268 11076
rect 24860 11024 24912 11076
rect 26700 11024 26752 11076
rect 20720 10956 20772 11008
rect 23572 10956 23624 11008
rect 24124 10956 24176 11008
rect 25412 10956 25464 11008
rect 27804 11024 27856 11076
rect 27712 10956 27764 11008
rect 28632 11024 28684 11076
rect 28724 11067 28776 11076
rect 28724 11033 28733 11067
rect 28733 11033 28767 11067
rect 28767 11033 28776 11067
rect 28724 11024 28776 11033
rect 30012 11067 30064 11076
rect 30012 11033 30021 11067
rect 30021 11033 30055 11067
rect 30055 11033 30064 11067
rect 30012 11024 30064 11033
rect 31300 11024 31352 11076
rect 47768 11024 47820 11076
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 1860 10616 1912 10668
rect 3056 10659 3108 10668
rect 3056 10625 3065 10659
rect 3065 10625 3099 10659
rect 3099 10625 3108 10659
rect 3056 10616 3108 10625
rect 6828 10752 6880 10804
rect 6920 10795 6972 10804
rect 6920 10761 6929 10795
rect 6929 10761 6963 10795
rect 6963 10761 6972 10795
rect 6920 10752 6972 10761
rect 11520 10752 11572 10804
rect 11704 10795 11756 10804
rect 11704 10761 11713 10795
rect 11713 10761 11747 10795
rect 11747 10761 11756 10795
rect 11704 10752 11756 10761
rect 9036 10684 9088 10736
rect 9680 10684 9732 10736
rect 10232 10727 10284 10736
rect 10232 10693 10241 10727
rect 10241 10693 10275 10727
rect 10275 10693 10284 10727
rect 10232 10684 10284 10693
rect 11060 10684 11112 10736
rect 14464 10752 14516 10804
rect 14556 10795 14608 10804
rect 14556 10761 14565 10795
rect 14565 10761 14599 10795
rect 14599 10761 14608 10795
rect 14556 10752 14608 10761
rect 18144 10752 18196 10804
rect 4988 10616 5040 10668
rect 5448 10616 5500 10668
rect 9404 10616 9456 10668
rect 1584 10548 1636 10600
rect 4804 10548 4856 10600
rect 6736 10548 6788 10600
rect 7104 10548 7156 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 7656 10548 7708 10600
rect 2964 10480 3016 10532
rect 5172 10480 5224 10532
rect 6920 10480 6972 10532
rect 2596 10455 2648 10464
rect 2596 10421 2605 10455
rect 2605 10421 2639 10455
rect 2639 10421 2648 10455
rect 2596 10412 2648 10421
rect 2780 10412 2832 10464
rect 5908 10412 5960 10464
rect 6828 10412 6880 10464
rect 8024 10591 8076 10600
rect 8024 10557 8033 10591
rect 8033 10557 8067 10591
rect 8067 10557 8076 10591
rect 8024 10548 8076 10557
rect 9128 10480 9180 10532
rect 8484 10412 8536 10464
rect 9772 10412 9824 10464
rect 10600 10548 10652 10600
rect 10968 10591 11020 10600
rect 10968 10557 10977 10591
rect 10977 10557 11011 10591
rect 11011 10557 11020 10591
rect 10968 10548 11020 10557
rect 11520 10616 11572 10668
rect 12808 10684 12860 10736
rect 14096 10684 14148 10736
rect 15200 10684 15252 10736
rect 16856 10684 16908 10736
rect 17408 10684 17460 10736
rect 19524 10752 19576 10804
rect 21272 10752 21324 10804
rect 22652 10752 22704 10804
rect 22836 10752 22888 10804
rect 29368 10752 29420 10804
rect 30012 10752 30064 10804
rect 15936 10616 15988 10668
rect 17500 10659 17552 10668
rect 17500 10625 17509 10659
rect 17509 10625 17543 10659
rect 17543 10625 17552 10659
rect 17500 10616 17552 10625
rect 20260 10684 20312 10736
rect 21732 10684 21784 10736
rect 22100 10684 22152 10736
rect 24124 10684 24176 10736
rect 25596 10684 25648 10736
rect 22836 10616 22888 10668
rect 23112 10659 23164 10668
rect 23112 10625 23121 10659
rect 23121 10625 23155 10659
rect 23155 10625 23164 10659
rect 23112 10616 23164 10625
rect 23940 10616 23992 10668
rect 24032 10616 24084 10668
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 12072 10548 12124 10600
rect 14372 10548 14424 10600
rect 14740 10548 14792 10600
rect 10876 10412 10928 10464
rect 11060 10412 11112 10464
rect 11888 10480 11940 10532
rect 11704 10412 11756 10464
rect 11980 10455 12032 10464
rect 11980 10421 11989 10455
rect 11989 10421 12023 10455
rect 12023 10421 12032 10455
rect 11980 10412 12032 10421
rect 13544 10480 13596 10532
rect 15936 10480 15988 10532
rect 18420 10548 18472 10600
rect 14556 10412 14608 10464
rect 14740 10412 14792 10464
rect 15108 10412 15160 10464
rect 16764 10412 16816 10464
rect 17040 10412 17092 10464
rect 22468 10548 22520 10600
rect 27436 10659 27488 10668
rect 27436 10625 27445 10659
rect 27445 10625 27479 10659
rect 27479 10625 27488 10659
rect 27436 10616 27488 10625
rect 28816 10659 28868 10668
rect 28816 10625 28825 10659
rect 28825 10625 28859 10659
rect 28859 10625 28868 10659
rect 28816 10616 28868 10625
rect 36084 10616 36136 10668
rect 19616 10480 19668 10532
rect 21180 10480 21232 10532
rect 20076 10412 20128 10464
rect 20720 10412 20772 10464
rect 20996 10412 21048 10464
rect 32588 10548 32640 10600
rect 24216 10480 24268 10532
rect 23848 10412 23900 10464
rect 28540 10480 28592 10532
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 2320 10208 2372 10260
rect 3148 10208 3200 10260
rect 8024 10208 8076 10260
rect 8116 10208 8168 10260
rect 11060 10208 11112 10260
rect 11244 10251 11296 10260
rect 11244 10217 11253 10251
rect 11253 10217 11287 10251
rect 11287 10217 11296 10251
rect 11244 10208 11296 10217
rect 11336 10208 11388 10260
rect 15292 10208 15344 10260
rect 15844 10208 15896 10260
rect 17960 10208 18012 10260
rect 18144 10208 18196 10260
rect 19432 10208 19484 10260
rect 19616 10208 19668 10260
rect 20168 10208 20220 10260
rect 20812 10208 20864 10260
rect 2228 10140 2280 10192
rect 2964 10140 3016 10192
rect 3240 10140 3292 10192
rect 3792 10140 3844 10192
rect 4068 10140 4120 10192
rect 4344 10140 4396 10192
rect 4068 9936 4120 9988
rect 5356 10004 5408 10056
rect 6736 10072 6788 10124
rect 6276 10004 6328 10056
rect 8208 10072 8260 10124
rect 7564 10004 7616 10056
rect 8852 10072 8904 10124
rect 9036 10072 9088 10124
rect 10784 10140 10836 10192
rect 11060 10072 11112 10124
rect 11336 10072 11388 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 13820 10183 13872 10192
rect 13820 10149 13829 10183
rect 13829 10149 13863 10183
rect 13863 10149 13872 10183
rect 13820 10140 13872 10149
rect 15936 10140 15988 10192
rect 18236 10140 18288 10192
rect 23848 10183 23900 10192
rect 23848 10149 23857 10183
rect 23857 10149 23891 10183
rect 23891 10149 23900 10183
rect 23848 10140 23900 10149
rect 14096 10072 14148 10124
rect 17500 10072 17552 10124
rect 17592 10072 17644 10124
rect 19432 10072 19484 10124
rect 24216 10072 24268 10124
rect 24676 10140 24728 10192
rect 8484 10004 8536 10056
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 8116 9936 8168 9988
rect 8392 9936 8444 9988
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2320 9868 2372 9877
rect 5448 9868 5500 9920
rect 7380 9868 7432 9920
rect 7748 9868 7800 9920
rect 8576 9868 8628 9920
rect 8852 9868 8904 9920
rect 9680 9868 9732 9920
rect 11888 9936 11940 9988
rect 12716 9868 12768 9920
rect 13176 9868 13228 9920
rect 13544 9868 13596 9920
rect 14740 9979 14792 9988
rect 14740 9945 14749 9979
rect 14749 9945 14783 9979
rect 14783 9945 14792 9979
rect 14740 9936 14792 9945
rect 15384 9936 15436 9988
rect 16948 9979 17000 9988
rect 16948 9945 16957 9979
rect 16957 9945 16991 9979
rect 16991 9945 17000 9979
rect 16948 9936 17000 9945
rect 18696 9936 18748 9988
rect 22744 10004 22796 10056
rect 23296 10004 23348 10056
rect 24032 10004 24084 10056
rect 25320 10004 25372 10056
rect 19708 9936 19760 9988
rect 21732 9936 21784 9988
rect 22284 9936 22336 9988
rect 30380 10072 30432 10124
rect 14096 9868 14148 9920
rect 14832 9868 14884 9920
rect 15476 9868 15528 9920
rect 17684 9868 17736 9920
rect 17960 9868 18012 9920
rect 19524 9868 19576 9920
rect 19892 9868 19944 9920
rect 20720 9868 20772 9920
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 22744 9911 22796 9920
rect 22744 9877 22753 9911
rect 22753 9877 22787 9911
rect 22787 9877 22796 9911
rect 22744 9868 22796 9877
rect 26700 9936 26752 9988
rect 33324 9936 33376 9988
rect 26056 9911 26108 9920
rect 26056 9877 26065 9911
rect 26065 9877 26099 9911
rect 26099 9877 26108 9911
rect 26056 9868 26108 9877
rect 26608 9911 26660 9920
rect 26608 9877 26617 9911
rect 26617 9877 26651 9911
rect 26651 9877 26660 9911
rect 26608 9868 26660 9877
rect 28448 9868 28500 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 1492 9664 1544 9716
rect 2688 9664 2740 9716
rect 3700 9664 3752 9716
rect 1952 9596 2004 9648
rect 2872 9596 2924 9648
rect 664 9528 716 9580
rect 848 9528 900 9580
rect 2228 9528 2280 9580
rect 3700 9528 3752 9580
rect 4252 9571 4304 9580
rect 4252 9537 4261 9571
rect 4261 9537 4295 9571
rect 4295 9537 4304 9571
rect 4252 9528 4304 9537
rect 5632 9596 5684 9648
rect 6460 9596 6512 9648
rect 6920 9664 6972 9716
rect 9404 9664 9456 9716
rect 9496 9664 9548 9716
rect 12072 9664 12124 9716
rect 12164 9664 12216 9716
rect 7380 9528 7432 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 8668 9596 8720 9648
rect 8852 9596 8904 9648
rect 10232 9596 10284 9648
rect 11336 9596 11388 9648
rect 11888 9596 11940 9648
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 11520 9528 11572 9580
rect 480 9460 532 9512
rect 5632 9460 5684 9512
rect 6828 9460 6880 9512
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 1400 9392 1452 9444
rect 3240 9392 3292 9444
rect 4068 9392 4120 9444
rect 5080 9392 5132 9444
rect 7104 9392 7156 9444
rect 9220 9460 9272 9512
rect 11152 9460 11204 9512
rect 12072 9460 12124 9512
rect 12532 9460 12584 9512
rect 13176 9460 13228 9512
rect 13360 9664 13412 9716
rect 13544 9664 13596 9716
rect 14464 9664 14516 9716
rect 16856 9664 16908 9716
rect 17316 9664 17368 9716
rect 14740 9639 14792 9648
rect 14740 9605 14749 9639
rect 14749 9605 14783 9639
rect 14783 9605 14792 9639
rect 14740 9596 14792 9605
rect 15384 9596 15436 9648
rect 17040 9596 17092 9648
rect 18696 9664 18748 9716
rect 22560 9664 22612 9716
rect 18604 9596 18656 9648
rect 19064 9596 19116 9648
rect 23572 9596 23624 9648
rect 28816 9664 28868 9716
rect 18420 9528 18472 9580
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 21456 9528 21508 9580
rect 27620 9596 27672 9648
rect 27712 9596 27764 9648
rect 32036 9596 32088 9648
rect 25228 9528 25280 9580
rect 25320 9528 25372 9580
rect 26332 9528 26384 9580
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 11520 9392 11572 9444
rect 940 9324 992 9376
rect 1860 9324 1912 9376
rect 2412 9324 2464 9376
rect 2688 9367 2740 9376
rect 2688 9333 2697 9367
rect 2697 9333 2731 9367
rect 2731 9333 2740 9367
rect 2688 9324 2740 9333
rect 4804 9324 4856 9376
rect 5264 9324 5316 9376
rect 5724 9324 5776 9376
rect 9772 9324 9824 9376
rect 10048 9324 10100 9376
rect 10140 9324 10192 9376
rect 13084 9392 13136 9444
rect 15844 9392 15896 9444
rect 16028 9392 16080 9444
rect 19340 9392 19392 9444
rect 21272 9460 21324 9512
rect 21640 9460 21692 9512
rect 23756 9392 23808 9444
rect 26148 9460 26200 9512
rect 31852 9460 31904 9512
rect 26240 9392 26292 9444
rect 12072 9324 12124 9376
rect 13820 9324 13872 9376
rect 14188 9367 14240 9376
rect 14188 9333 14197 9367
rect 14197 9333 14231 9367
rect 14231 9333 14240 9367
rect 14188 9324 14240 9333
rect 14556 9324 14608 9376
rect 17224 9324 17276 9376
rect 18144 9324 18196 9376
rect 20536 9324 20588 9376
rect 26792 9324 26844 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 1216 9120 1268 9172
rect 2228 9120 2280 9172
rect 3792 9163 3844 9172
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 6368 9120 6420 9172
rect 7564 9120 7616 9172
rect 10048 9120 10100 9172
rect 11060 9120 11112 9172
rect 15844 9120 15896 9172
rect 9772 9052 9824 9104
rect 10508 9052 10560 9104
rect 296 8984 348 9036
rect 1216 8984 1268 9036
rect 3792 8984 3844 9036
rect 7196 8984 7248 9036
rect 2412 8916 2464 8968
rect 2780 8959 2832 8968
rect 2780 8925 2789 8959
rect 2789 8925 2823 8959
rect 2823 8925 2832 8959
rect 2780 8916 2832 8925
rect 4712 8916 4764 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 5908 8916 5960 8968
rect 4344 8848 4396 8900
rect 7196 8848 7248 8900
rect 9404 8916 9456 8968
rect 10140 8916 10192 8968
rect 11336 8984 11388 9036
rect 11152 8916 11204 8968
rect 14096 9052 14148 9104
rect 14556 9052 14608 9104
rect 17868 9120 17920 9172
rect 18512 9120 18564 9172
rect 18788 9120 18840 9172
rect 20260 9120 20312 9172
rect 21364 9120 21416 9172
rect 26332 9163 26384 9172
rect 26332 9129 26341 9163
rect 26341 9129 26375 9163
rect 26375 9129 26384 9163
rect 26332 9120 26384 9129
rect 31300 9120 31352 9172
rect 12900 8984 12952 9036
rect 13360 8916 13412 8968
rect 14924 9027 14976 9036
rect 14924 8993 14933 9027
rect 14933 8993 14967 9027
rect 14967 8993 14976 9027
rect 14924 8984 14976 8993
rect 20904 9052 20956 9104
rect 16488 8984 16540 9036
rect 21824 9052 21876 9104
rect 22376 9052 22428 9104
rect 25044 9052 25096 9104
rect 27712 9052 27764 9104
rect 32772 9052 32824 9104
rect 40592 9052 40644 9104
rect 16028 8916 16080 8968
rect 17132 8959 17184 8968
rect 17132 8925 17141 8959
rect 17141 8925 17175 8959
rect 17175 8925 17184 8959
rect 17132 8916 17184 8925
rect 18788 8916 18840 8968
rect 20904 8959 20956 8968
rect 20904 8925 20913 8959
rect 20913 8925 20947 8959
rect 20947 8925 20956 8959
rect 20904 8916 20956 8925
rect 22008 8959 22060 8968
rect 22008 8925 22028 8959
rect 22028 8925 22060 8959
rect 29000 8984 29052 9036
rect 38476 8984 38528 9036
rect 22008 8916 22060 8925
rect 4712 8780 4764 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 5264 8823 5316 8832
rect 5264 8789 5273 8823
rect 5273 8789 5307 8823
rect 5307 8789 5316 8823
rect 5264 8780 5316 8789
rect 5356 8780 5408 8832
rect 6460 8780 6512 8832
rect 8392 8780 8444 8832
rect 8760 8780 8812 8832
rect 10232 8891 10284 8900
rect 10232 8857 10241 8891
rect 10241 8857 10275 8891
rect 10275 8857 10284 8891
rect 10232 8848 10284 8857
rect 10416 8848 10468 8900
rect 11060 8848 11112 8900
rect 11336 8780 11388 8832
rect 11888 8780 11940 8832
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 15108 8848 15160 8900
rect 12900 8780 12952 8832
rect 13360 8780 13412 8832
rect 13912 8780 13964 8832
rect 14924 8780 14976 8832
rect 15936 8823 15988 8832
rect 15936 8789 15945 8823
rect 15945 8789 15979 8823
rect 15979 8789 15988 8823
rect 15936 8780 15988 8789
rect 16028 8823 16080 8832
rect 16028 8789 16037 8823
rect 16037 8789 16071 8823
rect 16071 8789 16080 8823
rect 16028 8780 16080 8789
rect 17500 8780 17552 8832
rect 17868 8848 17920 8900
rect 19064 8848 19116 8900
rect 25688 8959 25740 8968
rect 25688 8925 25697 8959
rect 25697 8925 25731 8959
rect 25731 8925 25740 8959
rect 25688 8916 25740 8925
rect 20444 8780 20496 8832
rect 26240 8848 26292 8900
rect 27620 8916 27672 8968
rect 41328 8916 41380 8968
rect 25228 8823 25280 8832
rect 25228 8789 25237 8823
rect 25237 8789 25271 8823
rect 25271 8789 25280 8823
rect 25228 8780 25280 8789
rect 27712 8780 27764 8832
rect 28356 8780 28408 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 1584 8619 1636 8628
rect 1584 8585 1593 8619
rect 1593 8585 1627 8619
rect 1627 8585 1636 8619
rect 1584 8576 1636 8585
rect 1676 8619 1728 8628
rect 1676 8585 1685 8619
rect 1685 8585 1719 8619
rect 1719 8585 1728 8619
rect 1676 8576 1728 8585
rect 3976 8576 4028 8628
rect 5540 8576 5592 8628
rect 7012 8576 7064 8628
rect 2596 8508 2648 8560
rect 1584 8440 1636 8492
rect 7564 8508 7616 8560
rect 1952 8372 2004 8424
rect 2596 8372 2648 8424
rect 4896 8440 4948 8492
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 12164 8576 12216 8628
rect 18420 8576 18472 8628
rect 18788 8576 18840 8628
rect 20628 8619 20680 8628
rect 20628 8585 20637 8619
rect 20637 8585 20671 8619
rect 20671 8585 20680 8619
rect 20628 8576 20680 8585
rect 22468 8576 22520 8628
rect 23756 8619 23808 8628
rect 23756 8585 23765 8619
rect 23765 8585 23799 8619
rect 23799 8585 23808 8619
rect 23756 8576 23808 8585
rect 24124 8576 24176 8628
rect 10048 8508 10100 8560
rect 6368 8372 6420 8424
rect 7472 8372 7524 8424
rect 8576 8372 8628 8424
rect 8760 8483 8812 8492
rect 8760 8449 8769 8483
rect 8769 8449 8803 8483
rect 8803 8449 8812 8483
rect 8760 8440 8812 8449
rect 9220 8440 9272 8492
rect 10232 8440 10284 8492
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 12532 8508 12584 8560
rect 11060 8440 11112 8492
rect 9496 8372 9548 8424
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 2320 8304 2372 8356
rect 4068 8304 4120 8356
rect 1032 8236 1084 8288
rect 1952 8236 2004 8288
rect 7012 8304 7064 8356
rect 7748 8304 7800 8356
rect 10232 8304 10284 8356
rect 10692 8304 10744 8356
rect 10968 8415 11020 8424
rect 10968 8381 10977 8415
rect 10977 8381 11011 8415
rect 11011 8381 11020 8415
rect 10968 8372 11020 8381
rect 11060 8304 11112 8356
rect 5724 8236 5776 8288
rect 6828 8236 6880 8288
rect 9404 8279 9456 8288
rect 9404 8245 9413 8279
rect 9413 8245 9447 8279
rect 9447 8245 9456 8279
rect 9404 8236 9456 8245
rect 9680 8236 9732 8288
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 12072 8440 12124 8492
rect 12256 8372 12308 8424
rect 14556 8440 14608 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 11980 8347 12032 8356
rect 11980 8313 11989 8347
rect 11989 8313 12023 8347
rect 12023 8313 12032 8347
rect 11980 8304 12032 8313
rect 11336 8236 11388 8288
rect 12164 8236 12216 8288
rect 13544 8304 13596 8356
rect 15384 8372 15436 8424
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 18052 8415 18104 8424
rect 18052 8381 18061 8415
rect 18061 8381 18095 8415
rect 18095 8381 18104 8415
rect 18052 8372 18104 8381
rect 18972 8440 19024 8492
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 19340 8372 19392 8424
rect 19524 8372 19576 8424
rect 21732 8508 21784 8560
rect 25964 8576 26016 8628
rect 28356 8576 28408 8628
rect 36360 8576 36412 8628
rect 22744 8440 22796 8492
rect 23388 8440 23440 8492
rect 26516 8508 26568 8560
rect 29736 8440 29788 8492
rect 12716 8236 12768 8288
rect 12808 8236 12860 8288
rect 14280 8236 14332 8288
rect 16396 8236 16448 8288
rect 20996 8304 21048 8356
rect 27804 8372 27856 8424
rect 31024 8372 31076 8424
rect 32312 8304 32364 8356
rect 23940 8236 23992 8288
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 2412 8032 2464 8084
rect 4804 8032 4856 8084
rect 5080 8032 5132 8084
rect 5816 8032 5868 8084
rect 6092 8032 6144 8084
rect 7196 8032 7248 8084
rect 8300 8032 8352 8084
rect 8760 8032 8812 8084
rect 9680 8032 9732 8084
rect 9864 8075 9916 8084
rect 9864 8041 9873 8075
rect 9873 8041 9907 8075
rect 9907 8041 9916 8075
rect 9864 8032 9916 8041
rect 10048 8032 10100 8084
rect 11520 8032 11572 8084
rect 11704 8032 11756 8084
rect 13176 8032 13228 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 16764 8032 16816 8084
rect 17132 8032 17184 8084
rect 20904 8032 20956 8084
rect 23388 8032 23440 8084
rect 24400 8032 24452 8084
rect 1308 7964 1360 8016
rect 4344 7964 4396 8016
rect 2228 7828 2280 7880
rect 3516 7828 3568 7880
rect 3976 7828 4028 7880
rect 10968 7964 11020 8016
rect 11152 7964 11204 8016
rect 15200 7964 15252 8016
rect 4896 7760 4948 7812
rect 5264 7760 5316 7812
rect 6828 7828 6880 7880
rect 9588 7896 9640 7948
rect 10048 7828 10100 7880
rect 10324 7828 10376 7880
rect 10876 7896 10928 7948
rect 11060 7896 11112 7948
rect 13912 7896 13964 7948
rect 15936 7896 15988 7948
rect 16120 7896 16172 7948
rect 17868 7896 17920 7948
rect 25320 7964 25372 8016
rect 25504 8032 25556 8084
rect 39396 8032 39448 8084
rect 49056 7964 49108 8016
rect 11244 7828 11296 7880
rect 12164 7828 12216 7880
rect 13176 7828 13228 7880
rect 14924 7828 14976 7880
rect 15752 7828 15804 7880
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 18880 7828 18932 7880
rect 18972 7828 19024 7880
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 22192 7896 22244 7948
rect 24860 7939 24912 7948
rect 24860 7905 24869 7939
rect 24869 7905 24903 7939
rect 24903 7905 24912 7939
rect 24860 7896 24912 7905
rect 25596 7896 25648 7948
rect 21272 7828 21324 7880
rect 23112 7871 23164 7880
rect 23112 7837 23121 7871
rect 23121 7837 23155 7871
rect 23155 7837 23164 7871
rect 23112 7828 23164 7837
rect 24768 7828 24820 7880
rect 2780 7692 2832 7744
rect 12072 7760 12124 7812
rect 15200 7760 15252 7812
rect 16488 7760 16540 7812
rect 7564 7692 7616 7744
rect 10232 7692 10284 7744
rect 10600 7692 10652 7744
rect 10968 7692 11020 7744
rect 12348 7692 12400 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 15660 7692 15712 7744
rect 18512 7692 18564 7744
rect 24124 7692 24176 7744
rect 24860 7760 24912 7812
rect 25596 7760 25648 7812
rect 27804 7692 27856 7744
rect 38752 7692 38804 7744
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 4160 7488 4212 7540
rect 4436 7488 4488 7540
rect 4988 7531 5040 7540
rect 4988 7497 4997 7531
rect 4997 7497 5031 7531
rect 5031 7497 5040 7531
rect 4988 7488 5040 7497
rect 6552 7488 6604 7540
rect 10968 7488 11020 7540
rect 11060 7488 11112 7540
rect 12256 7488 12308 7540
rect 12440 7488 12492 7540
rect 1216 7420 1268 7472
rect 1584 7420 1636 7472
rect 2136 7420 2188 7472
rect 8392 7420 8444 7472
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 4068 7395 4120 7404
rect 4068 7361 4077 7395
rect 4077 7361 4111 7395
rect 4111 7361 4120 7395
rect 4068 7352 4120 7361
rect 4712 7352 4764 7404
rect 5264 7284 5316 7336
rect 7104 7284 7156 7336
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 7932 7352 7984 7404
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 3516 7216 3568 7268
rect 4712 7216 4764 7268
rect 5448 7216 5500 7268
rect 7932 7216 7984 7268
rect 4620 7148 4672 7200
rect 5540 7148 5592 7200
rect 6736 7148 6788 7200
rect 8300 7148 8352 7200
rect 10324 7284 10376 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 11152 7463 11204 7472
rect 11152 7429 11161 7463
rect 11161 7429 11195 7463
rect 11195 7429 11204 7463
rect 11152 7420 11204 7429
rect 12624 7420 12676 7472
rect 11244 7352 11296 7404
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 15292 7488 15344 7540
rect 16764 7488 16816 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 19984 7488 20036 7540
rect 21456 7531 21508 7540
rect 21456 7497 21465 7531
rect 21465 7497 21499 7531
rect 21499 7497 21508 7531
rect 21456 7488 21508 7497
rect 21548 7488 21600 7540
rect 23112 7488 23164 7540
rect 23756 7531 23808 7540
rect 23756 7497 23765 7531
rect 23765 7497 23799 7531
rect 23799 7497 23808 7531
rect 23756 7488 23808 7497
rect 25688 7488 25740 7540
rect 15108 7420 15160 7472
rect 19248 7420 19300 7472
rect 22284 7463 22336 7472
rect 22284 7429 22293 7463
rect 22293 7429 22327 7463
rect 22327 7429 22336 7463
rect 22284 7420 22336 7429
rect 22836 7420 22888 7472
rect 15200 7352 15252 7404
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 15384 7284 15436 7336
rect 9404 7216 9456 7268
rect 10968 7216 11020 7268
rect 11336 7259 11388 7268
rect 11336 7225 11345 7259
rect 11345 7225 11379 7259
rect 11379 7225 11388 7259
rect 11336 7216 11388 7225
rect 11520 7216 11572 7268
rect 16672 7352 16724 7404
rect 17132 7352 17184 7404
rect 18512 7352 18564 7404
rect 19800 7352 19852 7404
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 21916 7352 21968 7404
rect 29000 7420 29052 7472
rect 16120 7284 16172 7336
rect 24860 7284 24912 7336
rect 8944 7148 8996 7200
rect 12072 7148 12124 7200
rect 16672 7216 16724 7268
rect 17224 7216 17276 7268
rect 18972 7216 19024 7268
rect 24400 7259 24452 7268
rect 24400 7225 24409 7259
rect 24409 7225 24443 7259
rect 24443 7225 24452 7259
rect 24400 7216 24452 7225
rect 15660 7148 15712 7200
rect 17132 7148 17184 7200
rect 25780 7148 25832 7200
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 2596 6944 2648 6996
rect 5356 6944 5408 6996
rect 6368 6987 6420 6996
rect 6368 6953 6377 6987
rect 6377 6953 6411 6987
rect 6411 6953 6420 6987
rect 6368 6944 6420 6953
rect 7288 6944 7340 6996
rect 9220 6944 9272 6996
rect 13728 6944 13780 6996
rect 1124 6876 1176 6928
rect 2688 6876 2740 6928
rect 3700 6876 3752 6928
rect 1768 6808 1820 6860
rect 7196 6876 7248 6928
rect 10600 6876 10652 6928
rect 10692 6876 10744 6928
rect 15844 6944 15896 6996
rect 15936 6944 15988 6996
rect 14740 6876 14792 6928
rect 16304 6876 16356 6928
rect 7380 6808 7432 6860
rect 7748 6808 7800 6860
rect 2136 6740 2188 6792
rect 2596 6740 2648 6792
rect 3516 6740 3568 6792
rect 4252 6740 4304 6792
rect 4344 6740 4396 6792
rect 5264 6783 5316 6792
rect 5264 6749 5273 6783
rect 5273 6749 5307 6783
rect 5307 6749 5316 6783
rect 5264 6740 5316 6749
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6000 6740 6052 6792
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 10232 6808 10284 6860
rect 10784 6851 10836 6860
rect 10784 6817 10793 6851
rect 10793 6817 10827 6851
rect 10827 6817 10836 6851
rect 10784 6808 10836 6817
rect 10968 6808 11020 6860
rect 9036 6783 9088 6792
rect 9036 6749 9045 6783
rect 9045 6749 9079 6783
rect 9079 6749 9088 6783
rect 9036 6740 9088 6749
rect 11704 6740 11756 6792
rect 12532 6808 12584 6860
rect 12072 6740 12124 6792
rect 13452 6808 13504 6860
rect 14556 6851 14608 6860
rect 14556 6817 14565 6851
rect 14565 6817 14599 6851
rect 14599 6817 14608 6851
rect 14556 6808 14608 6817
rect 15936 6808 15988 6860
rect 16488 6808 16540 6860
rect 16580 6808 16632 6860
rect 17500 6808 17552 6860
rect 3240 6715 3292 6724
rect 3240 6681 3249 6715
rect 3249 6681 3283 6715
rect 3283 6681 3292 6715
rect 3240 6672 3292 6681
rect 7840 6672 7892 6724
rect 9680 6715 9732 6724
rect 9680 6681 9689 6715
rect 9689 6681 9723 6715
rect 9723 6681 9732 6715
rect 9680 6672 9732 6681
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 1952 6604 2004 6656
rect 3700 6604 3752 6656
rect 6460 6604 6512 6656
rect 9036 6604 9088 6656
rect 10232 6604 10284 6656
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 10692 6604 10744 6656
rect 10876 6604 10928 6656
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 15476 6783 15528 6792
rect 15476 6749 15485 6783
rect 15485 6749 15519 6783
rect 15519 6749 15528 6783
rect 15476 6740 15528 6749
rect 16764 6783 16816 6792
rect 16764 6749 16773 6783
rect 16773 6749 16807 6783
rect 16807 6749 16816 6783
rect 16764 6740 16816 6749
rect 13912 6672 13964 6724
rect 16028 6672 16080 6724
rect 16396 6672 16448 6724
rect 18512 6851 18564 6860
rect 18512 6817 18521 6851
rect 18521 6817 18555 6851
rect 18555 6817 18564 6851
rect 18512 6808 18564 6817
rect 20536 6944 20588 6996
rect 22284 6944 22336 6996
rect 22836 6944 22888 6996
rect 25320 6944 25372 6996
rect 26884 6944 26936 6996
rect 26884 6808 26936 6860
rect 19340 6740 19392 6792
rect 20812 6740 20864 6792
rect 21732 6672 21784 6724
rect 23020 6715 23072 6724
rect 23020 6681 23029 6715
rect 23029 6681 23063 6715
rect 23063 6681 23072 6715
rect 23020 6672 23072 6681
rect 23204 6715 23256 6724
rect 23204 6681 23213 6715
rect 23213 6681 23247 6715
rect 23247 6681 23256 6715
rect 23204 6672 23256 6681
rect 15200 6604 15252 6656
rect 17592 6604 17644 6656
rect 21180 6604 21232 6656
rect 24124 6604 24176 6656
rect 30472 6604 30524 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 3332 6400 3384 6452
rect 3976 6400 4028 6452
rect 4068 6400 4120 6452
rect 3792 6332 3844 6384
rect 4896 6443 4948 6452
rect 4896 6409 4905 6443
rect 4905 6409 4939 6443
rect 4939 6409 4948 6443
rect 4896 6400 4948 6409
rect 5632 6400 5684 6452
rect 1308 6264 1360 6316
rect 1952 6264 2004 6316
rect 2688 6196 2740 6248
rect 4068 6264 4120 6316
rect 5356 6307 5408 6316
rect 5356 6273 5365 6307
rect 5365 6273 5399 6307
rect 5399 6273 5408 6307
rect 5356 6264 5408 6273
rect 7748 6332 7800 6384
rect 9036 6332 9088 6384
rect 16764 6400 16816 6452
rect 17776 6400 17828 6452
rect 10692 6332 10744 6384
rect 3516 6128 3568 6180
rect 3976 6196 4028 6248
rect 6460 6196 6512 6248
rect 8300 6307 8352 6316
rect 8300 6273 8309 6307
rect 8309 6273 8343 6307
rect 8343 6273 8352 6307
rect 8300 6264 8352 6273
rect 8944 6196 8996 6248
rect 10968 6264 11020 6316
rect 12164 6264 12216 6316
rect 11060 6196 11112 6248
rect 16212 6332 16264 6384
rect 16304 6375 16356 6384
rect 16304 6341 16313 6375
rect 16313 6341 16347 6375
rect 16347 6341 16356 6375
rect 16304 6332 16356 6341
rect 16948 6332 17000 6384
rect 20812 6443 20864 6452
rect 20812 6409 20821 6443
rect 20821 6409 20855 6443
rect 20855 6409 20864 6443
rect 20812 6400 20864 6409
rect 23020 6400 23072 6452
rect 23296 6400 23348 6452
rect 26240 6400 26292 6452
rect 26884 6400 26936 6452
rect 33876 6400 33928 6452
rect 13728 6264 13780 6316
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 26056 6332 26108 6384
rect 16764 6196 16816 6248
rect 20996 6264 21048 6316
rect 21456 6307 21508 6316
rect 21456 6273 21465 6307
rect 21465 6273 21499 6307
rect 21499 6273 21508 6307
rect 21456 6264 21508 6273
rect 22192 6307 22244 6316
rect 22192 6273 22201 6307
rect 22201 6273 22235 6307
rect 22235 6273 22244 6307
rect 22192 6264 22244 6273
rect 22836 6307 22888 6316
rect 22836 6273 22845 6307
rect 22845 6273 22879 6307
rect 22879 6273 22888 6307
rect 22836 6264 22888 6273
rect 23296 6264 23348 6316
rect 25228 6196 25280 6248
rect 27620 6196 27672 6248
rect 43628 6196 43680 6248
rect 3332 6060 3384 6112
rect 4160 6128 4212 6180
rect 6368 6060 6420 6112
rect 6460 6103 6512 6112
rect 6460 6069 6469 6103
rect 6469 6069 6503 6103
rect 6503 6069 6512 6103
rect 6460 6060 6512 6069
rect 6736 6128 6788 6180
rect 14188 6128 14240 6180
rect 9864 6060 9916 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11704 6103 11756 6112
rect 11704 6069 11713 6103
rect 11713 6069 11747 6103
rect 11747 6069 11756 6103
rect 11704 6060 11756 6069
rect 12716 6060 12768 6112
rect 14556 6060 14608 6112
rect 14832 6060 14884 6112
rect 17132 6060 17184 6112
rect 18328 6128 18380 6180
rect 21548 6128 21600 6180
rect 23756 6128 23808 6180
rect 26148 6128 26200 6180
rect 42064 6128 42116 6180
rect 23296 6103 23348 6112
rect 23296 6069 23305 6103
rect 23305 6069 23339 6103
rect 23339 6069 23348 6103
rect 23296 6060 23348 6069
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 4436 5856 4488 5908
rect 5448 5899 5500 5908
rect 5448 5865 5457 5899
rect 5457 5865 5491 5899
rect 5491 5865 5500 5899
rect 5448 5856 5500 5865
rect 7380 5856 7432 5908
rect 10232 5856 10284 5908
rect 11612 5856 11664 5908
rect 12808 5856 12860 5908
rect 13728 5899 13780 5908
rect 13728 5865 13737 5899
rect 13737 5865 13771 5899
rect 13771 5865 13780 5899
rect 13728 5856 13780 5865
rect 756 5788 808 5840
rect 3332 5788 3384 5840
rect 3424 5831 3476 5840
rect 3424 5797 3433 5831
rect 3433 5797 3467 5831
rect 3467 5797 3476 5831
rect 3424 5788 3476 5797
rect 3700 5788 3752 5840
rect 2044 5720 2096 5772
rect 1308 5652 1360 5704
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 1860 5516 1912 5568
rect 3792 5652 3844 5704
rect 9312 5720 9364 5772
rect 9956 5720 10008 5772
rect 5540 5652 5592 5704
rect 7472 5652 7524 5704
rect 7932 5695 7984 5704
rect 7932 5661 7941 5695
rect 7941 5661 7975 5695
rect 7975 5661 7984 5695
rect 7932 5652 7984 5661
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 15292 5763 15344 5772
rect 15292 5729 15301 5763
rect 15301 5729 15335 5763
rect 15335 5729 15344 5763
rect 15292 5720 15344 5729
rect 16856 5720 16908 5772
rect 18604 5720 18656 5772
rect 23848 5856 23900 5908
rect 20996 5788 21048 5840
rect 21180 5831 21232 5840
rect 21180 5797 21189 5831
rect 21189 5797 21223 5831
rect 21223 5797 21232 5831
rect 21180 5788 21232 5797
rect 19708 5763 19760 5772
rect 19708 5729 19717 5763
rect 19717 5729 19751 5763
rect 19751 5729 19760 5763
rect 19708 5720 19760 5729
rect 30656 5788 30708 5840
rect 12440 5652 12492 5704
rect 4620 5584 4672 5636
rect 6552 5584 6604 5636
rect 4896 5516 4948 5568
rect 5172 5559 5224 5568
rect 5172 5525 5181 5559
rect 5181 5525 5215 5559
rect 5215 5525 5224 5559
rect 5172 5516 5224 5525
rect 8300 5516 8352 5568
rect 11796 5584 11848 5636
rect 12808 5584 12860 5636
rect 13912 5652 13964 5704
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 19156 5652 19208 5704
rect 20352 5652 20404 5704
rect 21180 5652 21232 5704
rect 12532 5516 12584 5568
rect 13544 5516 13596 5568
rect 15108 5516 15160 5568
rect 17316 5584 17368 5636
rect 27712 5720 27764 5772
rect 24952 5584 25004 5636
rect 23756 5516 23808 5568
rect 27068 5516 27120 5568
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 2412 5312 2464 5364
rect 3424 5312 3476 5364
rect 3884 5355 3936 5364
rect 3884 5321 3893 5355
rect 3893 5321 3927 5355
rect 3927 5321 3936 5355
rect 3884 5312 3936 5321
rect 5080 5312 5132 5364
rect 7196 5312 7248 5364
rect 7748 5312 7800 5364
rect 8944 5355 8996 5364
rect 8944 5321 8953 5355
rect 8953 5321 8987 5355
rect 8987 5321 8996 5355
rect 8944 5312 8996 5321
rect 11336 5312 11388 5364
rect 12072 5312 12124 5364
rect 12808 5355 12860 5364
rect 12808 5321 12817 5355
rect 12817 5321 12851 5355
rect 12851 5321 12860 5355
rect 12808 5312 12860 5321
rect 13452 5312 13504 5364
rect 2228 5244 2280 5296
rect 8392 5244 8444 5296
rect 9128 5244 9180 5296
rect 4528 5176 4580 5228
rect 5724 5176 5776 5228
rect 8208 5176 8260 5228
rect 8300 5219 8352 5228
rect 8300 5185 8309 5219
rect 8309 5185 8343 5219
rect 8343 5185 8352 5219
rect 8300 5176 8352 5185
rect 10140 5176 10192 5228
rect 10968 5244 11020 5296
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 17408 5312 17460 5364
rect 18328 5312 18380 5364
rect 21180 5312 21232 5364
rect 12440 5176 12492 5228
rect 12716 5176 12768 5228
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 14556 5219 14608 5228
rect 14556 5185 14565 5219
rect 14565 5185 14599 5219
rect 14599 5185 14608 5219
rect 14556 5176 14608 5185
rect 15844 5176 15896 5228
rect 19432 5244 19484 5296
rect 19616 5244 19668 5296
rect 29736 5312 29788 5364
rect 23664 5244 23716 5296
rect 24952 5287 25004 5296
rect 24952 5253 24961 5287
rect 24961 5253 24995 5287
rect 24995 5253 25004 5287
rect 24952 5244 25004 5253
rect 27528 5244 27580 5296
rect 16948 5176 17000 5228
rect 2964 5108 3016 5160
rect 664 5040 716 5092
rect 9220 5108 9272 5160
rect 10416 5108 10468 5160
rect 11704 5151 11756 5160
rect 11704 5117 11713 5151
rect 11713 5117 11747 5151
rect 11747 5117 11756 5151
rect 11704 5108 11756 5117
rect 13912 5108 13964 5160
rect 18696 5219 18748 5228
rect 18696 5185 18705 5219
rect 18705 5185 18739 5219
rect 18739 5185 18748 5219
rect 18696 5176 18748 5185
rect 19800 5176 19852 5228
rect 19984 5219 20036 5228
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 21272 5176 21324 5228
rect 22192 5218 22244 5228
rect 22192 5184 22236 5218
rect 22236 5184 22244 5218
rect 22192 5176 22244 5184
rect 23296 5176 23348 5228
rect 31760 5244 31812 5296
rect 18880 5108 18932 5160
rect 6368 5040 6420 5092
rect 1676 4972 1728 5024
rect 5448 4972 5500 5024
rect 6184 4972 6236 5024
rect 15660 5040 15712 5092
rect 24308 5108 24360 5160
rect 9312 4972 9364 5024
rect 12072 4972 12124 5024
rect 13820 4972 13872 5024
rect 14096 4972 14148 5024
rect 16304 5015 16356 5024
rect 16304 4981 16313 5015
rect 16313 4981 16347 5015
rect 16347 4981 16356 5015
rect 16304 4972 16356 4981
rect 18420 4972 18472 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 22560 4972 22612 5024
rect 25504 5040 25556 5092
rect 27068 4972 27120 5024
rect 27344 5151 27396 5160
rect 27344 5117 27353 5151
rect 27353 5117 27387 5151
rect 27387 5117 27396 5151
rect 27344 5108 27396 5117
rect 28908 5151 28960 5160
rect 28908 5117 28917 5151
rect 28917 5117 28951 5151
rect 28951 5117 28960 5151
rect 28908 5108 28960 5117
rect 29644 5151 29696 5160
rect 29644 5117 29653 5151
rect 29653 5117 29687 5151
rect 29687 5117 29696 5151
rect 29644 5108 29696 5117
rect 33508 5040 33560 5092
rect 30840 4972 30892 5024
rect 49424 4972 49476 5024
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 2780 4768 2832 4820
rect 4528 4768 4580 4820
rect 5356 4768 5408 4820
rect 7288 4768 7340 4820
rect 7472 4811 7524 4820
rect 7472 4777 7481 4811
rect 7481 4777 7515 4811
rect 7515 4777 7524 4811
rect 7472 4768 7524 4777
rect 8208 4768 8260 4820
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 1584 4700 1636 4752
rect 1308 4564 1360 4616
rect 1768 4564 1820 4616
rect 2964 4607 3016 4616
rect 2964 4573 2973 4607
rect 2973 4573 3007 4607
rect 3007 4573 3016 4607
rect 2964 4564 3016 4573
rect 3148 4607 3200 4616
rect 3148 4573 3157 4607
rect 3157 4573 3191 4607
rect 3191 4573 3200 4607
rect 3148 4564 3200 4573
rect 5724 4632 5776 4684
rect 7196 4632 7248 4684
rect 11428 4768 11480 4820
rect 12072 4811 12124 4820
rect 12072 4777 12081 4811
rect 12081 4777 12115 4811
rect 12115 4777 12124 4811
rect 12072 4768 12124 4777
rect 10876 4700 10928 4752
rect 14372 4768 14424 4820
rect 15108 4768 15160 4820
rect 16948 4768 17000 4820
rect 18604 4811 18656 4820
rect 18604 4777 18613 4811
rect 18613 4777 18647 4811
rect 18647 4777 18656 4811
rect 18604 4768 18656 4777
rect 18880 4768 18932 4820
rect 20996 4811 21048 4820
rect 20996 4777 21005 4811
rect 21005 4777 21039 4811
rect 21039 4777 21048 4811
rect 20996 4768 21048 4777
rect 22836 4768 22888 4820
rect 27344 4768 27396 4820
rect 31760 4768 31812 4820
rect 41420 4768 41472 4820
rect 16304 4700 16356 4752
rect 23756 4700 23808 4752
rect 29644 4700 29696 4752
rect 29736 4700 29788 4752
rect 34704 4700 34756 4752
rect 10968 4675 11020 4684
rect 10968 4641 10977 4675
rect 10977 4641 11011 4675
rect 11011 4641 11020 4675
rect 10968 4632 11020 4641
rect 11152 4632 11204 4684
rect 4620 4564 4672 4616
rect 5172 4607 5224 4616
rect 5172 4573 5181 4607
rect 5181 4573 5215 4607
rect 5215 4573 5224 4607
rect 5172 4564 5224 4573
rect 6276 4564 6328 4616
rect 6828 4607 6880 4616
rect 6828 4573 6837 4607
rect 6837 4573 6871 4607
rect 6871 4573 6880 4607
rect 6828 4564 6880 4573
rect 7012 4564 7064 4616
rect 9312 4607 9364 4616
rect 9312 4573 9321 4607
rect 9321 4573 9355 4607
rect 9355 4573 9364 4607
rect 9312 4564 9364 4573
rect 9404 4564 9456 4616
rect 12348 4564 12400 4616
rect 3516 4428 3568 4480
rect 5264 4428 5316 4480
rect 5908 4539 5960 4548
rect 5908 4505 5917 4539
rect 5917 4505 5951 4539
rect 5951 4505 5960 4539
rect 5908 4496 5960 4505
rect 6092 4539 6144 4548
rect 6092 4505 6101 4539
rect 6101 4505 6135 4539
rect 6135 4505 6144 4539
rect 6092 4496 6144 4505
rect 7564 4496 7616 4548
rect 6000 4428 6052 4480
rect 7472 4428 7524 4480
rect 12716 4564 12768 4616
rect 13728 4564 13780 4616
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 15660 4632 15712 4641
rect 19248 4632 19300 4684
rect 20720 4632 20772 4684
rect 21916 4675 21968 4684
rect 21916 4641 21925 4675
rect 21925 4641 21959 4675
rect 21959 4641 21968 4675
rect 21916 4632 21968 4641
rect 22560 4632 22612 4684
rect 27068 4675 27120 4684
rect 27068 4641 27077 4675
rect 27077 4641 27111 4675
rect 27111 4641 27120 4675
rect 27068 4632 27120 4641
rect 27160 4632 27212 4684
rect 30748 4632 30800 4684
rect 12624 4496 12676 4548
rect 14464 4496 14516 4548
rect 13636 4428 13688 4480
rect 13728 4428 13780 4480
rect 17408 4496 17460 4548
rect 17868 4564 17920 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 22192 4496 22244 4548
rect 20352 4428 20404 4480
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 23480 4564 23532 4616
rect 21364 4428 21416 4437
rect 27804 4428 27856 4480
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 3148 4224 3200 4276
rect 1952 4156 2004 4208
rect 1492 4088 1544 4140
rect 2320 4088 2372 4140
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 2780 4020 2832 4072
rect 5540 4156 5592 4208
rect 6184 4224 6236 4276
rect 7472 4156 7524 4208
rect 4620 4131 4672 4140
rect 4620 4097 4629 4131
rect 4629 4097 4663 4131
rect 4663 4097 4672 4131
rect 4620 4088 4672 4097
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 7196 4131 7248 4140
rect 7196 4097 7205 4131
rect 7205 4097 7239 4131
rect 7239 4097 7248 4131
rect 7196 4088 7248 4097
rect 7656 4020 7708 4072
rect 11520 4224 11572 4276
rect 11704 4224 11756 4276
rect 13728 4224 13780 4276
rect 17868 4224 17920 4276
rect 19248 4224 19300 4276
rect 9956 4156 10008 4208
rect 8852 4131 8904 4140
rect 8852 4097 8861 4131
rect 8861 4097 8895 4131
rect 8895 4097 8904 4131
rect 8852 4088 8904 4097
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 10048 4088 10100 4140
rect 11428 4088 11480 4140
rect 12072 4088 12124 4140
rect 12164 4088 12216 4140
rect 14096 4156 14148 4208
rect 14280 4156 14332 4208
rect 13360 4088 13412 4140
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 14648 4131 14700 4140
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 14740 4088 14792 4140
rect 15292 4088 15344 4140
rect 15476 4088 15528 4140
rect 25136 4224 25188 4276
rect 9312 4020 9364 4029
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 11336 4020 11388 4072
rect 17132 4020 17184 4072
rect 20076 4020 20128 4072
rect 20628 4131 20680 4140
rect 20628 4097 20637 4131
rect 20637 4097 20671 4131
rect 20671 4097 20680 4131
rect 20628 4088 20680 4097
rect 20904 4020 20956 4072
rect 22836 4156 22888 4208
rect 9956 3952 10008 4004
rect 13452 3952 13504 4004
rect 13728 3952 13780 4004
rect 31208 3952 31260 4004
rect 2872 3884 2924 3936
rect 3516 3927 3568 3936
rect 3516 3893 3525 3927
rect 3525 3893 3559 3927
rect 3559 3893 3568 3927
rect 3516 3884 3568 3893
rect 8760 3884 8812 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 9496 3884 9548 3936
rect 12532 3884 12584 3936
rect 15292 3927 15344 3936
rect 15292 3893 15301 3927
rect 15301 3893 15335 3927
rect 15335 3893 15344 3927
rect 15292 3884 15344 3893
rect 15476 3884 15528 3936
rect 16120 3884 16172 3936
rect 19524 3927 19576 3936
rect 19524 3893 19533 3927
rect 19533 3893 19567 3927
rect 19567 3893 19576 3927
rect 19524 3884 19576 3893
rect 19892 3927 19944 3936
rect 19892 3893 19901 3927
rect 19901 3893 19935 3927
rect 19935 3893 19944 3927
rect 19892 3884 19944 3893
rect 21640 3884 21692 3936
rect 23480 3884 23532 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 2320 3723 2372 3732
rect 2320 3689 2329 3723
rect 2329 3689 2363 3723
rect 2363 3689 2372 3723
rect 2320 3680 2372 3689
rect 3976 3680 4028 3732
rect 2780 3612 2832 3664
rect 8668 3680 8720 3732
rect 9680 3680 9732 3732
rect 12164 3680 12216 3732
rect 13544 3680 13596 3732
rect 11336 3612 11388 3664
rect 18512 3680 18564 3732
rect 19892 3680 19944 3732
rect 21640 3680 21692 3732
rect 14556 3655 14608 3664
rect 14556 3621 14565 3655
rect 14565 3621 14599 3655
rect 14599 3621 14608 3655
rect 14556 3612 14608 3621
rect 15384 3612 15436 3664
rect 15752 3655 15804 3664
rect 15752 3621 15761 3655
rect 15761 3621 15795 3655
rect 15795 3621 15804 3655
rect 15752 3612 15804 3621
rect 15936 3655 15988 3664
rect 15936 3621 15945 3655
rect 15945 3621 15979 3655
rect 15979 3621 15988 3655
rect 15936 3612 15988 3621
rect 17132 3612 17184 3664
rect 21364 3612 21416 3664
rect 22100 3612 22152 3664
rect 28724 3612 28776 3664
rect 848 3544 900 3596
rect 9404 3544 9456 3596
rect 9772 3544 9824 3596
rect 1676 3519 1728 3528
rect 1676 3485 1685 3519
rect 1685 3485 1719 3519
rect 1719 3485 1728 3519
rect 1676 3476 1728 3485
rect 2780 3519 2832 3528
rect 2780 3485 2789 3519
rect 2789 3485 2823 3519
rect 2823 3485 2832 3519
rect 2780 3476 2832 3485
rect 1400 3408 1452 3460
rect 6000 3519 6052 3528
rect 6000 3485 6009 3519
rect 6009 3485 6043 3519
rect 6043 3485 6052 3519
rect 6000 3476 6052 3485
rect 6920 3476 6972 3528
rect 8300 3408 8352 3460
rect 8576 3451 8628 3460
rect 8576 3417 8585 3451
rect 8585 3417 8619 3451
rect 8619 3417 8628 3451
rect 8576 3408 8628 3417
rect 9496 3519 9548 3528
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9496 3476 9548 3485
rect 11888 3519 11940 3528
rect 11888 3485 11897 3519
rect 11897 3485 11931 3519
rect 11931 3485 11940 3519
rect 11888 3476 11940 3485
rect 9680 3408 9732 3460
rect 3884 3340 3936 3392
rect 4068 3340 4120 3392
rect 5816 3340 5868 3392
rect 11980 3408 12032 3460
rect 19524 3544 19576 3596
rect 21088 3544 21140 3596
rect 12348 3519 12400 3528
rect 12348 3485 12357 3519
rect 12357 3485 12391 3519
rect 12391 3485 12400 3519
rect 12348 3476 12400 3485
rect 14648 3476 14700 3528
rect 10508 3340 10560 3392
rect 15108 3451 15160 3460
rect 15108 3417 15117 3451
rect 15117 3417 15151 3451
rect 15151 3417 15160 3451
rect 15108 3408 15160 3417
rect 15752 3476 15804 3528
rect 17040 3476 17092 3528
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 17684 3476 17736 3528
rect 18420 3408 18472 3460
rect 17224 3340 17276 3392
rect 17684 3340 17736 3392
rect 18696 3340 18748 3392
rect 18880 3408 18932 3460
rect 28908 3476 28960 3528
rect 44088 3476 44140 3528
rect 27068 3408 27120 3460
rect 46756 3408 46808 3460
rect 19340 3340 19392 3392
rect 19800 3340 19852 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 9220 3068 9272 3120
rect 12072 3136 12124 3188
rect 15108 3136 15160 3188
rect 17592 3136 17644 3188
rect 17868 3136 17920 3188
rect 20812 3179 20864 3188
rect 20812 3145 20821 3179
rect 20821 3145 20855 3179
rect 20855 3145 20864 3179
rect 20812 3136 20864 3145
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 3884 3000 3936 3052
rect 8484 3000 8536 3052
rect 10600 3000 10652 3052
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 12164 3000 12216 3052
rect 1584 2975 1636 2984
rect 1584 2941 1593 2975
rect 1593 2941 1627 2975
rect 1627 2941 1636 2975
rect 1584 2932 1636 2941
rect 3332 2864 3384 2916
rect 3884 2864 3936 2916
rect 4068 2864 4120 2916
rect 9864 2932 9916 2984
rect 14832 3111 14884 3120
rect 14832 3077 14841 3111
rect 14841 3077 14875 3111
rect 14875 3077 14884 3111
rect 14832 3068 14884 3077
rect 15016 3111 15068 3120
rect 15016 3077 15025 3111
rect 15025 3077 15059 3111
rect 15059 3077 15068 3111
rect 15016 3068 15068 3077
rect 19892 3068 19944 3120
rect 22744 3068 22796 3120
rect 12716 3000 12768 3052
rect 13084 3043 13136 3052
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13544 3043 13596 3052
rect 13544 3009 13553 3043
rect 13553 3009 13587 3043
rect 13587 3009 13596 3043
rect 13544 3000 13596 3009
rect 17132 3000 17184 3052
rect 18420 3000 18472 3052
rect 18512 3043 18564 3052
rect 18512 3009 18521 3043
rect 18521 3009 18555 3043
rect 18555 3009 18564 3043
rect 18512 3000 18564 3009
rect 22192 3043 22244 3052
rect 22192 3009 22201 3043
rect 22201 3009 22235 3043
rect 22235 3009 22244 3043
rect 22192 3000 22244 3009
rect 15936 2932 15988 2984
rect 4160 2839 4212 2848
rect 4160 2805 4169 2839
rect 4169 2805 4203 2839
rect 4203 2805 4212 2839
rect 4160 2796 4212 2805
rect 8852 2864 8904 2916
rect 16396 2907 16448 2916
rect 16396 2873 16405 2907
rect 16405 2873 16439 2907
rect 16439 2873 16448 2907
rect 16396 2864 16448 2873
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 14188 2839 14240 2848
rect 14188 2805 14197 2839
rect 14197 2805 14231 2839
rect 14231 2805 14240 2839
rect 14188 2796 14240 2805
rect 15384 2839 15436 2848
rect 15384 2805 15393 2839
rect 15393 2805 15427 2839
rect 15427 2805 15436 2839
rect 15384 2796 15436 2805
rect 15936 2839 15988 2848
rect 15936 2805 15945 2839
rect 15945 2805 15979 2839
rect 15979 2805 15988 2839
rect 15936 2796 15988 2805
rect 20812 2796 20864 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 2044 2592 2096 2644
rect 5540 2592 5592 2644
rect 8300 2592 8352 2644
rect 13544 2592 13596 2644
rect 14004 2592 14056 2644
rect 15200 2592 15252 2644
rect 15936 2592 15988 2644
rect 16948 2635 17000 2644
rect 16948 2601 16957 2635
rect 16957 2601 16991 2635
rect 16991 2601 17000 2635
rect 16948 2592 17000 2601
rect 17592 2635 17644 2644
rect 17592 2601 17601 2635
rect 17601 2601 17635 2635
rect 17635 2601 17644 2635
rect 17592 2592 17644 2601
rect 17684 2592 17736 2644
rect 22008 2635 22060 2644
rect 22008 2601 22017 2635
rect 22017 2601 22051 2635
rect 22051 2601 22060 2635
rect 22008 2592 22060 2601
rect 22560 2635 22612 2644
rect 22560 2601 22569 2635
rect 22569 2601 22603 2635
rect 22603 2601 22612 2635
rect 22560 2592 22612 2601
rect 23388 2592 23440 2644
rect 25504 2635 25556 2644
rect 25504 2601 25513 2635
rect 25513 2601 25547 2635
rect 25547 2601 25556 2635
rect 25504 2592 25556 2601
rect 27804 2592 27856 2644
rect 30840 2635 30892 2644
rect 30840 2601 30849 2635
rect 30849 2601 30883 2635
rect 30883 2601 30892 2635
rect 30840 2592 30892 2601
rect 33508 2635 33560 2644
rect 33508 2601 33517 2635
rect 33517 2601 33551 2635
rect 33551 2601 33560 2635
rect 33508 2592 33560 2601
rect 1124 2524 1176 2576
rect 664 2456 716 2508
rect 3332 2456 3384 2508
rect 1308 2388 1360 2440
rect 1768 2388 1820 2440
rect 4068 2456 4120 2508
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 6184 2456 6236 2508
rect 6736 2456 6788 2508
rect 9404 2456 9456 2508
rect 4344 2431 4396 2440
rect 4344 2397 4353 2431
rect 4353 2397 4387 2431
rect 4387 2397 4396 2431
rect 4344 2388 4396 2397
rect 14188 2524 14240 2576
rect 15016 2524 15068 2576
rect 18420 2524 18472 2576
rect 12072 2456 12124 2508
rect 14648 2456 14700 2508
rect 15200 2388 15252 2440
rect 4896 2252 4948 2304
rect 12624 2320 12676 2372
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9036 2252 9088 2261
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 14372 2295 14424 2304
rect 14372 2261 14381 2295
rect 14381 2261 14415 2295
rect 14415 2261 14424 2295
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16396 2456 16448 2508
rect 19432 2567 19484 2576
rect 19432 2533 19441 2567
rect 19441 2533 19475 2567
rect 19475 2533 19484 2567
rect 19432 2524 19484 2533
rect 32404 2524 32456 2576
rect 16488 2388 16540 2440
rect 17776 2431 17828 2440
rect 17776 2397 17785 2431
rect 17785 2397 17819 2431
rect 17819 2397 17828 2431
rect 17776 2388 17828 2397
rect 36360 2499 36412 2508
rect 36360 2465 36369 2499
rect 36369 2465 36403 2499
rect 36403 2465 36412 2499
rect 36360 2456 36412 2465
rect 19432 2388 19484 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 22560 2388 22612 2440
rect 25412 2388 25464 2440
rect 28356 2431 28408 2440
rect 28356 2397 28365 2431
rect 28365 2397 28399 2431
rect 28399 2397 28408 2431
rect 28356 2388 28408 2397
rect 30748 2388 30800 2440
rect 33416 2388 33468 2440
rect 36084 2431 36136 2440
rect 36084 2397 36093 2431
rect 36093 2397 36127 2431
rect 36127 2397 36136 2431
rect 36084 2388 36136 2397
rect 14372 2252 14424 2261
rect 18788 2295 18840 2304
rect 18788 2261 18797 2295
rect 18797 2261 18831 2295
rect 18831 2261 18840 2295
rect 18788 2252 18840 2261
rect 18972 2295 19024 2304
rect 18972 2261 18981 2295
rect 18981 2261 19015 2295
rect 19015 2261 19024 2295
rect 20720 2363 20772 2372
rect 20720 2329 20729 2363
rect 20729 2329 20763 2363
rect 20763 2329 20772 2363
rect 20720 2320 20772 2329
rect 20904 2320 20956 2372
rect 28724 2320 28776 2372
rect 18972 2252 19024 2261
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 2872 2048 2924 2100
rect 11520 2048 11572 2100
rect 9036 1980 9088 2032
rect 15200 2048 15252 2100
rect 18788 2048 18840 2100
rect 19616 2048 19668 2100
rect 11704 1980 11756 2032
rect 22100 1980 22152 2032
rect 4160 1912 4212 1964
rect 17776 1912 17828 1964
rect 3424 1844 3476 1896
rect 15384 1844 15436 1896
rect 16488 1844 16540 1896
rect 17500 1844 17552 1896
rect 20904 1844 20956 1896
rect 3608 1776 3660 1828
rect 4344 1640 4396 1692
rect 11888 1708 11940 1760
rect 18972 1708 19024 1760
rect 10968 1640 11020 1692
rect 20720 1640 20772 1692
rect 1584 1572 1636 1624
rect 11152 1572 11204 1624
rect 3332 1504 3384 1556
rect 14372 1504 14424 1556
rect 10324 1436 10376 1488
rect 19340 1436 19392 1488
rect 572 1300 624 1352
rect 11060 1368 11112 1420
rect 16488 1368 16540 1420
rect 11336 1300 11388 1352
rect 5632 1232 5684 1284
rect 11704 1232 11756 1284
rect 22192 1300 22244 1352
rect 25320 1232 25372 1284
rect 13636 1164 13688 1216
rect 21456 1164 21508 1216
rect 22100 1164 22152 1216
rect 22468 1164 22520 1216
rect 35440 1164 35492 1216
rect 15752 1096 15804 1148
rect 25964 1096 26016 1148
rect 3700 1028 3752 1080
rect 18696 1028 18748 1080
rect 4804 960 4856 1012
rect 20352 960 20404 1012
rect 4712 892 4764 944
rect 17868 892 17920 944
rect 3976 824 4028 876
rect 21180 824 21232 876
rect 6644 756 6696 808
rect 16488 756 16540 808
rect 6368 688 6420 740
rect 34980 688 35032 740
rect 1492 552 1544 604
rect 21272 552 21324 604
rect 3516 484 3568 536
rect 18788 484 18840 536
rect 2228 416 2280 468
rect 15476 416 15528 468
rect 3792 212 3844 264
rect 18880 212 18932 264
rect 5908 144 5960 196
rect 20812 144 20864 196
<< metal2 >>
rect 1308 26376 1360 26382
rect 1308 26318 1360 26324
rect 2226 26330 2282 27000
rect 572 26308 624 26314
rect 572 26250 624 26256
rect 388 22568 440 22574
rect 388 22510 440 22516
rect 296 13932 348 13938
rect 296 13874 348 13880
rect 308 9042 336 13874
rect 400 13258 428 22510
rect 480 18896 532 18902
rect 480 18838 532 18844
rect 388 13252 440 13258
rect 388 13194 440 13200
rect 388 11620 440 11626
rect 388 11562 440 11568
rect 296 9036 348 9042
rect 296 8978 348 8984
rect 400 2774 428 11562
rect 492 9518 520 18838
rect 584 13326 612 26250
rect 848 24404 900 24410
rect 848 24346 900 24352
rect 756 23792 808 23798
rect 756 23734 808 23740
rect 664 19440 716 19446
rect 664 19382 716 19388
rect 676 15094 704 19382
rect 664 15088 716 15094
rect 664 15030 716 15036
rect 572 13320 624 13326
rect 572 13262 624 13268
rect 572 11552 624 11558
rect 572 11494 624 11500
rect 480 9512 532 9518
rect 480 9454 532 9460
rect 584 4978 612 11494
rect 664 9580 716 9586
rect 664 9522 716 9528
rect 676 5098 704 9522
rect 768 5846 796 23734
rect 860 9586 888 24346
rect 1124 20460 1176 20466
rect 1124 20402 1176 20408
rect 1032 19848 1084 19854
rect 1032 19790 1084 19796
rect 940 15428 992 15434
rect 940 15370 992 15376
rect 952 11898 980 15370
rect 940 11892 992 11898
rect 940 11834 992 11840
rect 848 9580 900 9586
rect 848 9522 900 9528
rect 938 9480 994 9489
rect 860 9438 938 9466
rect 756 5840 808 5846
rect 756 5782 808 5788
rect 664 5092 716 5098
rect 664 5034 716 5040
rect 584 4950 704 4978
rect 400 2746 612 2774
rect 584 1358 612 2746
rect 676 2514 704 4950
rect 860 3602 888 9438
rect 938 9415 994 9424
rect 940 9376 992 9382
rect 940 9318 992 9324
rect 848 3596 900 3602
rect 848 3538 900 3544
rect 664 2508 716 2514
rect 664 2450 716 2456
rect 952 1873 980 9318
rect 1044 8294 1072 19790
rect 1136 15706 1164 20402
rect 1320 17882 1348 26318
rect 2226 26302 2544 26330
rect 2226 26200 2282 26302
rect 2044 25628 2096 25634
rect 2044 25570 2096 25576
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1768 24064 1820 24070
rect 1768 24006 1820 24012
rect 1780 23866 1808 24006
rect 1768 23860 1820 23866
rect 1768 23802 1820 23808
rect 1872 23118 1900 25162
rect 1952 23588 2004 23594
rect 1952 23530 2004 23536
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1492 22092 1544 22098
rect 1492 22034 1544 22040
rect 1400 20392 1452 20398
rect 1504 20369 1532 22034
rect 1584 22024 1636 22030
rect 1584 21966 1636 21972
rect 1400 20334 1452 20340
rect 1490 20360 1546 20369
rect 1412 19145 1440 20334
rect 1490 20295 1546 20304
rect 1492 19916 1544 19922
rect 1492 19858 1544 19864
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1400 18828 1452 18834
rect 1400 18770 1452 18776
rect 1412 17921 1440 18770
rect 1504 18737 1532 19858
rect 1490 18728 1546 18737
rect 1490 18663 1546 18672
rect 1596 18612 1624 21966
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1688 20913 1716 21490
rect 1674 20904 1730 20913
rect 1674 20839 1730 20848
rect 1504 18584 1624 18612
rect 1398 17912 1454 17921
rect 1308 17876 1360 17882
rect 1398 17847 1454 17856
rect 1308 17818 1360 17824
rect 1216 17740 1268 17746
rect 1216 17682 1268 17688
rect 1228 17105 1256 17682
rect 1400 17536 1452 17542
rect 1400 17478 1452 17484
rect 1308 17128 1360 17134
rect 1214 17096 1270 17105
rect 1308 17070 1360 17076
rect 1214 17031 1270 17040
rect 1320 16697 1348 17070
rect 1306 16688 1362 16697
rect 1306 16623 1362 16632
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1320 16289 1348 16458
rect 1306 16280 1362 16289
rect 1306 16215 1362 16224
rect 1412 16164 1440 17478
rect 1228 16136 1440 16164
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 1122 13424 1178 13433
rect 1122 13359 1178 13368
rect 1136 12782 1164 13359
rect 1124 12776 1176 12782
rect 1124 12718 1176 12724
rect 1032 8288 1084 8294
rect 1032 8230 1084 8236
rect 1136 6934 1164 12718
rect 1228 9178 1256 16136
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15881 1348 15982
rect 1306 15872 1362 15881
rect 1306 15807 1362 15816
rect 1308 15564 1360 15570
rect 1308 15506 1360 15512
rect 1320 15473 1348 15506
rect 1306 15464 1362 15473
rect 1306 15399 1362 15408
rect 1306 15056 1362 15065
rect 1306 14991 1362 15000
rect 1320 14958 1348 14991
rect 1308 14952 1360 14958
rect 1308 14894 1360 14900
rect 1306 14648 1362 14657
rect 1306 14583 1362 14592
rect 1320 14482 1348 14583
rect 1308 14476 1360 14482
rect 1308 14418 1360 14424
rect 1306 14240 1362 14249
rect 1306 14175 1362 14184
rect 1320 13870 1348 14175
rect 1504 13938 1532 18584
rect 1584 17876 1636 17882
rect 1584 17818 1636 17824
rect 1596 13977 1624 17818
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1780 16574 1808 17138
rect 1780 16546 1900 16574
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1780 14890 1808 16050
rect 1872 15978 1900 16546
rect 1860 15972 1912 15978
rect 1860 15914 1912 15920
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1768 14884 1820 14890
rect 1768 14826 1820 14832
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1582 13968 1638 13977
rect 1492 13932 1544 13938
rect 1582 13903 1584 13912
rect 1492 13874 1544 13880
rect 1636 13903 1638 13912
rect 1584 13874 1636 13880
rect 1308 13864 1360 13870
rect 1308 13806 1360 13812
rect 1780 13716 1808 14554
rect 1504 13688 1808 13716
rect 1398 12200 1454 12209
rect 1398 12135 1454 12144
rect 1308 11824 1360 11830
rect 1308 11766 1360 11772
rect 1216 9172 1268 9178
rect 1216 9114 1268 9120
rect 1216 9036 1268 9042
rect 1216 8978 1268 8984
rect 1228 7585 1256 8978
rect 1320 8022 1348 11766
rect 1412 11218 1440 12135
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1504 11098 1532 13688
rect 1584 13320 1636 13326
rect 1582 13288 1584 13297
rect 1636 13288 1638 13297
rect 1582 13223 1638 13232
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1412 11070 1532 11098
rect 1412 9450 1440 11070
rect 1596 10810 1624 12038
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1596 10606 1624 10746
rect 1584 10600 1636 10606
rect 1584 10542 1636 10548
rect 1688 9874 1716 12718
rect 1780 11121 1808 13126
rect 1872 12238 1900 15438
rect 1964 13190 1992 23530
rect 2056 22642 2084 25570
rect 2136 25560 2188 25566
rect 2136 25502 2188 25508
rect 2044 22636 2096 22642
rect 2044 22578 2096 22584
rect 2044 21004 2096 21010
rect 2044 20946 2096 20952
rect 2056 19553 2084 20946
rect 2042 19544 2098 19553
rect 2042 19479 2098 19488
rect 2148 19378 2176 25502
rect 2226 24304 2282 24313
rect 2226 24239 2282 24248
rect 2240 24206 2268 24239
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2228 22568 2280 22574
rect 2228 22510 2280 22516
rect 2240 21185 2268 22510
rect 2226 21176 2282 21185
rect 2226 21111 2282 21120
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2136 19372 2188 19378
rect 2136 19314 2188 19320
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18329 2084 19246
rect 2136 19168 2188 19174
rect 2136 19110 2188 19116
rect 2042 18320 2098 18329
rect 2042 18255 2098 18264
rect 2044 18216 2096 18222
rect 2044 18158 2096 18164
rect 2056 17513 2084 18158
rect 2042 17504 2098 17513
rect 2042 17439 2098 17448
rect 2148 14618 2176 19110
rect 2136 14612 2188 14618
rect 2136 14554 2188 14560
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 2056 13394 2084 13767
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 2148 12628 2176 13874
rect 2056 12600 2176 12628
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1766 11112 1822 11121
rect 1766 11047 1822 11056
rect 1766 10840 1822 10849
rect 1766 10775 1822 10784
rect 1596 9846 1716 9874
rect 1492 9716 1544 9722
rect 1492 9658 1544 9664
rect 1400 9444 1452 9450
rect 1400 9386 1452 9392
rect 1398 9344 1454 9353
rect 1398 9279 1454 9288
rect 1308 8016 1360 8022
rect 1308 7958 1360 7964
rect 1214 7576 1270 7585
rect 1214 7511 1270 7520
rect 1216 7472 1268 7478
rect 1216 7414 1268 7420
rect 1124 6928 1176 6934
rect 1124 6870 1176 6876
rect 1228 2774 1256 7414
rect 1308 6316 1360 6322
rect 1308 6258 1360 6264
rect 1320 6089 1348 6258
rect 1306 6080 1362 6089
rect 1306 6015 1362 6024
rect 1308 5704 1360 5710
rect 1306 5672 1308 5681
rect 1360 5672 1362 5681
rect 1306 5607 1362 5616
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1320 4622 1348 5199
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1412 4026 1440 9279
rect 1504 8514 1532 9658
rect 1596 8809 1624 9846
rect 1674 9616 1730 9625
rect 1674 9551 1730 9560
rect 1582 8800 1638 8809
rect 1582 8735 1638 8744
rect 1596 8634 1624 8735
rect 1688 8634 1716 9551
rect 1584 8628 1636 8634
rect 1584 8570 1636 8576
rect 1676 8628 1728 8634
rect 1676 8570 1728 8576
rect 1780 8514 1808 10775
rect 1872 10674 1900 12038
rect 1952 11756 2004 11762
rect 1952 11698 2004 11704
rect 1964 10849 1992 11698
rect 1950 10840 2006 10849
rect 1950 10775 2006 10784
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1950 10568 2006 10577
rect 1950 10503 2006 10512
rect 1964 9897 1992 10503
rect 1950 9888 2006 9897
rect 1950 9823 2006 9832
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1504 8498 1624 8514
rect 1504 8492 1636 8498
rect 1504 8486 1584 8492
rect 1584 8434 1636 8440
rect 1688 8486 1808 8514
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1504 7546 1532 8191
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1596 7478 1624 8434
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1490 4856 1546 4865
rect 1490 4791 1546 4800
rect 1504 4146 1532 4791
rect 1596 4758 1624 5646
rect 1688 5386 1716 8486
rect 1872 8412 1900 9318
rect 1964 8430 1992 9590
rect 1780 8384 1900 8412
rect 1952 8424 2004 8430
rect 1780 6866 1808 8384
rect 1952 8366 2004 8372
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1766 6760 1822 6769
rect 1766 6695 1822 6704
rect 1780 6662 1808 6695
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1872 5574 1900 7346
rect 1964 6662 1992 8230
rect 1952 6656 2004 6662
rect 1952 6598 2004 6604
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1688 5358 1900 5386
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1584 4752 1636 4758
rect 1584 4694 1636 4700
rect 1492 4140 1544 4146
rect 1492 4082 1544 4088
rect 1412 3998 1532 4026
rect 1400 3460 1452 3466
rect 1400 3402 1452 3408
rect 1136 2746 1256 2774
rect 1136 2582 1164 2746
rect 1124 2576 1176 2582
rect 1124 2518 1176 2524
rect 1308 2440 1360 2446
rect 1306 2408 1308 2417
rect 1360 2408 1362 2417
rect 1306 2343 1362 2352
rect 938 1864 994 1873
rect 938 1799 994 1808
rect 572 1352 624 1358
rect 572 1294 624 1300
rect 1412 800 1440 3402
rect 1398 0 1454 800
rect 1504 610 1532 3998
rect 1688 3534 1716 4966
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 1584 2984 1636 2990
rect 1584 2926 1636 2932
rect 1596 2825 1624 2926
rect 1582 2816 1638 2825
rect 1582 2751 1638 2760
rect 1596 1630 1624 2751
rect 1780 2446 1808 4558
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1584 1624 1636 1630
rect 1584 1566 1636 1572
rect 1872 1465 1900 5358
rect 1964 4214 1992 6258
rect 2056 5778 2084 12600
rect 2240 12442 2268 20878
rect 2424 18970 2452 23598
rect 2516 21418 2544 26302
rect 2870 26200 2926 27000
rect 3514 26200 3570 27000
rect 4158 26200 4214 27000
rect 4802 26330 4858 27000
rect 4802 26302 5120 26330
rect 4802 26200 4858 26302
rect 2778 24440 2834 24449
rect 2778 24375 2834 24384
rect 2792 23662 2820 24375
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2596 23520 2648 23526
rect 2596 23462 2648 23468
rect 2504 21412 2556 21418
rect 2504 21354 2556 21360
rect 2608 20874 2636 23462
rect 2884 23322 2912 26200
rect 3330 25256 3386 25265
rect 3330 25191 3386 25200
rect 3344 24886 3372 25191
rect 3332 24880 3384 24886
rect 3332 24822 3384 24828
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 3528 24274 3556 26200
rect 3884 25764 3936 25770
rect 3884 25706 3936 25712
rect 3516 24268 3568 24274
rect 3516 24210 3568 24216
rect 3516 24064 3568 24070
rect 3516 24006 3568 24012
rect 3698 24032 3754 24041
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 2872 23316 2924 23322
rect 2872 23258 2924 23264
rect 2780 23044 2832 23050
rect 2780 22986 2832 22992
rect 2792 22250 2820 22986
rect 3330 22536 3386 22545
rect 3330 22471 3386 22480
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 2700 22222 2820 22250
rect 3344 22234 3372 22471
rect 3424 22432 3476 22438
rect 3424 22374 3476 22380
rect 3332 22228 3384 22234
rect 2700 21593 2728 22222
rect 3332 22170 3384 22176
rect 3332 22092 3384 22098
rect 3332 22034 3384 22040
rect 3344 22001 3372 22034
rect 3330 21992 3386 22001
rect 3330 21927 3386 21936
rect 3332 21888 3384 21894
rect 3332 21830 3384 21836
rect 2686 21584 2742 21593
rect 2686 21519 2742 21528
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2792 19961 2820 21422
rect 3344 21321 3372 21830
rect 3330 21312 3386 21321
rect 2950 21244 3258 21253
rect 3330 21247 3386 21256
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 2778 19952 2834 19961
rect 2778 19887 2834 19896
rect 3436 19854 3464 22374
rect 3424 19848 3476 19854
rect 2594 19816 2650 19825
rect 3424 19790 3476 19796
rect 2594 19751 2650 19760
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2424 16658 2452 18906
rect 2504 17604 2556 17610
rect 2504 17546 2556 17552
rect 2412 16652 2464 16658
rect 2412 16594 2464 16600
rect 2320 15564 2372 15570
rect 2320 15506 2372 15512
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2228 12164 2280 12170
rect 2228 12106 2280 12112
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2148 7478 2176 11086
rect 2240 10198 2268 12106
rect 2332 11354 2360 15506
rect 2412 15360 2464 15366
rect 2412 15302 2464 15308
rect 2424 12374 2452 15302
rect 2412 12368 2464 12374
rect 2412 12310 2464 12316
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2320 11348 2372 11354
rect 2320 11290 2372 11296
rect 2424 11286 2452 12174
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2320 10260 2372 10266
rect 2320 10202 2372 10208
rect 2228 10192 2280 10198
rect 2332 10169 2360 10202
rect 2228 10134 2280 10140
rect 2318 10160 2374 10169
rect 2318 10095 2374 10104
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2240 9178 2268 9522
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2240 7970 2268 9114
rect 2332 8362 2360 9862
rect 2424 9382 2452 11086
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2320 8356 2372 8362
rect 2320 8298 2372 8304
rect 2318 8120 2374 8129
rect 2424 8090 2452 8910
rect 2318 8055 2320 8064
rect 2372 8055 2374 8064
rect 2412 8084 2464 8090
rect 2320 8026 2372 8032
rect 2412 8026 2464 8032
rect 2410 7984 2466 7993
rect 2240 7942 2360 7970
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2136 7472 2188 7478
rect 2136 7414 2188 7420
rect 2136 6792 2188 6798
rect 2134 6760 2136 6769
rect 2188 6760 2190 6769
rect 2134 6695 2190 6704
rect 2044 5772 2096 5778
rect 2044 5714 2096 5720
rect 2240 5302 2268 7822
rect 2228 5296 2280 5302
rect 2228 5238 2280 5244
rect 2332 5148 2360 7942
rect 2410 7919 2466 7928
rect 2424 5370 2452 7919
rect 2516 7546 2544 17546
rect 2608 11898 2636 19751
rect 3424 19712 3476 19718
rect 3424 19654 3476 19660
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2780 17876 2832 17882
rect 2780 17818 2832 17824
rect 2792 16574 2820 17818
rect 2700 16546 2820 16574
rect 2700 15026 2728 16546
rect 2884 16402 2912 19246
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 3436 18834 3464 19654
rect 3424 18828 3476 18834
rect 3424 18770 3476 18776
rect 3436 18426 3464 18770
rect 3528 18766 3556 24006
rect 3698 23967 3754 23976
rect 3608 23248 3660 23254
rect 3606 23216 3608 23225
rect 3660 23216 3662 23225
rect 3606 23151 3662 23160
rect 3606 22128 3662 22137
rect 3606 22063 3662 22072
rect 3620 21554 3648 22063
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3608 21140 3660 21146
rect 3608 21082 3660 21088
rect 3620 18834 3648 21082
rect 3712 19786 3740 23967
rect 3896 23168 3924 25706
rect 4066 25664 4122 25673
rect 4066 25599 4122 25608
rect 4080 25090 4108 25599
rect 4068 25084 4120 25090
rect 4068 25026 4120 25032
rect 3974 24848 4030 24857
rect 3974 24783 4030 24792
rect 3988 24410 4016 24783
rect 3976 24404 4028 24410
rect 3976 24346 4028 24352
rect 4172 23730 4200 26200
rect 4802 25120 4858 25129
rect 4802 25055 4858 25064
rect 4528 25016 4580 25022
rect 4528 24958 4580 24964
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 4066 23624 4122 23633
rect 4122 23582 4476 23610
rect 4066 23559 4122 23568
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 3896 23140 4016 23168
rect 3882 23080 3938 23089
rect 3882 23015 3938 23024
rect 3790 22808 3846 22817
rect 3790 22743 3846 22752
rect 3804 21146 3832 22743
rect 3792 21140 3844 21146
rect 3792 21082 3844 21088
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 3804 20777 3832 20946
rect 3790 20768 3846 20777
rect 3790 20703 3846 20712
rect 3792 20596 3844 20602
rect 3792 20538 3844 20544
rect 3804 20058 3832 20538
rect 3792 20052 3844 20058
rect 3792 19994 3844 20000
rect 3700 19780 3752 19786
rect 3700 19722 3752 19728
rect 3700 19440 3752 19446
rect 3700 19382 3752 19388
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3516 18760 3568 18766
rect 3516 18702 3568 18708
rect 3608 18624 3660 18630
rect 3608 18566 3660 18572
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3620 18329 3648 18566
rect 3606 18320 3662 18329
rect 3332 18284 3384 18290
rect 3606 18255 3662 18264
rect 3332 18226 3384 18232
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 2792 16374 2912 16402
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2792 14822 2820 16374
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 2950 15739 3258 15748
rect 2872 15700 2924 15706
rect 2872 15642 2924 15648
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2780 14816 2832 14822
rect 2780 14758 2832 14764
rect 2700 14498 2728 14758
rect 2700 14470 2820 14498
rect 2792 11914 2820 14470
rect 2884 13161 2912 15642
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3344 13274 3372 18226
rect 3606 17776 3662 17785
rect 3606 17711 3608 17720
rect 3660 17711 3662 17720
rect 3608 17682 3660 17688
rect 3424 16720 3476 16726
rect 3422 16688 3424 16697
rect 3608 16720 3660 16726
rect 3476 16688 3478 16697
rect 3422 16623 3478 16632
rect 3528 16680 3608 16708
rect 3422 15464 3478 15473
rect 3422 15399 3424 15408
rect 3476 15399 3478 15408
rect 3424 15370 3476 15376
rect 3424 14816 3476 14822
rect 3424 14758 3476 14764
rect 3436 13394 3464 14758
rect 3528 14618 3556 16680
rect 3608 16662 3660 16668
rect 3608 15632 3660 15638
rect 3606 15600 3608 15609
rect 3660 15600 3662 15609
rect 3606 15535 3662 15544
rect 3608 15428 3660 15434
rect 3608 15370 3660 15376
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3620 14414 3648 15370
rect 3712 15201 3740 19382
rect 3896 18222 3924 23015
rect 3988 22166 4016 23140
rect 4068 22568 4120 22574
rect 4068 22510 4120 22516
rect 3976 22160 4028 22166
rect 3976 22102 4028 22108
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 3988 21593 4016 21966
rect 3974 21584 4030 21593
rect 3974 21519 4030 21528
rect 4080 21162 4108 22510
rect 4172 21486 4200 23258
rect 4344 22228 4396 22234
rect 4344 22170 4396 22176
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4160 21480 4212 21486
rect 4160 21422 4212 21428
rect 3988 21134 4108 21162
rect 3988 20618 4016 21134
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 4080 20942 4108 20975
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3988 20590 4108 20618
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3988 20233 4016 20402
rect 3974 20224 4030 20233
rect 3974 20159 4030 20168
rect 3988 19446 4016 20159
rect 3976 19440 4028 19446
rect 3976 19382 4028 19388
rect 3884 18216 3936 18222
rect 4080 18193 4108 20590
rect 4264 20534 4292 22102
rect 4252 20528 4304 20534
rect 4252 20470 4304 20476
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3884 18158 3936 18164
rect 4066 18184 4122 18193
rect 4066 18119 4122 18128
rect 3884 17672 3936 17678
rect 3884 17614 3936 17620
rect 3896 16969 3924 17614
rect 4172 17134 4200 19722
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 4264 17610 4292 19654
rect 4356 19446 4384 22170
rect 4448 21622 4476 23582
rect 4540 22778 4568 24958
rect 4816 24206 4844 25055
rect 4896 24880 4948 24886
rect 4896 24822 4948 24828
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4724 23497 4752 24142
rect 4710 23488 4766 23497
rect 4710 23423 4766 23432
rect 4528 22772 4580 22778
rect 4528 22714 4580 22720
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4436 21616 4488 21622
rect 4436 21558 4488 21564
rect 4528 20392 4580 20398
rect 4528 20334 4580 20340
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4344 17672 4396 17678
rect 4342 17640 4344 17649
rect 4396 17640 4398 17649
rect 4252 17604 4304 17610
rect 4342 17575 4398 17584
rect 4252 17546 4304 17552
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3882 16960 3938 16969
rect 3882 16895 3938 16904
rect 3792 16652 3844 16658
rect 3792 16594 3844 16600
rect 3698 15192 3754 15201
rect 3698 15127 3754 15136
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3608 14272 3660 14278
rect 3606 14240 3608 14249
rect 3660 14240 3662 14249
rect 3606 14175 3662 14184
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3516 13864 3568 13870
rect 3514 13832 3516 13841
rect 3568 13832 3570 13841
rect 3514 13767 3570 13776
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3514 13288 3570 13297
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 3252 13025 3280 13262
rect 3344 13246 3464 13274
rect 2870 13016 2926 13025
rect 2870 12951 2926 12960
rect 3238 13016 3294 13025
rect 3238 12951 3294 12960
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2700 11886 2820 11914
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2608 11218 2636 11494
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2596 10464 2648 10470
rect 2596 10406 2648 10412
rect 2608 8566 2636 10406
rect 2700 9722 2728 11886
rect 2780 11756 2832 11762
rect 2780 11698 2832 11704
rect 2792 11014 2820 11698
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2688 9376 2740 9382
rect 2688 9318 2740 9324
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 2596 8424 2648 8430
rect 2596 8366 2648 8372
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2608 7154 2636 8366
rect 2516 7126 2636 7154
rect 2412 5364 2464 5370
rect 2412 5306 2464 5312
rect 2148 5120 2360 5148
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2148 2774 2176 5120
rect 2320 4140 2372 4146
rect 2320 4082 2372 4088
rect 2332 3738 2360 4082
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 2516 2774 2544 7126
rect 2700 7018 2728 9318
rect 2792 9092 2820 10406
rect 2884 9654 2912 12951
rect 3252 12918 3280 12951
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3344 12345 3372 12650
rect 3330 12336 3386 12345
rect 3330 12271 3386 12280
rect 3238 11792 3294 11801
rect 3238 11727 3294 11736
rect 3332 11756 3384 11762
rect 3252 11694 3280 11727
rect 3332 11698 3384 11704
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 2962 10840 3018 10849
rect 2962 10775 3018 10784
rect 2976 10538 3004 10775
rect 3056 10668 3108 10674
rect 3056 10610 3108 10616
rect 3068 10577 3096 10610
rect 3054 10568 3110 10577
rect 2964 10532 3016 10538
rect 3054 10503 3110 10512
rect 2964 10474 3016 10480
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 3148 10260 3200 10266
rect 3148 10202 3200 10208
rect 2964 10192 3016 10198
rect 3160 10169 3188 10202
rect 3240 10192 3292 10198
rect 2964 10134 3016 10140
rect 3146 10160 3202 10169
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 2976 9489 3004 10134
rect 3240 10134 3292 10140
rect 3146 10095 3202 10104
rect 2962 9480 3018 9489
rect 3252 9450 3280 10134
rect 2962 9415 3018 9424
rect 3240 9444 3292 9450
rect 3240 9386 3292 9392
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 2792 9064 3004 9092
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2792 7750 2820 8910
rect 2976 8401 3004 9064
rect 2962 8392 3018 8401
rect 2962 8327 3018 8336
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 2608 7002 2728 7018
rect 2596 6996 2728 7002
rect 2648 6990 2728 6996
rect 2596 6938 2648 6944
rect 2688 6928 2740 6934
rect 2740 6886 2820 6914
rect 2688 6870 2740 6876
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 5545 2636 6734
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2594 5536 2650 5545
rect 2594 5471 2650 5480
rect 2700 4729 2728 6190
rect 2792 4826 2820 6886
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3252 6497 3280 6666
rect 3238 6488 3294 6497
rect 3344 6458 3372 11698
rect 3238 6423 3294 6432
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3332 6112 3384 6118
rect 3332 6054 3384 6060
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3344 5846 3372 6054
rect 3436 5846 3464 13246
rect 3514 13223 3570 13232
rect 3528 13190 3556 13223
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3516 12640 3568 12646
rect 3516 12582 3568 12588
rect 3528 11354 3556 12582
rect 3620 11762 3648 14010
rect 3712 12986 3740 14962
rect 3804 13802 3832 16594
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3974 15056 4030 15065
rect 3974 14991 4030 15000
rect 3988 14958 4016 14991
rect 4080 14958 4108 15302
rect 3976 14952 4028 14958
rect 3882 14920 3938 14929
rect 3976 14894 4028 14900
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 3882 14855 3938 14864
rect 3896 14006 3924 14855
rect 3884 14000 3936 14006
rect 3884 13942 3936 13948
rect 3792 13796 3844 13802
rect 3792 13738 3844 13744
rect 3976 13728 4028 13734
rect 3790 13696 3846 13705
rect 3976 13670 4028 13676
rect 3790 13631 3846 13640
rect 3804 13530 3832 13631
rect 3792 13524 3844 13530
rect 3792 13466 3844 13472
rect 3790 13424 3846 13433
rect 3790 13359 3846 13368
rect 3884 13388 3936 13394
rect 3700 12980 3752 12986
rect 3700 12922 3752 12928
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3712 12073 3740 12786
rect 3698 12064 3754 12073
rect 3698 11999 3754 12008
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3804 11642 3832 13359
rect 3884 13330 3936 13336
rect 3896 12646 3924 13330
rect 3884 12640 3936 12646
rect 3884 12582 3936 12588
rect 3882 12472 3938 12481
rect 3882 12407 3938 12416
rect 3620 11614 3832 11642
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3516 11144 3568 11150
rect 3516 11086 3568 11092
rect 3528 7886 3556 11086
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3514 7712 3570 7721
rect 3514 7647 3570 7656
rect 3528 7274 3556 7647
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 6633 3556 6734
rect 3514 6624 3570 6633
rect 3514 6559 3570 6568
rect 3516 6180 3568 6186
rect 3516 6122 3568 6128
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 2962 5264 3018 5273
rect 2962 5199 3018 5208
rect 2976 5166 3004 5199
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 2686 4720 2742 4729
rect 2686 4655 2742 4664
rect 3146 4720 3202 4729
rect 3146 4655 3202 4664
rect 3160 4622 3188 4655
rect 2964 4616 3016 4622
rect 2962 4584 2964 4593
rect 3148 4616 3200 4622
rect 3016 4584 3018 4593
rect 3148 4558 3200 4564
rect 2962 4519 3018 4528
rect 3160 4282 3188 4558
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2792 3670 2820 4014
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 2056 2746 2176 2774
rect 2240 2746 2544 2774
rect 2056 2650 2084 2746
rect 2044 2644 2096 2650
rect 2044 2586 2096 2592
rect 1858 1456 1914 1465
rect 1858 1391 1914 1400
rect 1492 604 1544 610
rect 1492 546 1544 552
rect 2240 474 2268 2746
rect 2792 2553 2820 3470
rect 2778 2544 2834 2553
rect 2778 2479 2834 2488
rect 2884 2106 2912 3878
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3068 3058 3096 3431
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3344 2922 3372 5782
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 3330 2680 3386 2689
rect 3330 2615 3386 2624
rect 3344 2514 3372 2615
rect 3332 2508 3384 2514
rect 3332 2450 3384 2456
rect 3436 2394 3464 5306
rect 3528 4486 3556 6122
rect 3620 5250 3648 11614
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3712 9722 3740 11494
rect 3790 11248 3846 11257
rect 3790 11183 3846 11192
rect 3804 10198 3832 11183
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3700 9716 3752 9722
rect 3700 9658 3752 9664
rect 3790 9616 3846 9625
rect 3700 9580 3752 9586
rect 3790 9551 3846 9560
rect 3700 9522 3752 9528
rect 3712 6934 3740 9522
rect 3804 9178 3832 9551
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3700 6928 3752 6934
rect 3700 6870 3752 6876
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3712 5846 3740 6598
rect 3804 6390 3832 8978
rect 3792 6384 3844 6390
rect 3792 6326 3844 6332
rect 3790 6080 3846 6089
rect 3790 6015 3846 6024
rect 3700 5840 3752 5846
rect 3700 5782 3752 5788
rect 3804 5710 3832 6015
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3896 5370 3924 12407
rect 3988 8634 4016 13670
rect 4080 12714 4108 14894
rect 4264 14793 4292 17138
rect 4448 15162 4476 19790
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4250 14784 4306 14793
rect 4250 14719 4306 14728
rect 4540 14074 4568 20334
rect 4632 19378 4660 22170
rect 4908 22094 4936 24822
rect 4988 23588 5040 23594
rect 4988 23530 5040 23536
rect 4816 22066 4936 22094
rect 4816 19938 4844 22066
rect 4724 19910 4844 19938
rect 4620 19372 4672 19378
rect 4620 19314 4672 19320
rect 4620 16448 4672 16454
rect 4620 16390 4672 16396
rect 4528 14068 4580 14074
rect 4528 14010 4580 14016
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 4172 13326 4200 13942
rect 4250 13560 4306 13569
rect 4250 13495 4252 13504
rect 4304 13495 4306 13504
rect 4344 13524 4396 13530
rect 4252 13466 4304 13472
rect 4344 13466 4396 13472
rect 4160 13320 4212 13326
rect 4356 13308 4384 13466
rect 4160 13262 4212 13268
rect 4264 13280 4384 13308
rect 4172 12986 4200 13262
rect 4160 12980 4212 12986
rect 4160 12922 4212 12928
rect 4172 12850 4200 12922
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4172 12458 4200 12582
rect 4080 12430 4200 12458
rect 4264 12442 4292 13280
rect 4632 13172 4660 16390
rect 4724 16182 4752 19910
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4816 17746 4844 19722
rect 4894 19136 4950 19145
rect 4894 19071 4950 19080
rect 4804 17740 4856 17746
rect 4804 17682 4856 17688
rect 4712 16176 4764 16182
rect 4712 16118 4764 16124
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4724 14958 4752 15982
rect 4816 15570 4844 17682
rect 4804 15564 4856 15570
rect 4804 15506 4856 15512
rect 4712 14952 4764 14958
rect 4712 14894 4764 14900
rect 4724 14113 4752 14894
rect 4816 14414 4844 15506
rect 4908 15502 4936 19071
rect 5000 16590 5028 23530
rect 5092 22574 5120 26302
rect 5264 26240 5316 26246
rect 5446 26200 5502 27000
rect 6090 26200 6146 27000
rect 6734 26330 6790 27000
rect 6734 26302 6868 26330
rect 6734 26200 6790 26302
rect 5264 26182 5316 26188
rect 5276 23186 5304 26182
rect 5460 23662 5488 26200
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5448 23656 5500 23662
rect 5448 23598 5500 23604
rect 5356 23588 5408 23594
rect 5356 23530 5408 23536
rect 5264 23180 5316 23186
rect 5264 23122 5316 23128
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5172 17604 5224 17610
rect 5172 17546 5224 17552
rect 4988 16584 5040 16590
rect 4988 16526 5040 16532
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 5000 14346 5028 15846
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 5092 14482 5120 14758
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 4988 14340 5040 14346
rect 4988 14282 5040 14288
rect 5184 14226 5212 17546
rect 5276 16454 5304 20334
rect 5368 18034 5396 23530
rect 5538 22672 5594 22681
rect 5538 22607 5594 22616
rect 5552 21962 5580 22607
rect 5540 21956 5592 21962
rect 5540 21898 5592 21904
rect 5736 21690 5764 24890
rect 6104 23186 6132 26200
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6182 25528 6238 25537
rect 6182 25463 6238 25472
rect 6092 23180 6144 23186
rect 6092 23122 6144 23128
rect 6196 23118 6224 25463
rect 6552 24812 6604 24818
rect 6552 24754 6604 24760
rect 6564 24206 6592 24754
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6184 23112 6236 23118
rect 6184 23054 6236 23060
rect 6656 22574 6684 25774
rect 6736 25152 6788 25158
rect 6736 25094 6788 25100
rect 6748 23730 6776 25094
rect 6736 23724 6788 23730
rect 6736 23666 6788 23672
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6000 22500 6052 22506
rect 6000 22442 6052 22448
rect 5816 21888 5868 21894
rect 5816 21830 5868 21836
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5828 21593 5856 21830
rect 5814 21584 5870 21593
rect 5632 21548 5684 21554
rect 5814 21519 5870 21528
rect 5632 21490 5684 21496
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5460 19360 5488 21286
rect 5540 20800 5592 20806
rect 5644 20777 5672 21490
rect 5816 20868 5868 20874
rect 5816 20810 5868 20816
rect 5724 20800 5776 20806
rect 5540 20742 5592 20748
rect 5630 20768 5686 20777
rect 5552 20505 5580 20742
rect 5724 20742 5776 20748
rect 5630 20703 5686 20712
rect 5538 20496 5594 20505
rect 5538 20431 5594 20440
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5644 19718 5672 20402
rect 5736 20262 5764 20742
rect 5724 20256 5776 20262
rect 5724 20198 5776 20204
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5724 19508 5776 19514
rect 5724 19450 5776 19456
rect 5460 19332 5672 19360
rect 5368 18006 5580 18034
rect 5264 16448 5316 16454
rect 5264 16390 5316 16396
rect 5552 15201 5580 18006
rect 5644 15314 5672 19332
rect 5736 18630 5764 19450
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5828 18358 5856 20810
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5920 20369 5948 20742
rect 5906 20360 5962 20369
rect 5906 20295 5962 20304
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5816 18352 5868 18358
rect 5816 18294 5868 18300
rect 5920 18222 5948 20198
rect 6012 18766 6040 22442
rect 6840 22094 6868 26302
rect 7378 26200 7434 27000
rect 7748 26988 7800 26994
rect 7748 26930 7800 26936
rect 7104 25288 7156 25294
rect 7104 25230 7156 25236
rect 7012 22094 7064 22098
rect 6840 22092 7064 22094
rect 6840 22066 7012 22092
rect 7012 22034 7064 22040
rect 6920 22024 6972 22030
rect 7024 22003 7052 22034
rect 6920 21966 6972 21972
rect 6828 21888 6880 21894
rect 6828 21830 6880 21836
rect 6276 21616 6328 21622
rect 6276 21558 6328 21564
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6196 19922 6224 20878
rect 6184 19916 6236 19922
rect 6184 19858 6236 19864
rect 6184 19712 6236 19718
rect 6184 19654 6236 19660
rect 6196 19514 6224 19654
rect 6184 19508 6236 19514
rect 6184 19450 6236 19456
rect 6092 19236 6144 19242
rect 6092 19178 6144 19184
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6104 18601 6132 19178
rect 6090 18592 6146 18601
rect 6090 18527 6146 18536
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 6092 18216 6144 18222
rect 6092 18158 6144 18164
rect 5736 17066 5764 18158
rect 5920 17134 5948 18158
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 5908 17128 5960 17134
rect 5908 17070 5960 17076
rect 5724 17060 5776 17066
rect 5724 17002 5776 17008
rect 5816 16516 5868 16522
rect 5816 16458 5868 16464
rect 5644 15286 5764 15314
rect 5538 15192 5594 15201
rect 5736 15162 5764 15286
rect 5538 15127 5594 15136
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4908 14198 5212 14226
rect 4710 14104 4766 14113
rect 4710 14039 4766 14048
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4356 13144 4660 13172
rect 4252 12436 4304 12442
rect 4080 11150 4108 12430
rect 4252 12378 4304 12384
rect 4356 12322 4384 13144
rect 4436 12912 4488 12918
rect 4436 12854 4488 12860
rect 4264 12294 4384 12322
rect 4264 11558 4292 12294
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4066 10432 4122 10441
rect 4066 10367 4122 10376
rect 4080 10198 4108 10367
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 4080 9450 4108 9930
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3988 6712 4016 7822
rect 4080 7410 4108 8298
rect 4172 7546 4200 11018
rect 4356 10198 4384 12174
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4342 10024 4398 10033
rect 4342 9959 4398 9968
rect 4250 9616 4306 9625
rect 4250 9551 4252 9560
rect 4304 9551 4306 9560
rect 4252 9522 4304 9528
rect 4356 8906 4384 9959
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4250 8528 4306 8537
rect 4250 8463 4306 8472
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4264 6798 4292 8463
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4356 6798 4384 7958
rect 4448 7546 4476 12854
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 8129 4568 12106
rect 4632 12102 4660 12582
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4526 8120 4582 8129
rect 4526 8055 4582 8064
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4632 7206 4660 11630
rect 4724 8974 4752 13670
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4816 12238 4844 12922
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 11218 4844 12174
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4802 11112 4858 11121
rect 4802 11047 4858 11056
rect 4816 10606 4844 11047
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 4816 9382 4844 10542
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 8968 4764 8974
rect 4908 8922 4936 14198
rect 4986 14104 5042 14113
rect 4986 14039 4988 14048
rect 5040 14039 5042 14048
rect 4988 14010 5040 14016
rect 5000 13394 5028 14010
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 4988 13388 5040 13394
rect 4988 13330 5040 13336
rect 5000 12594 5028 13330
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5092 12889 5120 13194
rect 5078 12880 5134 12889
rect 5078 12815 5134 12824
rect 5184 12646 5212 13398
rect 5276 13394 5304 14758
rect 5368 13734 5396 14894
rect 5552 14822 5580 15030
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5724 14476 5776 14482
rect 5724 14418 5776 14424
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5356 13728 5408 13734
rect 5356 13670 5408 13676
rect 5460 13410 5488 14214
rect 5552 14006 5580 14214
rect 5540 14000 5592 14006
rect 5540 13942 5592 13948
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5368 13382 5488 13410
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5172 12640 5224 12646
rect 5078 12608 5134 12617
rect 5000 12566 5078 12594
rect 5172 12582 5224 12588
rect 5078 12543 5134 12552
rect 5172 12368 5224 12374
rect 5078 12336 5134 12345
rect 5172 12310 5224 12316
rect 5078 12271 5134 12280
rect 4986 12200 5042 12209
rect 4986 12135 5042 12144
rect 5000 12102 5028 12135
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 5000 11694 5028 12038
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4712 8910 4764 8916
rect 4816 8894 4936 8922
rect 4712 8832 4764 8838
rect 4712 8774 4764 8780
rect 4724 7410 4752 8774
rect 4816 8090 4844 8894
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8498 4936 8774
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 5000 8344 5028 10610
rect 5092 9489 5120 12271
rect 5184 11937 5212 12310
rect 5170 11928 5226 11937
rect 5170 11863 5226 11872
rect 5276 11830 5304 12922
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 5184 10538 5212 11698
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5172 10532 5224 10538
rect 5172 10474 5224 10480
rect 5078 9480 5134 9489
rect 5276 9466 5304 11630
rect 5368 10690 5396 13382
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12374 5488 13126
rect 5644 12730 5672 14282
rect 5736 12986 5764 14418
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5552 12702 5672 12730
rect 5448 12368 5500 12374
rect 5448 12310 5500 12316
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5460 11898 5488 12174
rect 5448 11892 5500 11898
rect 5448 11834 5500 11840
rect 5368 10674 5488 10690
rect 5368 10668 5500 10674
rect 5368 10662 5448 10668
rect 5448 10610 5500 10616
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5078 9415 5080 9424
rect 5132 9415 5134 9424
rect 5184 9438 5304 9466
rect 5080 9386 5132 9392
rect 5000 8316 5120 8344
rect 4986 8256 5042 8265
rect 4986 8191 5042 8200
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4802 7984 4858 7993
rect 4802 7919 4858 7928
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4434 7032 4490 7041
rect 4434 6967 4490 6976
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 3988 6684 4108 6712
rect 4080 6458 4108 6684
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 4068 6452 4120 6458
rect 4068 6394 4120 6400
rect 3988 6254 4016 6394
rect 4158 6352 4214 6361
rect 4068 6316 4120 6322
rect 4158 6287 4214 6296
rect 4068 6258 4120 6264
rect 3976 6248 4028 6254
rect 3976 6190 4028 6196
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3620 5222 3924 5250
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3698 4448 3754 4457
rect 3698 4383 3754 4392
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 3058 3556 3878
rect 3606 3632 3662 3641
rect 3606 3567 3662 3576
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3344 2366 3464 2394
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 3344 1562 3372 2366
rect 3514 2000 3570 2009
rect 3514 1935 3570 1944
rect 3424 1896 3476 1902
rect 3424 1838 3476 1844
rect 3436 1601 3464 1838
rect 3422 1592 3478 1601
rect 3332 1556 3384 1562
rect 3422 1527 3478 1536
rect 3332 1498 3384 1504
rect 3528 542 3556 1935
rect 3620 1834 3648 3567
rect 3608 1828 3660 1834
rect 3608 1770 3660 1776
rect 3712 1086 3740 4383
rect 3790 4040 3846 4049
rect 3790 3975 3846 3984
rect 3700 1080 3752 1086
rect 3700 1022 3752 1028
rect 3516 536 3568 542
rect 3516 478 3568 484
rect 2228 468 2280 474
rect 2228 410 2280 416
rect 3804 270 3832 3975
rect 3896 3618 3924 5222
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3988 3738 4016 4082
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 3896 3590 4016 3618
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3058 3924 3334
rect 3884 3052 3936 3058
rect 3884 2994 3936 3000
rect 3884 2916 3936 2922
rect 3884 2858 3936 2864
rect 3896 921 3924 2858
rect 3882 912 3938 921
rect 3988 882 4016 3590
rect 4080 3398 4108 6258
rect 4172 6186 4200 6287
rect 4160 6180 4212 6186
rect 4160 6122 4212 6128
rect 4448 5914 4476 6967
rect 4618 6352 4674 6361
rect 4618 6287 4674 6296
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4632 5642 4660 6287
rect 4620 5636 4672 5642
rect 4620 5578 4672 5584
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4540 4826 4568 5170
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4632 4146 4660 4558
rect 4620 4140 4672 4146
rect 4620 4082 4672 4088
rect 4068 3392 4120 3398
rect 4068 3334 4120 3340
rect 4066 3224 4122 3233
rect 4066 3159 4122 3168
rect 4080 2922 4108 3159
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 3882 847 3938 856
rect 3976 876 4028 882
rect 3976 818 4028 824
rect 4080 800 4108 2450
rect 4172 1970 4200 2790
rect 4344 2440 4396 2446
rect 4344 2382 4396 2388
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4356 1698 4384 2382
rect 4344 1692 4396 1698
rect 4344 1634 4396 1640
rect 4724 950 4752 7210
rect 4816 1018 4844 7919
rect 4896 7812 4948 7818
rect 4896 7754 4948 7760
rect 4908 6458 4936 7754
rect 5000 7546 5028 8191
rect 5092 8090 5120 8316
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 5078 7984 5134 7993
rect 5078 7919 5134 7928
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 2310 4936 5510
rect 5092 5370 5120 7919
rect 5184 5574 5212 9438
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 8838 5304 9318
rect 5368 8838 5396 9998
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5276 7818 5304 8774
rect 5264 7812 5316 7818
rect 5264 7754 5316 7760
rect 5354 7440 5410 7449
rect 5354 7375 5410 7384
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5276 6798 5304 7278
rect 5368 7154 5396 7375
rect 5460 7274 5488 9862
rect 5552 8634 5580 12702
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5644 11830 5672 12582
rect 5736 11830 5764 12786
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5724 11824 5776 11830
rect 5724 11766 5776 11772
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 9648 5684 9654
rect 5630 9616 5632 9625
rect 5684 9616 5686 9625
rect 5630 9551 5686 9560
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9058 5672 9454
rect 5736 9382 5764 11630
rect 5828 11354 5856 16458
rect 6012 16153 6040 18022
rect 6104 16454 6132 18158
rect 6196 17678 6224 19450
rect 6288 18834 6316 21558
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20641 6500 20810
rect 6564 20777 6592 21286
rect 6840 21010 6868 21830
rect 6932 21185 6960 21966
rect 7116 21690 7144 25230
rect 7392 24274 7420 26200
rect 7564 25900 7616 25906
rect 7564 25842 7616 25848
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7380 24064 7432 24070
rect 7380 24006 7432 24012
rect 7288 23248 7340 23254
rect 7288 23190 7340 23196
rect 7104 21684 7156 21690
rect 7104 21626 7156 21632
rect 7104 21480 7156 21486
rect 7104 21422 7156 21428
rect 7012 21412 7064 21418
rect 7012 21354 7064 21360
rect 6918 21176 6974 21185
rect 6918 21111 6974 21120
rect 6828 21004 6880 21010
rect 6828 20946 6880 20952
rect 6550 20768 6606 20777
rect 6550 20703 6606 20712
rect 6458 20632 6514 20641
rect 6458 20567 6514 20576
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6552 20324 6604 20330
rect 6552 20266 6604 20272
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6564 19922 6592 20266
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6460 19712 6512 19718
rect 6460 19654 6512 19660
rect 6368 19440 6420 19446
rect 6368 19382 6420 19388
rect 6380 18902 6408 19382
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6276 18828 6328 18834
rect 6276 18770 6328 18776
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 5998 16144 6054 16153
rect 5998 16079 6054 16088
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 12594 6040 14758
rect 6104 13530 6132 16390
rect 6196 15366 6224 17614
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6380 15706 6408 17138
rect 6472 17105 6500 19654
rect 6564 19378 6592 19858
rect 6748 19718 6776 20266
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6736 19712 6788 19718
rect 6840 19689 6868 19722
rect 6736 19654 6788 19660
rect 6826 19680 6882 19689
rect 6748 19514 6776 19654
rect 6826 19615 6882 19624
rect 6736 19508 6788 19514
rect 6736 19450 6788 19456
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6552 17808 6604 17814
rect 6552 17750 6604 17756
rect 6564 17202 6592 17750
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6458 17096 6514 17105
rect 6458 17031 6514 17040
rect 6460 16516 6512 16522
rect 6460 16458 6512 16464
rect 6368 15700 6420 15706
rect 6368 15642 6420 15648
rect 6276 15632 6328 15638
rect 6276 15574 6328 15580
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6288 14618 6316 15574
rect 6276 14612 6328 14618
rect 6276 14554 6328 14560
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 14006 6408 14214
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6288 13734 6316 13874
rect 6276 13728 6328 13734
rect 6276 13670 6328 13676
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 5920 12566 6040 12594
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5920 10554 5948 12566
rect 5998 12472 6054 12481
rect 5998 12407 6054 12416
rect 6012 11937 6040 12407
rect 5998 11928 6054 11937
rect 5998 11863 6054 11872
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 5828 10526 5948 10554
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5644 9030 5764 9058
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5540 7200 5592 7206
rect 5368 7126 5488 7154
rect 5540 7142 5592 7148
rect 5356 6996 5408 7002
rect 5356 6938 5408 6944
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5368 6322 5396 6938
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5460 6202 5488 7126
rect 5552 6304 5580 7142
rect 5644 6458 5672 8910
rect 5736 8294 5764 9030
rect 5828 8401 5856 10526
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 8974 5948 10406
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5814 8392 5870 8401
rect 5814 8327 5870 8336
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5736 6361 5764 6734
rect 5722 6352 5778 6361
rect 5552 6276 5672 6304
rect 5722 6287 5778 6296
rect 5368 6174 5488 6202
rect 5538 6216 5594 6225
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5170 5400 5226 5409
rect 5080 5364 5132 5370
rect 5170 5335 5226 5344
rect 5080 5306 5132 5312
rect 5184 4622 5212 5335
rect 5368 4826 5396 6174
rect 5538 6151 5594 6160
rect 5446 5944 5502 5953
rect 5446 5879 5448 5888
rect 5500 5879 5502 5888
rect 5448 5850 5500 5856
rect 5552 5710 5580 6151
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5356 4820 5408 4826
rect 5356 4762 5408 4768
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5264 4480 5316 4486
rect 5264 4422 5316 4428
rect 5276 3097 5304 4422
rect 5354 4176 5410 4185
rect 5354 4111 5356 4120
rect 5408 4111 5410 4120
rect 5356 4082 5408 4088
rect 5262 3088 5318 3097
rect 5262 3023 5318 3032
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4804 1012 4856 1018
rect 4804 954 4856 960
rect 4712 944 4764 950
rect 4712 886 4764 892
rect 3792 264 3844 270
rect 3792 206 3844 212
rect 4066 0 4122 800
rect 5460 785 5488 4966
rect 5538 4720 5594 4729
rect 5538 4655 5594 4664
rect 5552 4214 5580 4655
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5552 2650 5580 4150
rect 5540 2644 5592 2650
rect 5540 2586 5592 2592
rect 5644 1290 5672 6276
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 4690 5764 5170
rect 5724 4684 5776 4690
rect 5724 4626 5776 4632
rect 5828 3641 5856 8026
rect 6012 6798 6040 11766
rect 6104 8090 6132 12718
rect 6196 12170 6224 12854
rect 6288 12850 6316 13330
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6380 12481 6408 13942
rect 6366 12472 6422 12481
rect 6276 12436 6328 12442
rect 6366 12407 6422 12416
rect 6276 12378 6328 12384
rect 6288 12345 6316 12378
rect 6274 12336 6330 12345
rect 6274 12271 6330 12280
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6196 11150 6224 12106
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6274 11928 6330 11937
rect 6274 11863 6330 11872
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6288 10146 6316 11863
rect 6196 10118 6316 10146
rect 6092 8084 6144 8090
rect 6092 8026 6144 8032
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6090 6080 6146 6089
rect 6090 6015 6146 6024
rect 6104 5681 6132 6015
rect 6090 5672 6146 5681
rect 6090 5607 6146 5616
rect 6196 5114 6224 10118
rect 6276 10056 6328 10062
rect 6276 9998 6328 10004
rect 6288 5137 6316 9998
rect 6380 9178 6408 12038
rect 6472 9654 6500 16458
rect 6642 16144 6698 16153
rect 6552 16108 6604 16114
rect 6642 16079 6644 16088
rect 6552 16050 6604 16056
rect 6696 16079 6698 16088
rect 6644 16050 6696 16056
rect 6564 15994 6592 16050
rect 6564 15966 6684 15994
rect 6552 15428 6604 15434
rect 6552 15370 6604 15376
rect 6564 14346 6592 15370
rect 6656 14618 6684 15966
rect 6748 15502 6776 18906
rect 6826 18048 6882 18057
rect 6826 17983 6882 17992
rect 6840 17542 6868 17983
rect 6932 17746 6960 20402
rect 7024 20398 7052 21354
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7116 19938 7144 21422
rect 7024 19910 7144 19938
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6828 17536 6880 17542
rect 6828 17478 6880 17484
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 17134 6960 17478
rect 6828 17128 6880 17134
rect 6828 17070 6880 17076
rect 6920 17128 6972 17134
rect 6920 17070 6972 17076
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 6840 15434 6868 17070
rect 6932 16833 6960 17070
rect 6918 16824 6974 16833
rect 6918 16759 6974 16768
rect 7024 16640 7052 19910
rect 7104 19780 7156 19786
rect 7104 19722 7156 19728
rect 7116 18086 7144 19722
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7208 17728 7236 19450
rect 7300 18222 7328 23190
rect 7392 21894 7420 24006
rect 7380 21888 7432 21894
rect 7380 21830 7432 21836
rect 7392 18970 7420 21830
rect 7380 18964 7432 18970
rect 7380 18906 7432 18912
rect 7484 18358 7512 24346
rect 7576 22642 7604 25842
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7576 21078 7604 21422
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7576 19689 7604 20878
rect 7562 19680 7618 19689
rect 7562 19615 7618 19624
rect 7576 19446 7604 19615
rect 7668 19514 7696 23462
rect 7760 22642 7788 26930
rect 8022 26330 8078 27000
rect 8666 26330 8722 27000
rect 7852 26302 8078 26330
rect 7852 23186 7880 26302
rect 8022 26200 8078 26302
rect 8588 26302 8722 26330
rect 8300 25696 8352 25702
rect 8300 25638 8352 25644
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7932 23656 7984 23662
rect 7984 23604 8156 23610
rect 7932 23598 8156 23604
rect 7944 23594 8156 23598
rect 7944 23588 8168 23594
rect 7944 23582 8116 23588
rect 8116 23530 8168 23536
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7840 23180 7892 23186
rect 7840 23122 7892 23128
rect 7944 23066 7972 23462
rect 8024 23316 8076 23322
rect 8024 23258 8076 23264
rect 8036 23118 8064 23258
rect 7852 23038 7972 23066
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7748 22636 7800 22642
rect 7748 22578 7800 22584
rect 7852 21010 7880 23038
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 8024 21480 8076 21486
rect 8024 21422 8076 21428
rect 7840 21004 7892 21010
rect 7840 20946 7892 20952
rect 8036 20913 8064 21422
rect 8022 20904 8078 20913
rect 8022 20839 8078 20848
rect 7840 20800 7892 20806
rect 7840 20742 7892 20748
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 19440 7616 19446
rect 7564 19382 7616 19388
rect 7564 18624 7616 18630
rect 7564 18566 7616 18572
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7380 18352 7432 18358
rect 7380 18294 7432 18300
rect 7472 18352 7524 18358
rect 7472 18294 7524 18300
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7208 17700 7328 17728
rect 7194 17640 7250 17649
rect 7194 17575 7250 17584
rect 7208 17202 7236 17575
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 7196 16652 7248 16658
rect 7024 16612 7196 16640
rect 6920 16448 6972 16454
rect 6920 16390 6972 16396
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6828 15020 6880 15026
rect 6828 14962 6880 14968
rect 6736 14816 6788 14822
rect 6736 14758 6788 14764
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6642 14376 6698 14385
rect 6552 14340 6604 14346
rect 6642 14311 6698 14320
rect 6552 14282 6604 14288
rect 6550 14104 6606 14113
rect 6550 14039 6606 14048
rect 6564 13802 6592 14039
rect 6656 14006 6684 14311
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6656 13258 6684 13670
rect 6644 13252 6696 13258
rect 6644 13194 6696 13200
rect 6748 13025 6776 14758
rect 6734 13016 6790 13025
rect 6840 12986 6868 14962
rect 6932 14074 6960 16390
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 7024 15065 7052 15370
rect 7010 15056 7066 15065
rect 7010 14991 7066 15000
rect 7116 14958 7144 16612
rect 7196 16594 7248 16600
rect 7300 16454 7328 17700
rect 7288 16448 7340 16454
rect 7288 16390 7340 16396
rect 7196 15360 7248 15366
rect 7196 15302 7248 15308
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7208 14822 7236 15302
rect 7300 14940 7328 16390
rect 7392 15065 7420 18294
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7484 17785 7512 17818
rect 7470 17776 7526 17785
rect 7470 17711 7526 17720
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7378 15056 7434 15065
rect 7378 14991 7434 15000
rect 7300 14912 7420 14940
rect 7196 14816 7248 14822
rect 7102 14784 7158 14793
rect 7196 14758 7248 14764
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7102 14719 7158 14728
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6734 12951 6790 12960
rect 6828 12980 6880 12986
rect 6828 12922 6880 12928
rect 6550 12880 6606 12889
rect 6550 12815 6552 12824
rect 6604 12815 6606 12824
rect 6552 12786 6604 12792
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6642 12608 6698 12617
rect 6564 11014 6592 12582
rect 6642 12543 6698 12552
rect 6656 12434 6684 12543
rect 6656 12406 6868 12434
rect 6736 12368 6788 12374
rect 6736 12310 6788 12316
rect 6748 12073 6776 12310
rect 6734 12064 6790 12073
rect 6734 11999 6790 12008
rect 6840 11830 6868 12406
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6550 10840 6606 10849
rect 6550 10775 6606 10784
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6564 9353 6592 10775
rect 6748 10606 6776 11562
rect 6840 10810 6868 11630
rect 6920 11552 6972 11558
rect 6920 11494 6972 11500
rect 6932 10810 6960 11494
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6920 10532 6972 10538
rect 6920 10474 6972 10480
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6734 10296 6790 10305
rect 6734 10231 6790 10240
rect 6748 10130 6776 10231
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6642 9616 6698 9625
rect 6840 9602 6868 10406
rect 6932 9722 6960 10474
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6840 9574 6960 9602
rect 6642 9551 6698 9560
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 6656 9217 6684 9551
rect 6828 9512 6880 9518
rect 6826 9480 6828 9489
rect 6880 9480 6882 9489
rect 6826 9415 6882 9424
rect 6642 9208 6698 9217
rect 6368 9172 6420 9178
rect 6642 9143 6698 9152
rect 6368 9114 6420 9120
rect 6460 8832 6512 8838
rect 6460 8774 6512 8780
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6380 7002 6408 8366
rect 6368 6996 6420 7002
rect 6368 6938 6420 6944
rect 6472 6662 6500 8774
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6564 7546 6592 8434
rect 6642 8392 6698 8401
rect 6642 8327 6698 8336
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6460 6248 6512 6254
rect 6460 6190 6512 6196
rect 6472 6118 6500 6190
rect 6368 6112 6420 6118
rect 6366 6080 6368 6089
rect 6460 6112 6512 6118
rect 6420 6080 6422 6089
rect 6460 6054 6512 6060
rect 6366 6015 6422 6024
rect 6012 5086 6224 5114
rect 6274 5128 6330 5137
rect 5908 4548 5960 4554
rect 5908 4490 5960 4496
rect 5814 3632 5870 3641
rect 5814 3567 5870 3576
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 2514 5856 3334
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5828 2417 5856 2450
rect 5814 2408 5870 2417
rect 5814 2343 5870 2352
rect 5632 1284 5684 1290
rect 5632 1226 5684 1232
rect 5446 776 5502 785
rect 5446 711 5502 720
rect 5920 202 5948 4490
rect 6012 4486 6040 5086
rect 6274 5063 6330 5072
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6184 5024 6236 5030
rect 6184 4966 6236 4972
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5998 3904 6054 3913
rect 5998 3839 6054 3848
rect 6012 3534 6040 3839
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6104 1329 6132 4490
rect 6196 4282 6224 4966
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4276 6236 4282
rect 6184 4218 6236 4224
rect 6288 2774 6316 4558
rect 6196 2746 6316 2774
rect 6196 2514 6224 2746
rect 6184 2508 6236 2514
rect 6184 2450 6236 2456
rect 6090 1320 6146 1329
rect 6090 1255 6146 1264
rect 6380 746 6408 5034
rect 6472 4865 6500 6054
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5545 6592 5578
rect 6550 5536 6606 5545
rect 6550 5471 6606 5480
rect 6458 4856 6514 4865
rect 6458 4791 6514 4800
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6564 4049 6592 4082
rect 6550 4040 6606 4049
rect 6550 3975 6606 3984
rect 6656 814 6684 8327
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7886 6868 8230
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6826 7712 6882 7721
rect 6826 7647 6882 7656
rect 6736 7200 6788 7206
rect 6734 7168 6736 7177
rect 6788 7168 6790 7177
rect 6734 7103 6790 7112
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6748 6186 6776 6695
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6840 4622 6868 7647
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6932 3534 6960 9574
rect 7024 8634 7052 13194
rect 7116 11286 7144 14719
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7208 13870 7236 14486
rect 7300 14385 7328 14758
rect 7286 14376 7342 14385
rect 7286 14311 7342 14320
rect 7392 14260 7420 14912
rect 7300 14249 7420 14260
rect 7286 14240 7420 14249
rect 7342 14232 7420 14240
rect 7286 14175 7342 14184
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 7194 13288 7250 13297
rect 7194 13223 7250 13232
rect 7208 12850 7236 13223
rect 7300 13025 7328 14175
rect 7484 13841 7512 17070
rect 7576 15978 7604 18566
rect 7668 17338 7696 18566
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7654 16688 7710 16697
rect 7654 16623 7710 16632
rect 7668 16046 7696 16623
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7564 15972 7616 15978
rect 7564 15914 7616 15920
rect 7668 15745 7696 15982
rect 7760 15978 7788 19654
rect 7852 19310 7880 20742
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 8116 20256 8168 20262
rect 8116 20198 8168 20204
rect 8128 19990 8156 20198
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 7840 19304 7892 19310
rect 7840 19246 7892 19252
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7852 18630 7880 18906
rect 7932 18896 7984 18902
rect 7932 18838 7984 18844
rect 7944 18698 7972 18838
rect 8312 18834 8340 25638
rect 8392 24880 8444 24886
rect 8392 24822 8444 24828
rect 8404 22438 8432 24822
rect 8482 23488 8538 23497
rect 8482 23423 8538 23432
rect 8496 22522 8524 23423
rect 8588 22710 8616 26302
rect 8666 26200 8722 26302
rect 9310 26200 9366 27000
rect 9496 26648 9548 26654
rect 9496 26590 9548 26596
rect 8944 25968 8996 25974
rect 8944 25910 8996 25916
rect 8576 22704 8628 22710
rect 8576 22646 8628 22652
rect 8668 22568 8720 22574
rect 8496 22494 8616 22522
rect 8668 22510 8720 22516
rect 8392 22432 8444 22438
rect 8392 22374 8444 22380
rect 8404 22094 8432 22374
rect 8404 22066 8524 22094
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8404 21486 8432 21898
rect 8392 21480 8444 21486
rect 8392 21422 8444 21428
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 8404 19961 8432 20198
rect 8390 19952 8446 19961
rect 8390 19887 8446 19896
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 8022 18728 8078 18737
rect 7932 18692 7984 18698
rect 8022 18663 8024 18672
rect 7932 18634 7984 18640
rect 8076 18663 8078 18672
rect 8024 18634 8076 18640
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7852 17921 7880 18566
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 7932 18352 7984 18358
rect 7932 18294 7984 18300
rect 7944 18154 7972 18294
rect 8208 18216 8260 18222
rect 8114 18184 8170 18193
rect 7932 18148 7984 18154
rect 8208 18158 8260 18164
rect 8114 18119 8170 18128
rect 7932 18090 7984 18096
rect 8128 18086 8156 18119
rect 8116 18080 8168 18086
rect 8116 18022 8168 18028
rect 7838 17912 7894 17921
rect 7838 17847 7894 17856
rect 8220 17785 8248 18158
rect 8298 17912 8354 17921
rect 8298 17847 8354 17856
rect 8206 17776 8262 17785
rect 8206 17711 8262 17720
rect 7840 17536 7892 17542
rect 7840 17478 7892 17484
rect 7852 16697 7880 17478
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8036 16833 8064 17274
rect 8208 17128 8260 17134
rect 8206 17096 8208 17105
rect 8260 17096 8262 17105
rect 8206 17031 8262 17040
rect 8022 16824 8078 16833
rect 8022 16759 8078 16768
rect 8116 16720 8168 16726
rect 7838 16688 7894 16697
rect 8116 16662 8168 16668
rect 7838 16623 7894 16632
rect 8128 16561 8156 16662
rect 8312 16561 8340 17847
rect 8114 16552 8170 16561
rect 8114 16487 8170 16496
rect 8298 16552 8354 16561
rect 8298 16487 8354 16496
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 7748 15972 7800 15978
rect 7748 15914 7800 15920
rect 7654 15736 7710 15745
rect 7654 15671 7710 15680
rect 7654 15600 7710 15609
rect 7576 15544 7654 15552
rect 7576 15524 7656 15544
rect 7576 14278 7604 15524
rect 7708 15535 7710 15544
rect 7656 15506 7708 15512
rect 7654 15192 7710 15201
rect 7654 15127 7656 15136
rect 7708 15127 7710 15136
rect 7656 15098 7708 15104
rect 7656 15020 7708 15026
rect 7656 14962 7708 14968
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7562 14104 7618 14113
rect 7562 14039 7618 14048
rect 7576 13938 7604 14039
rect 7668 13977 7696 14962
rect 7760 14074 7788 15914
rect 7852 14618 7880 16390
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 8312 16130 8340 16390
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8220 16102 8340 16130
rect 7944 15609 7972 16050
rect 7930 15600 7986 15609
rect 7930 15535 7986 15544
rect 7930 15464 7986 15473
rect 7930 15399 7932 15408
rect 7984 15399 7986 15408
rect 7932 15370 7984 15376
rect 8220 15348 8248 16102
rect 8220 15320 8340 15348
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7944 14498 7972 15098
rect 8036 14929 8064 15098
rect 8312 15042 8340 15320
rect 8220 15014 8340 15042
rect 8022 14920 8078 14929
rect 8022 14855 8024 14864
rect 8076 14855 8078 14864
rect 8024 14826 8076 14832
rect 7852 14470 7972 14498
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7654 13968 7710 13977
rect 7564 13932 7616 13938
rect 7654 13903 7710 13912
rect 7564 13874 7616 13880
rect 7656 13864 7708 13870
rect 7470 13832 7526 13841
rect 7656 13806 7708 13812
rect 7470 13767 7526 13776
rect 7668 13716 7696 13806
rect 7576 13688 7696 13716
rect 7852 13705 7880 14470
rect 7930 14376 7986 14385
rect 7930 14311 7932 14320
rect 7984 14311 7986 14320
rect 7932 14282 7984 14288
rect 8220 14260 8248 15014
rect 8220 14232 8340 14260
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 7838 13696 7894 13705
rect 7378 13560 7434 13569
rect 7378 13495 7434 13504
rect 7392 13161 7420 13495
rect 7378 13152 7434 13161
rect 7378 13087 7434 13096
rect 7286 13016 7342 13025
rect 7286 12951 7342 12960
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7288 12368 7340 12374
rect 7288 12310 7340 12316
rect 7104 11280 7156 11286
rect 7104 11222 7156 11228
rect 7196 11212 7248 11218
rect 7196 11154 7248 11160
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 7116 10985 7144 11018
rect 7102 10976 7158 10985
rect 7102 10911 7158 10920
rect 7208 10606 7236 11154
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7116 9625 7144 10542
rect 7102 9616 7158 9625
rect 7102 9551 7158 9560
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7012 8356 7064 8362
rect 7012 8298 7064 8304
rect 7024 4622 7052 8298
rect 7116 7342 7144 9386
rect 7208 9042 7236 10542
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7208 8090 7236 8842
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7300 7721 7328 12310
rect 7472 12232 7524 12238
rect 7470 12200 7472 12209
rect 7524 12200 7526 12209
rect 7470 12135 7526 12144
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7392 11150 7420 11290
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7380 9920 7432 9926
rect 7378 9888 7380 9897
rect 7432 9888 7434 9897
rect 7378 9823 7434 9832
rect 7380 9580 7432 9586
rect 7380 9522 7432 9528
rect 7392 7857 7420 9522
rect 7484 8430 7512 11766
rect 7576 11354 7604 13688
rect 7838 13631 7894 13640
rect 7656 13252 7708 13258
rect 7656 13194 7708 13200
rect 7668 12918 7696 13194
rect 7748 13184 7800 13190
rect 8036 13172 8064 14010
rect 8312 13954 8340 14232
rect 8404 14074 8432 18770
rect 8496 14414 8524 22066
rect 8588 20262 8616 22494
rect 8680 21350 8708 22510
rect 8760 21888 8812 21894
rect 8758 21856 8760 21865
rect 8812 21856 8814 21865
rect 8758 21791 8814 21800
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8680 20398 8708 21286
rect 8668 20392 8720 20398
rect 8668 20334 8720 20340
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8588 18193 8616 19994
rect 8680 19922 8708 20334
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8680 19786 8708 19858
rect 8668 19780 8720 19786
rect 8668 19722 8720 19728
rect 8956 19334 8984 25910
rect 9220 25492 9272 25498
rect 9220 25434 9272 25440
rect 9128 24064 9180 24070
rect 9128 24006 9180 24012
rect 9140 23798 9168 24006
rect 9128 23792 9180 23798
rect 9128 23734 9180 23740
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22273 9076 22918
rect 9034 22264 9090 22273
rect 9034 22199 9090 22208
rect 9034 21992 9090 22001
rect 9034 21927 9036 21936
rect 9088 21927 9090 21936
rect 9036 21898 9088 21904
rect 9034 20632 9090 20641
rect 9034 20567 9090 20576
rect 9048 20058 9076 20567
rect 9036 20052 9088 20058
rect 9036 19994 9088 20000
rect 9232 19854 9260 25434
rect 9324 24342 9352 26200
rect 9312 24336 9364 24342
rect 9312 24278 9364 24284
rect 9508 23118 9536 26590
rect 9954 26200 10010 27000
rect 10232 26920 10284 26926
rect 10232 26862 10284 26868
rect 9862 25256 9918 25265
rect 9862 25191 9918 25200
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9678 23760 9734 23769
rect 9678 23695 9734 23704
rect 9692 23526 9720 23695
rect 9680 23520 9732 23526
rect 9784 23497 9812 24142
rect 9876 23730 9904 25191
rect 9864 23724 9916 23730
rect 9864 23666 9916 23672
rect 9968 23662 9996 26200
rect 10048 25084 10100 25090
rect 10048 25026 10100 25032
rect 9956 23656 10008 23662
rect 9956 23598 10008 23604
rect 9680 23462 9732 23468
rect 9770 23488 9826 23497
rect 9770 23423 9826 23432
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9404 22976 9456 22982
rect 9404 22918 9456 22924
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9324 21729 9352 21830
rect 9310 21720 9366 21729
rect 9310 21655 9366 21664
rect 9416 21622 9444 22918
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9770 22128 9826 22137
rect 9770 22063 9826 22072
rect 9680 21888 9732 21894
rect 9680 21830 9732 21836
rect 9404 21616 9456 21622
rect 9404 21558 9456 21564
rect 9416 21010 9444 21558
rect 9586 21448 9642 21457
rect 9586 21383 9588 21392
rect 9640 21383 9642 21392
rect 9588 21354 9640 21360
rect 9404 21004 9456 21010
rect 9404 20946 9456 20952
rect 9692 20777 9720 21830
rect 9678 20768 9734 20777
rect 9678 20703 9734 20712
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9140 19514 9168 19654
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 8680 19306 8984 19334
rect 8574 18184 8630 18193
rect 8574 18119 8630 18128
rect 8680 18086 8708 19306
rect 9128 19304 9180 19310
rect 9128 19246 9180 19252
rect 8944 19168 8996 19174
rect 8942 19136 8944 19145
rect 8996 19136 8998 19145
rect 8942 19071 8998 19080
rect 9140 18986 9168 19246
rect 8944 18964 8996 18970
rect 8944 18906 8996 18912
rect 9048 18958 9168 18986
rect 8760 18624 8812 18630
rect 8760 18566 8812 18572
rect 8852 18624 8904 18630
rect 8852 18566 8904 18572
rect 8772 18086 8800 18566
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8668 18080 8720 18086
rect 8668 18022 8720 18028
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8588 17338 8616 18022
rect 8576 17332 8628 17338
rect 8576 17274 8628 17280
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8588 16833 8616 17138
rect 8574 16824 8630 16833
rect 8574 16759 8630 16768
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8588 16425 8616 16662
rect 8680 16436 8708 18022
rect 8772 16658 8800 18022
rect 8864 17610 8892 18566
rect 8956 18290 8984 18906
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 8956 17610 8984 18226
rect 8852 17604 8904 17610
rect 8852 17546 8904 17552
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8850 17232 8906 17241
rect 8850 17167 8906 17176
rect 8760 16652 8812 16658
rect 8760 16594 8812 16600
rect 8760 16448 8812 16454
rect 8574 16416 8630 16425
rect 8680 16408 8760 16436
rect 8760 16390 8812 16396
rect 8574 16351 8630 16360
rect 8666 16280 8722 16289
rect 8666 16215 8668 16224
rect 8720 16215 8722 16224
rect 8668 16186 8720 16192
rect 8772 16017 8800 16390
rect 8758 16008 8814 16017
rect 8758 15943 8814 15952
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8574 15192 8630 15201
rect 8772 15162 8800 15846
rect 8574 15127 8630 15136
rect 8760 15156 8812 15162
rect 8588 14958 8616 15127
rect 8760 15098 8812 15104
rect 8576 14952 8628 14958
rect 8576 14894 8628 14900
rect 8760 14816 8812 14822
rect 8760 14758 8812 14764
rect 8668 14544 8720 14550
rect 8668 14486 8720 14492
rect 8484 14408 8536 14414
rect 8482 14376 8484 14385
rect 8536 14376 8538 14385
rect 8482 14311 8538 14320
rect 8482 14104 8538 14113
rect 8392 14068 8444 14074
rect 8482 14039 8538 14048
rect 8392 14010 8444 14016
rect 8220 13926 8340 13954
rect 8392 13932 8444 13938
rect 8220 13433 8248 13926
rect 8496 13920 8524 14039
rect 8444 13892 8524 13920
rect 8576 13932 8628 13938
rect 8392 13874 8444 13880
rect 8576 13874 8628 13880
rect 8206 13424 8262 13433
rect 8206 13359 8262 13368
rect 7748 13126 7800 13132
rect 7852 13144 8064 13172
rect 8220 13172 8248 13359
rect 8220 13144 8340 13172
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7564 11348 7616 11354
rect 7564 11290 7616 11296
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10062 7604 10950
rect 7668 10606 7696 12718
rect 7760 11218 7788 13126
rect 7852 12374 7880 13144
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 8024 12912 8076 12918
rect 8312 12866 8340 13144
rect 8024 12854 8076 12860
rect 7840 12368 7892 12374
rect 7840 12310 7892 12316
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11642 7880 12174
rect 8036 12102 8064 12854
rect 8220 12838 8340 12866
rect 8220 12617 8248 12838
rect 8206 12608 8262 12617
rect 8588 12594 8616 13874
rect 8206 12543 8262 12552
rect 8496 12566 8616 12594
rect 8496 12424 8524 12566
rect 8404 12396 8524 12424
rect 8576 12436 8628 12442
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 8404 11914 8432 12396
rect 8576 12378 8628 12384
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8312 11886 8432 11914
rect 7852 11614 7972 11642
rect 7840 11552 7892 11558
rect 7840 11494 7892 11500
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7852 11150 7880 11494
rect 7840 11144 7892 11150
rect 7944 11121 7972 11614
rect 7840 11086 7892 11092
rect 7930 11112 7986 11121
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7656 10600 7708 10606
rect 7656 10542 7708 10548
rect 7564 10056 7616 10062
rect 7760 10010 7788 10950
rect 7564 9998 7616 10004
rect 7668 9982 7788 10010
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9489 7604 9522
rect 7562 9480 7618 9489
rect 7562 9415 7618 9424
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7576 8566 7604 9114
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7378 7848 7434 7857
rect 7378 7783 7434 7792
rect 7564 7744 7616 7750
rect 7286 7712 7342 7721
rect 7564 7686 7616 7692
rect 7286 7647 7342 7656
rect 7104 7336 7156 7342
rect 7104 7278 7156 7284
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7208 5370 7236 6870
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7300 4826 7328 6938
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 5914 7420 6802
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7484 4826 7512 5646
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7208 4146 7236 4626
rect 7576 4554 7604 7686
rect 7564 4548 7616 4554
rect 7564 4490 7616 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7484 4214 7512 4422
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7668 4078 7696 9982
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 8362 7788 9862
rect 7748 8356 7800 8362
rect 7748 8298 7800 8304
rect 7852 7410 7880 11086
rect 7930 11047 7986 11056
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 8312 10792 8340 11886
rect 8496 11830 8524 12038
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8588 11626 8616 12378
rect 8576 11620 8628 11626
rect 8576 11562 8628 11568
rect 8574 11384 8630 11393
rect 8574 11319 8630 11328
rect 8588 11218 8616 11319
rect 8576 11212 8628 11218
rect 8576 11154 8628 11160
rect 8484 11144 8536 11150
rect 8220 10764 8340 10792
rect 8404 11104 8484 11132
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8036 10266 8064 10542
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 8128 9994 8156 10202
rect 8220 10130 8248 10764
rect 8298 10704 8354 10713
rect 8298 10639 8354 10648
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 9988 8168 9994
rect 8116 9930 8168 9936
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 8312 8090 8340 10639
rect 8404 10441 8432 11104
rect 8484 11086 8536 11092
rect 8574 10840 8630 10849
rect 8574 10775 8630 10784
rect 8484 10464 8536 10470
rect 8390 10432 8446 10441
rect 8484 10406 8536 10412
rect 8390 10367 8446 10376
rect 8496 10062 8524 10406
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 9217 8432 9930
rect 8496 9518 8524 9998
rect 8588 9926 8616 10775
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8680 9654 8708 14486
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8404 7478 8432 8774
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7944 7274 7972 7346
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7760 6633 7788 6802
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 7746 6624 7802 6633
rect 7746 6559 7802 6568
rect 7746 6488 7802 6497
rect 7746 6423 7802 6432
rect 7760 6390 7788 6423
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7852 5817 7880 6666
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7930 6352 7986 6361
rect 8312 6322 8340 7142
rect 8390 6488 8446 6497
rect 8390 6423 8446 6432
rect 7930 6287 7986 6296
rect 8300 6316 8352 6322
rect 7838 5808 7894 5817
rect 7838 5743 7894 5752
rect 7944 5710 7972 6287
rect 8300 6258 8352 6264
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7746 5400 7802 5409
rect 7950 5403 8258 5412
rect 7746 5335 7748 5344
rect 7800 5335 7802 5344
rect 7748 5306 7800 5312
rect 8312 5234 8340 5510
rect 8404 5302 8432 6423
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8220 4826 8248 5170
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 8300 3460 8352 3466
rect 8300 3402 8352 3408
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 8312 2650 8340 3402
rect 8496 3058 8524 9454
rect 8772 8922 8800 14758
rect 8864 10441 8892 17167
rect 9048 16522 9076 18958
rect 9128 18760 9180 18766
rect 9128 18702 9180 18708
rect 9220 18760 9272 18766
rect 9220 18702 9272 18708
rect 9140 17746 9168 18702
rect 9232 18057 9260 18702
rect 9218 18048 9274 18057
rect 9218 17983 9274 17992
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 9232 17610 9260 17983
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9220 17604 9272 17610
rect 9220 17546 9272 17552
rect 9036 16516 9088 16522
rect 9036 16458 9088 16464
rect 9036 16244 9088 16250
rect 9036 16186 9088 16192
rect 9048 15745 9076 16186
rect 9034 15736 9090 15745
rect 9034 15671 9090 15680
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15094 8984 15302
rect 8944 15088 8996 15094
rect 8944 15030 8996 15036
rect 9048 14822 9076 15370
rect 9036 14816 9088 14822
rect 9036 14758 9088 14764
rect 8944 14408 8996 14414
rect 8944 14350 8996 14356
rect 9034 14376 9090 14385
rect 8956 13977 8984 14350
rect 9034 14311 9090 14320
rect 8942 13968 8998 13977
rect 8942 13903 8998 13912
rect 8942 13424 8998 13433
rect 8942 13359 8998 13368
rect 8956 12782 8984 13359
rect 8944 12776 8996 12782
rect 8944 12718 8996 12724
rect 8956 11150 8984 12718
rect 9048 12442 9076 14311
rect 9036 12436 9088 12442
rect 9036 12378 9088 12384
rect 9036 12096 9088 12102
rect 9036 12038 9088 12044
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8850 10432 8906 10441
rect 8850 10367 8906 10376
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9926 8892 10066
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 8864 9654 8892 9862
rect 8852 9648 8904 9654
rect 8850 9616 8852 9625
rect 8904 9616 8906 9625
rect 8850 9551 8906 9560
rect 8680 8894 8800 8922
rect 8576 8424 8628 8430
rect 8576 8366 8628 8372
rect 8588 6866 8616 8366
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8680 3738 8708 8894
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8850 8800 8906 8809
rect 8772 8498 8800 8774
rect 8850 8735 8906 8744
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8772 4026 8800 8026
rect 8864 6225 8892 8735
rect 8956 7206 8984 11086
rect 9048 10742 9076 12038
rect 9140 11762 9168 17546
rect 9324 17241 9352 20198
rect 9404 20052 9456 20058
rect 9404 19994 9456 20000
rect 9416 18698 9444 19994
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9496 19508 9548 19514
rect 9496 19450 9548 19456
rect 9508 19417 9536 19450
rect 9494 19408 9550 19417
rect 9494 19343 9550 19352
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9508 18601 9536 19110
rect 9494 18592 9550 18601
rect 9494 18527 9550 18536
rect 9600 18358 9628 19790
rect 9692 19281 9720 20198
rect 9678 19272 9734 19281
rect 9678 19207 9734 19216
rect 9588 18352 9640 18358
rect 9588 18294 9640 18300
rect 9404 18284 9456 18290
rect 9404 18226 9456 18232
rect 9416 17785 9444 18226
rect 9784 18057 9812 22063
rect 9968 21078 9996 22374
rect 9956 21072 10008 21078
rect 9956 21014 10008 21020
rect 9968 20618 9996 21014
rect 10060 21010 10088 25026
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10152 20806 10180 24074
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 9968 20590 10180 20618
rect 9956 20324 10008 20330
rect 9956 20266 10008 20272
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 9876 18465 9904 19246
rect 9968 18902 9996 20266
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9862 18456 9918 18465
rect 9862 18391 9918 18400
rect 9770 18048 9826 18057
rect 9770 17983 9826 17992
rect 9402 17776 9458 17785
rect 9402 17711 9458 17720
rect 9496 17740 9548 17746
rect 9496 17682 9548 17688
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 9508 17134 9536 17682
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9324 16726 9352 17070
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9312 16720 9364 16726
rect 9218 16688 9274 16697
rect 9312 16662 9364 16668
rect 9218 16623 9274 16632
rect 9232 16250 9260 16623
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9232 15910 9260 16186
rect 9324 16028 9352 16662
rect 9416 16289 9444 16730
rect 9586 16688 9642 16697
rect 9876 16674 9904 17274
rect 9968 16998 9996 17614
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9954 16688 10010 16697
rect 9876 16646 9954 16674
rect 9586 16623 9642 16632
rect 9954 16623 9956 16632
rect 9600 16590 9628 16623
rect 10008 16623 10010 16632
rect 9956 16594 10008 16600
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9588 16584 9640 16590
rect 9588 16526 9640 16532
rect 9402 16280 9458 16289
rect 9508 16250 9536 16526
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9402 16215 9458 16224
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9588 16040 9640 16046
rect 9324 16000 9588 16028
rect 9220 15904 9272 15910
rect 9220 15846 9272 15852
rect 9324 15502 9352 16000
rect 9588 15982 9640 15988
rect 9692 15978 9720 16390
rect 9680 15972 9732 15978
rect 9680 15914 9732 15920
rect 9496 15632 9548 15638
rect 9864 15632 9916 15638
rect 9496 15574 9548 15580
rect 9692 15592 9864 15620
rect 9404 15564 9456 15570
rect 9404 15506 9456 15512
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9416 15201 9444 15506
rect 9402 15192 9458 15201
rect 9402 15127 9458 15136
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 13394 9260 14962
rect 9404 14612 9456 14618
rect 9404 14554 9456 14560
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9232 12646 9260 13330
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9324 11830 9352 13806
rect 9416 13190 9444 14554
rect 9508 13433 9536 15574
rect 9692 15450 9720 15592
rect 9864 15574 9916 15580
rect 9600 15422 9720 15450
rect 9600 15366 9628 15422
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9600 14958 9628 15302
rect 9588 14952 9640 14958
rect 9588 14894 9640 14900
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9494 13424 9550 13433
rect 9494 13359 9550 13368
rect 9496 13320 9548 13326
rect 9496 13262 9548 13268
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9404 12912 9456 12918
rect 9404 12854 9456 12860
rect 9416 12238 9444 12854
rect 9508 12442 9536 13262
rect 9600 13025 9628 14350
rect 9692 14074 9720 15302
rect 9862 15192 9918 15201
rect 9862 15127 9918 15136
rect 9876 15026 9904 15127
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9680 14068 9732 14074
rect 9680 14010 9732 14016
rect 9678 13968 9734 13977
rect 9678 13903 9734 13912
rect 9586 13016 9642 13025
rect 9586 12951 9642 12960
rect 9692 12918 9720 13903
rect 9784 13433 9812 14758
rect 9770 13424 9826 13433
rect 9770 13359 9826 13368
rect 9770 13152 9826 13161
rect 9770 13087 9826 13096
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9496 12436 9548 12442
rect 9496 12378 9548 12384
rect 9600 12345 9628 12650
rect 9784 12458 9812 13087
rect 9876 12782 9904 14758
rect 9968 14385 9996 16594
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9954 14376 10010 14385
rect 9954 14311 10010 14320
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9968 12646 9996 13398
rect 10060 13326 10088 15846
rect 10152 13870 10180 20590
rect 10244 17338 10272 26862
rect 10598 26330 10654 27000
rect 10520 26302 10654 26330
rect 10520 23186 10548 26302
rect 10598 26200 10654 26302
rect 11242 26200 11298 27000
rect 11886 26200 11942 27000
rect 12530 26200 12586 27000
rect 13174 26200 13230 27000
rect 13280 26302 13492 26330
rect 11060 24880 11112 24886
rect 11058 24848 11060 24857
rect 11112 24848 11114 24857
rect 11058 24783 11114 24792
rect 10874 24032 10930 24041
rect 10874 23967 10930 23976
rect 10598 23896 10654 23905
rect 10598 23831 10654 23840
rect 10508 23180 10560 23186
rect 10508 23122 10560 23128
rect 10506 22128 10562 22137
rect 10416 22092 10468 22098
rect 10506 22063 10562 22072
rect 10416 22034 10468 22040
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10336 21554 10364 21898
rect 10324 21548 10376 21554
rect 10324 21490 10376 21496
rect 10428 20262 10456 22034
rect 10520 21486 10548 22063
rect 10508 21480 10560 21486
rect 10508 21422 10560 21428
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10520 20874 10548 21014
rect 10508 20868 10560 20874
rect 10508 20810 10560 20816
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10416 20256 10468 20262
rect 10416 20198 10468 20204
rect 10322 19816 10378 19825
rect 10322 19751 10324 19760
rect 10376 19751 10378 19760
rect 10324 19722 10376 19728
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10336 18630 10364 19314
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10336 17134 10364 18566
rect 10520 17513 10548 20402
rect 10612 19514 10640 23831
rect 10690 23624 10746 23633
rect 10690 23559 10746 23568
rect 10704 22030 10732 23559
rect 10784 22976 10836 22982
rect 10784 22918 10836 22924
rect 10796 22710 10824 22918
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10888 22094 10916 23967
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 10796 22066 10916 22094
rect 10692 22024 10744 22030
rect 10692 21966 10744 21972
rect 10796 20618 10824 22066
rect 10968 21480 11020 21486
rect 10968 21422 11020 21428
rect 10704 20602 10824 20618
rect 10692 20596 10824 20602
rect 10744 20590 10824 20596
rect 10692 20538 10744 20544
rect 10704 19514 10732 20538
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 10980 20482 11008 21422
rect 11072 20602 11100 22986
rect 11164 22642 11192 23054
rect 11152 22636 11204 22642
rect 11152 22578 11204 22584
rect 11256 22098 11284 26200
rect 11428 24404 11480 24410
rect 11428 24346 11480 24352
rect 11440 24154 11468 24346
rect 11532 24274 11652 24290
rect 11520 24268 11652 24274
rect 11572 24262 11652 24268
rect 11520 24210 11572 24216
rect 11440 24126 11560 24154
rect 11428 23044 11480 23050
rect 11428 22986 11480 22992
rect 11440 22681 11468 22986
rect 11426 22672 11482 22681
rect 11426 22607 11482 22616
rect 11336 22432 11388 22438
rect 11336 22374 11388 22380
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11244 22092 11296 22098
rect 11244 22034 11296 22040
rect 11152 21888 11204 21894
rect 11152 21830 11204 21836
rect 11060 20596 11112 20602
rect 11060 20538 11112 20544
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10796 19786 10824 20334
rect 10784 19780 10836 19786
rect 10784 19722 10836 19728
rect 10600 19508 10652 19514
rect 10600 19450 10652 19456
rect 10692 19508 10744 19514
rect 10692 19450 10744 19456
rect 10784 19304 10836 19310
rect 10782 19272 10784 19281
rect 10836 19272 10838 19281
rect 10782 19207 10838 19216
rect 10796 19009 10824 19207
rect 10782 19000 10838 19009
rect 10782 18935 10838 18944
rect 10598 18728 10654 18737
rect 10598 18663 10600 18672
rect 10652 18663 10654 18672
rect 10600 18634 10652 18640
rect 10888 18426 10916 20470
rect 10980 20454 11100 20482
rect 11072 20398 11100 20454
rect 11060 20392 11112 20398
rect 11060 20334 11112 20340
rect 11164 18850 11192 21830
rect 11348 21729 11376 22374
rect 11334 21720 11390 21729
rect 11334 21655 11390 21664
rect 11244 20800 11296 20806
rect 11336 20800 11388 20806
rect 11244 20742 11296 20748
rect 11334 20768 11336 20777
rect 11388 20768 11390 20777
rect 11072 18822 11192 18850
rect 11072 18630 11100 18822
rect 11152 18692 11204 18698
rect 11152 18634 11204 18640
rect 11060 18624 11112 18630
rect 11060 18566 11112 18572
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10690 18320 10746 18329
rect 10690 18255 10692 18264
rect 10744 18255 10746 18264
rect 10692 18226 10744 18232
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10612 17746 10640 18158
rect 10600 17740 10652 17746
rect 10600 17682 10652 17688
rect 10600 17536 10652 17542
rect 10506 17504 10562 17513
rect 10600 17478 10652 17484
rect 10506 17439 10562 17448
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10324 16992 10376 16998
rect 10322 16960 10324 16969
rect 10416 16992 10468 16998
rect 10376 16960 10378 16969
rect 10416 16934 10468 16940
rect 10322 16895 10378 16904
rect 10336 16658 10364 16895
rect 10324 16652 10376 16658
rect 10324 16594 10376 16600
rect 10336 16017 10364 16594
rect 10322 16008 10378 16017
rect 10322 15943 10378 15952
rect 10230 15736 10286 15745
rect 10230 15671 10286 15680
rect 10244 14618 10272 15671
rect 10428 15094 10456 16934
rect 10520 16454 10548 17439
rect 10612 17270 10640 17478
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10508 16448 10560 16454
rect 10508 16390 10560 16396
rect 10612 16182 10640 17070
rect 10784 17060 10836 17066
rect 10784 17002 10836 17008
rect 10690 16280 10746 16289
rect 10690 16215 10746 16224
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 10612 16046 10640 16118
rect 10600 16040 10652 16046
rect 10600 15982 10652 15988
rect 10506 15192 10562 15201
rect 10612 15162 10640 15982
rect 10704 15366 10732 16215
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10506 15127 10562 15136
rect 10600 15156 10652 15162
rect 10416 15088 10468 15094
rect 10416 15030 10468 15036
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10232 14612 10284 14618
rect 10232 14554 10284 14560
rect 10140 13864 10192 13870
rect 10140 13806 10192 13812
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10048 13320 10100 13326
rect 10048 13262 10100 13268
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 9956 12640 10008 12646
rect 9956 12582 10008 12588
rect 9784 12430 9996 12458
rect 9586 12336 9642 12345
rect 9968 12306 9996 12430
rect 9586 12271 9642 12280
rect 9956 12300 10008 12306
rect 9956 12242 10008 12248
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 10060 12170 10088 13126
rect 10152 12850 10180 13670
rect 10244 12918 10272 14554
rect 10428 13190 10456 14894
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10048 12164 10100 12170
rect 10152 12152 10180 12582
rect 10152 12124 10272 12152
rect 10048 12106 10100 12112
rect 9404 12096 9456 12102
rect 9404 12038 9456 12044
rect 9772 12096 9824 12102
rect 9824 12073 9904 12084
rect 9824 12064 9918 12073
rect 9824 12056 9862 12064
rect 9772 12038 9824 12044
rect 9312 11824 9364 11830
rect 9312 11766 9364 11772
rect 9128 11756 9180 11762
rect 9128 11698 9180 11704
rect 9128 11620 9180 11626
rect 9128 11562 9180 11568
rect 9036 10736 9088 10742
rect 9036 10678 9088 10684
rect 9048 10130 9076 10678
rect 9140 10538 9168 11562
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 9034 10024 9090 10033
rect 9034 9959 9090 9968
rect 9048 8537 9076 9959
rect 9140 8809 9168 10474
rect 9232 9518 9260 11086
rect 9220 9512 9272 9518
rect 9220 9454 9272 9460
rect 9126 8800 9182 8809
rect 9126 8735 9182 8744
rect 9034 8528 9090 8537
rect 9034 8463 9090 8472
rect 9220 8492 9272 8498
rect 9220 8434 9272 8440
rect 9126 8256 9182 8265
rect 9126 8191 9182 8200
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9036 6792 9088 6798
rect 9034 6760 9036 6769
rect 9088 6760 9090 6769
rect 9034 6695 9090 6704
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6390 9076 6598
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 8944 6248 8996 6254
rect 8850 6216 8906 6225
rect 8944 6190 8996 6196
rect 9034 6216 9090 6225
rect 8850 6151 8906 6160
rect 8864 4146 8892 6151
rect 8956 5370 8984 6190
rect 9034 6151 9090 6160
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9048 4593 9076 6151
rect 9140 5302 9168 8191
rect 9232 7002 9260 8434
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9324 5778 9352 11222
rect 9416 11082 9444 12038
rect 9862 11999 9918 12008
rect 9588 11892 9640 11898
rect 9588 11834 9640 11840
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9404 10668 9456 10674
rect 9404 10610 9456 10616
rect 9416 10033 9444 10610
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9508 9722 9536 10950
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9416 8974 9444 9658
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9496 8424 9548 8430
rect 9496 8366 9548 8372
rect 9404 8288 9456 8294
rect 9404 8230 9456 8236
rect 9416 7274 9444 8230
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9508 5624 9536 8366
rect 9600 7954 9628 11834
rect 9680 11756 9732 11762
rect 9680 11698 9732 11704
rect 9692 10742 9720 11698
rect 10244 11370 10272 12124
rect 9968 11342 10272 11370
rect 9968 11218 9996 11342
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 10048 11144 10100 11150
rect 10048 11086 10100 11092
rect 10060 10985 10088 11086
rect 9862 10976 9918 10985
rect 9862 10911 9918 10920
rect 10046 10976 10102 10985
rect 10046 10911 10102 10920
rect 9680 10736 9732 10742
rect 9680 10678 9732 10684
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10033 9812 10406
rect 9770 10024 9826 10033
rect 9770 9959 9826 9968
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9692 9674 9720 9862
rect 9692 9646 9812 9674
rect 9784 9382 9812 9646
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9772 9104 9824 9110
rect 9772 9046 9824 9052
rect 9678 8664 9734 8673
rect 9678 8599 9734 8608
rect 9692 8294 9720 8599
rect 9680 8288 9732 8294
rect 9680 8230 9732 8236
rect 9692 8090 9720 8230
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9588 7948 9640 7954
rect 9588 7890 9640 7896
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9692 6361 9720 6666
rect 9678 6352 9734 6361
rect 9678 6287 9734 6296
rect 9784 5710 9812 9046
rect 9876 8673 9904 10911
rect 10232 10736 10284 10742
rect 10232 10678 10284 10684
rect 9954 10296 10010 10305
rect 9954 10231 10010 10240
rect 9862 8664 9918 8673
rect 9862 8599 9918 8608
rect 9862 8528 9918 8537
rect 9862 8463 9918 8472
rect 9876 8090 9904 8463
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9508 5596 9720 5624
rect 9128 5296 9180 5302
rect 9128 5238 9180 5244
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9034 4584 9090 4593
rect 9034 4519 9090 4528
rect 8852 4140 8904 4146
rect 8852 4082 8904 4088
rect 8772 3998 8892 4026
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8668 3732 8720 3738
rect 8668 3674 8720 3680
rect 8574 3496 8630 3505
rect 8574 3431 8576 3440
rect 8628 3431 8630 3440
rect 8576 3402 8628 3408
rect 8484 3052 8536 3058
rect 8484 2994 8536 3000
rect 8772 2961 8800 3878
rect 8758 2952 8814 2961
rect 8864 2922 8892 3998
rect 8758 2887 8814 2896
rect 8852 2916 8904 2922
rect 8852 2858 8904 2864
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6644 808 6696 814
rect 6748 800 6776 2450
rect 9048 2310 9076 4519
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 9048 2038 9076 2246
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 9140 921 9168 3878
rect 9232 3126 9260 5102
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9324 4622 9352 4966
rect 9402 4856 9458 4865
rect 9402 4791 9458 4800
rect 9416 4622 9444 4791
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9692 4536 9720 5596
rect 9692 4508 9812 4536
rect 9678 4448 9734 4457
rect 9678 4383 9734 4392
rect 9312 4072 9364 4078
rect 9310 4040 9312 4049
rect 9364 4040 9366 4049
rect 9310 3975 9366 3984
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9220 3120 9272 3126
rect 9220 3062 9272 3068
rect 9416 2774 9444 3538
rect 9508 3534 9536 3878
rect 9692 3738 9720 4383
rect 9680 3732 9732 3738
rect 9680 3674 9732 3680
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9692 3466 9720 3674
rect 9784 3602 9812 4508
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9876 2990 9904 6054
rect 9968 5778 9996 10231
rect 10244 9654 10272 10678
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10060 9178 10088 9318
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10152 8974 10180 9318
rect 10230 9208 10286 9217
rect 10230 9143 10286 9152
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 10060 8566 10088 8599
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 10048 8424 10100 8430
rect 10046 8392 10048 8401
rect 10100 8392 10102 8401
rect 10046 8327 10102 8336
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7886 10088 8026
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10046 7168 10102 7177
rect 10046 7103 10102 7112
rect 9956 5772 10008 5778
rect 9956 5714 10008 5720
rect 9954 5128 10010 5137
rect 9954 5063 10010 5072
rect 9968 4826 9996 5063
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9968 4010 9996 4150
rect 10060 4146 10088 7103
rect 10152 5234 10180 8910
rect 10244 8906 10272 9143
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10244 8498 10272 8842
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10232 8356 10284 8362
rect 10232 8298 10284 8304
rect 10244 7750 10272 8298
rect 10336 7886 10364 12582
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10428 10577 10456 12242
rect 10414 10568 10470 10577
rect 10414 10503 10470 10512
rect 10428 9761 10456 10503
rect 10414 9752 10470 9761
rect 10414 9687 10470 9696
rect 10414 9616 10470 9625
rect 10414 9551 10470 9560
rect 10428 8906 10456 9551
rect 10520 9110 10548 15127
rect 10600 15098 10652 15104
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 14822 10640 14894
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14346 10640 14758
rect 10690 14648 10746 14657
rect 10690 14583 10746 14592
rect 10704 14414 10732 14583
rect 10692 14408 10744 14414
rect 10692 14350 10744 14356
rect 10600 14340 10652 14346
rect 10600 14282 10652 14288
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10612 13394 10640 13670
rect 10600 13388 10652 13394
rect 10600 13330 10652 13336
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10612 12238 10640 12718
rect 10704 12646 10732 14214
rect 10796 13161 10824 17002
rect 10888 16658 10916 18158
rect 10980 17882 11008 18158
rect 10968 17876 11020 17882
rect 10968 17818 11020 17824
rect 10968 17332 11020 17338
rect 10968 17274 11020 17280
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10876 16516 10928 16522
rect 10876 16458 10928 16464
rect 10888 15994 10916 16458
rect 10980 16250 11008 17274
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11072 16794 11100 17138
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11058 16688 11114 16697
rect 11058 16623 11060 16632
rect 11112 16623 11114 16632
rect 11060 16594 11112 16600
rect 10968 16244 11020 16250
rect 10968 16186 11020 16192
rect 11060 16176 11112 16182
rect 11058 16144 11060 16153
rect 11112 16144 11114 16153
rect 11058 16079 11114 16088
rect 10888 15966 11100 15994
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10980 14793 11008 14962
rect 10966 14784 11022 14793
rect 10966 14719 11022 14728
rect 10968 14476 11020 14482
rect 10888 14436 10968 14464
rect 10888 14385 10916 14436
rect 10968 14418 11020 14424
rect 10874 14376 10930 14385
rect 10874 14311 10930 14320
rect 10888 13258 10916 14311
rect 11072 14113 11100 15966
rect 11164 15473 11192 18634
rect 11150 15464 11206 15473
rect 11150 15399 11206 15408
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 11164 14006 11192 15302
rect 11256 14929 11284 20742
rect 11334 20703 11390 20712
rect 11440 20398 11468 22374
rect 11532 20806 11560 24126
rect 11520 20800 11572 20806
rect 11520 20742 11572 20748
rect 11428 20392 11480 20398
rect 11428 20334 11480 20340
rect 11336 19712 11388 19718
rect 11336 19654 11388 19660
rect 11348 18630 11376 19654
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11334 18320 11390 18329
rect 11334 18255 11390 18264
rect 11348 17785 11376 18255
rect 11334 17776 11390 17785
rect 11334 17711 11390 17720
rect 11440 16810 11468 20334
rect 11624 19553 11652 24262
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11716 23497 11744 24006
rect 11808 23798 11836 24006
rect 11796 23792 11848 23798
rect 11796 23734 11848 23740
rect 11702 23488 11758 23497
rect 11702 23423 11758 23432
rect 11900 23186 11928 26200
rect 11978 25392 12034 25401
rect 11978 25327 12034 25336
rect 11796 23180 11848 23186
rect 11796 23122 11848 23128
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 11808 23089 11836 23122
rect 11794 23080 11850 23089
rect 11992 23032 12020 25327
rect 12072 25084 12124 25090
rect 12072 25026 12124 25032
rect 11794 23015 11850 23024
rect 11900 23004 12020 23032
rect 11900 22488 11928 23004
rect 11978 22944 12034 22953
rect 11978 22879 12034 22888
rect 11992 22710 12020 22879
rect 11980 22704 12032 22710
rect 11980 22646 12032 22652
rect 11900 22460 12020 22488
rect 11888 22160 11940 22166
rect 11888 22102 11940 22108
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11716 19854 11744 20742
rect 11794 20496 11850 20505
rect 11794 20431 11796 20440
rect 11848 20431 11850 20440
rect 11796 20402 11848 20408
rect 11704 19848 11756 19854
rect 11704 19790 11756 19796
rect 11610 19544 11666 19553
rect 11610 19479 11666 19488
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11532 18426 11560 19314
rect 11612 19236 11664 19242
rect 11612 19178 11664 19184
rect 11520 18420 11572 18426
rect 11520 18362 11572 18368
rect 11624 18358 11652 19178
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11612 18352 11664 18358
rect 11610 18320 11612 18329
rect 11664 18320 11666 18329
rect 11610 18255 11666 18264
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 11532 17649 11560 17682
rect 11518 17640 11574 17649
rect 11518 17575 11520 17584
rect 11572 17575 11574 17584
rect 11520 17546 11572 17552
rect 11348 16782 11468 16810
rect 11348 15502 11376 16782
rect 11426 16280 11482 16289
rect 11426 16215 11428 16224
rect 11480 16215 11482 16224
rect 11428 16186 11480 16192
rect 11518 16144 11574 16153
rect 11518 16079 11574 16088
rect 11428 16040 11480 16046
rect 11428 15982 11480 15988
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11242 14920 11298 14929
rect 11242 14855 11298 14864
rect 11152 14000 11204 14006
rect 11152 13942 11204 13948
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10782 13152 10838 13161
rect 10782 13087 10838 13096
rect 10784 12912 10836 12918
rect 10784 12854 10836 12860
rect 10692 12640 10744 12646
rect 10692 12582 10744 12588
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10692 12096 10744 12102
rect 10692 12038 10744 12044
rect 10612 11257 10640 12038
rect 10598 11248 10654 11257
rect 10598 11183 10654 11192
rect 10600 10600 10652 10606
rect 10600 10542 10652 10548
rect 10612 10033 10640 10542
rect 10598 10024 10654 10033
rect 10598 9959 10654 9968
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10428 8294 10456 8842
rect 10704 8362 10732 12038
rect 10796 11286 10824 12854
rect 10980 12434 11008 13738
rect 11060 13728 11112 13734
rect 11060 13670 11112 13676
rect 11072 12782 11100 13670
rect 11150 13560 11206 13569
rect 11150 13495 11206 13504
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 10980 12406 11100 12434
rect 10876 12368 10928 12374
rect 10876 12310 10928 12316
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10796 10198 10824 11086
rect 10888 10470 10916 12310
rect 10968 11824 11020 11830
rect 10968 11766 11020 11772
rect 10980 11393 11008 11766
rect 10966 11384 11022 11393
rect 10966 11319 11022 11328
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10980 10606 11008 11086
rect 11072 10742 11100 12406
rect 11164 11286 11192 13495
rect 11256 12345 11284 13874
rect 11348 13802 11376 15438
rect 11440 15337 11468 15982
rect 11426 15328 11482 15337
rect 11426 15263 11482 15272
rect 11428 14340 11480 14346
rect 11428 14282 11480 14288
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 13546 11376 13738
rect 11440 13705 11468 14282
rect 11426 13696 11482 13705
rect 11426 13631 11482 13640
rect 11348 13518 11468 13546
rect 11336 12844 11388 12850
rect 11336 12786 11388 12792
rect 11242 12336 11298 12345
rect 11242 12271 11298 12280
rect 11242 11792 11298 11801
rect 11242 11727 11244 11736
rect 11296 11727 11298 11736
rect 11244 11698 11296 11704
rect 11242 11384 11298 11393
rect 11242 11319 11298 11328
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 11256 11098 11284 11319
rect 11164 11070 11284 11098
rect 11060 10736 11112 10742
rect 11060 10678 11112 10684
rect 10968 10600 11020 10606
rect 11164 10577 11192 11070
rect 10968 10542 11020 10548
rect 11150 10568 11206 10577
rect 11150 10503 11206 10512
rect 10876 10464 10928 10470
rect 10876 10406 10928 10412
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 11072 10266 11100 10406
rect 11242 10296 11298 10305
rect 11060 10260 11112 10266
rect 11348 10266 11376 12786
rect 11440 12073 11468 13518
rect 11532 13326 11560 16079
rect 11624 13734 11652 17682
rect 11716 17202 11744 18770
rect 11808 17746 11836 20402
rect 11900 19786 11928 22102
rect 11992 20942 12020 22460
rect 12084 21690 12112 25026
rect 12254 24712 12310 24721
rect 12254 24647 12310 24656
rect 12348 24676 12400 24682
rect 12268 23798 12296 24647
rect 12348 24618 12400 24624
rect 12360 23798 12388 24618
rect 12544 24290 12572 26200
rect 13188 26160 13216 26200
rect 13280 26160 13308 26302
rect 13188 26132 13308 26160
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12452 24262 12572 24290
rect 12452 24070 12480 24262
rect 12532 24200 12584 24206
rect 12530 24168 12532 24177
rect 12584 24168 12586 24177
rect 12530 24103 12586 24112
rect 12440 24064 12492 24070
rect 12440 24006 12492 24012
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12348 23792 12400 23798
rect 12544 23780 12572 24006
rect 12348 23734 12400 23740
rect 12452 23752 12572 23780
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 19440 12032 19446
rect 11980 19382 12032 19388
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11900 17814 11928 19314
rect 11992 19310 12020 19382
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11888 17808 11940 17814
rect 11888 17750 11940 17756
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11794 17368 11850 17377
rect 11794 17303 11850 17312
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11716 15366 11744 17138
rect 11808 16454 11836 17303
rect 11992 17270 12020 18566
rect 12084 17814 12112 19654
rect 12072 17808 12124 17814
rect 12072 17750 12124 17756
rect 11980 17264 12032 17270
rect 11980 17206 12032 17212
rect 11992 16998 12020 17206
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11980 16448 12032 16454
rect 11980 16390 12032 16396
rect 11992 16182 12020 16390
rect 11980 16176 12032 16182
rect 11980 16118 12032 16124
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 11796 15904 11848 15910
rect 11848 15864 12020 15892
rect 11796 15846 11848 15852
rect 11888 15428 11940 15434
rect 11888 15370 11940 15376
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11716 14657 11744 15098
rect 11796 14816 11848 14822
rect 11794 14784 11796 14793
rect 11848 14784 11850 14793
rect 11794 14719 11850 14728
rect 11702 14648 11758 14657
rect 11702 14583 11758 14592
rect 11796 14408 11848 14414
rect 11900 14385 11928 15370
rect 11992 15337 12020 15864
rect 11978 15328 12034 15337
rect 11978 15263 12034 15272
rect 11796 14350 11848 14356
rect 11886 14376 11942 14385
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11520 13320 11572 13326
rect 11520 13262 11572 13268
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11532 12646 11560 12786
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11624 12442 11652 13466
rect 11808 13394 11836 14350
rect 11886 14311 11942 14320
rect 12084 14260 12112 16050
rect 11992 14232 12112 14260
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 13433 11928 13670
rect 11886 13424 11942 13433
rect 11796 13388 11848 13394
rect 11886 13359 11942 13368
rect 11796 13330 11848 13336
rect 11888 13252 11940 13258
rect 11888 13194 11940 13200
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11704 12912 11756 12918
rect 11702 12880 11704 12889
rect 11756 12880 11758 12889
rect 11702 12815 11758 12824
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11612 12436 11664 12442
rect 11612 12378 11664 12384
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11426 12064 11482 12073
rect 11532 12050 11560 12174
rect 11532 12022 11652 12050
rect 11426 11999 11482 12008
rect 11428 11892 11480 11898
rect 11428 11834 11480 11840
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11440 11801 11468 11834
rect 11426 11792 11482 11801
rect 11426 11727 11482 11736
rect 11532 11529 11560 11834
rect 11518 11520 11574 11529
rect 11518 11455 11574 11464
rect 11518 11248 11574 11257
rect 11428 11212 11480 11218
rect 11518 11183 11574 11192
rect 11428 11154 11480 11160
rect 11242 10231 11244 10240
rect 11060 10202 11112 10208
rect 11296 10231 11298 10240
rect 11336 10260 11388 10266
rect 11244 10202 11296 10208
rect 11336 10202 11388 10208
rect 10784 10192 10836 10198
rect 10784 10134 10836 10140
rect 10796 9674 10824 10134
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10796 9646 10916 9674
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10796 8945 10824 9522
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10796 8401 10824 8434
rect 10782 8392 10838 8401
rect 10692 8356 10744 8362
rect 10782 8327 10838 8336
rect 10692 8298 10744 8304
rect 10428 8266 10548 8294
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10324 7336 10376 7342
rect 10324 7278 10376 7284
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10244 6769 10272 6802
rect 10230 6760 10286 6769
rect 10230 6695 10286 6704
rect 10232 6656 10284 6662
rect 10230 6624 10232 6633
rect 10284 6624 10286 6633
rect 10230 6559 10286 6568
rect 10230 5944 10286 5953
rect 10230 5879 10232 5888
rect 10284 5879 10286 5888
rect 10232 5850 10284 5856
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9416 2746 9536 2774
rect 9508 2689 9536 2746
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9126 912 9182 921
rect 9126 847 9182 856
rect 9416 800 9444 2450
rect 10336 1494 10364 7278
rect 10428 5166 10456 7346
rect 10520 6780 10548 8266
rect 10598 8256 10654 8265
rect 10598 8191 10654 8200
rect 10612 7750 10640 8191
rect 10888 7954 10916 9646
rect 11072 9178 11100 10066
rect 11150 9752 11206 9761
rect 11150 9687 11206 9696
rect 11164 9518 11192 9687
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 10980 9030 11192 9058
rect 10980 8537 11008 9030
rect 11164 8974 11192 9030
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10966 8528 11022 8537
rect 11072 8498 11100 8842
rect 11150 8800 11206 8809
rect 11150 8735 11206 8744
rect 10966 8463 11022 8472
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 8424 11020 8430
rect 10968 8366 11020 8372
rect 10980 8022 11008 8366
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10968 8016 11020 8022
rect 10968 7958 11020 7964
rect 11072 7954 11100 8298
rect 11164 8022 11192 8735
rect 11256 8537 11284 10202
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11348 9654 11376 10066
rect 11336 9648 11388 9654
rect 11336 9590 11388 9596
rect 11334 9208 11390 9217
rect 11334 9143 11390 9152
rect 11348 9042 11376 9143
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11242 8528 11298 8537
rect 11242 8463 11298 8472
rect 11348 8294 11376 8774
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 10600 7744 10652 7750
rect 10600 7686 10652 7692
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10612 6934 10640 7686
rect 10980 7546 11008 7686
rect 11072 7546 11100 7890
rect 11244 7880 11296 7886
rect 11244 7822 11296 7828
rect 11334 7848 11390 7857
rect 11150 7712 11206 7721
rect 11150 7647 11206 7656
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7478 11192 7647
rect 11256 7585 11284 7822
rect 11334 7783 11390 7792
rect 11242 7576 11298 7585
rect 11242 7511 11298 7520
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11244 7404 11296 7410
rect 11244 7346 11296 7352
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 6934 10732 7278
rect 10968 7268 11020 7274
rect 10968 7210 11020 7216
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10692 6928 10744 6934
rect 10692 6870 10744 6876
rect 10980 6866 11008 7210
rect 10784 6860 10836 6866
rect 10784 6802 10836 6808
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10520 6752 10640 6780
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10520 3398 10548 6598
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10612 3058 10640 6752
rect 10692 6656 10744 6662
rect 10692 6598 10744 6604
rect 10704 6390 10732 6598
rect 10796 6497 10824 6802
rect 10874 6760 10930 6769
rect 10874 6695 10930 6704
rect 10888 6662 10916 6695
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10782 6488 10838 6497
rect 10782 6423 10838 6432
rect 10692 6384 10744 6390
rect 10692 6326 10744 6332
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10888 4758 10916 5646
rect 10980 5302 11008 6258
rect 11060 6248 11112 6254
rect 11060 6190 11112 6196
rect 11072 5545 11100 6190
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11058 5536 11114 5545
rect 11058 5471 11114 5480
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 10966 5128 11022 5137
rect 10966 5063 11022 5072
rect 10876 4752 10928 4758
rect 10876 4694 10928 4700
rect 10980 4690 11008 5063
rect 11164 4690 11192 6054
rect 10968 4684 11020 4690
rect 10968 4626 11020 4632
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 11152 4072 11204 4078
rect 11150 4040 11152 4049
rect 11204 4040 11206 4049
rect 11150 3975 11206 3984
rect 10874 3224 10930 3233
rect 10874 3159 10930 3168
rect 10888 3058 10916 3159
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11256 2774 11284 7346
rect 11348 7274 11376 7783
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11348 6225 11376 7210
rect 11334 6216 11390 6225
rect 11334 6151 11390 6160
rect 11334 5672 11390 5681
rect 11334 5607 11390 5616
rect 11348 5370 11376 5607
rect 11336 5364 11388 5370
rect 11336 5306 11388 5312
rect 11440 4826 11468 11154
rect 11532 10810 11560 11183
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10130 11560 10610
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11532 9586 11560 10066
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11520 9444 11572 9450
rect 11520 9386 11572 9392
rect 11532 9217 11560 9386
rect 11518 9208 11574 9217
rect 11518 9143 11574 9152
rect 11518 8936 11574 8945
rect 11518 8871 11574 8880
rect 11532 8498 11560 8871
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11532 7274 11560 8026
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11624 7154 11652 12022
rect 11716 11694 11744 12718
rect 11808 12617 11836 12922
rect 11794 12608 11850 12617
rect 11794 12543 11850 12552
rect 11900 12458 11928 13194
rect 11992 12986 12020 14232
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 12084 13258 12112 13670
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11808 12430 11928 12458
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11808 11540 11836 12430
rect 11980 12232 12032 12238
rect 11980 12174 12032 12180
rect 11888 12164 11940 12170
rect 11888 12106 11940 12112
rect 11900 11898 11928 12106
rect 11992 11898 12020 12174
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12084 11830 12112 12922
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11716 11512 11836 11540
rect 11716 10810 11744 11512
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11702 10568 11758 10577
rect 11702 10503 11758 10512
rect 11716 10470 11744 10503
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11702 9344 11758 9353
rect 11702 9279 11758 9288
rect 11716 8090 11744 9279
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11532 7126 11652 7154
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11532 4282 11560 7126
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11716 6118 11744 6734
rect 11704 6112 11756 6118
rect 11704 6054 11756 6060
rect 11610 5944 11666 5953
rect 11610 5879 11612 5888
rect 11664 5879 11666 5888
rect 11612 5850 11664 5856
rect 11716 5681 11744 6054
rect 11702 5672 11758 5681
rect 11808 5642 11836 11018
rect 11900 10538 11928 11698
rect 12176 11218 12204 23462
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12268 21622 12296 22578
rect 12256 21616 12308 21622
rect 12256 21558 12308 21564
rect 12256 21480 12308 21486
rect 12254 21448 12256 21457
rect 12308 21448 12310 21457
rect 12254 21383 12310 21392
rect 12360 21332 12388 23598
rect 12452 22488 12480 23752
rect 12636 23712 12664 25978
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12544 23684 12664 23712
rect 13360 23724 13412 23730
rect 12544 22817 12572 23684
rect 13360 23666 13412 23672
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 13372 23361 13400 23666
rect 13358 23352 13414 23361
rect 12624 23316 12676 23322
rect 13358 23287 13414 23296
rect 12624 23258 12676 23264
rect 12530 22808 12586 22817
rect 12530 22743 12586 22752
rect 12544 22710 12572 22743
rect 12532 22704 12584 22710
rect 12532 22646 12584 22652
rect 12452 22460 12572 22488
rect 12438 22400 12494 22409
rect 12438 22335 12494 22344
rect 12268 21304 12388 21332
rect 12268 20482 12296 21304
rect 12452 21162 12480 22335
rect 12544 22030 12572 22460
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12544 21321 12572 21966
rect 12530 21312 12586 21321
rect 12530 21247 12586 21256
rect 12360 21134 12480 21162
rect 12360 20602 12388 21134
rect 12348 20596 12400 20602
rect 12348 20538 12400 20544
rect 12268 20454 12388 20482
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12268 18222 12296 19246
rect 12360 18902 12388 20454
rect 12440 19372 12492 19378
rect 12636 19360 12664 23258
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12714 22264 12770 22273
rect 12714 22199 12770 22208
rect 12728 22166 12756 22199
rect 12716 22160 12768 22166
rect 12716 22102 12768 22108
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12728 20890 12756 21490
rect 12820 21010 12848 23122
rect 12992 23044 13044 23050
rect 12992 22986 13044 22992
rect 13360 23044 13412 23050
rect 13360 22986 13412 22992
rect 12898 22808 12954 22817
rect 12898 22743 12954 22752
rect 12912 22545 12940 22743
rect 13004 22710 13032 22986
rect 12992 22704 13044 22710
rect 12992 22646 13044 22652
rect 12898 22536 12954 22545
rect 12898 22471 12954 22480
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12808 21004 12860 21010
rect 12808 20946 12860 20952
rect 12728 20862 12940 20890
rect 12912 20534 12940 20862
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12992 20392 13044 20398
rect 12990 20360 12992 20369
rect 13044 20360 13046 20369
rect 12990 20295 13046 20304
rect 12714 20224 12770 20233
rect 12714 20159 12770 20168
rect 12728 19825 12756 20159
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 13176 19916 13228 19922
rect 13176 19858 13228 19864
rect 12714 19816 12770 19825
rect 12714 19751 12770 19760
rect 12808 19780 12860 19786
rect 12808 19722 12860 19728
rect 12636 19332 12756 19360
rect 12440 19314 12492 19320
rect 12452 18970 12480 19314
rect 12622 19272 12678 19281
rect 12622 19207 12678 19216
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12452 18358 12480 18906
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12256 18216 12308 18222
rect 12256 18158 12308 18164
rect 12544 17921 12572 19110
rect 12636 18970 12664 19207
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12728 18873 12756 19332
rect 12714 18864 12770 18873
rect 12714 18799 12770 18808
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12530 17912 12586 17921
rect 12530 17847 12586 17856
rect 12348 17740 12400 17746
rect 12348 17682 12400 17688
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12268 15162 12296 17478
rect 12360 15201 12388 17682
rect 12532 17604 12584 17610
rect 12452 17564 12532 17592
rect 12452 15910 12480 17564
rect 12532 17546 12584 17552
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12636 17134 12664 17478
rect 12624 17128 12676 17134
rect 12624 17070 12676 17076
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12530 16416 12586 16425
rect 12530 16351 12586 16360
rect 12440 15904 12492 15910
rect 12440 15846 12492 15852
rect 12544 15609 12572 16351
rect 12530 15600 12586 15609
rect 12530 15535 12586 15544
rect 12636 15434 12664 16934
rect 12624 15428 12676 15434
rect 12624 15370 12676 15376
rect 12532 15360 12584 15366
rect 12532 15302 12584 15308
rect 12544 15201 12572 15302
rect 12346 15192 12402 15201
rect 12256 15156 12308 15162
rect 12346 15127 12402 15136
rect 12530 15192 12586 15201
rect 12530 15127 12586 15136
rect 12256 15098 12308 15104
rect 12440 15020 12492 15026
rect 12440 14962 12492 14968
rect 12452 14618 12480 14962
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12544 14618 12572 14894
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 12544 13977 12572 14554
rect 12636 14346 12664 15370
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12530 13968 12586 13977
rect 12530 13903 12586 13912
rect 12532 13796 12584 13802
rect 12636 13784 12664 14282
rect 12584 13756 12664 13784
rect 12532 13738 12584 13744
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 11830 12296 13330
rect 12636 13258 12664 13756
rect 12728 13530 12756 18702
rect 12820 17882 12848 19722
rect 13188 19281 13216 19858
rect 13174 19272 13230 19281
rect 13174 19207 13230 19216
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 13372 18465 13400 22986
rect 13464 22098 13492 26302
rect 13818 26200 13874 27000
rect 14462 26200 14518 27000
rect 14740 26376 14792 26382
rect 14740 26318 14792 26324
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13636 24880 13688 24886
rect 13636 24822 13688 24828
rect 13542 24304 13598 24313
rect 13542 24239 13598 24248
rect 13556 23322 13584 24239
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13544 23180 13596 23186
rect 13544 23122 13596 23128
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13556 21962 13584 23122
rect 13544 21956 13596 21962
rect 13544 21898 13596 21904
rect 13556 21486 13584 21898
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13544 21344 13596 21350
rect 13544 21286 13596 21292
rect 13556 20398 13584 21286
rect 13544 20392 13596 20398
rect 13544 20334 13596 20340
rect 13452 19916 13504 19922
rect 13452 19858 13504 19864
rect 13464 19718 13492 19858
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13556 19446 13584 20334
rect 13544 19440 13596 19446
rect 13544 19382 13596 19388
rect 13648 18970 13676 24822
rect 13740 24750 13768 24890
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13832 24138 13860 26200
rect 14188 26172 14240 26178
rect 14188 26114 14240 26120
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 13910 24304 13966 24313
rect 13910 24239 13966 24248
rect 13820 24132 13872 24138
rect 13820 24074 13872 24080
rect 13924 23798 13952 24239
rect 13912 23792 13964 23798
rect 13912 23734 13964 23740
rect 13912 23520 13964 23526
rect 13912 23462 13964 23468
rect 13924 23254 13952 23462
rect 13912 23248 13964 23254
rect 13912 23190 13964 23196
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22137 13768 22918
rect 14016 22794 14044 24550
rect 14200 24070 14228 26114
rect 14476 24342 14504 26200
rect 14556 25560 14608 25566
rect 14556 25502 14608 25508
rect 14464 24336 14516 24342
rect 14464 24278 14516 24284
rect 14372 24268 14424 24274
rect 14372 24210 14424 24216
rect 14278 24168 14334 24177
rect 14278 24103 14334 24112
rect 14292 24070 14320 24103
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14280 24064 14332 24070
rect 14280 24006 14332 24012
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 14096 23248 14148 23254
rect 14096 23190 14148 23196
rect 14108 22953 14136 23190
rect 14094 22944 14150 22953
rect 14094 22879 14150 22888
rect 14016 22766 14136 22794
rect 14004 22432 14056 22438
rect 14004 22374 14056 22380
rect 13726 22128 13782 22137
rect 13782 22086 13860 22114
rect 13726 22063 13782 22072
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13740 19961 13768 21422
rect 13832 20369 13860 22086
rect 13818 20360 13874 20369
rect 13818 20295 13874 20304
rect 14016 20233 14044 22374
rect 14108 20534 14136 22766
rect 14096 20528 14148 20534
rect 14096 20470 14148 20476
rect 14002 20224 14058 20233
rect 14002 20159 14058 20168
rect 14096 19984 14148 19990
rect 13726 19952 13782 19961
rect 14096 19926 14148 19932
rect 13726 19887 13782 19896
rect 13820 19848 13872 19854
rect 13818 19816 13820 19825
rect 13872 19816 13874 19825
rect 13818 19751 13874 19760
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13636 18964 13688 18970
rect 13636 18906 13688 18912
rect 13358 18456 13414 18465
rect 12900 18420 12952 18426
rect 13358 18391 13414 18400
rect 12900 18362 12952 18368
rect 12912 18086 12940 18362
rect 12900 18080 12952 18086
rect 13372 18057 13400 18391
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 12900 18022 12952 18028
rect 13358 18048 13414 18057
rect 12950 17980 13258 17989
rect 13358 17983 13414 17992
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12808 17876 12860 17882
rect 12808 17818 12860 17824
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13280 16980 13308 17478
rect 13464 16998 13492 18158
rect 13740 17954 13768 19654
rect 13820 19236 13872 19242
rect 13820 19178 13872 19184
rect 13556 17926 13768 17954
rect 13452 16992 13504 16998
rect 13280 16952 13400 16980
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 13372 16794 13400 16952
rect 13452 16934 13504 16940
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 12992 16652 13044 16658
rect 12992 16594 13044 16600
rect 13004 16250 13032 16594
rect 13268 16584 13320 16590
rect 13360 16584 13412 16590
rect 13268 16526 13320 16532
rect 13358 16552 13360 16561
rect 13412 16552 13414 16561
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12900 16176 12952 16182
rect 12898 16144 12900 16153
rect 12952 16144 12954 16153
rect 12898 16079 12954 16088
rect 13280 15994 13308 16526
rect 13358 16487 13414 16496
rect 13358 16144 13414 16153
rect 13358 16079 13360 16088
rect 13412 16079 13414 16088
rect 13360 16050 13412 16056
rect 13280 15966 13400 15994
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 13268 15496 13320 15502
rect 13268 15438 13320 15444
rect 13176 15428 13228 15434
rect 13176 15370 13228 15376
rect 13188 15094 13216 15370
rect 13176 15088 13228 15094
rect 13176 15030 13228 15036
rect 13280 14822 13308 15438
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12806 14648 12862 14657
rect 12950 14651 13258 14660
rect 12862 14592 12940 14600
rect 12806 14583 12940 14592
rect 12820 14572 12940 14583
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12532 13184 12584 13190
rect 12532 13126 12584 13132
rect 12348 12300 12400 12306
rect 12348 12242 12400 12248
rect 12360 11898 12388 12242
rect 12438 11928 12494 11937
rect 12348 11892 12400 11898
rect 12438 11863 12440 11872
rect 12348 11834 12400 11840
rect 12492 11863 12494 11872
rect 12440 11834 12492 11840
rect 12256 11824 12308 11830
rect 12256 11766 12308 11772
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 11218 12296 11630
rect 12164 11212 12216 11218
rect 12164 11154 12216 11160
rect 12256 11212 12308 11218
rect 12256 11154 12308 11160
rect 11980 11008 12032 11014
rect 11980 10950 12032 10956
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11992 10470 12020 10950
rect 12072 10600 12124 10606
rect 12072 10542 12124 10548
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11992 10169 12020 10406
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 12084 10033 12112 10542
rect 12162 10296 12218 10305
rect 12162 10231 12218 10240
rect 12070 10024 12126 10033
rect 11888 9988 11940 9994
rect 12070 9959 12126 9968
rect 11888 9930 11940 9936
rect 11900 9654 11928 9930
rect 12176 9722 12204 10231
rect 12072 9716 12124 9722
rect 11992 9664 12072 9674
rect 11992 9658 12124 9664
rect 12164 9716 12216 9722
rect 12164 9658 12216 9664
rect 11888 9648 11940 9654
rect 11886 9616 11888 9625
rect 11992 9646 12112 9658
rect 11940 9616 11942 9625
rect 11886 9551 11942 9560
rect 11992 9194 12020 9646
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 9382 12112 9454
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 11992 9166 12112 9194
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11702 5607 11758 5616
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11702 5264 11758 5273
rect 11702 5199 11758 5208
rect 11716 5166 11744 5199
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11716 4282 11744 5102
rect 11520 4276 11572 4282
rect 11520 4218 11572 4224
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11428 4140 11480 4146
rect 11428 4082 11480 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11348 3670 11376 4014
rect 11336 3664 11388 3670
rect 11336 3606 11388 3612
rect 11440 2774 11468 4082
rect 11900 3534 11928 8774
rect 11992 8362 12020 9007
rect 12084 8838 12112 9166
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12176 8634 12204 9658
rect 12164 8628 12216 8634
rect 12164 8570 12216 8576
rect 12268 8514 12296 11154
rect 12360 9761 12388 11698
rect 12440 11552 12492 11558
rect 12440 11494 12492 11500
rect 12452 11354 12480 11494
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12440 11008 12492 11014
rect 12440 10950 12492 10956
rect 12346 9752 12402 9761
rect 12346 9687 12402 9696
rect 12452 9636 12480 10950
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12176 8486 12296 8514
rect 12360 9608 12480 9636
rect 12544 9625 12572 13126
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 12636 12306 12664 12650
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12530 9616 12586 9625
rect 11980 8356 12032 8362
rect 11980 8298 12032 8304
rect 12084 7970 12112 8434
rect 12176 8294 12204 8486
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12162 8120 12218 8129
rect 12162 8055 12218 8064
rect 11992 7942 12112 7970
rect 11888 3528 11940 3534
rect 11888 3470 11940 3476
rect 11992 3466 12020 7942
rect 12176 7886 12204 8055
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 7206 12112 7754
rect 12162 7712 12218 7721
rect 12162 7647 12218 7656
rect 12176 7313 12204 7647
rect 12268 7546 12296 8366
rect 12360 7750 12388 9608
rect 12530 9551 12586 9560
rect 12532 9512 12584 9518
rect 12438 9480 12494 9489
rect 12532 9454 12584 9460
rect 12438 9415 12494 9424
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12452 7698 12480 9415
rect 12544 8566 12572 9454
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12452 7670 12572 7698
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12162 7304 12218 7313
rect 12162 7239 12218 7248
rect 12072 7200 12124 7206
rect 12072 7142 12124 7148
rect 12162 7168 12218 7177
rect 12162 7103 12218 7112
rect 12072 6792 12124 6798
rect 12070 6760 12072 6769
rect 12124 6760 12126 6769
rect 12070 6695 12126 6704
rect 12084 5370 12112 6695
rect 12176 6322 12204 7103
rect 12452 6769 12480 7482
rect 12544 6866 12572 7670
rect 12636 7478 12664 12038
rect 12728 11014 12756 12786
rect 12820 12102 12848 14214
rect 12912 13870 12940 14572
rect 13372 14414 13400 15966
rect 13360 14408 13412 14414
rect 13360 14350 13412 14356
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12900 13864 12952 13870
rect 12900 13806 12952 13812
rect 13096 13734 13124 14214
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13280 13802 13308 14010
rect 13268 13796 13320 13802
rect 13268 13738 13320 13744
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13096 12714 13124 13126
rect 13280 12782 13308 13398
rect 13360 12912 13412 12918
rect 13360 12854 13412 12860
rect 13268 12776 13320 12782
rect 13174 12744 13230 12753
rect 13084 12708 13136 12714
rect 13268 12718 13320 12724
rect 13372 12714 13400 12854
rect 13174 12679 13176 12688
rect 13084 12650 13136 12656
rect 13228 12679 13230 12688
rect 13360 12708 13412 12714
rect 13176 12650 13228 12656
rect 13360 12650 13412 12656
rect 13464 12594 13492 16934
rect 13372 12566 13492 12594
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11286 12848 11698
rect 12912 11626 12940 12242
rect 12900 11620 12952 11626
rect 12900 11562 12952 11568
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 13280 11121 13308 11290
rect 13266 11112 13322 11121
rect 12808 11076 12860 11082
rect 13266 11047 13322 11056
rect 12808 11018 12860 11024
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12820 10742 12848 11018
rect 12808 10736 12860 10742
rect 12728 10696 12808 10724
rect 12728 9926 12756 10696
rect 12808 10678 12860 10684
rect 12806 10432 12862 10441
rect 12806 10367 12862 10376
rect 12820 10248 12848 10367
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12820 10220 13032 10248
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 13004 9674 13032 10220
rect 13372 10180 13400 12566
rect 13556 12442 13584 17926
rect 13728 17740 13780 17746
rect 13728 17682 13780 17688
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13648 16658 13676 16934
rect 13636 16652 13688 16658
rect 13636 16594 13688 16600
rect 13740 16289 13768 17682
rect 13832 16658 13860 19178
rect 13912 18964 13964 18970
rect 13912 18906 13964 18912
rect 13924 18737 13952 18906
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13910 18728 13966 18737
rect 13910 18663 13966 18672
rect 13912 18284 13964 18290
rect 13912 18226 13964 18232
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13924 16522 13952 18226
rect 14016 16969 14044 18838
rect 14108 17338 14136 19926
rect 14200 19122 14228 23258
rect 14384 23225 14412 24210
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14476 23866 14504 24142
rect 14464 23860 14516 23866
rect 14464 23802 14516 23808
rect 14370 23216 14426 23225
rect 14370 23151 14426 23160
rect 14280 22976 14332 22982
rect 14384 22953 14412 23151
rect 14280 22918 14332 22924
rect 14370 22944 14426 22953
rect 14292 22545 14320 22918
rect 14568 22930 14596 25502
rect 14646 23216 14702 23225
rect 14752 23186 14780 26318
rect 15106 26200 15162 27000
rect 15750 26200 15806 27000
rect 16394 26330 16450 27000
rect 17038 26602 17094 27000
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 17038 26574 17356 26602
rect 16132 26302 16450 26330
rect 14832 25560 14884 25566
rect 14832 25502 14884 25508
rect 14646 23151 14702 23160
rect 14740 23180 14792 23186
rect 14660 23118 14688 23151
rect 14740 23122 14792 23128
rect 14648 23112 14700 23118
rect 14648 23054 14700 23060
rect 14740 22976 14792 22982
rect 14568 22902 14688 22930
rect 14740 22918 14792 22924
rect 14370 22879 14426 22888
rect 14556 22636 14608 22642
rect 14556 22578 14608 22584
rect 14278 22536 14334 22545
rect 14278 22471 14334 22480
rect 14280 22024 14332 22030
rect 14280 21966 14332 21972
rect 14292 19990 14320 21966
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14372 21412 14424 21418
rect 14372 21354 14424 21360
rect 14384 21146 14412 21354
rect 14372 21140 14424 21146
rect 14372 21082 14424 21088
rect 14372 20936 14424 20942
rect 14372 20878 14424 20884
rect 14384 20505 14412 20878
rect 14476 20534 14504 21490
rect 14464 20528 14516 20534
rect 14370 20496 14426 20505
rect 14464 20470 14516 20476
rect 14370 20431 14426 20440
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14372 19848 14424 19854
rect 14278 19816 14334 19825
rect 14372 19790 14424 19796
rect 14278 19751 14334 19760
rect 14292 19242 14320 19751
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14200 19094 14320 19122
rect 14186 18184 14242 18193
rect 14186 18119 14242 18128
rect 14200 17338 14228 18119
rect 14292 17513 14320 19094
rect 14384 18834 14412 19790
rect 14476 19718 14504 20470
rect 14464 19712 14516 19718
rect 14464 19654 14516 19660
rect 14462 18864 14518 18873
rect 14372 18828 14424 18834
rect 14462 18799 14464 18808
rect 14372 18770 14424 18776
rect 14516 18799 14518 18808
rect 14464 18770 14516 18776
rect 14384 18358 14412 18770
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 14384 17921 14412 18022
rect 14370 17912 14426 17921
rect 14568 17882 14596 22578
rect 14660 22094 14688 22902
rect 14752 22234 14780 22918
rect 14844 22642 14872 25502
rect 15016 25356 15068 25362
rect 15016 25298 15068 25304
rect 15028 24041 15056 25298
rect 15014 24032 15070 24041
rect 15014 23967 15070 23976
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14936 23497 14964 23666
rect 14922 23488 14978 23497
rect 14922 23423 14978 23432
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 14832 22432 14884 22438
rect 14830 22400 14832 22409
rect 14884 22400 14886 22409
rect 14830 22335 14886 22344
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14660 22066 14780 22094
rect 14648 22024 14700 22030
rect 14648 21966 14700 21972
rect 14660 21010 14688 21966
rect 14648 21004 14700 21010
rect 14648 20946 14700 20952
rect 14648 20868 14700 20874
rect 14648 20810 14700 20816
rect 14660 20097 14688 20810
rect 14646 20088 14702 20097
rect 14646 20023 14702 20032
rect 14648 19780 14700 19786
rect 14648 19722 14700 19728
rect 14660 19689 14688 19722
rect 14646 19680 14702 19689
rect 14646 19615 14702 19624
rect 14646 18728 14702 18737
rect 14646 18663 14702 18672
rect 14660 18426 14688 18663
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14370 17847 14426 17856
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14568 17678 14596 17818
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14372 17536 14424 17542
rect 14278 17504 14334 17513
rect 14372 17478 14424 17484
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14646 17504 14702 17513
rect 14278 17439 14334 17448
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14188 17332 14240 17338
rect 14188 17274 14240 17280
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14096 16992 14148 16998
rect 14002 16960 14058 16969
rect 14096 16934 14148 16940
rect 14002 16895 14058 16904
rect 14108 16776 14136 16934
rect 14016 16748 14136 16776
rect 13912 16516 13964 16522
rect 13912 16458 13964 16464
rect 14016 16454 14044 16748
rect 14292 16590 14320 17138
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14280 16448 14332 16454
rect 14280 16390 14332 16396
rect 13726 16280 13782 16289
rect 13726 16215 13782 16224
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13636 15088 13688 15094
rect 13634 15056 13636 15065
rect 13688 15056 13690 15065
rect 13634 14991 13690 15000
rect 13636 14816 13688 14822
rect 13832 14793 13860 15846
rect 13924 15450 13952 15982
rect 14016 15745 14044 16390
rect 14002 15736 14058 15745
rect 14002 15671 14058 15680
rect 14016 15570 14044 15671
rect 14108 15609 14136 16390
rect 14292 16182 14320 16390
rect 14384 16250 14412 17478
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 14280 16176 14332 16182
rect 14476 16130 14504 17478
rect 14646 17439 14702 17448
rect 14660 17218 14688 17439
rect 14752 17320 14780 22066
rect 14844 21486 14872 22170
rect 14936 22137 14964 22578
rect 14922 22128 14978 22137
rect 15120 22098 15148 26200
rect 15658 24440 15714 24449
rect 15658 24375 15714 24384
rect 15290 23760 15346 23769
rect 15290 23695 15346 23704
rect 15304 23594 15332 23695
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 14922 22063 14978 22072
rect 15108 22092 15160 22098
rect 14936 22001 14964 22063
rect 15108 22034 15160 22040
rect 15212 22030 15240 23530
rect 15474 23488 15530 23497
rect 15474 23423 15530 23432
rect 15488 23118 15516 23423
rect 15476 23112 15528 23118
rect 15396 23060 15476 23066
rect 15396 23054 15528 23060
rect 15396 23038 15516 23054
rect 15200 22024 15252 22030
rect 14922 21992 14978 22001
rect 14922 21927 14978 21936
rect 15198 21992 15200 22001
rect 15252 21992 15254 22001
rect 15198 21927 15254 21936
rect 15396 21865 15424 23038
rect 15566 22944 15622 22953
rect 15566 22879 15622 22888
rect 15476 22568 15528 22574
rect 15476 22510 15528 22516
rect 15382 21856 15438 21865
rect 15382 21791 15438 21800
rect 15108 21616 15160 21622
rect 15106 21584 15108 21593
rect 15160 21584 15162 21593
rect 15106 21519 15162 21528
rect 14832 21480 14884 21486
rect 14832 21422 14884 21428
rect 15108 21480 15160 21486
rect 15108 21422 15160 21428
rect 14924 21344 14976 21350
rect 14924 21286 14976 21292
rect 15120 21298 15148 21422
rect 15384 21344 15436 21350
rect 14832 20868 14884 20874
rect 14832 20810 14884 20816
rect 14844 20641 14872 20810
rect 14830 20632 14886 20641
rect 14830 20567 14886 20576
rect 14830 20224 14886 20233
rect 14830 20159 14886 20168
rect 14844 19310 14872 20159
rect 14936 19378 14964 21286
rect 15120 21270 15240 21298
rect 15384 21286 15436 21292
rect 15108 21140 15160 21146
rect 15108 21082 15160 21088
rect 15120 21049 15148 21082
rect 15106 21040 15162 21049
rect 15212 21010 15240 21270
rect 15106 20975 15162 20984
rect 15200 21004 15252 21010
rect 15200 20946 15252 20952
rect 15198 19952 15254 19961
rect 15198 19887 15254 19896
rect 15292 19916 15344 19922
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14832 19304 14884 19310
rect 14832 19246 14884 19252
rect 14844 18970 14872 19246
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14844 17882 14872 18906
rect 14936 18086 14964 19314
rect 15016 18692 15068 18698
rect 15016 18634 15068 18640
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14830 17776 14886 17785
rect 14936 17746 14964 18022
rect 14830 17711 14886 17720
rect 14924 17740 14976 17746
rect 14844 17513 14872 17711
rect 14924 17682 14976 17688
rect 14830 17504 14886 17513
rect 14830 17439 14886 17448
rect 14832 17332 14884 17338
rect 14752 17292 14832 17320
rect 14832 17274 14884 17280
rect 14738 17232 14794 17241
rect 14660 17190 14738 17218
rect 14738 17167 14794 17176
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14832 17128 14884 17134
rect 14832 17070 14884 17076
rect 14660 16402 14688 17070
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14752 16697 14780 16730
rect 14738 16688 14794 16697
rect 14738 16623 14794 16632
rect 14752 16522 14780 16623
rect 14740 16516 14792 16522
rect 14740 16458 14792 16464
rect 14660 16374 14780 16402
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14280 16118 14332 16124
rect 14384 16102 14504 16130
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 14094 15600 14150 15609
rect 14004 15564 14056 15570
rect 14094 15535 14150 15544
rect 14004 15506 14056 15512
rect 13924 15422 14044 15450
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13636 14758 13688 14764
rect 13818 14784 13874 14793
rect 13648 13938 13676 14758
rect 13818 14719 13874 14728
rect 13924 14618 13952 14962
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13726 14512 13782 14521
rect 13726 14447 13782 14456
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13636 13728 13688 13734
rect 13636 13670 13688 13676
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13544 12300 13596 12306
rect 13464 12260 13544 12288
rect 13464 11914 13492 12260
rect 13544 12242 13596 12248
rect 13648 12186 13676 13670
rect 13556 12158 13676 12186
rect 13556 12073 13584 12158
rect 13636 12096 13688 12102
rect 13542 12064 13598 12073
rect 13636 12038 13688 12044
rect 13542 11999 13598 12008
rect 13464 11886 13584 11914
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13280 10152 13400 10180
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13004 9646 13124 9674
rect 13096 9450 13124 9646
rect 13188 9518 13216 9862
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 13280 9364 13308 10152
rect 13360 9716 13412 9722
rect 13360 9658 13412 9664
rect 13372 9432 13400 9658
rect 13464 9500 13492 11766
rect 13556 11354 13584 11886
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13542 11248 13598 11257
rect 13542 11183 13598 11192
rect 13556 10538 13584 11183
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13556 9722 13584 9862
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13464 9472 13584 9500
rect 13372 9404 13492 9432
rect 13280 9336 13400 9364
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 13372 9160 13400 9336
rect 13280 9132 13400 9160
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12912 8838 12940 8978
rect 13280 8945 13308 9132
rect 13464 9092 13492 9404
rect 13372 9064 13492 9092
rect 13372 8974 13400 9064
rect 13556 9024 13584 9472
rect 13464 8996 13584 9024
rect 13360 8968 13412 8974
rect 13266 8936 13322 8945
rect 13360 8910 13412 8916
rect 13266 8871 13322 8880
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12808 8288 12860 8294
rect 12808 8230 12860 8236
rect 12624 7472 12676 7478
rect 12624 7414 12676 7420
rect 12532 6860 12584 6866
rect 12532 6802 12584 6808
rect 12438 6760 12494 6769
rect 12438 6695 12494 6704
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12728 6202 12756 8230
rect 12636 6174 12756 6202
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12452 5386 12480 5646
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12268 5358 12480 5386
rect 12072 5024 12124 5030
rect 12072 4966 12124 4972
rect 12084 4826 12112 4966
rect 12072 4820 12124 4826
rect 12072 4762 12124 4768
rect 12084 4146 12112 4762
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12164 4140 12216 4146
rect 12164 4082 12216 4088
rect 12176 3738 12204 4082
rect 12164 3732 12216 3738
rect 12164 3674 12216 3680
rect 12268 3618 12296 5358
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12348 4616 12400 4622
rect 12452 4570 12480 5170
rect 12400 4564 12480 4570
rect 12348 4558 12480 4564
rect 12360 4542 12480 4558
rect 12438 4312 12494 4321
rect 12438 4247 12494 4256
rect 12176 3590 12296 3618
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12084 2938 12112 3130
rect 12176 3058 12204 3590
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12164 3052 12216 3058
rect 12164 2994 12216 3000
rect 12360 2938 12388 3470
rect 12084 2910 12388 2938
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11072 2746 11284 2774
rect 11348 2746 11468 2774
rect 10966 1864 11022 1873
rect 10966 1799 11022 1808
rect 10980 1698 11008 1799
rect 10968 1692 11020 1698
rect 10968 1634 11020 1640
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 11072 1426 11100 2746
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 1630 11192 2246
rect 11152 1624 11204 1630
rect 11152 1566 11204 1572
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 11348 1358 11376 2746
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 2106 11560 2246
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11704 2032 11756 2038
rect 11704 1974 11756 1980
rect 11336 1352 11388 1358
rect 11336 1294 11388 1300
rect 11716 1290 11744 1974
rect 11900 1766 11928 2790
rect 12452 2689 12480 4247
rect 12544 3942 12572 5510
rect 12636 4554 12664 6174
rect 12716 6112 12768 6118
rect 12714 6080 12716 6089
rect 12768 6080 12770 6089
rect 12714 6015 12770 6024
rect 12820 5914 12848 8230
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 13188 7886 13216 8026
rect 13176 7880 13228 7886
rect 13176 7822 13228 7828
rect 12898 7576 12954 7585
rect 12898 7511 12954 7520
rect 12912 7342 12940 7511
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12714 5808 12770 5817
rect 12714 5743 12770 5752
rect 12728 5234 12756 5743
rect 12808 5636 12860 5642
rect 12808 5578 12860 5584
rect 12820 5370 12848 5578
rect 12808 5364 12860 5370
rect 12808 5306 12860 5312
rect 13372 5234 13400 8774
rect 13464 6866 13492 8996
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13556 8537 13584 8871
rect 13542 8528 13598 8537
rect 13542 8463 13598 8472
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 6860 13504 6866
rect 13452 6802 13504 6808
rect 13450 6760 13506 6769
rect 13450 6695 13506 6704
rect 13464 5370 13492 6695
rect 13556 5574 13584 8298
rect 13648 6633 13676 12038
rect 13740 8090 13768 14447
rect 13912 14408 13964 14414
rect 13912 14350 13964 14356
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13832 12646 13860 14282
rect 13924 13002 13952 14350
rect 14016 13190 14044 15422
rect 14096 15360 14148 15366
rect 14096 15302 14148 15308
rect 14108 15162 14136 15302
rect 14200 15162 14228 15846
rect 14292 15706 14320 15846
rect 14280 15700 14332 15706
rect 14280 15642 14332 15648
rect 14278 15464 14334 15473
rect 14278 15399 14334 15408
rect 14096 15156 14148 15162
rect 14096 15098 14148 15104
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14108 13734 14136 15098
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 14200 14482 14228 14962
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 14096 13728 14148 13734
rect 14096 13670 14148 13676
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13924 12974 14044 13002
rect 13910 12880 13966 12889
rect 13910 12815 13966 12824
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13924 11937 13952 12815
rect 13910 11928 13966 11937
rect 13910 11863 13966 11872
rect 13818 11792 13874 11801
rect 13818 11727 13874 11736
rect 13832 11354 13860 11727
rect 13912 11688 13964 11694
rect 13912 11630 13964 11636
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13818 11248 13874 11257
rect 13818 11183 13820 11192
rect 13872 11183 13874 11192
rect 13820 11154 13872 11160
rect 13820 11008 13872 11014
rect 13818 10976 13820 10985
rect 13872 10976 13874 10985
rect 13818 10911 13874 10920
rect 13818 10840 13874 10849
rect 13818 10775 13874 10784
rect 13832 10198 13860 10775
rect 13820 10192 13872 10198
rect 13818 10160 13820 10169
rect 13872 10160 13874 10169
rect 13818 10095 13874 10104
rect 13818 10024 13874 10033
rect 13818 9959 13874 9968
rect 13832 9382 13860 9959
rect 13820 9376 13872 9382
rect 13820 9318 13872 9324
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 13740 7002 13768 7239
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13634 6624 13690 6633
rect 13634 6559 13690 6568
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 5914 13768 6258
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13452 5364 13504 5370
rect 13452 5306 13504 5312
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13832 5030 13860 9318
rect 13924 8838 13952 11630
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13910 8120 13966 8129
rect 13910 8055 13966 8064
rect 13924 7954 13952 8055
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13924 5710 13952 6666
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13912 5160 13964 5166
rect 13912 5102 13964 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13818 4584 13874 4593
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12728 3058 12756 4558
rect 13740 4486 13768 4558
rect 13818 4519 13874 4528
rect 13636 4480 13688 4486
rect 13636 4422 13688 4428
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 13372 3233 13400 4082
rect 13452 4004 13504 4010
rect 13452 3946 13504 3952
rect 13082 3224 13138 3233
rect 13082 3159 13138 3168
rect 13358 3224 13414 3233
rect 13358 3159 13414 3168
rect 13096 3058 13124 3159
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12624 2848 12676 2854
rect 13360 2848 13412 2854
rect 12624 2790 12676 2796
rect 13358 2816 13360 2825
rect 13412 2816 13414 2825
rect 12438 2680 12494 2689
rect 12438 2615 12494 2624
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11704 1284 11756 1290
rect 11704 1226 11756 1232
rect 12084 800 12112 2450
rect 12636 2378 12664 2790
rect 12950 2748 13258 2757
rect 13358 2751 13414 2760
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13464 2689 13492 3946
rect 13556 3738 13584 4082
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13544 3052 13596 3058
rect 13544 2994 13596 3000
rect 13450 2680 13506 2689
rect 13556 2650 13584 2994
rect 13450 2615 13506 2624
rect 13544 2644 13596 2650
rect 13544 2586 13596 2592
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 13648 1222 13676 4422
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13740 4010 13768 4218
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13832 2666 13860 4519
rect 13740 2638 13860 2666
rect 13740 1873 13768 2638
rect 13726 1864 13782 1873
rect 13726 1799 13782 1808
rect 13636 1216 13688 1222
rect 13924 1193 13952 5102
rect 14016 2650 14044 12974
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14200 11529 14228 11834
rect 14186 11520 14242 11529
rect 14186 11455 14242 11464
rect 14188 11280 14240 11286
rect 14188 11222 14240 11228
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14108 10130 14136 10678
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14096 9920 14148 9926
rect 14094 9888 14096 9897
rect 14148 9888 14150 9897
rect 14094 9823 14150 9832
rect 14200 9466 14228 11222
rect 14108 9438 14228 9466
rect 14108 9110 14136 9438
rect 14188 9376 14240 9382
rect 14186 9344 14188 9353
rect 14240 9344 14242 9353
rect 14186 9279 14242 9288
rect 14096 9104 14148 9110
rect 14096 9046 14148 9052
rect 14094 8528 14150 8537
rect 14094 8463 14150 8472
rect 14108 6633 14136 8463
rect 14186 8392 14242 8401
rect 14186 8327 14242 8336
rect 14094 6624 14150 6633
rect 14094 6559 14150 6568
rect 14200 6186 14228 8327
rect 14292 8294 14320 15399
rect 14384 14822 14412 16102
rect 14462 16008 14518 16017
rect 14462 15943 14464 15952
rect 14516 15943 14518 15952
rect 14464 15914 14516 15920
rect 14462 15736 14518 15745
rect 14462 15671 14518 15680
rect 14476 14958 14504 15671
rect 14660 15502 14688 16186
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14556 15428 14608 15434
rect 14556 15370 14608 15376
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14568 14482 14596 15370
rect 14660 14822 14688 15438
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14556 14476 14608 14482
rect 14556 14418 14608 14424
rect 14648 14408 14700 14414
rect 14648 14350 14700 14356
rect 14660 14006 14688 14350
rect 14648 14000 14700 14006
rect 14648 13942 14700 13948
rect 14660 13394 14688 13942
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14648 13252 14700 13258
rect 14648 13194 14700 13200
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14476 12918 14504 13126
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 11898 14412 12582
rect 14568 12434 14596 12718
rect 14476 12406 14596 12434
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 14370 11792 14426 11801
rect 14370 11727 14426 11736
rect 14384 11082 14412 11727
rect 14476 11354 14504 12406
rect 14554 11792 14610 11801
rect 14554 11727 14610 11736
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14568 11286 14596 11727
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 14372 11076 14424 11082
rect 14372 11018 14424 11024
rect 14384 10713 14412 11018
rect 14476 10810 14504 11086
rect 14554 10976 14610 10985
rect 14554 10911 14610 10920
rect 14568 10810 14596 10911
rect 14464 10804 14516 10810
rect 14464 10746 14516 10752
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14370 10704 14426 10713
rect 14370 10639 14426 10648
rect 14372 10600 14424 10606
rect 14372 10542 14424 10548
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 14292 7449 14320 7686
rect 14278 7440 14334 7449
rect 14278 7375 14334 7384
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4214 14136 4966
rect 14292 4214 14320 5646
rect 14384 4826 14412 10542
rect 14476 10062 14504 10746
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 10056 14516 10062
rect 14568 10033 14596 10406
rect 14464 9998 14516 10004
rect 14554 10024 14610 10033
rect 14476 9722 14504 9998
rect 14554 9959 14610 9968
rect 14464 9716 14516 9722
rect 14464 9658 14516 9664
rect 14556 9376 14608 9382
rect 14556 9318 14608 9324
rect 14568 9110 14596 9318
rect 14556 9104 14608 9110
rect 14556 9046 14608 9052
rect 14660 8616 14688 13194
rect 14752 12617 14780 16374
rect 14844 15162 14872 17070
rect 15028 16658 15056 18634
rect 15108 18420 15160 18426
rect 15212 18408 15240 19887
rect 15292 19858 15344 19864
rect 15304 19689 15332 19858
rect 15290 19680 15346 19689
rect 15290 19615 15346 19624
rect 15304 19378 15332 19615
rect 15292 19372 15344 19378
rect 15292 19314 15344 19320
rect 15292 18624 15344 18630
rect 15292 18566 15344 18572
rect 15396 18578 15424 21286
rect 15488 20466 15516 22510
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15580 20369 15608 22879
rect 15672 20874 15700 24375
rect 15764 23798 15792 26200
rect 15844 25016 15896 25022
rect 15844 24958 15896 24964
rect 15752 23792 15804 23798
rect 15752 23734 15804 23740
rect 15856 23361 15884 24958
rect 15936 23792 15988 23798
rect 15936 23734 15988 23740
rect 15842 23352 15898 23361
rect 15842 23287 15898 23296
rect 15948 22094 15976 23734
rect 16132 22710 16160 26302
rect 16394 26200 16450 26302
rect 16212 25628 16264 25634
rect 16212 25570 16264 25576
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16120 22500 16172 22506
rect 16120 22442 16172 22448
rect 15856 22066 15976 22094
rect 15752 21480 15804 21486
rect 15752 21422 15804 21428
rect 15764 21146 15792 21422
rect 15752 21140 15804 21146
rect 15752 21082 15804 21088
rect 15856 20992 15884 22066
rect 15934 21720 15990 21729
rect 15934 21655 15990 21664
rect 15948 21554 15976 21655
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16132 21486 16160 22442
rect 16224 22114 16252 25570
rect 16396 25152 16448 25158
rect 16396 25094 16448 25100
rect 16304 24744 16356 24750
rect 16304 24686 16356 24692
rect 16316 24562 16344 24686
rect 16408 24664 16436 25094
rect 16488 25016 16540 25022
rect 16488 24958 16540 24964
rect 16500 24857 16528 24958
rect 16486 24848 16542 24857
rect 16486 24783 16542 24792
rect 16408 24636 16620 24664
rect 16316 24534 16528 24562
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16316 22234 16344 23802
rect 16394 23624 16450 23633
rect 16394 23559 16450 23568
rect 16304 22228 16356 22234
rect 16304 22170 16356 22176
rect 16224 22086 16344 22114
rect 16212 21888 16264 21894
rect 16212 21830 16264 21836
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 15764 20964 15884 20992
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15566 20360 15622 20369
rect 15566 20295 15622 20304
rect 15660 20256 15712 20262
rect 15660 20198 15712 20204
rect 15672 19922 15700 20198
rect 15660 19916 15712 19922
rect 15660 19858 15712 19864
rect 15764 19802 15792 20964
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 15844 20868 15896 20874
rect 15844 20810 15896 20816
rect 15580 19774 15792 19802
rect 15476 19712 15528 19718
rect 15476 19654 15528 19660
rect 15488 18698 15516 19654
rect 15476 18692 15528 18698
rect 15476 18634 15528 18640
rect 15160 18380 15240 18408
rect 15108 18362 15160 18368
rect 15304 18290 15332 18566
rect 15396 18550 15516 18578
rect 15200 18284 15252 18290
rect 15200 18226 15252 18232
rect 15292 18284 15344 18290
rect 15292 18226 15344 18232
rect 15106 17776 15162 17785
rect 15106 17711 15162 17720
rect 15120 17270 15148 17711
rect 15212 17377 15240 18226
rect 15384 18216 15436 18222
rect 15382 18184 15384 18193
rect 15436 18184 15438 18193
rect 15382 18119 15438 18128
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15198 17368 15254 17377
rect 15198 17303 15254 17312
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 14924 16516 14976 16522
rect 14924 16458 14976 16464
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 14936 13938 14964 16458
rect 15304 16454 15332 17818
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15396 16833 15424 17002
rect 15382 16824 15438 16833
rect 15382 16759 15438 16768
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 15028 15706 15056 15914
rect 15016 15700 15068 15706
rect 15016 15642 15068 15648
rect 15028 14958 15056 15642
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 15028 13394 15056 13806
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15016 13388 15068 13394
rect 15016 13330 15068 13336
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14738 12608 14794 12617
rect 14738 12543 14794 12552
rect 14740 12436 14792 12442
rect 14740 12378 14792 12384
rect 14752 10606 14780 12378
rect 14844 11014 14872 12854
rect 14936 12306 14964 13330
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14936 11626 14964 11698
rect 14924 11620 14976 11626
rect 14924 11562 14976 11568
rect 14922 11248 14978 11257
rect 14922 11183 14978 11192
rect 14936 11082 14964 11183
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9994 14780 10406
rect 14740 9988 14792 9994
rect 14740 9930 14792 9936
rect 14844 9926 14872 10950
rect 14832 9920 14884 9926
rect 14832 9862 14884 9868
rect 14740 9648 14792 9654
rect 14738 9616 14740 9625
rect 14792 9616 14794 9625
rect 14738 9551 14794 9560
rect 14660 8588 14780 8616
rect 14646 8528 14702 8537
rect 14556 8492 14608 8498
rect 14646 8463 14648 8472
rect 14556 8434 14608 8440
rect 14700 8463 14702 8472
rect 14648 8434 14700 8440
rect 14568 6866 14596 8434
rect 14752 6934 14780 8588
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14556 6860 14608 6866
rect 14556 6802 14608 6808
rect 14844 6118 14872 9862
rect 14922 9208 14978 9217
rect 14922 9143 14978 9152
rect 14936 9042 14964 9143
rect 15028 9058 15056 12038
rect 15120 10470 15148 15370
rect 15212 13938 15240 16050
rect 15488 14657 15516 18550
rect 15580 16794 15608 19774
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 15672 19145 15700 19654
rect 15658 19136 15714 19145
rect 15658 19071 15714 19080
rect 15672 17202 15700 19071
rect 15856 18850 15884 20810
rect 16132 20806 16160 20878
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16132 20505 16160 20742
rect 16118 20496 16174 20505
rect 16118 20431 16174 20440
rect 16224 20448 16252 21830
rect 16316 21729 16344 22086
rect 16302 21720 16358 21729
rect 16302 21655 16358 21664
rect 16304 21344 16356 21350
rect 16302 21312 16304 21321
rect 16356 21312 16358 21321
rect 16302 21247 16358 21256
rect 16316 21010 16344 21247
rect 16408 21078 16436 23559
rect 16500 23497 16528 24534
rect 16486 23488 16542 23497
rect 16486 23423 16542 23432
rect 16592 22794 16620 24636
rect 16868 24614 16896 26522
rect 17038 26200 17094 26574
rect 17224 26512 17276 26518
rect 17224 26454 17276 26460
rect 17040 25628 17092 25634
rect 17040 25570 17092 25576
rect 16948 25288 17000 25294
rect 16948 25230 17000 25236
rect 16960 25090 16988 25230
rect 16948 25084 17000 25090
rect 16948 25026 17000 25032
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16948 24608 17000 24614
rect 16948 24550 17000 24556
rect 16960 24426 16988 24550
rect 16672 24404 16724 24410
rect 16672 24346 16724 24352
rect 16868 24398 16988 24426
rect 16684 23905 16712 24346
rect 16868 24342 16896 24398
rect 16856 24336 16908 24342
rect 16856 24278 16908 24284
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 16764 24132 16816 24138
rect 16764 24074 16816 24080
rect 16670 23896 16726 23905
rect 16670 23831 16726 23840
rect 16500 22766 16620 22794
rect 16500 22114 16528 22766
rect 16580 22636 16632 22642
rect 16580 22578 16632 22584
rect 16592 22234 16620 22578
rect 16670 22264 16726 22273
rect 16580 22228 16632 22234
rect 16670 22199 16726 22208
rect 16580 22170 16632 22176
rect 16500 22086 16620 22114
rect 16592 22001 16620 22086
rect 16578 21992 16634 22001
rect 16578 21927 16634 21936
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16396 21072 16448 21078
rect 16396 21014 16448 21020
rect 16304 21004 16356 21010
rect 16304 20946 16356 20952
rect 16500 20924 16528 21490
rect 16580 21140 16632 21146
rect 16580 21082 16632 21088
rect 16592 20942 16620 21082
rect 16408 20896 16528 20924
rect 16580 20936 16632 20942
rect 16408 20534 16436 20896
rect 16580 20878 16632 20884
rect 16684 20754 16712 22199
rect 16776 22166 16804 24074
rect 16868 23186 16896 24142
rect 17052 23905 17080 25570
rect 17132 24608 17184 24614
rect 17132 24550 17184 24556
rect 17038 23896 17094 23905
rect 17038 23831 17094 23840
rect 17038 23760 17094 23769
rect 17038 23695 17094 23704
rect 16856 23180 16908 23186
rect 16856 23122 16908 23128
rect 16868 22574 16896 23122
rect 16856 22568 16908 22574
rect 16856 22510 16908 22516
rect 16764 22160 16816 22166
rect 16762 22128 16764 22137
rect 16816 22128 16818 22137
rect 16868 22098 16896 22510
rect 16762 22063 16818 22072
rect 16856 22092 16908 22098
rect 16856 22034 16908 22040
rect 16764 21480 16816 21486
rect 16764 21422 16816 21428
rect 16776 20913 16804 21422
rect 16762 20904 16818 20913
rect 16868 20874 16896 22034
rect 16762 20839 16818 20848
rect 16856 20868 16908 20874
rect 16856 20810 16908 20816
rect 16500 20726 16712 20754
rect 16948 20800 17000 20806
rect 16948 20742 17000 20748
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16304 20460 16356 20466
rect 16224 20420 16304 20448
rect 16304 20402 16356 20408
rect 16500 20398 16528 20726
rect 16578 20632 16634 20641
rect 16578 20567 16634 20576
rect 16856 20596 16908 20602
rect 16488 20392 16540 20398
rect 16488 20334 16540 20340
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 16118 20224 16174 20233
rect 16118 20159 16174 20168
rect 16132 19310 16160 20159
rect 16302 19544 16358 19553
rect 16302 19479 16358 19488
rect 16316 19446 16344 19479
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 15936 19304 15988 19310
rect 15936 19246 15988 19252
rect 16028 19304 16080 19310
rect 16028 19246 16080 19252
rect 16120 19304 16172 19310
rect 16120 19246 16172 19252
rect 15764 18834 15884 18850
rect 15752 18828 15884 18834
rect 15804 18822 15884 18828
rect 15752 18770 15804 18776
rect 15752 18624 15804 18630
rect 15752 18566 15804 18572
rect 15764 18222 15792 18566
rect 15752 18216 15804 18222
rect 15752 18158 15804 18164
rect 15750 18048 15806 18057
rect 15750 17983 15806 17992
rect 15764 17490 15792 17983
rect 15856 17746 15884 18822
rect 15844 17740 15896 17746
rect 15844 17682 15896 17688
rect 15844 17604 15896 17610
rect 15948 17592 15976 19246
rect 16040 18329 16068 19246
rect 16118 19000 16174 19009
rect 16118 18935 16174 18944
rect 16132 18601 16160 18935
rect 16224 18902 16252 19382
rect 16212 18896 16264 18902
rect 16212 18838 16264 18844
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 16118 18592 16174 18601
rect 16118 18527 16174 18536
rect 16026 18320 16082 18329
rect 16132 18290 16160 18527
rect 16026 18255 16082 18264
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16132 17728 16160 18226
rect 16224 18057 16252 18226
rect 16210 18048 16266 18057
rect 16210 17983 16266 17992
rect 16316 17882 16344 18634
rect 16408 18601 16436 20266
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16500 20097 16528 20198
rect 16486 20088 16542 20097
rect 16486 20023 16542 20032
rect 16486 19408 16542 19417
rect 16486 19343 16542 19352
rect 16394 18592 16450 18601
rect 16394 18527 16450 18536
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 15896 17564 15976 17592
rect 16040 17700 16160 17728
rect 15844 17546 15896 17552
rect 15764 17462 15884 17490
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15566 15872 15622 15881
rect 15566 15807 15622 15816
rect 15474 14648 15530 14657
rect 15474 14583 15530 14592
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15290 14376 15346 14385
rect 15290 14311 15346 14320
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15212 12374 15240 12786
rect 15200 12368 15252 12374
rect 15200 12310 15252 12316
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15212 10742 15240 12106
rect 15304 11937 15332 14311
rect 15290 11928 15346 11937
rect 15290 11863 15346 11872
rect 15292 11824 15344 11830
rect 15292 11766 15344 11772
rect 15396 11778 15424 14418
rect 15580 13802 15608 15807
rect 15764 15706 15792 17070
rect 15856 16794 15884 17462
rect 16040 17218 16068 17700
rect 16120 17604 16172 17610
rect 16120 17546 16172 17552
rect 15948 17190 16068 17218
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15658 15464 15714 15473
rect 15658 15399 15660 15408
rect 15712 15399 15714 15408
rect 15660 15370 15712 15376
rect 15672 14346 15700 15370
rect 15764 15065 15792 15642
rect 15750 15056 15806 15065
rect 15750 14991 15806 15000
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15672 13326 15700 14282
rect 15856 14278 15884 16730
rect 15948 16590 15976 17190
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 15936 16584 15988 16590
rect 15936 16526 15988 16532
rect 15936 16040 15988 16046
rect 15936 15982 15988 15988
rect 15844 14272 15896 14278
rect 15844 14214 15896 14220
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15660 13320 15712 13326
rect 15660 13262 15712 13268
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15474 12064 15530 12073
rect 15474 11999 15530 12008
rect 15488 11898 15516 11999
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15304 11064 15332 11766
rect 15396 11750 15516 11778
rect 15384 11076 15436 11082
rect 15304 11036 15384 11064
rect 15384 11018 15436 11024
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15292 10260 15344 10266
rect 15292 10202 15344 10208
rect 14924 9036 14976 9042
rect 15028 9030 15240 9058
rect 14924 8978 14976 8984
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14936 7886 14964 8774
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 14568 5234 14596 6054
rect 14556 5228 14608 5234
rect 14556 5170 14608 5176
rect 14372 4820 14424 4826
rect 14372 4762 14424 4768
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14280 4208 14332 4214
rect 14280 4150 14332 4156
rect 14476 3346 14504 4490
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14554 3768 14610 3777
rect 14554 3703 14610 3712
rect 14568 3670 14596 3703
rect 14556 3664 14608 3670
rect 14556 3606 14608 3612
rect 14660 3534 14688 4082
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14476 3318 14688 3346
rect 14188 2848 14240 2854
rect 14188 2790 14240 2796
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14200 2582 14228 2790
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 14660 2514 14688 3318
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14200 1465 14228 2246
rect 14384 1562 14412 2246
rect 14372 1556 14424 1562
rect 14372 1498 14424 1504
rect 14186 1456 14242 1465
rect 14186 1391 14242 1400
rect 13636 1158 13688 1164
rect 13910 1184 13966 1193
rect 13910 1119 13966 1128
rect 14752 800 14780 4082
rect 14832 3120 14884 3126
rect 14830 3088 14832 3097
rect 14884 3088 14886 3097
rect 14830 3023 14886 3032
rect 14936 2564 14964 7822
rect 15120 7478 15148 8842
rect 15212 8022 15240 9030
rect 15200 8016 15252 8022
rect 15200 7958 15252 7964
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15212 7410 15240 7754
rect 15304 7546 15332 10202
rect 15396 9994 15424 11018
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9654 15424 9930
rect 15488 9926 15516 11750
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15384 8424 15436 8430
rect 15580 8412 15608 12582
rect 15660 12368 15712 12374
rect 15660 12310 15712 12316
rect 15672 11626 15700 12310
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15436 8384 15608 8412
rect 15384 8366 15436 8372
rect 15764 7886 15792 13806
rect 15842 13424 15898 13433
rect 15842 13359 15898 13368
rect 15856 12714 15884 13359
rect 15948 13172 15976 15982
rect 16040 15162 16068 17070
rect 16132 16697 16160 17546
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16118 16688 16174 16697
rect 16118 16623 16174 16632
rect 16120 16584 16172 16590
rect 16224 16561 16252 17070
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16304 16584 16356 16590
rect 16120 16526 16172 16532
rect 16210 16552 16266 16561
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16028 13184 16080 13190
rect 15948 13144 16028 13172
rect 16028 13126 16080 13132
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11937 15884 12038
rect 15842 11928 15898 11937
rect 15842 11863 15898 11872
rect 15948 11778 15976 12786
rect 16040 11898 16068 13126
rect 16028 11892 16080 11898
rect 16028 11834 16080 11840
rect 16132 11801 16160 16526
rect 16304 16526 16356 16532
rect 16210 16487 16266 16496
rect 16316 15994 16344 16526
rect 16224 15966 16344 15994
rect 16224 13161 16252 15966
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16316 15065 16344 15846
rect 16408 15638 16436 16594
rect 16396 15632 16448 15638
rect 16396 15574 16448 15580
rect 16500 15162 16528 19343
rect 16592 18970 16620 20567
rect 16856 20538 16908 20544
rect 16868 20233 16896 20538
rect 16960 20330 16988 20742
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 16854 20224 16910 20233
rect 16854 20159 16910 20168
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16776 19174 16804 19858
rect 16868 19689 16896 19994
rect 16948 19848 17000 19854
rect 16948 19790 17000 19796
rect 16854 19680 16910 19689
rect 16854 19615 16910 19624
rect 16960 19553 16988 19790
rect 16946 19544 17002 19553
rect 16946 19479 17002 19488
rect 17052 19334 17080 23695
rect 17144 22094 17172 24550
rect 17236 22982 17264 26454
rect 17224 22976 17276 22982
rect 17224 22918 17276 22924
rect 17236 22710 17264 22918
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17144 22066 17264 22094
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17144 21457 17172 21490
rect 17130 21448 17186 21457
rect 17130 21383 17186 21392
rect 17130 21176 17186 21185
rect 17130 21111 17186 21120
rect 17144 20233 17172 21111
rect 17236 20913 17264 22066
rect 17328 21486 17356 26574
rect 17682 26200 17738 27000
rect 17776 26580 17828 26586
rect 17776 26522 17828 26528
rect 17592 26104 17644 26110
rect 17592 26046 17644 26052
rect 17500 25424 17552 25430
rect 17500 25366 17552 25372
rect 17512 22234 17540 25366
rect 17604 23798 17632 26046
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17696 23050 17724 26200
rect 17788 23186 17816 26522
rect 18326 26200 18382 27000
rect 18880 26444 18932 26450
rect 18880 26386 18932 26392
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 17880 24750 17908 25842
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 17960 24880 18012 24886
rect 17960 24822 18012 24828
rect 17868 24744 17920 24750
rect 17868 24686 17920 24692
rect 17972 24614 18000 24822
rect 17960 24608 18012 24614
rect 17960 24550 18012 24556
rect 18156 24342 18184 24890
rect 18144 24336 18196 24342
rect 18144 24278 18196 24284
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23848 17908 24006
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17880 23820 18000 23848
rect 17776 23180 17828 23186
rect 17776 23122 17828 23128
rect 17972 23089 18000 23820
rect 18340 23662 18368 26200
rect 18696 25356 18748 25362
rect 18696 25298 18748 25304
rect 18512 24880 18564 24886
rect 18512 24822 18564 24828
rect 18420 24132 18472 24138
rect 18420 24074 18472 24080
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18236 23588 18288 23594
rect 18236 23530 18288 23536
rect 17958 23080 18014 23089
rect 17684 23044 17736 23050
rect 17958 23015 18014 23024
rect 18248 23032 18276 23530
rect 18432 23050 18460 24074
rect 18524 23730 18552 24822
rect 18602 24712 18658 24721
rect 18602 24647 18658 24656
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18420 23044 18472 23050
rect 18248 23004 18368 23032
rect 17684 22986 17736 22992
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17500 22228 17552 22234
rect 17500 22170 17552 22176
rect 17960 22228 18012 22234
rect 17960 22170 18012 22176
rect 17500 22092 17552 22098
rect 17972 22094 18000 22170
rect 17500 22034 17552 22040
rect 17696 22066 18000 22094
rect 18052 22092 18104 22098
rect 17406 21856 17462 21865
rect 17406 21791 17462 21800
rect 17316 21480 17368 21486
rect 17316 21422 17368 21428
rect 17316 21072 17368 21078
rect 17316 21014 17368 21020
rect 17222 20904 17278 20913
rect 17222 20839 17278 20848
rect 17328 20602 17356 21014
rect 17420 20942 17448 21791
rect 17512 21486 17540 22034
rect 17696 21962 17724 22066
rect 18052 22034 18104 22040
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17592 21888 17644 21894
rect 18064 21876 18092 22034
rect 17592 21830 17644 21836
rect 17880 21848 18092 21876
rect 17500 21480 17552 21486
rect 17500 21422 17552 21428
rect 17500 21004 17552 21010
rect 17500 20946 17552 20952
rect 17408 20936 17460 20942
rect 17408 20878 17460 20884
rect 17408 20800 17460 20806
rect 17406 20768 17408 20777
rect 17460 20768 17462 20777
rect 17406 20703 17462 20712
rect 17316 20596 17368 20602
rect 17316 20538 17368 20544
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17130 20224 17186 20233
rect 17130 20159 17186 20168
rect 17236 20097 17264 20402
rect 17408 20324 17460 20330
rect 17408 20266 17460 20272
rect 17222 20088 17278 20097
rect 17222 20023 17278 20032
rect 17420 19854 17448 20266
rect 17316 19848 17368 19854
rect 16868 19306 17080 19334
rect 17236 19808 17316 19836
rect 17236 19334 17264 19808
rect 17316 19790 17368 19796
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17512 19802 17540 20946
rect 17604 20602 17632 21830
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17682 20632 17738 20641
rect 17592 20596 17644 20602
rect 17682 20567 17738 20576
rect 17592 20538 17644 20544
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17604 20058 17632 20402
rect 17696 20262 17724 20567
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 17682 20088 17738 20097
rect 17592 20052 17644 20058
rect 17788 20058 17816 21490
rect 17880 21078 17908 21848
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17958 21448 18014 21457
rect 17958 21383 17960 21392
rect 18012 21383 18014 21392
rect 17960 21354 18012 21360
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 18340 20534 18368 23004
rect 18420 22986 18472 22992
rect 18432 22710 18460 22986
rect 18616 22930 18644 24647
rect 18708 23594 18736 25298
rect 18786 24304 18842 24313
rect 18786 24239 18842 24248
rect 18800 24070 18828 24239
rect 18788 24064 18840 24070
rect 18786 24032 18788 24041
rect 18840 24032 18842 24041
rect 18786 23967 18842 23976
rect 18788 23656 18840 23662
rect 18788 23598 18840 23604
rect 18696 23588 18748 23594
rect 18696 23530 18748 23536
rect 18800 23526 18828 23598
rect 18788 23520 18840 23526
rect 18892 23508 18920 26386
rect 18970 26200 19026 27000
rect 19064 26444 19116 26450
rect 19064 26386 19116 26392
rect 18984 24274 19012 26200
rect 19076 26178 19104 26386
rect 19352 26302 19564 26330
rect 19064 26172 19116 26178
rect 19064 26114 19116 26120
rect 19352 24290 19380 26302
rect 19536 26160 19564 26302
rect 19614 26200 19670 27000
rect 19708 26920 19760 26926
rect 19708 26862 19760 26868
rect 19628 26160 19656 26200
rect 19536 26132 19656 26160
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 19168 24262 19380 24290
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 19076 23866 19104 24006
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 18984 23610 19012 23802
rect 19168 23798 19196 24262
rect 19616 24200 19668 24206
rect 19616 24142 19668 24148
rect 19524 24132 19576 24138
rect 19524 24074 19576 24080
rect 19536 23798 19564 24074
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19156 23656 19208 23662
rect 18984 23604 19156 23610
rect 18984 23598 19208 23604
rect 18984 23582 19196 23598
rect 18892 23480 19288 23508
rect 18788 23462 18840 23468
rect 19062 23352 19118 23361
rect 19062 23287 19118 23296
rect 18524 22902 18644 22930
rect 18972 22976 19024 22982
rect 18972 22918 19024 22924
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18432 21622 18460 22646
rect 18420 21616 18472 21622
rect 18420 21558 18472 21564
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18432 20777 18460 20878
rect 18418 20768 18474 20777
rect 18418 20703 18474 20712
rect 18144 20528 18196 20534
rect 18144 20470 18196 20476
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17868 20324 17920 20330
rect 17868 20266 17920 20272
rect 17682 20023 17738 20032
rect 17776 20052 17828 20058
rect 17592 19994 17644 20000
rect 17696 19990 17724 20023
rect 17776 19994 17828 20000
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17880 19922 17908 20266
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17512 19786 17816 19802
rect 17512 19780 17828 19786
rect 17512 19774 17776 19780
rect 17408 19712 17460 19718
rect 17408 19654 17460 19660
rect 17236 19306 17356 19334
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16580 18828 16632 18834
rect 16580 18770 16632 18776
rect 16592 18329 16620 18770
rect 16578 18320 16634 18329
rect 16578 18255 16634 18264
rect 16580 18216 16632 18222
rect 16580 18158 16632 18164
rect 16592 17882 16620 18158
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16302 15056 16358 15065
rect 16592 15026 16620 17818
rect 16684 15706 16712 19110
rect 16762 18864 16818 18873
rect 16762 18799 16818 18808
rect 16776 18698 16804 18799
rect 16764 18692 16816 18698
rect 16764 18634 16816 18640
rect 16868 18578 16896 19306
rect 17038 19136 17094 19145
rect 17038 19071 17094 19080
rect 17052 18766 17080 19071
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17130 18864 17186 18873
rect 17130 18799 17186 18808
rect 17040 18760 17092 18766
rect 17040 18702 17092 18708
rect 16776 18550 16896 18578
rect 16776 18154 16804 18550
rect 16854 18456 16910 18465
rect 16854 18391 16910 18400
rect 16764 18148 16816 18154
rect 16764 18090 16816 18096
rect 16868 17542 16896 18391
rect 17144 18290 17172 18799
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17132 18148 17184 18154
rect 17132 18090 17184 18096
rect 17038 18048 17094 18057
rect 17038 17983 17094 17992
rect 16856 17536 16908 17542
rect 16856 17478 16908 17484
rect 16868 17218 16896 17478
rect 16868 17202 16988 17218
rect 16868 17196 17000 17202
rect 16868 17190 16948 17196
rect 16948 17138 17000 17144
rect 16764 16992 16816 16998
rect 16764 16934 16816 16940
rect 16856 16992 16908 16998
rect 16856 16934 16908 16940
rect 16672 15700 16724 15706
rect 16672 15642 16724 15648
rect 16670 15600 16726 15609
rect 16670 15535 16726 15544
rect 16302 14991 16358 15000
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16684 14929 16712 15535
rect 16776 15366 16804 16934
rect 16868 16726 16896 16934
rect 16856 16720 16908 16726
rect 16856 16662 16908 16668
rect 16856 16040 16908 16046
rect 16908 16000 16988 16028
rect 16856 15982 16908 15988
rect 16854 15600 16910 15609
rect 16854 15535 16910 15544
rect 16868 15434 16896 15535
rect 16960 15502 16988 16000
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16856 15428 16908 15434
rect 16856 15370 16908 15376
rect 16764 15360 16816 15366
rect 16764 15302 16816 15308
rect 16854 15328 16910 15337
rect 16854 15263 16910 15272
rect 16764 15156 16816 15162
rect 16764 15098 16816 15104
rect 16486 14920 16542 14929
rect 16670 14920 16726 14929
rect 16542 14878 16620 14906
rect 16486 14855 16542 14864
rect 16302 14512 16358 14521
rect 16302 14447 16358 14456
rect 16316 13682 16344 14447
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16486 14240 16542 14249
rect 16408 13870 16436 14214
rect 16486 14175 16542 14184
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 16316 13654 16436 13682
rect 16302 13560 16358 13569
rect 16302 13495 16304 13504
rect 16356 13495 16358 13504
rect 16304 13466 16356 13472
rect 16210 13152 16266 13161
rect 16210 13087 16266 13096
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16224 12050 16252 12718
rect 16316 12617 16344 13466
rect 16302 12608 16358 12617
rect 16302 12543 16358 12552
rect 16408 12434 16436 13654
rect 16500 13530 16528 14175
rect 16592 13954 16620 14878
rect 16670 14855 16726 14864
rect 16670 14104 16726 14113
rect 16670 14039 16672 14048
rect 16724 14039 16726 14048
rect 16672 14010 16724 14016
rect 16592 13926 16712 13954
rect 16684 13705 16712 13926
rect 16670 13696 16726 13705
rect 16670 13631 16726 13640
rect 16578 13560 16634 13569
rect 16488 13524 16540 13530
rect 16776 13546 16804 15098
rect 16868 13569 16896 15263
rect 16960 14482 16988 15438
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16684 13530 16804 13546
rect 16578 13495 16634 13504
rect 16672 13524 16804 13530
rect 16488 13466 16540 13472
rect 16592 13410 16620 13495
rect 16724 13518 16804 13524
rect 16854 13560 16910 13569
rect 16854 13495 16910 13504
rect 16672 13466 16724 13472
rect 16500 13382 16620 13410
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16672 13388 16724 13394
rect 16500 13258 16528 13382
rect 16672 13330 16724 13336
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16486 13152 16542 13161
rect 16486 13087 16542 13096
rect 16500 12986 16528 13087
rect 16488 12980 16540 12986
rect 16488 12922 16540 12928
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16500 12646 16528 12718
rect 16488 12640 16540 12646
rect 16488 12582 16540 12588
rect 16408 12406 16528 12434
rect 16500 12345 16528 12406
rect 16486 12336 16542 12345
rect 16486 12271 16542 12280
rect 16403 12164 16455 12170
rect 16455 12124 16528 12152
rect 16403 12106 16455 12112
rect 16224 12022 16436 12050
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16304 11892 16356 11898
rect 16304 11834 16356 11840
rect 16118 11792 16174 11801
rect 15844 11756 15896 11762
rect 15948 11750 16068 11778
rect 15844 11698 15896 11704
rect 15856 10266 15884 11698
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 10674 15976 11630
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15936 10532 15988 10538
rect 15936 10474 15988 10480
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 10198 15976 10474
rect 15936 10192 15988 10198
rect 15936 10134 15988 10140
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15856 9178 15884 9386
rect 15844 9172 15896 9178
rect 15844 9114 15896 9120
rect 15948 8922 15976 10134
rect 16040 9450 16068 11750
rect 16118 11727 16174 11736
rect 16120 11212 16172 11218
rect 16120 11154 16172 11160
rect 16028 9444 16080 9450
rect 16028 9386 16080 9392
rect 15856 8894 15976 8922
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15752 7880 15804 7886
rect 15752 7822 15804 7828
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15292 7540 15344 7546
rect 15292 7482 15344 7488
rect 15672 7410 15700 7686
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15384 7336 15436 7342
rect 15384 7278 15436 7284
rect 15200 6792 15252 6798
rect 15198 6760 15200 6769
rect 15252 6760 15254 6769
rect 15198 6695 15254 6704
rect 15200 6656 15252 6662
rect 15200 6598 15252 6604
rect 15108 5568 15160 5574
rect 15108 5510 15160 5516
rect 15120 4826 15148 5510
rect 15212 5370 15240 6598
rect 15292 5772 15344 5778
rect 15292 5714 15344 5720
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15304 4146 15332 5714
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15014 4040 15070 4049
rect 15014 3975 15070 3984
rect 15028 3126 15056 3975
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 3641 15332 3878
rect 15396 3670 15424 7278
rect 15660 7200 15712 7206
rect 15660 7142 15712 7148
rect 15476 6792 15528 6798
rect 15474 6760 15476 6769
rect 15528 6760 15530 6769
rect 15474 6695 15530 6704
rect 15672 6322 15700 7142
rect 15856 7002 15884 8894
rect 16040 8838 16068 8910
rect 15936 8832 15988 8838
rect 15936 8774 15988 8780
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15948 7954 15976 8774
rect 16132 8344 16160 11154
rect 16040 8316 16160 8344
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 15750 6624 15806 6633
rect 15750 6559 15806 6568
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15660 5092 15712 5098
rect 15660 5034 15712 5040
rect 15672 4690 15700 5034
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15488 3942 15516 4082
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15384 3664 15436 3670
rect 15290 3632 15346 3641
rect 15384 3606 15436 3612
rect 15290 3567 15346 3576
rect 15108 3460 15160 3466
rect 15108 3402 15160 3408
rect 15120 3194 15148 3402
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15384 2848 15436 2854
rect 15384 2790 15436 2796
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15016 2576 15068 2582
rect 14936 2536 15016 2564
rect 15016 2518 15068 2524
rect 15212 2446 15240 2586
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15212 1193 15240 2042
rect 15396 1902 15424 2790
rect 15384 1896 15436 1902
rect 15384 1838 15436 1844
rect 15198 1184 15254 1193
rect 15198 1119 15254 1128
rect 6644 750 6696 756
rect 6368 740 6420 746
rect 6368 682 6420 688
rect 5908 196 5960 202
rect 5908 138 5960 144
rect 6734 0 6790 800
rect 9402 0 9458 800
rect 12070 0 12126 800
rect 14738 0 14794 800
rect 15488 474 15516 3878
rect 15764 3670 15792 6559
rect 15856 5234 15884 6938
rect 15948 6866 15976 6938
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 16040 6730 16068 8316
rect 16118 8256 16174 8265
rect 16118 8191 16174 8200
rect 16132 7954 16160 8191
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 15934 5808 15990 5817
rect 15934 5743 15990 5752
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15948 3670 15976 5743
rect 16132 3942 16160 7278
rect 16224 6390 16252 11834
rect 16316 7698 16344 11834
rect 16408 11762 16436 12022
rect 16396 11756 16448 11762
rect 16396 11698 16448 11704
rect 16394 11384 16450 11393
rect 16394 11319 16450 11328
rect 16408 8673 16436 11319
rect 16500 9674 16528 12124
rect 16592 12102 16620 13194
rect 16684 12102 16712 13330
rect 16776 12918 16804 13398
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16764 12912 16816 12918
rect 16764 12854 16816 12860
rect 16868 12306 16896 13330
rect 16960 12986 16988 14282
rect 17052 13938 17080 17983
rect 17144 17270 17172 18090
rect 17236 17882 17264 18906
rect 17224 17876 17276 17882
rect 17224 17818 17276 17824
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17224 17264 17276 17270
rect 17224 17206 17276 17212
rect 17132 16720 17184 16726
rect 17132 16662 17184 16668
rect 17144 16289 17172 16662
rect 17130 16280 17186 16289
rect 17130 16215 17186 16224
rect 17236 16182 17264 17206
rect 17224 16176 17276 16182
rect 17224 16118 17276 16124
rect 17132 16040 17184 16046
rect 17132 15982 17184 15988
rect 17144 15473 17172 15982
rect 17130 15464 17186 15473
rect 17130 15399 17186 15408
rect 17328 15162 17356 19306
rect 17420 17678 17448 19654
rect 17498 19544 17554 19553
rect 17498 19479 17554 19488
rect 17512 19310 17540 19479
rect 17604 19378 17632 19774
rect 17776 19722 17828 19728
rect 17972 19700 18000 20334
rect 18156 20330 18184 20470
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18524 20262 18552 22902
rect 18604 22772 18656 22778
rect 18604 22714 18656 22720
rect 18616 21010 18644 22714
rect 18694 22128 18750 22137
rect 18694 22063 18750 22072
rect 18708 21729 18736 22063
rect 18694 21720 18750 21729
rect 18694 21655 18750 21664
rect 18880 21616 18932 21622
rect 18878 21584 18880 21593
rect 18932 21584 18934 21593
rect 18878 21519 18934 21528
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18984 20942 19012 22918
rect 19076 21622 19104 23287
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 19064 21480 19116 21486
rect 19168 21457 19196 21830
rect 19064 21422 19116 21428
rect 19154 21448 19210 21457
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 19076 20874 19104 21422
rect 19154 21383 19210 21392
rect 19154 21176 19210 21185
rect 19154 21111 19210 21120
rect 19064 20868 19116 20874
rect 19064 20810 19116 20816
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 17880 19672 18000 19700
rect 18512 19712 18564 19718
rect 18510 19680 18512 19689
rect 18564 19680 18566 19689
rect 17880 19666 17908 19672
rect 17788 19638 17908 19666
rect 17788 19553 17816 19638
rect 17950 19612 18258 19621
rect 18510 19615 18566 19624
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17774 19544 17830 19553
rect 17950 19547 18258 19556
rect 18616 19553 18644 20402
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 17774 19479 17830 19488
rect 18602 19544 18658 19553
rect 18800 19514 18828 20334
rect 18602 19479 18658 19488
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 17776 19440 17828 19446
rect 17774 19408 17776 19417
rect 17828 19408 17830 19417
rect 17592 19372 17644 19378
rect 17774 19343 17830 19352
rect 18340 19378 18460 19394
rect 18340 19372 18472 19378
rect 18340 19366 18420 19372
rect 17592 19314 17644 19320
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17960 19304 18012 19310
rect 18236 19304 18288 19310
rect 18012 19264 18236 19292
rect 17960 19246 18012 19252
rect 18236 19246 18288 19252
rect 17696 19122 17724 19246
rect 17604 19094 17724 19122
rect 17868 19168 17920 19174
rect 17920 19128 18000 19156
rect 17868 19110 17920 19116
rect 17972 19122 18000 19128
rect 18340 19122 18368 19366
rect 18420 19314 18472 19320
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18696 19236 18748 19242
rect 18696 19178 18748 19184
rect 17972 19094 18368 19122
rect 18602 19136 18658 19145
rect 17500 18896 17552 18902
rect 17500 18838 17552 18844
rect 17512 18329 17540 18838
rect 17604 18601 17632 19094
rect 18602 19071 18658 19080
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 18156 18924 18552 18952
rect 17590 18592 17646 18601
rect 17590 18527 17646 18536
rect 17696 18465 17724 18906
rect 18050 18864 18106 18873
rect 17776 18828 17828 18834
rect 18156 18850 18184 18924
rect 18106 18834 18184 18850
rect 18234 18864 18290 18873
rect 18106 18828 18196 18834
rect 18106 18822 18144 18828
rect 18050 18799 18106 18808
rect 17776 18770 17828 18776
rect 18234 18799 18290 18808
rect 18144 18770 18196 18776
rect 17682 18456 17738 18465
rect 17682 18391 17738 18400
rect 17788 18340 17816 18770
rect 17868 18692 17920 18698
rect 17868 18634 17920 18640
rect 17880 18408 17908 18634
rect 18248 18630 18276 18799
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17880 18380 18000 18408
rect 17498 18320 17554 18329
rect 17498 18255 17554 18264
rect 17696 18312 17816 18340
rect 17972 18329 18000 18380
rect 17958 18320 18014 18329
rect 17696 17814 17724 18312
rect 17868 18284 17920 18290
rect 17958 18255 18014 18264
rect 18144 18284 18196 18290
rect 17868 18226 17920 18232
rect 18144 18226 18196 18232
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 17776 17740 17828 17746
rect 17776 17682 17828 17688
rect 17408 17672 17460 17678
rect 17408 17614 17460 17620
rect 17500 17604 17552 17610
rect 17500 17546 17552 17552
rect 17512 17338 17540 17546
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17512 16504 17540 17274
rect 17604 17066 17632 17478
rect 17592 17060 17644 17066
rect 17592 17002 17644 17008
rect 17788 16697 17816 17682
rect 17880 17610 17908 18226
rect 18156 17814 18184 18226
rect 18432 18086 18460 18566
rect 18524 18465 18552 18924
rect 18510 18456 18566 18465
rect 18510 18391 18566 18400
rect 18420 18080 18472 18086
rect 18420 18022 18472 18028
rect 18420 17876 18472 17882
rect 18420 17818 18472 17824
rect 18144 17808 18196 17814
rect 18144 17750 18196 17756
rect 18144 17672 18196 17678
rect 18196 17632 18368 17660
rect 18144 17614 18196 17620
rect 17868 17604 17920 17610
rect 17868 17546 17920 17552
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 18340 17338 18368 17632
rect 18432 17354 18460 17818
rect 18616 17513 18644 19071
rect 18708 17954 18736 19178
rect 18800 18873 18828 19246
rect 18786 18864 18842 18873
rect 18786 18799 18842 18808
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18800 18057 18828 18566
rect 18786 18048 18842 18057
rect 18786 17983 18842 17992
rect 18708 17926 18828 17954
rect 18602 17504 18658 17513
rect 18602 17439 18658 17448
rect 18328 17332 18380 17338
rect 18432 17326 18644 17354
rect 18328 17274 18380 17280
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17774 16688 17830 16697
rect 17774 16623 17830 16632
rect 17880 16590 17908 17206
rect 18510 16960 18566 16969
rect 18510 16895 18566 16904
rect 18418 16824 18474 16833
rect 18418 16759 18474 16768
rect 17868 16584 17920 16590
rect 17868 16526 17920 16532
rect 17684 16516 17736 16522
rect 17512 16476 17684 16504
rect 17684 16458 17736 16464
rect 17406 16416 17462 16425
rect 17406 16351 17462 16360
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 17420 14929 17448 16351
rect 17590 16280 17646 16289
rect 17590 16215 17646 16224
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17130 14920 17186 14929
rect 17406 14920 17462 14929
rect 17130 14855 17132 14864
rect 17184 14855 17186 14864
rect 17328 14878 17406 14906
rect 17132 14826 17184 14832
rect 17328 14346 17356 14878
rect 17406 14855 17462 14864
rect 17316 14340 17368 14346
rect 17316 14282 17368 14288
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 12442 16988 12582
rect 17052 12442 17080 13466
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16856 12164 16908 12170
rect 16856 12106 16908 12112
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11892 16632 11898
rect 16684 11880 16712 12038
rect 16632 11852 16712 11880
rect 16580 11834 16632 11840
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16672 11552 16724 11558
rect 16672 11494 16724 11500
rect 16500 9646 16620 9674
rect 16486 9208 16542 9217
rect 16486 9143 16542 9152
rect 16500 9042 16528 9143
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16394 8664 16450 8673
rect 16394 8599 16450 8608
rect 16396 8288 16448 8294
rect 16396 8230 16448 8236
rect 16408 7886 16436 8230
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16488 7812 16540 7818
rect 16488 7754 16540 7760
rect 16316 7670 16436 7698
rect 16304 6928 16356 6934
rect 16304 6870 16356 6876
rect 16316 6390 16344 6870
rect 16408 6730 16436 7670
rect 16500 6866 16528 7754
rect 16592 6866 16620 9646
rect 16684 7410 16712 11494
rect 16776 11082 16804 11630
rect 16764 11076 16816 11082
rect 16764 11018 16816 11024
rect 16868 11014 16896 12106
rect 17040 11620 17092 11626
rect 17040 11562 17092 11568
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16960 11121 16988 11290
rect 16946 11112 17002 11121
rect 16946 11047 17002 11056
rect 16856 11008 16908 11014
rect 16908 10968 16988 10996
rect 16856 10950 16908 10956
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16764 10464 16816 10470
rect 16764 10406 16816 10412
rect 16776 8090 16804 10406
rect 16868 9722 16896 10678
rect 16960 10112 16988 10968
rect 17052 10470 17080 11562
rect 17040 10464 17092 10470
rect 17040 10406 17092 10412
rect 16960 10084 17080 10112
rect 16948 9988 17000 9994
rect 16948 9930 17000 9936
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16868 9518 16896 9658
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 8084 16816 8090
rect 16764 8026 16816 8032
rect 16762 7576 16818 7585
rect 16762 7511 16764 7520
rect 16816 7511 16818 7520
rect 16764 7482 16816 7488
rect 16672 7404 16724 7410
rect 16672 7346 16724 7352
rect 16672 7268 16724 7274
rect 16672 7210 16724 7216
rect 16488 6860 16540 6866
rect 16488 6802 16540 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16684 6497 16712 7210
rect 16764 6792 16816 6798
rect 16764 6734 16816 6740
rect 16670 6488 16726 6497
rect 16776 6458 16804 6734
rect 16670 6423 16726 6432
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16212 6384 16264 6390
rect 16212 6326 16264 6332
rect 16304 6384 16356 6390
rect 16304 6326 16356 6332
rect 16764 6248 16816 6254
rect 16764 6190 16816 6196
rect 16776 5216 16804 6190
rect 16868 5778 16896 9454
rect 16960 6390 16988 9930
rect 17052 9654 17080 10084
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 17144 9058 17172 14010
rect 17316 14000 17368 14006
rect 17236 13960 17316 13988
rect 17236 12458 17264 13960
rect 17316 13942 17368 13948
rect 17420 13682 17448 14282
rect 17512 14278 17540 15982
rect 17604 15609 17632 16215
rect 17696 16182 17724 16458
rect 18328 16448 18380 16454
rect 18328 16390 18380 16396
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17590 15600 17646 15609
rect 17590 15535 17646 15544
rect 17696 15434 17724 16118
rect 18340 15638 18368 16390
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17696 15337 17724 15370
rect 17682 15328 17738 15337
rect 17682 15263 17738 15272
rect 17696 14346 17724 15263
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 18432 15201 18460 16759
rect 18524 16454 18552 16895
rect 18512 16448 18564 16454
rect 18616 16425 18644 17326
rect 18694 16552 18750 16561
rect 18694 16487 18750 16496
rect 18512 16390 18564 16396
rect 18602 16416 18658 16425
rect 18524 16130 18552 16390
rect 18602 16351 18658 16360
rect 18602 16144 18658 16153
rect 18524 16102 18602 16130
rect 18602 16079 18658 16088
rect 18708 15366 18736 16487
rect 18800 15745 18828 17926
rect 18892 17610 18920 20742
rect 18970 20496 19026 20505
rect 18970 20431 18972 20440
rect 19024 20431 19026 20440
rect 18972 20402 19024 20408
rect 19076 20398 19104 20810
rect 19064 20392 19116 20398
rect 19064 20334 19116 20340
rect 18972 20324 19024 20330
rect 18972 20266 19024 20272
rect 18984 18465 19012 20266
rect 19168 20262 19196 21111
rect 19156 20256 19208 20262
rect 19156 20198 19208 20204
rect 19260 20058 19288 23480
rect 19628 22817 19656 24142
rect 19720 23905 19748 26862
rect 20076 26240 20128 26246
rect 20258 26200 20314 27000
rect 20536 26648 20588 26654
rect 20536 26590 20588 26596
rect 20076 26182 20128 26188
rect 19892 25152 19944 25158
rect 19892 25094 19944 25100
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19800 24608 19852 24614
rect 19800 24550 19852 24556
rect 19706 23896 19762 23905
rect 19706 23831 19762 23840
rect 19614 22808 19670 22817
rect 19614 22743 19670 22752
rect 19616 22568 19668 22574
rect 19616 22510 19668 22516
rect 19708 22568 19760 22574
rect 19708 22510 19760 22516
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 19444 22137 19472 22170
rect 19430 22128 19486 22137
rect 19628 22098 19656 22510
rect 19430 22063 19486 22072
rect 19616 22092 19668 22098
rect 19616 22034 19668 22040
rect 19432 21888 19484 21894
rect 19338 21856 19394 21865
rect 19616 21888 19668 21894
rect 19484 21848 19616 21876
rect 19432 21830 19484 21836
rect 19616 21830 19668 21836
rect 19338 21791 19394 21800
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19248 20052 19300 20058
rect 19248 19994 19300 20000
rect 19064 19916 19116 19922
rect 19064 19858 19116 19864
rect 19076 19417 19104 19858
rect 19168 19446 19196 19994
rect 19156 19440 19208 19446
rect 19062 19408 19118 19417
rect 19156 19382 19208 19388
rect 19062 19343 19118 19352
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 19154 18728 19210 18737
rect 18970 18456 19026 18465
rect 18970 18391 19026 18400
rect 18972 18284 19024 18290
rect 18972 18226 19024 18232
rect 18984 17678 19012 18226
rect 18972 17672 19024 17678
rect 18972 17614 19024 17620
rect 18880 17604 18932 17610
rect 18880 17546 18932 17552
rect 18970 16824 19026 16833
rect 18970 16759 19026 16768
rect 18984 16658 19012 16759
rect 18880 16652 18932 16658
rect 18880 16594 18932 16600
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18786 15736 18842 15745
rect 18786 15671 18842 15680
rect 18800 15570 18828 15671
rect 18788 15564 18840 15570
rect 18788 15506 18840 15512
rect 18512 15360 18564 15366
rect 18510 15328 18512 15337
rect 18696 15360 18748 15366
rect 18564 15328 18566 15337
rect 18510 15263 18566 15272
rect 18694 15328 18696 15337
rect 18748 15328 18750 15337
rect 18694 15263 18750 15272
rect 18418 15192 18474 15201
rect 18236 15156 18288 15162
rect 18418 15127 18474 15136
rect 18236 15098 18288 15104
rect 18248 14890 18276 15098
rect 18788 14952 18840 14958
rect 18788 14894 18840 14900
rect 18052 14884 18104 14890
rect 18052 14826 18104 14832
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18512 14884 18564 14890
rect 18512 14826 18564 14832
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17500 14272 17552 14278
rect 17500 14214 17552 14220
rect 17696 14006 17724 14282
rect 18064 14278 18092 14826
rect 18052 14272 18104 14278
rect 18524 14249 18552 14826
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18602 14512 18658 14521
rect 18602 14447 18658 14456
rect 18052 14214 18104 14220
rect 18510 14240 18566 14249
rect 17950 14172 18258 14181
rect 18510 14175 18566 14184
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 18052 14068 18104 14074
rect 17972 14028 18052 14056
rect 17684 14000 17736 14006
rect 17684 13942 17736 13948
rect 17972 13682 18000 14028
rect 18052 14010 18104 14016
rect 18616 13802 18644 14447
rect 18708 14414 18736 14758
rect 18800 14618 18828 14894
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18694 13832 18750 13841
rect 18604 13796 18656 13802
rect 18694 13767 18750 13776
rect 18604 13738 18656 13744
rect 18708 13734 18736 13767
rect 17328 13654 17448 13682
rect 17512 13654 18000 13682
rect 18144 13728 18196 13734
rect 18144 13670 18196 13676
rect 18696 13728 18748 13734
rect 18696 13670 18748 13676
rect 17328 13530 17356 13654
rect 17512 13546 17540 13654
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 17420 13518 17540 13546
rect 17316 13320 17368 13326
rect 17316 13262 17368 13268
rect 17328 12850 17356 13262
rect 17420 12968 17448 13518
rect 17592 13388 17644 13394
rect 17512 13348 17592 13376
rect 17512 13172 17540 13348
rect 18156 13376 18184 13670
rect 18708 13546 18736 13670
rect 18616 13518 18736 13546
rect 18512 13456 18564 13462
rect 18432 13416 18512 13444
rect 18236 13388 18288 13394
rect 18156 13348 18236 13376
rect 17592 13330 17644 13336
rect 18236 13330 18288 13336
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17512 13144 17724 13172
rect 17788 13161 17816 13262
rect 18432 13240 18460 13416
rect 18616 13444 18644 13518
rect 18616 13416 18690 13444
rect 18512 13398 18564 13404
rect 18662 13410 18690 13416
rect 18662 13394 18736 13410
rect 18662 13388 18748 13394
rect 18662 13382 18696 13388
rect 18696 13330 18748 13336
rect 18694 13288 18750 13297
rect 18432 13212 18644 13240
rect 18694 13223 18696 13232
rect 17868 13184 17920 13190
rect 17696 12968 17724 13144
rect 17774 13152 17830 13161
rect 17868 13126 17920 13132
rect 17774 13087 17830 13096
rect 17776 12980 17828 12986
rect 17420 12940 17540 12968
rect 17696 12940 17776 12968
rect 17512 12900 17540 12940
rect 17776 12922 17828 12928
rect 17512 12872 17724 12900
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17236 12430 17448 12458
rect 17420 11812 17448 12430
rect 17500 11824 17552 11830
rect 17420 11784 17500 11812
rect 17500 11766 17552 11772
rect 17604 11778 17632 12650
rect 17696 11898 17724 12872
rect 17880 12866 17908 13126
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 18616 12968 18644 13212
rect 18748 13223 18750 13232
rect 18696 13194 18748 13200
rect 17788 12838 17908 12866
rect 18432 12940 18644 12968
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 17788 12073 17816 12838
rect 17868 12776 17920 12782
rect 17868 12718 17920 12724
rect 17774 12064 17830 12073
rect 17774 11999 17830 12008
rect 17684 11892 17736 11898
rect 17880 11880 17908 12718
rect 17958 12472 18014 12481
rect 18142 12472 18198 12481
rect 17958 12407 18014 12416
rect 18064 12430 18142 12458
rect 17972 12084 18000 12407
rect 18064 12374 18092 12430
rect 18142 12407 18198 12416
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 18236 12096 18288 12102
rect 17972 12056 18236 12084
rect 18236 12038 18288 12044
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 18328 11892 18380 11898
rect 17880 11852 18000 11880
rect 17684 11834 17736 11840
rect 17604 11750 17816 11778
rect 17592 11688 17644 11694
rect 17592 11630 17644 11636
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17420 11218 17448 11494
rect 17408 11212 17460 11218
rect 17460 11172 17540 11200
rect 17408 11154 17460 11160
rect 17408 10736 17460 10742
rect 17408 10678 17460 10684
rect 17420 9897 17448 10678
rect 17512 10674 17540 11172
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17512 10130 17540 10610
rect 17604 10130 17632 11630
rect 17788 11354 17816 11750
rect 17868 11620 17920 11626
rect 17868 11562 17920 11568
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17880 11218 17908 11562
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17972 11098 18000 11852
rect 18328 11834 18380 11840
rect 17880 11070 18000 11098
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17592 10124 17644 10130
rect 17592 10066 17644 10072
rect 17684 9920 17736 9926
rect 17406 9888 17462 9897
rect 17684 9862 17736 9868
rect 17774 9888 17830 9897
rect 17406 9823 17462 9832
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17052 9030 17172 9058
rect 16948 6384 17000 6390
rect 16948 6326 17000 6332
rect 16856 5772 16908 5778
rect 16856 5714 16908 5720
rect 16948 5228 17000 5234
rect 16776 5188 16948 5216
rect 16948 5170 17000 5176
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4758 16344 4966
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16304 4752 16356 4758
rect 16304 4694 16356 4700
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15752 3664 15804 3670
rect 15752 3606 15804 3612
rect 15936 3664 15988 3670
rect 15936 3606 15988 3612
rect 15764 3534 15792 3606
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15948 2990 15976 3606
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15948 2650 15976 2790
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16408 2514 16436 2858
rect 16960 2650 16988 4762
rect 17052 3534 17080 9030
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17144 8090 17172 8910
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17144 7206 17172 7346
rect 17236 7274 17264 9318
rect 17224 7268 17276 7274
rect 17224 7210 17276 7216
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17132 6112 17184 6118
rect 17184 6072 17264 6100
rect 17132 6054 17184 6060
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17144 3670 17172 4014
rect 17132 3664 17184 3670
rect 17132 3606 17184 3612
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17144 3058 17172 3606
rect 17236 3398 17264 6072
rect 17328 5642 17356 9658
rect 17406 9480 17462 9489
rect 17406 9415 17462 9424
rect 17420 8498 17448 9415
rect 17498 9344 17554 9353
rect 17498 9279 17554 9288
rect 17512 8838 17540 9279
rect 17590 9208 17646 9217
rect 17590 9143 17646 9152
rect 17604 8945 17632 9143
rect 17590 8936 17646 8945
rect 17590 8871 17646 8880
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17512 6866 17540 8774
rect 17590 7712 17646 7721
rect 17590 7647 17646 7656
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17604 6662 17632 7647
rect 17592 6656 17644 6662
rect 17592 6598 17644 6604
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17420 5250 17448 5306
rect 17420 5222 17540 5250
rect 17314 4720 17370 4729
rect 17314 4655 17370 4664
rect 17328 4457 17356 4655
rect 17408 4548 17460 4554
rect 17408 4490 17460 4496
rect 17314 4448 17370 4457
rect 17314 4383 17370 4392
rect 17224 3392 17276 3398
rect 17224 3334 17276 3340
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 16948 2644 17000 2650
rect 16948 2586 17000 2592
rect 16396 2508 16448 2514
rect 16396 2450 16448 2456
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 16488 2440 16540 2446
rect 16488 2382 16540 2388
rect 15764 1154 15792 2382
rect 16500 1902 16528 2382
rect 16488 1896 16540 1902
rect 16488 1838 16540 1844
rect 16488 1420 16540 1426
rect 16488 1362 16540 1368
rect 15752 1148 15804 1154
rect 15752 1090 15804 1096
rect 16500 814 16528 1362
rect 16488 808 16540 814
rect 17420 800 17448 4490
rect 17512 1902 17540 5222
rect 17696 3534 17724 9862
rect 17774 9823 17830 9832
rect 17788 6458 17816 9823
rect 17880 9674 17908 11070
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18156 10266 18184 10746
rect 18234 10296 18290 10305
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 18144 10260 18196 10266
rect 18234 10231 18290 10240
rect 18144 10202 18196 10208
rect 17972 9926 18000 10202
rect 18248 10198 18276 10231
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 17960 9920 18012 9926
rect 17960 9862 18012 9868
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17880 9646 18184 9674
rect 18156 9382 18184 9646
rect 18144 9376 18196 9382
rect 17866 9344 17922 9353
rect 18144 9318 18196 9324
rect 17866 9279 17922 9288
rect 17880 9178 17908 9279
rect 17868 9172 17920 9178
rect 17868 9114 17920 9120
rect 17866 8936 17922 8945
rect 17866 8871 17868 8880
rect 17920 8871 17922 8880
rect 17868 8842 17920 8848
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 18052 8424 18104 8430
rect 18050 8392 18052 8401
rect 18104 8392 18106 8401
rect 18050 8327 18106 8336
rect 17868 7948 17920 7954
rect 17868 7890 17920 7896
rect 17776 6452 17828 6458
rect 17776 6394 17828 6400
rect 17880 6338 17908 7890
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 18340 7546 18368 11834
rect 18432 10606 18460 12940
rect 18604 12844 18656 12850
rect 18708 12832 18736 12951
rect 18656 12804 18736 12832
rect 18604 12786 18656 12792
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18512 12232 18564 12238
rect 18512 12174 18564 12180
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18420 9580 18472 9586
rect 18420 9522 18472 9528
rect 18432 8634 18460 9522
rect 18524 9500 18552 12174
rect 18616 12073 18644 12242
rect 18602 12064 18658 12073
rect 18602 11999 18658 12008
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18616 9654 18644 11222
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 18708 9994 18736 11018
rect 18800 10520 18828 14554
rect 18892 13870 18920 16594
rect 18972 16448 19024 16454
rect 18970 16416 18972 16425
rect 19024 16416 19026 16425
rect 18970 16351 19026 16360
rect 18972 16244 19024 16250
rect 18972 16186 19024 16192
rect 18984 16046 19012 16186
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 19076 15978 19104 18702
rect 19154 18663 19210 18672
rect 19168 18630 19196 18663
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19156 18216 19208 18222
rect 19156 18158 19208 18164
rect 19248 18216 19300 18222
rect 19248 18158 19300 18164
rect 19168 17241 19196 18158
rect 19260 18057 19288 18158
rect 19246 18048 19302 18057
rect 19246 17983 19302 17992
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19154 17232 19210 17241
rect 19154 17167 19210 17176
rect 19168 17066 19196 17167
rect 19156 17060 19208 17066
rect 19156 17002 19208 17008
rect 19260 16810 19288 17546
rect 19168 16782 19288 16810
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 18984 14056 19012 15642
rect 19076 14958 19104 15914
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 19076 14346 19104 14894
rect 19064 14340 19116 14346
rect 19064 14282 19116 14288
rect 18984 14028 19104 14056
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18892 13376 18920 13806
rect 18892 13348 19012 13376
rect 18878 13288 18934 13297
rect 18878 13223 18934 13232
rect 18892 12986 18920 13223
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18892 12481 18920 12650
rect 18878 12472 18934 12481
rect 18878 12407 18880 12416
rect 18932 12407 18934 12416
rect 18880 12378 18932 12384
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18892 11393 18920 11834
rect 18878 11384 18934 11393
rect 18878 11319 18934 11328
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18892 10985 18920 11086
rect 18878 10976 18934 10985
rect 18878 10911 18934 10920
rect 18800 10492 18920 10520
rect 18786 10024 18842 10033
rect 18696 9988 18748 9994
rect 18786 9959 18842 9968
rect 18696 9930 18748 9936
rect 18708 9722 18736 9930
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18524 9472 18736 9500
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18524 7750 18552 9114
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18326 7304 18382 7313
rect 18326 7239 18382 7248
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 18340 6361 18368 7239
rect 18524 6866 18552 7346
rect 18512 6860 18564 6866
rect 18512 6802 18564 6808
rect 17788 6310 17908 6338
rect 18326 6352 18382 6361
rect 17788 4162 17816 6310
rect 18326 6287 18382 6296
rect 18328 6180 18380 6186
rect 18328 6122 18380 6128
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 18340 5370 18368 6122
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18328 5364 18380 5370
rect 18328 5306 18380 5312
rect 18326 5128 18382 5137
rect 18326 5063 18382 5072
rect 17868 4616 17920 4622
rect 17868 4558 17920 4564
rect 17880 4282 17908 4558
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 17868 4276 17920 4282
rect 17868 4218 17920 4224
rect 17788 4134 18000 4162
rect 17972 3754 18000 4134
rect 18340 3913 18368 5063
rect 18420 5024 18472 5030
rect 18420 4966 18472 4972
rect 18326 3904 18382 3913
rect 18326 3839 18382 3848
rect 17972 3726 18368 3754
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17604 3194 17632 3470
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17696 2650 17724 3334
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17592 2644 17644 2650
rect 17592 2586 17644 2592
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17604 2553 17632 2586
rect 17590 2544 17646 2553
rect 17590 2479 17646 2488
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17788 1970 17816 2382
rect 17776 1964 17828 1970
rect 17776 1906 17828 1912
rect 17500 1896 17552 1902
rect 17500 1838 17552 1844
rect 17880 950 17908 3130
rect 18340 2774 18368 3726
rect 18432 3466 18460 4966
rect 18616 4826 18644 5714
rect 18708 5234 18736 9472
rect 18800 9178 18828 9959
rect 18788 9172 18840 9178
rect 18788 9114 18840 9120
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18800 8634 18828 8910
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18892 7886 18920 10492
rect 18984 8498 19012 13348
rect 19076 9761 19104 14028
rect 19168 13530 19196 16782
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19260 15978 19288 16662
rect 19248 15972 19300 15978
rect 19248 15914 19300 15920
rect 19352 15706 19380 21791
rect 19720 21350 19748 22510
rect 19812 22166 19840 24550
rect 19800 22160 19852 22166
rect 19904 22137 19932 25094
rect 19800 22102 19852 22108
rect 19890 22128 19946 22137
rect 19890 22063 19946 22072
rect 19708 21344 19760 21350
rect 19708 21286 19760 21292
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19522 20904 19578 20913
rect 19444 20602 19472 20878
rect 19996 20874 20024 25094
rect 20088 24206 20116 26182
rect 20272 24954 20300 26200
rect 20260 24948 20312 24954
rect 20260 24890 20312 24896
rect 20352 24608 20404 24614
rect 20352 24550 20404 24556
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 20076 23520 20128 23526
rect 20076 23462 20128 23468
rect 20088 23186 20116 23462
rect 20076 23180 20128 23186
rect 20076 23122 20128 23128
rect 20074 22808 20130 22817
rect 20074 22743 20130 22752
rect 20088 22710 20116 22743
rect 20076 22704 20128 22710
rect 20076 22646 20128 22652
rect 20088 22409 20116 22646
rect 20074 22400 20130 22409
rect 20074 22335 20130 22344
rect 20076 22092 20128 22098
rect 20076 22034 20128 22040
rect 19522 20839 19578 20848
rect 19984 20868 20036 20874
rect 19432 20596 19484 20602
rect 19432 20538 19484 20544
rect 19432 20460 19484 20466
rect 19432 20402 19484 20408
rect 19444 18766 19472 20402
rect 19536 19922 19564 20839
rect 19984 20810 20036 20816
rect 19614 20768 19670 20777
rect 19614 20703 19670 20712
rect 19524 19916 19576 19922
rect 19524 19858 19576 19864
rect 19628 19854 19656 20703
rect 20088 19922 20116 22034
rect 20180 21146 20208 24142
rect 20364 23594 20392 24550
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22545 20300 22986
rect 20258 22536 20314 22545
rect 20258 22471 20314 22480
rect 20364 22438 20392 23530
rect 20352 22432 20404 22438
rect 20352 22374 20404 22380
rect 20260 22024 20312 22030
rect 20352 22024 20404 22030
rect 20260 21966 20312 21972
rect 20350 21992 20352 22001
rect 20404 21992 20406 22001
rect 20272 21554 20300 21966
rect 20350 21927 20406 21936
rect 20260 21548 20312 21554
rect 20260 21490 20312 21496
rect 20260 21344 20312 21350
rect 20260 21286 20312 21292
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 20272 19854 20300 21286
rect 20548 20398 20576 26590
rect 20902 26200 20958 27000
rect 21546 26200 21602 27000
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 20812 25492 20864 25498
rect 20812 25434 20864 25440
rect 20824 25226 20852 25434
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20628 24268 20680 24274
rect 20628 24210 20680 24216
rect 20640 23050 20668 24210
rect 20628 23044 20680 23050
rect 20628 22986 20680 22992
rect 20640 22710 20668 22986
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20640 21962 20668 22646
rect 20732 22098 20760 24890
rect 20812 24880 20864 24886
rect 20812 24822 20864 24828
rect 20720 22092 20772 22098
rect 20720 22034 20772 22040
rect 20628 21956 20680 21962
rect 20628 21898 20680 21904
rect 20640 21622 20668 21898
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20720 20800 20772 20806
rect 20720 20742 20772 20748
rect 20732 20618 20760 20742
rect 20640 20590 20760 20618
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20640 20058 20668 20590
rect 20628 20052 20680 20058
rect 20628 19994 20680 20000
rect 20720 20052 20772 20058
rect 20720 19994 20772 20000
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19432 18624 19484 18630
rect 19432 18566 19484 18572
rect 19444 17542 19472 18566
rect 19536 18329 19564 19110
rect 19522 18320 19578 18329
rect 19522 18255 19524 18264
rect 19576 18255 19578 18264
rect 19524 18226 19576 18232
rect 19524 18148 19576 18154
rect 19524 18090 19576 18096
rect 19432 17536 19484 17542
rect 19432 17478 19484 17484
rect 19430 16416 19486 16425
rect 19430 16351 19486 16360
rect 19444 16250 19472 16351
rect 19432 16244 19484 16250
rect 19432 16186 19484 16192
rect 19432 16108 19484 16114
rect 19432 16050 19484 16056
rect 19340 15700 19392 15706
rect 19340 15642 19392 15648
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19156 13524 19208 13530
rect 19156 13466 19208 13472
rect 19156 13388 19208 13394
rect 19156 13330 19208 13336
rect 19168 12866 19196 13330
rect 19260 13297 19288 15438
rect 19444 14464 19472 16050
rect 19536 15337 19564 18090
rect 19628 18057 19656 19314
rect 19614 18048 19670 18057
rect 19614 17983 19670 17992
rect 19614 17776 19670 17785
rect 19614 17711 19670 17720
rect 19628 17542 19656 17711
rect 19616 17536 19668 17542
rect 19616 17478 19668 17484
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19522 15328 19578 15337
rect 19522 15263 19578 15272
rect 19352 14436 19472 14464
rect 19246 13288 19302 13297
rect 19352 13258 19380 14436
rect 19524 14408 19576 14414
rect 19524 14350 19576 14356
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19246 13223 19302 13232
rect 19340 13252 19392 13258
rect 19340 13194 19392 13200
rect 19338 13152 19394 13161
rect 19338 13087 19394 13096
rect 19168 12838 19288 12866
rect 19156 12776 19208 12782
rect 19156 12718 19208 12724
rect 19062 9752 19118 9761
rect 19062 9687 19118 9696
rect 19064 9648 19116 9654
rect 19064 9590 19116 9596
rect 19076 8906 19104 9590
rect 19064 8900 19116 8906
rect 19064 8842 19116 8848
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18972 7880 19024 7886
rect 18972 7822 19024 7828
rect 18984 7274 19012 7822
rect 18972 7268 19024 7274
rect 18972 7210 19024 7216
rect 19168 5710 19196 12718
rect 19260 11937 19288 12838
rect 19246 11928 19302 11937
rect 19246 11863 19302 11872
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19260 7478 19288 11630
rect 19352 9450 19380 13087
rect 19444 11150 19472 14282
rect 19536 13870 19564 14350
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19628 13394 19656 17138
rect 19720 16658 19748 19314
rect 19812 18358 19840 19722
rect 19984 19168 20036 19174
rect 19984 19110 20036 19116
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19798 17776 19854 17785
rect 19798 17711 19854 17720
rect 19812 17270 19840 17711
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19720 15502 19748 16594
rect 19904 15706 19932 18906
rect 19996 18834 20024 19110
rect 20272 18834 20300 19790
rect 20536 19780 20588 19786
rect 20536 19722 20588 19728
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 19984 18828 20036 18834
rect 19984 18770 20036 18776
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 19996 18222 20024 18770
rect 20258 18728 20314 18737
rect 20258 18663 20314 18672
rect 19984 18216 20036 18222
rect 19984 18158 20036 18164
rect 20076 18080 20128 18086
rect 19982 18048 20038 18057
rect 20076 18022 20128 18028
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 19982 17983 20038 17992
rect 19996 17785 20024 17983
rect 19982 17776 20038 17785
rect 19982 17711 20038 17720
rect 19996 16454 20024 17711
rect 20088 16794 20116 18022
rect 20180 17134 20208 18022
rect 20272 17542 20300 18663
rect 20364 18578 20392 19450
rect 20442 18592 20498 18601
rect 20364 18550 20442 18578
rect 20442 18527 20498 18536
rect 20442 18320 20498 18329
rect 20442 18255 20498 18264
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 20364 17354 20392 18022
rect 20272 17326 20392 17354
rect 20168 17128 20220 17134
rect 20168 17070 20220 17076
rect 20272 16998 20300 17326
rect 20352 17264 20404 17270
rect 20352 17206 20404 17212
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19984 16448 20036 16454
rect 19984 16390 20036 16396
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19892 15700 19944 15706
rect 19892 15642 19944 15648
rect 19890 15600 19946 15609
rect 19890 15535 19946 15544
rect 19708 15496 19760 15502
rect 19708 15438 19760 15444
rect 19708 14952 19760 14958
rect 19708 14894 19760 14900
rect 19720 14482 19748 14894
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19904 14362 19932 15535
rect 19996 14958 20024 15846
rect 20088 15570 20116 15846
rect 20166 15600 20222 15609
rect 20076 15564 20128 15570
rect 20166 15535 20168 15544
rect 20076 15506 20128 15512
rect 20220 15535 20222 15544
rect 20168 15506 20220 15512
rect 20272 15314 20300 16934
rect 20088 15286 20300 15314
rect 19984 14952 20036 14958
rect 19984 14894 20036 14900
rect 20088 14385 20116 15286
rect 20258 14784 20314 14793
rect 20258 14719 20314 14728
rect 20272 14482 20300 14719
rect 20260 14476 20312 14482
rect 20260 14418 20312 14424
rect 20074 14376 20130 14385
rect 19812 14113 19840 14350
rect 19904 14334 20024 14362
rect 19892 14272 19944 14278
rect 19892 14214 19944 14220
rect 19798 14104 19854 14113
rect 19798 14039 19800 14048
rect 19852 14039 19854 14048
rect 19800 14010 19852 14016
rect 19798 13696 19854 13705
rect 19798 13631 19854 13640
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19708 13320 19760 13326
rect 19708 13262 19760 13268
rect 19524 13184 19576 13190
rect 19524 13126 19576 13132
rect 19536 12850 19564 13126
rect 19616 12912 19668 12918
rect 19616 12854 19668 12860
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19628 12102 19656 12854
rect 19720 12850 19748 13262
rect 19812 13025 19840 13631
rect 19798 13016 19854 13025
rect 19798 12951 19854 12960
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19616 12096 19668 12102
rect 19616 12038 19668 12044
rect 19536 11694 19564 12038
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19524 11688 19576 11694
rect 19524 11630 19576 11636
rect 19628 11626 19656 11698
rect 19616 11620 19668 11626
rect 19616 11562 19668 11568
rect 19628 11336 19656 11562
rect 19720 11558 19748 12786
rect 19800 12096 19852 12102
rect 19800 12038 19852 12044
rect 19812 11558 19840 12038
rect 19708 11552 19760 11558
rect 19708 11494 19760 11500
rect 19800 11552 19852 11558
rect 19800 11494 19852 11500
rect 19536 11308 19656 11336
rect 19432 11144 19484 11150
rect 19432 11086 19484 11092
rect 19444 10266 19472 11086
rect 19536 11082 19564 11308
rect 19720 11218 19748 11494
rect 19616 11212 19668 11218
rect 19616 11154 19668 11160
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19628 11082 19656 11154
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19536 10810 19564 11018
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19616 10532 19668 10538
rect 19616 10474 19668 10480
rect 19628 10266 19656 10474
rect 19432 10260 19484 10266
rect 19432 10202 19484 10208
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19432 10124 19484 10130
rect 19432 10066 19484 10072
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 19352 6798 19380 8366
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19338 6216 19394 6225
rect 19338 6151 19394 6160
rect 19246 5808 19302 5817
rect 19246 5743 19302 5752
rect 19156 5704 19208 5710
rect 19156 5646 19208 5652
rect 18696 5228 18748 5234
rect 18696 5170 18748 5176
rect 18880 5160 18932 5166
rect 18880 5102 18932 5108
rect 18892 5001 18920 5102
rect 18878 4992 18934 5001
rect 18878 4927 18934 4936
rect 18892 4826 18920 4927
rect 18604 4820 18656 4826
rect 18604 4762 18656 4768
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 19260 4690 19288 5743
rect 19248 4684 19300 4690
rect 19248 4626 19300 4632
rect 19260 4282 19288 4626
rect 19248 4276 19300 4282
rect 19248 4218 19300 4224
rect 19352 4049 19380 6151
rect 19444 5302 19472 10066
rect 19720 9994 19748 11154
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19536 8430 19564 9862
rect 19614 9344 19670 9353
rect 19614 9279 19670 9288
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19628 5302 19656 9279
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7177 19748 7822
rect 19812 7410 19840 11494
rect 19904 9926 19932 14214
rect 19996 13954 20024 14334
rect 20074 14311 20130 14320
rect 20272 14074 20300 14418
rect 20260 14068 20312 14074
rect 20260 14010 20312 14016
rect 19996 13926 20208 13954
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19996 12238 20024 13806
rect 20088 12646 20116 13806
rect 20180 12646 20208 13926
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20168 12640 20220 12646
rect 20168 12582 20220 12588
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 20088 10470 20116 12582
rect 20272 12186 20300 13738
rect 20364 12442 20392 17206
rect 20456 15450 20484 18255
rect 20548 18057 20576 19722
rect 20640 19689 20668 19994
rect 20626 19680 20682 19689
rect 20626 19615 20682 19624
rect 20732 18766 20760 19994
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20534 18048 20590 18057
rect 20534 17983 20590 17992
rect 20640 17746 20668 18566
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20534 16960 20590 16969
rect 20534 16895 20590 16904
rect 20548 15638 20576 16895
rect 20640 16708 20668 17478
rect 20732 17338 20760 17575
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20824 16810 20852 24822
rect 20916 24274 20944 26200
rect 21272 25900 21324 25906
rect 21272 25842 21324 25848
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20916 23186 20944 23598
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20916 20602 20944 23122
rect 21008 22953 21036 23666
rect 21100 22982 21128 25434
rect 21088 22976 21140 22982
rect 20994 22944 21050 22953
rect 21088 22918 21140 22924
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 20994 22879 21050 22888
rect 21008 22574 21036 22879
rect 20996 22568 21048 22574
rect 20996 22510 21048 22516
rect 20996 21616 21048 21622
rect 21088 21616 21140 21622
rect 20996 21558 21048 21564
rect 21086 21584 21088 21593
rect 21140 21584 21142 21593
rect 21008 20874 21036 21558
rect 21086 21519 21142 21528
rect 21086 21176 21142 21185
rect 21086 21111 21142 21120
rect 21100 21078 21128 21111
rect 21088 21072 21140 21078
rect 21088 21014 21140 21020
rect 20996 20868 21048 20874
rect 20996 20810 21048 20816
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 20916 18834 20944 20538
rect 21008 19786 21036 20810
rect 21086 20360 21142 20369
rect 21086 20295 21142 20304
rect 20996 19780 21048 19786
rect 20996 19722 21048 19728
rect 21008 19446 21036 19722
rect 20996 19440 21048 19446
rect 20996 19382 21048 19388
rect 20994 19136 21050 19145
rect 20994 19071 21050 19080
rect 20904 18828 20956 18834
rect 20904 18770 20956 18776
rect 21008 18329 21036 19071
rect 21100 18737 21128 20295
rect 21192 19718 21220 22918
rect 21284 22817 21312 25842
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21376 23798 21404 24754
rect 21456 24336 21508 24342
rect 21456 24278 21508 24284
rect 21364 23792 21416 23798
rect 21364 23734 21416 23740
rect 21270 22808 21326 22817
rect 21270 22743 21326 22752
rect 21272 22228 21324 22234
rect 21272 22170 21324 22176
rect 21284 21350 21312 22170
rect 21362 22128 21418 22137
rect 21468 22098 21496 24278
rect 21560 24274 21588 26200
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21744 22409 21772 26930
rect 22190 26330 22246 27000
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 22190 26302 22784 26330
rect 22112 25922 22140 26250
rect 22190 26200 22246 26302
rect 22376 26240 22428 26246
rect 22376 26182 22428 26188
rect 22112 25894 22232 25922
rect 22100 25696 22152 25702
rect 22100 25638 22152 25644
rect 22112 25294 22140 25638
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 21916 25220 21968 25226
rect 21916 25162 21968 25168
rect 21824 22976 21876 22982
rect 21824 22918 21876 22924
rect 21730 22400 21786 22409
rect 21730 22335 21786 22344
rect 21730 22264 21786 22273
rect 21730 22199 21786 22208
rect 21638 22128 21694 22137
rect 21362 22063 21418 22072
rect 21456 22092 21508 22098
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21376 20874 21404 22063
rect 21638 22063 21694 22072
rect 21456 22034 21508 22040
rect 21454 21856 21510 21865
rect 21454 21791 21510 21800
rect 21468 21321 21496 21791
rect 21652 21486 21680 22063
rect 21640 21480 21692 21486
rect 21640 21422 21692 21428
rect 21640 21344 21692 21350
rect 21454 21312 21510 21321
rect 21640 21286 21692 21292
rect 21454 21247 21510 21256
rect 21364 20868 21416 20874
rect 21364 20810 21416 20816
rect 21272 20800 21324 20806
rect 21272 20742 21324 20748
rect 21284 20466 21312 20742
rect 21272 20460 21324 20466
rect 21272 20402 21324 20408
rect 21468 20398 21496 21247
rect 21546 20632 21602 20641
rect 21546 20567 21602 20576
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21454 20088 21510 20097
rect 21454 20023 21510 20032
rect 21180 19712 21232 19718
rect 21180 19654 21232 19660
rect 21468 19514 21496 20023
rect 21456 19508 21508 19514
rect 21456 19450 21508 19456
rect 21272 19440 21324 19446
rect 21272 19382 21324 19388
rect 21086 18728 21142 18737
rect 21086 18663 21142 18672
rect 20994 18320 21050 18329
rect 20994 18255 21050 18264
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 16998 20944 17478
rect 21192 17270 21220 17818
rect 21284 17610 21312 19382
rect 21364 19304 21416 19310
rect 21364 19246 21416 19252
rect 21272 17604 21324 17610
rect 21272 17546 21324 17552
rect 21180 17264 21232 17270
rect 21180 17206 21232 17212
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20824 16782 21312 16810
rect 20720 16720 20772 16726
rect 20640 16680 20720 16708
rect 20720 16662 20772 16668
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20628 16040 20680 16046
rect 20628 15982 20680 15988
rect 20536 15632 20588 15638
rect 20534 15600 20536 15609
rect 20588 15600 20590 15609
rect 20534 15535 20590 15544
rect 20456 15422 20576 15450
rect 20444 15360 20496 15366
rect 20444 15302 20496 15308
rect 20352 12436 20404 12442
rect 20352 12378 20404 12384
rect 20272 12158 20392 12186
rect 20260 12096 20312 12102
rect 20260 12038 20312 12044
rect 20166 11928 20222 11937
rect 20272 11898 20300 12038
rect 20166 11863 20222 11872
rect 20260 11892 20312 11898
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 20180 10418 20208 11863
rect 20260 11834 20312 11840
rect 20364 11830 20392 12158
rect 20352 11824 20404 11830
rect 20352 11766 20404 11772
rect 20260 11212 20312 11218
rect 20260 11154 20312 11160
rect 20272 10742 20300 11154
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20180 10390 20300 10418
rect 19982 10296 20038 10305
rect 19982 10231 20038 10240
rect 20168 10260 20220 10266
rect 19996 10033 20024 10231
rect 20168 10202 20220 10208
rect 19982 10024 20038 10033
rect 19982 9959 20038 9968
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 19996 7546 20024 8434
rect 19984 7540 20036 7546
rect 19984 7482 20036 7488
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19706 7168 19762 7177
rect 19706 7103 19762 7112
rect 19706 6760 19762 6769
rect 19706 6695 19762 6704
rect 19720 5778 19748 6695
rect 19708 5772 19760 5778
rect 19708 5714 19760 5720
rect 19432 5296 19484 5302
rect 19432 5238 19484 5244
rect 19616 5296 19668 5302
rect 19616 5238 19668 5244
rect 19982 5264 20038 5273
rect 19800 5228 19852 5234
rect 19982 5199 19984 5208
rect 19800 5170 19852 5176
rect 20036 5199 20038 5208
rect 19984 5170 20036 5176
rect 19338 4040 19394 4049
rect 19338 3975 19394 3984
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18432 3058 18460 3402
rect 18524 3058 18552 3674
rect 19536 3602 19564 3878
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 18880 3460 18932 3466
rect 18880 3402 18932 3408
rect 18696 3392 18748 3398
rect 18696 3334 18748 3340
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18340 2746 18460 2774
rect 18432 2582 18460 2746
rect 18420 2576 18472 2582
rect 18420 2518 18472 2524
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18708 1086 18736 3334
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18800 2106 18828 2246
rect 18788 2100 18840 2106
rect 18788 2042 18840 2048
rect 18696 1080 18748 1086
rect 18696 1022 18748 1028
rect 17868 944 17920 950
rect 17868 886 17920 892
rect 16488 750 16540 756
rect 15476 468 15528 474
rect 15476 410 15528 416
rect 17406 0 17462 800
rect 18800 542 18828 2042
rect 18788 536 18840 542
rect 18788 478 18840 484
rect 18892 270 18920 3402
rect 19812 3398 19840 5170
rect 20076 4072 20128 4078
rect 20076 4014 20128 4020
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19904 3738 19932 3878
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18984 1766 19012 2246
rect 18972 1760 19024 1766
rect 18972 1702 19024 1708
rect 19352 1494 19380 3334
rect 19904 3126 19932 3674
rect 19892 3120 19944 3126
rect 19892 3062 19944 3068
rect 19432 2576 19484 2582
rect 19432 2518 19484 2524
rect 19444 2446 19472 2518
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19628 2106 19656 2382
rect 19616 2100 19668 2106
rect 19616 2042 19668 2048
rect 19340 1488 19392 1494
rect 19340 1430 19392 1436
rect 20088 800 20116 4014
rect 20180 2553 20208 10202
rect 20272 9178 20300 10390
rect 20350 10296 20406 10305
rect 20350 10231 20406 10240
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20364 6882 20392 10231
rect 20456 8838 20484 15302
rect 20548 14521 20576 15422
rect 20640 15162 20668 15982
rect 20904 15564 20956 15570
rect 20904 15506 20956 15512
rect 20812 15428 20864 15434
rect 20812 15370 20864 15376
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20628 14816 20680 14822
rect 20680 14776 20760 14804
rect 20628 14758 20680 14764
rect 20534 14512 20590 14521
rect 20534 14447 20590 14456
rect 20548 13394 20576 14447
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20536 13252 20588 13258
rect 20536 13194 20588 13200
rect 20548 9382 20576 13194
rect 20640 12073 20668 13942
rect 20732 13705 20760 14776
rect 20824 14074 20852 15370
rect 20916 14074 20944 15506
rect 21008 15094 21036 16594
rect 21180 16040 21232 16046
rect 21180 15982 21232 15988
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20904 14068 20956 14074
rect 20904 14010 20956 14016
rect 20902 13968 20958 13977
rect 20902 13903 20958 13912
rect 20812 13796 20864 13802
rect 20812 13738 20864 13744
rect 20718 13696 20774 13705
rect 20718 13631 20774 13640
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20626 12064 20682 12073
rect 20626 11999 20682 12008
rect 20628 11756 20680 11762
rect 20628 11698 20680 11704
rect 20640 11286 20668 11698
rect 20732 11558 20760 12378
rect 20824 12356 20852 13738
rect 20916 12617 20944 13903
rect 21008 13258 21036 15030
rect 21100 14890 21128 15302
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 21100 13841 21128 13874
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21192 13138 21220 15982
rect 21008 13110 21220 13138
rect 20902 12608 20958 12617
rect 20902 12543 20958 12552
rect 20824 12328 20944 12356
rect 20720 11552 20772 11558
rect 20916 11529 20944 12328
rect 21008 11898 21036 13110
rect 21284 13002 21312 16782
rect 21376 14482 21404 19246
rect 21468 17066 21496 19450
rect 21456 17060 21508 17066
rect 21456 17002 21508 17008
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 21468 16114 21496 16662
rect 21560 16590 21588 20567
rect 21652 20534 21680 21286
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21640 20324 21692 20330
rect 21640 20266 21692 20272
rect 21652 19009 21680 20266
rect 21638 19000 21694 19009
rect 21638 18935 21694 18944
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21652 17202 21680 17614
rect 21640 17196 21692 17202
rect 21640 17138 21692 17144
rect 21744 16658 21772 22199
rect 21836 20913 21864 22918
rect 21822 20904 21878 20913
rect 21822 20839 21878 20848
rect 21824 20800 21876 20806
rect 21824 20742 21876 20748
rect 21836 20641 21864 20742
rect 21822 20632 21878 20641
rect 21822 20567 21878 20576
rect 21824 20528 21876 20534
rect 21824 20470 21876 20476
rect 21836 19258 21864 20470
rect 21928 19514 21956 25162
rect 22006 23488 22062 23497
rect 22006 23423 22062 23432
rect 22020 22545 22048 23423
rect 22006 22536 22062 22545
rect 22006 22471 22062 22480
rect 22100 22160 22152 22166
rect 22100 22102 22152 22108
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 21350 22048 21490
rect 22008 21344 22060 21350
rect 22008 21286 22060 21292
rect 22008 20460 22060 20466
rect 22008 20402 22060 20408
rect 22020 20058 22048 20402
rect 22008 20052 22060 20058
rect 22008 19994 22060 20000
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 22112 19334 22140 22102
rect 22204 20777 22232 25894
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22296 24206 22324 25638
rect 22284 24200 22336 24206
rect 22284 24142 22336 24148
rect 22284 23860 22336 23866
rect 22284 23802 22336 23808
rect 22296 23186 22324 23802
rect 22388 23662 22416 26182
rect 22560 25288 22612 25294
rect 22560 25230 22612 25236
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22466 24984 22522 24993
rect 22466 24919 22522 24928
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22480 23361 22508 24919
rect 22572 24886 22600 25230
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22560 24744 22612 24750
rect 22560 24686 22612 24692
rect 22572 24274 22600 24686
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22560 23792 22612 23798
rect 22560 23734 22612 23740
rect 22466 23352 22522 23361
rect 22466 23287 22522 23296
rect 22284 23180 22336 23186
rect 22284 23122 22336 23128
rect 22296 22642 22324 23122
rect 22466 22808 22522 22817
rect 22466 22743 22522 22752
rect 22284 22636 22336 22642
rect 22284 22578 22336 22584
rect 22282 22264 22338 22273
rect 22282 22199 22338 22208
rect 22296 21418 22324 22199
rect 22480 22137 22508 22743
rect 22466 22128 22522 22137
rect 22466 22063 22522 22072
rect 22376 21480 22428 21486
rect 22376 21422 22428 21428
rect 22284 21412 22336 21418
rect 22284 21354 22336 21360
rect 22190 20768 22246 20777
rect 22190 20703 22246 20712
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22204 20466 22232 20538
rect 22192 20460 22244 20466
rect 22192 20402 22244 20408
rect 22296 19990 22324 21354
rect 22284 19984 22336 19990
rect 22284 19926 22336 19932
rect 22388 19836 22416 21422
rect 22572 20942 22600 23734
rect 22664 23186 22692 25230
rect 22756 24154 22784 26302
rect 22834 26200 22890 27000
rect 22928 26852 22980 26858
rect 22928 26794 22980 26800
rect 23388 26852 23440 26858
rect 23388 26794 23440 26800
rect 22848 24954 22876 26200
rect 22836 24948 22888 24954
rect 22836 24890 22888 24896
rect 22940 24857 22968 26794
rect 23400 26246 23428 26794
rect 23478 26330 23534 27000
rect 23478 26302 23888 26330
rect 23388 26240 23440 26246
rect 23478 26200 23534 26302
rect 23388 26182 23440 26188
rect 23388 25084 23440 25090
rect 23388 25026 23440 25032
rect 22926 24848 22982 24857
rect 22926 24783 22982 24792
rect 22836 24744 22888 24750
rect 22836 24686 22888 24692
rect 22848 24290 22876 24686
rect 23400 24585 23428 25026
rect 23480 25016 23532 25022
rect 23480 24958 23532 24964
rect 23386 24576 23442 24585
rect 22950 24508 23258 24517
rect 23386 24511 23442 24520
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22848 24262 22968 24290
rect 22756 24126 22876 24154
rect 22744 23656 22796 23662
rect 22744 23598 22796 23604
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22652 22432 22704 22438
rect 22652 22374 22704 22380
rect 22664 22234 22692 22374
rect 22652 22228 22704 22234
rect 22652 22170 22704 22176
rect 22756 22098 22784 23598
rect 22652 22092 22704 22098
rect 22652 22034 22704 22040
rect 22744 22092 22796 22098
rect 22744 22034 22796 22040
rect 22560 20936 22612 20942
rect 22560 20878 22612 20884
rect 22560 20800 22612 20806
rect 22560 20742 22612 20748
rect 22468 20392 22520 20398
rect 22468 20334 22520 20340
rect 22296 19808 22416 19836
rect 22112 19306 22232 19334
rect 21836 19230 22140 19258
rect 22008 18284 22060 18290
rect 22008 18226 22060 18232
rect 21822 18048 21878 18057
rect 21822 17983 21878 17992
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21468 14482 21496 16050
rect 21640 15972 21692 15978
rect 21640 15914 21692 15920
rect 21652 15366 21680 15914
rect 21640 15360 21692 15366
rect 21640 15302 21692 15308
rect 21548 15156 21600 15162
rect 21548 15098 21600 15104
rect 21560 14550 21588 15098
rect 21548 14544 21600 14550
rect 21548 14486 21600 14492
rect 21364 14476 21416 14482
rect 21364 14418 21416 14424
rect 21456 14476 21508 14482
rect 21456 14418 21508 14424
rect 21364 14272 21416 14278
rect 21364 14214 21416 14220
rect 21192 12974 21312 13002
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21192 11762 21220 12974
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20720 11494 20772 11500
rect 20902 11520 20958 11529
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20732 11014 20760 11494
rect 20902 11455 20958 11464
rect 20720 11008 20772 11014
rect 20720 10950 20772 10956
rect 20720 10464 20772 10470
rect 20772 10424 20852 10452
rect 20720 10406 20772 10412
rect 20824 10266 20852 10424
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20444 8832 20496 8838
rect 20444 8774 20496 8780
rect 20640 8634 20668 9522
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 7002 20576 7346
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20364 6854 20668 6882
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 4486 20392 5646
rect 20352 4480 20404 4486
rect 20352 4422 20404 4428
rect 20166 2544 20222 2553
rect 20166 2479 20222 2488
rect 20364 1018 20392 4422
rect 20640 4146 20668 6854
rect 20732 4690 20760 9862
rect 20916 9110 20944 11455
rect 20996 10464 21048 10470
rect 20996 10406 21048 10412
rect 21100 10418 21128 11630
rect 21376 11608 21404 14214
rect 21548 14068 21600 14074
rect 21548 14010 21600 14016
rect 21454 13968 21510 13977
rect 21454 13903 21456 13912
rect 21508 13903 21510 13912
rect 21456 13874 21508 13880
rect 21560 13462 21588 14010
rect 21548 13456 21600 13462
rect 21548 13398 21600 13404
rect 21548 12912 21600 12918
rect 21548 12854 21600 12860
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21284 11580 21404 11608
rect 21180 11076 21232 11082
rect 21180 11018 21232 11024
rect 21192 10538 21220 11018
rect 21284 10810 21312 11580
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21272 10804 21324 10810
rect 21272 10746 21324 10752
rect 21180 10532 21232 10538
rect 21180 10474 21232 10480
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20916 8090 20944 8910
rect 21008 8362 21036 10406
rect 21100 10390 21220 10418
rect 21086 9208 21142 9217
rect 21086 9143 21142 9152
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20824 6458 20852 6734
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 21008 5846 21036 6258
rect 20996 5840 21048 5846
rect 20996 5782 21048 5788
rect 21008 4826 21036 5782
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 20720 4684 20772 4690
rect 20720 4626 20772 4632
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20916 4078 20944 4558
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20810 3632 20866 3641
rect 21100 3602 21128 9143
rect 21192 7698 21220 10390
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21284 9518 21312 9862
rect 21272 9512 21324 9518
rect 21272 9454 21324 9460
rect 21284 7886 21312 9454
rect 21376 9178 21404 11018
rect 21468 9586 21496 12582
rect 21560 11898 21588 12854
rect 21652 12442 21680 15302
rect 21732 14816 21784 14822
rect 21730 14784 21732 14793
rect 21784 14784 21786 14793
rect 21730 14719 21786 14728
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 21744 14074 21772 14214
rect 21732 14068 21784 14074
rect 21732 14010 21784 14016
rect 21836 13376 21864 17983
rect 22020 17814 22048 18226
rect 22008 17808 22060 17814
rect 22008 17750 22060 17756
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21928 15434 21956 16458
rect 22020 15570 22048 17614
rect 22112 17218 22140 19230
rect 22204 17882 22232 19306
rect 22192 17876 22244 17882
rect 22192 17818 22244 17824
rect 22190 17504 22246 17513
rect 22190 17439 22246 17448
rect 22204 17338 22232 17439
rect 22192 17332 22244 17338
rect 22192 17274 22244 17280
rect 22112 17190 22232 17218
rect 22098 17096 22154 17105
rect 22098 17031 22100 17040
rect 22152 17031 22154 17040
rect 22100 17002 22152 17008
rect 22100 16652 22152 16658
rect 22100 16594 22152 16600
rect 22112 16114 22140 16594
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 21916 15428 21968 15434
rect 21916 15370 21968 15376
rect 21916 14884 21968 14890
rect 21916 14826 21968 14832
rect 21928 14634 21956 14826
rect 21928 14606 22140 14634
rect 21916 14476 21968 14482
rect 21968 14436 22048 14464
rect 21916 14418 21968 14424
rect 21916 14272 21968 14278
rect 21916 14214 21968 14220
rect 21928 13938 21956 14214
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 22020 13802 22048 14436
rect 22112 14414 22140 14606
rect 22100 14408 22152 14414
rect 22100 14350 22152 14356
rect 22008 13796 22060 13802
rect 22008 13738 22060 13744
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 21744 13348 21864 13376
rect 21744 12442 21772 13348
rect 21928 13274 21956 13466
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 21928 13246 22048 13274
rect 22020 12850 22048 13246
rect 22008 12844 22060 12850
rect 22008 12786 22060 12792
rect 21914 12608 21970 12617
rect 21914 12543 21970 12552
rect 21640 12436 21692 12442
rect 21640 12378 21692 12384
rect 21732 12436 21784 12442
rect 21732 12378 21784 12384
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21640 12096 21692 12102
rect 21640 12038 21692 12044
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 21456 9580 21508 9586
rect 21456 9522 21508 9528
rect 21652 9518 21680 12038
rect 21744 11626 21772 12106
rect 21824 12096 21876 12102
rect 21824 12038 21876 12044
rect 21836 11694 21864 12038
rect 21928 11937 21956 12543
rect 21914 11928 21970 11937
rect 21914 11863 21970 11872
rect 22112 11830 22140 13330
rect 22204 13326 22232 17190
rect 22296 16522 22324 19808
rect 22376 19712 22428 19718
rect 22376 19654 22428 19660
rect 22388 19553 22416 19654
rect 22374 19544 22430 19553
rect 22374 19479 22430 19488
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22388 18970 22416 19314
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22480 18272 22508 20334
rect 22572 18601 22600 20742
rect 22664 19417 22692 22034
rect 22744 21888 22796 21894
rect 22744 21830 22796 21836
rect 22756 21321 22784 21830
rect 22742 21312 22798 21321
rect 22742 21247 22798 21256
rect 22744 20800 22796 20806
rect 22744 20742 22796 20748
rect 22756 20398 22784 20742
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22848 20346 22876 24126
rect 22940 23662 22968 24262
rect 23296 23792 23348 23798
rect 23296 23734 23348 23740
rect 22928 23656 22980 23662
rect 22928 23598 22980 23604
rect 22950 23420 23258 23429
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23308 23186 23336 23734
rect 23388 23588 23440 23594
rect 23388 23530 23440 23536
rect 23296 23180 23348 23186
rect 23296 23122 23348 23128
rect 23308 23050 23336 23122
rect 23296 23044 23348 23050
rect 23296 22986 23348 22992
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 23124 21418 23152 22102
rect 23308 21690 23336 22986
rect 23400 22710 23428 23530
rect 23388 22704 23440 22710
rect 23388 22646 23440 22652
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 23400 21486 23428 22646
rect 23492 22574 23520 24958
rect 23754 23352 23810 23361
rect 23860 23322 23888 26302
rect 24122 26200 24178 27000
rect 24766 26330 24822 27000
rect 24228 26302 24822 26330
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23754 23287 23810 23296
rect 23848 23316 23900 23322
rect 23664 23112 23716 23118
rect 23664 23054 23716 23060
rect 23676 22710 23704 23054
rect 23664 22704 23716 22710
rect 23664 22646 23716 22652
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23662 22400 23718 22409
rect 23662 22335 23718 22344
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23388 21480 23440 21486
rect 23584 21468 23612 21966
rect 23676 21622 23704 22335
rect 23664 21616 23716 21622
rect 23664 21558 23716 21564
rect 23664 21480 23716 21486
rect 23388 21422 23440 21428
rect 23492 21440 23664 21468
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23296 21412 23348 21418
rect 23296 21354 23348 21360
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23204 20936 23256 20942
rect 23204 20878 23256 20884
rect 23216 20806 23244 20878
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 22848 20318 22968 20346
rect 22940 20262 22968 20318
rect 22836 20256 22888 20262
rect 22742 20224 22798 20233
rect 22836 20198 22888 20204
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22742 20159 22798 20168
rect 22756 19553 22784 20159
rect 22742 19544 22798 19553
rect 22742 19479 22798 19488
rect 22650 19408 22706 19417
rect 22650 19343 22706 19352
rect 22664 19174 22692 19343
rect 22744 19304 22796 19310
rect 22744 19246 22796 19252
rect 22848 19258 22876 20198
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23112 19984 23164 19990
rect 23112 19926 23164 19932
rect 23124 19417 23152 19926
rect 23308 19514 23336 21354
rect 23492 21298 23520 21440
rect 23664 21422 23716 21428
rect 23768 21332 23796 23287
rect 23848 23258 23900 23264
rect 23952 22574 23980 25162
rect 24136 23254 24164 26200
rect 24124 23248 24176 23254
rect 24124 23190 24176 23196
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24136 22817 24164 22918
rect 24122 22808 24178 22817
rect 24122 22743 24178 22752
rect 23940 22568 23992 22574
rect 23940 22510 23992 22516
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 23940 22092 23992 22098
rect 23400 21270 23520 21298
rect 23676 21304 23796 21332
rect 23860 22052 23940 22080
rect 23400 20788 23428 21270
rect 23478 21176 23534 21185
rect 23478 21111 23480 21120
rect 23532 21111 23534 21120
rect 23572 21140 23624 21146
rect 23480 21082 23532 21088
rect 23572 21082 23624 21088
rect 23584 21010 23612 21082
rect 23572 21004 23624 21010
rect 23572 20946 23624 20952
rect 23572 20868 23624 20874
rect 23676 20856 23704 21304
rect 23624 20828 23704 20856
rect 23754 20904 23810 20913
rect 23754 20839 23810 20848
rect 23572 20810 23624 20816
rect 23480 20800 23532 20806
rect 23400 20760 23480 20788
rect 23480 20742 23532 20748
rect 23570 20632 23626 20641
rect 23570 20567 23572 20576
rect 23624 20567 23626 20576
rect 23572 20538 23624 20544
rect 23572 20460 23624 20466
rect 23572 20402 23624 20408
rect 23388 20324 23440 20330
rect 23388 20266 23440 20272
rect 23296 19508 23348 19514
rect 23296 19450 23348 19456
rect 22926 19408 22982 19417
rect 22926 19343 22928 19352
rect 22980 19343 22982 19352
rect 23110 19408 23166 19417
rect 23110 19343 23166 19352
rect 22928 19314 22980 19320
rect 22652 19168 22704 19174
rect 22652 19110 22704 19116
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22558 18592 22614 18601
rect 22558 18527 22614 18536
rect 22558 18456 22614 18465
rect 22558 18391 22614 18400
rect 22388 18244 22508 18272
rect 22284 16516 22336 16522
rect 22284 16458 22336 16464
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22296 15978 22324 16118
rect 22284 15972 22336 15978
rect 22284 15914 22336 15920
rect 22284 15564 22336 15570
rect 22284 15506 22336 15512
rect 22296 15026 22324 15506
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22296 14482 22324 14962
rect 22284 14476 22336 14482
rect 22284 14418 22336 14424
rect 22284 14340 22336 14346
rect 22284 14282 22336 14288
rect 22296 14074 22324 14282
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22192 13320 22244 13326
rect 22192 13262 22244 13268
rect 22204 12986 22232 13262
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22388 12866 22416 18244
rect 22468 18148 22520 18154
rect 22468 18090 22520 18096
rect 22480 17882 22508 18090
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22480 17338 22508 17478
rect 22468 17332 22520 17338
rect 22468 17274 22520 17280
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22480 16658 22508 17070
rect 22572 16794 22600 18391
rect 22664 18358 22692 18634
rect 22756 18630 22784 19246
rect 22848 19230 23336 19258
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22744 18624 22796 18630
rect 22744 18566 22796 18572
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22756 17105 22784 18566
rect 22742 17096 22798 17105
rect 22742 17031 22798 17040
rect 22744 16992 22796 16998
rect 22744 16934 22796 16940
rect 22560 16788 22612 16794
rect 22560 16730 22612 16736
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22756 16522 22784 16934
rect 22848 16708 22876 19110
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 23308 18442 23336 19230
rect 23400 18970 23428 20266
rect 23480 19508 23532 19514
rect 23480 19450 23532 19456
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23308 18414 23428 18442
rect 23296 18352 23348 18358
rect 23296 18294 23348 18300
rect 23112 18284 23164 18290
rect 23112 18226 23164 18232
rect 23124 18086 23152 18226
rect 23112 18080 23164 18086
rect 23112 18022 23164 18028
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23202 17776 23258 17785
rect 23202 17711 23258 17720
rect 23216 17338 23244 17711
rect 23204 17332 23256 17338
rect 23204 17274 23256 17280
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22848 16680 23060 16708
rect 22744 16516 22796 16522
rect 22744 16458 22796 16464
rect 22468 16448 22520 16454
rect 22468 16390 22520 16396
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22480 14278 22508 16390
rect 22650 16280 22706 16289
rect 22650 16215 22706 16224
rect 22560 15904 22612 15910
rect 22560 15846 22612 15852
rect 22572 15434 22600 15846
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22560 14952 22612 14958
rect 22560 14894 22612 14900
rect 22572 14618 22600 14894
rect 22560 14612 22612 14618
rect 22560 14554 22612 14560
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22468 14068 22520 14074
rect 22468 14010 22520 14016
rect 22480 13977 22508 14010
rect 22560 14000 22612 14006
rect 22466 13968 22522 13977
rect 22664 13977 22692 16215
rect 22744 16040 22796 16046
rect 22744 15982 22796 15988
rect 22756 14074 22784 15982
rect 22744 14068 22796 14074
rect 22744 14010 22796 14016
rect 22560 13942 22612 13948
rect 22650 13968 22706 13977
rect 22466 13903 22522 13912
rect 22572 13841 22600 13942
rect 22650 13903 22706 13912
rect 22558 13832 22614 13841
rect 22558 13767 22614 13776
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22560 13456 22612 13462
rect 22560 13398 22612 13404
rect 22204 12838 22416 12866
rect 22008 11824 22060 11830
rect 22008 11766 22060 11772
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 21824 11688 21876 11694
rect 21824 11630 21876 11636
rect 21732 11620 21784 11626
rect 21732 11562 21784 11568
rect 21744 10742 21772 11562
rect 21732 10736 21784 10742
rect 21732 10678 21784 10684
rect 21744 9994 21772 10678
rect 21732 9988 21784 9994
rect 21732 9930 21784 9936
rect 21640 9512 21692 9518
rect 21640 9454 21692 9460
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21836 9110 21864 11630
rect 21916 11212 21968 11218
rect 21916 11154 21968 11160
rect 21824 9104 21876 9110
rect 21824 9046 21876 9052
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21192 7670 21312 7698
rect 21180 6656 21232 6662
rect 21180 6598 21232 6604
rect 21192 5846 21220 6598
rect 21284 6202 21312 7670
rect 21454 7576 21510 7585
rect 21454 7511 21456 7520
rect 21508 7511 21510 7520
rect 21548 7540 21600 7546
rect 21456 7482 21508 7488
rect 21548 7482 21600 7488
rect 21468 6322 21496 7482
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21284 6174 21496 6202
rect 21560 6186 21588 7482
rect 21744 6730 21772 8502
rect 21928 7410 21956 11154
rect 22020 10588 22048 11766
rect 22098 11656 22154 11665
rect 22098 11591 22100 11600
rect 22152 11591 22154 11600
rect 22100 11562 22152 11568
rect 22112 10742 22140 11562
rect 22100 10736 22152 10742
rect 22100 10678 22152 10684
rect 22020 10560 22140 10588
rect 22006 9072 22062 9081
rect 22006 9007 22062 9016
rect 22020 8974 22048 9007
rect 22008 8968 22060 8974
rect 22008 8910 22060 8916
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21732 6724 21784 6730
rect 21732 6666 21784 6672
rect 21180 5840 21232 5846
rect 21180 5782 21232 5788
rect 21192 5710 21220 5782
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21192 5370 21220 5646
rect 21180 5364 21232 5370
rect 21180 5306 21232 5312
rect 21272 5228 21324 5234
rect 21272 5170 21324 5176
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 20810 3567 20866 3576
rect 21088 3596 21140 3602
rect 20824 3194 20852 3567
rect 21088 3538 21140 3544
rect 20812 3188 20864 3194
rect 20812 3130 20864 3136
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20732 1698 20760 2314
rect 20720 1692 20772 1698
rect 20720 1634 20772 1640
rect 20352 1012 20404 1018
rect 20352 954 20404 960
rect 18880 264 18932 270
rect 18880 206 18932 212
rect 20074 0 20130 800
rect 20824 202 20852 2790
rect 20904 2372 20956 2378
rect 20904 2314 20956 2320
rect 20916 1902 20944 2314
rect 20904 1896 20956 1902
rect 20904 1838 20956 1844
rect 21192 882 21220 4966
rect 21180 876 21232 882
rect 21180 818 21232 824
rect 21284 610 21312 5170
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21376 3670 21404 4422
rect 21364 3664 21416 3670
rect 21364 3606 21416 3612
rect 21468 1222 21496 6174
rect 21548 6180 21600 6186
rect 21548 6122 21600 6128
rect 21914 4720 21970 4729
rect 21914 4655 21916 4664
rect 21968 4655 21970 4664
rect 21916 4626 21968 4632
rect 21640 3936 21692 3942
rect 21640 3878 21692 3884
rect 21652 3738 21680 3878
rect 22112 3777 22140 10560
rect 22204 7954 22232 12838
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22284 12708 22336 12714
rect 22284 12650 22336 12656
rect 22296 12617 22324 12650
rect 22282 12608 22338 12617
rect 22282 12543 22338 12552
rect 22284 11688 22336 11694
rect 22284 11630 22336 11636
rect 22296 11286 22324 11630
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22282 10160 22338 10169
rect 22282 10095 22338 10104
rect 22296 9994 22324 10095
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22282 9752 22338 9761
rect 22282 9687 22338 9696
rect 22296 8922 22324 9687
rect 22388 9110 22416 12718
rect 22468 12708 22520 12714
rect 22468 12650 22520 12656
rect 22480 12434 22508 12650
rect 22572 12646 22600 13398
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22480 12406 22600 12434
rect 22480 11762 22508 12406
rect 22572 12306 22600 12406
rect 22560 12300 22612 12306
rect 22560 12242 22612 12248
rect 22560 12164 22612 12170
rect 22560 12106 22612 12112
rect 22468 11756 22520 11762
rect 22468 11698 22520 11704
rect 22480 11218 22508 11698
rect 22468 11212 22520 11218
rect 22468 11154 22520 11160
rect 22468 10600 22520 10606
rect 22468 10542 22520 10548
rect 22376 9104 22428 9110
rect 22376 9046 22428 9052
rect 22296 8894 22416 8922
rect 22192 7948 22244 7954
rect 22192 7890 22244 7896
rect 22284 7472 22336 7478
rect 22284 7414 22336 7420
rect 22296 7002 22324 7414
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 22190 6896 22246 6905
rect 22190 6831 22246 6840
rect 22204 6322 22232 6831
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22204 4554 22232 5170
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 22098 3768 22154 3777
rect 21640 3732 21692 3738
rect 22098 3703 22154 3712
rect 21640 3674 21692 3680
rect 22100 3664 22152 3670
rect 22100 3606 22152 3612
rect 22006 2680 22062 2689
rect 22006 2615 22008 2624
rect 22060 2615 22062 2624
rect 22008 2586 22060 2592
rect 22112 2038 22140 3606
rect 22192 3052 22244 3058
rect 22192 2994 22244 3000
rect 22100 2032 22152 2038
rect 22100 1974 22152 1980
rect 22204 1358 22232 2994
rect 22388 2774 22416 8894
rect 22480 8634 22508 10542
rect 22572 9722 22600 12106
rect 22664 10810 22692 13670
rect 22756 11218 22784 13738
rect 22848 13512 22876 16390
rect 23032 15910 23060 16680
rect 23308 16590 23336 18294
rect 23400 18170 23428 18414
rect 23492 18272 23520 19450
rect 23584 19417 23612 20402
rect 23664 20256 23716 20262
rect 23664 20198 23716 20204
rect 23570 19408 23626 19417
rect 23570 19343 23626 19352
rect 23572 19168 23624 19174
rect 23676 19145 23704 20198
rect 23768 20097 23796 20839
rect 23754 20088 23810 20097
rect 23754 20023 23810 20032
rect 23860 19718 23888 22052
rect 23940 22034 23992 22040
rect 23940 21684 23992 21690
rect 23940 21626 23992 21632
rect 23952 21010 23980 21626
rect 24136 21434 24164 22510
rect 24044 21406 24164 21434
rect 23940 21004 23992 21010
rect 23940 20946 23992 20952
rect 23940 20528 23992 20534
rect 23940 20470 23992 20476
rect 23848 19712 23900 19718
rect 23848 19654 23900 19660
rect 23572 19110 23624 19116
rect 23662 19136 23718 19145
rect 23584 18986 23612 19110
rect 23662 19071 23718 19080
rect 23584 18958 23704 18986
rect 23572 18896 23624 18902
rect 23572 18838 23624 18844
rect 23584 18766 23612 18838
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23584 18340 23612 18702
rect 23676 18630 23704 18958
rect 23860 18834 23888 19654
rect 23848 18828 23900 18834
rect 23848 18770 23900 18776
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 18465 23888 18566
rect 23846 18456 23902 18465
rect 23846 18391 23902 18400
rect 23848 18352 23900 18358
rect 23584 18312 23704 18340
rect 23676 18306 23704 18312
rect 23676 18300 23848 18306
rect 23676 18294 23900 18300
rect 23676 18278 23888 18294
rect 23492 18244 23612 18272
rect 23400 18142 23520 18170
rect 23492 18086 23520 18142
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23400 17678 23428 18022
rect 23388 17672 23440 17678
rect 23388 17614 23440 17620
rect 23584 17524 23612 18244
rect 23952 17898 23980 20470
rect 24044 18057 24072 21406
rect 24124 21344 24176 21350
rect 24124 21286 24176 21292
rect 24136 20942 24164 21286
rect 24124 20936 24176 20942
rect 24124 20878 24176 20884
rect 24136 20602 24164 20878
rect 24124 20596 24176 20602
rect 24124 20538 24176 20544
rect 24124 19508 24176 19514
rect 24124 19450 24176 19456
rect 24136 19378 24164 19450
rect 24124 19372 24176 19378
rect 24124 19314 24176 19320
rect 24122 18320 24178 18329
rect 24122 18255 24178 18264
rect 24030 18048 24086 18057
rect 24030 17983 24086 17992
rect 24136 17921 24164 18255
rect 24122 17912 24178 17921
rect 23952 17870 24072 17898
rect 23664 17672 23716 17678
rect 23756 17672 23808 17678
rect 23664 17614 23716 17620
rect 23754 17640 23756 17649
rect 23808 17640 23810 17649
rect 23400 17496 23612 17524
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23202 16416 23258 16425
rect 23202 16351 23258 16360
rect 23216 16114 23244 16351
rect 23400 16182 23428 17496
rect 23676 17082 23704 17614
rect 23754 17575 23810 17584
rect 23768 17338 23796 17575
rect 23848 17536 23900 17542
rect 23846 17504 23848 17513
rect 23900 17504 23902 17513
rect 23846 17439 23902 17448
rect 23756 17332 23808 17338
rect 23756 17274 23808 17280
rect 23756 17196 23808 17202
rect 23808 17156 23888 17184
rect 23756 17138 23808 17144
rect 23676 17066 23796 17082
rect 23664 17060 23796 17066
rect 23716 17054 23796 17060
rect 23664 17002 23716 17008
rect 23480 16992 23532 16998
rect 23480 16934 23532 16940
rect 23492 16250 23520 16934
rect 23570 16824 23626 16833
rect 23570 16759 23572 16768
rect 23624 16759 23626 16768
rect 23664 16788 23716 16794
rect 23572 16730 23624 16736
rect 23664 16730 23716 16736
rect 23570 16280 23626 16289
rect 23480 16244 23532 16250
rect 23570 16215 23626 16224
rect 23480 16186 23532 16192
rect 23388 16176 23440 16182
rect 23388 16118 23440 16124
rect 23584 16114 23612 16215
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 23124 15910 23152 16050
rect 23020 15904 23072 15910
rect 23020 15846 23072 15852
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23216 14929 23244 15438
rect 23388 15360 23440 15366
rect 23388 15302 23440 15308
rect 23296 14952 23348 14958
rect 23202 14920 23258 14929
rect 23296 14894 23348 14900
rect 23202 14855 23258 14864
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 23308 14482 23336 14894
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23296 14340 23348 14346
rect 23296 14282 23348 14288
rect 22928 14272 22980 14278
rect 22928 14214 22980 14220
rect 23112 14272 23164 14278
rect 23112 14214 23164 14220
rect 22940 13734 22968 14214
rect 23124 13870 23152 14214
rect 23112 13864 23164 13870
rect 23112 13806 23164 13812
rect 23308 13802 23336 14282
rect 23296 13796 23348 13802
rect 23296 13738 23348 13744
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22848 13484 23152 13512
rect 23124 13326 23152 13484
rect 23112 13320 23164 13326
rect 23112 13262 23164 13268
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 22848 12102 22876 13194
rect 23308 12918 23336 13194
rect 23296 12912 23348 12918
rect 23296 12854 23348 12860
rect 23296 12776 23348 12782
rect 23296 12718 23348 12724
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 23308 12434 23336 12718
rect 23216 12406 23336 12434
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 23020 11824 23072 11830
rect 22834 11792 22890 11801
rect 23020 11766 23072 11772
rect 22834 11727 22890 11736
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22652 10804 22704 10810
rect 22652 10746 22704 10752
rect 22756 10062 22784 11154
rect 22848 10810 22876 11727
rect 23032 11540 23060 11766
rect 23216 11665 23244 12406
rect 23294 12336 23350 12345
rect 23294 12271 23350 12280
rect 23308 11801 23336 12271
rect 23294 11792 23350 11801
rect 23294 11727 23350 11736
rect 23202 11656 23258 11665
rect 23202 11591 23258 11600
rect 23032 11512 23336 11540
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 23308 11098 23336 11512
rect 23400 11218 23428 15302
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23492 14074 23520 14418
rect 23480 14068 23532 14074
rect 23480 14010 23532 14016
rect 23572 14068 23624 14074
rect 23572 14010 23624 14016
rect 23480 13728 23532 13734
rect 23480 13670 23532 13676
rect 23492 13394 23520 13670
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23480 13184 23532 13190
rect 23480 13126 23532 13132
rect 23388 11212 23440 11218
rect 23388 11154 23440 11160
rect 23492 11098 23520 13126
rect 23584 11150 23612 14010
rect 23676 13190 23704 16730
rect 23768 16436 23796 17054
rect 23860 16590 23888 17156
rect 23940 16652 23992 16658
rect 23940 16594 23992 16600
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23768 16408 23888 16436
rect 23756 15360 23808 15366
rect 23756 15302 23808 15308
rect 23768 14278 23796 15302
rect 23860 15094 23888 16408
rect 23952 16250 23980 16594
rect 23940 16244 23992 16250
rect 23940 16186 23992 16192
rect 23940 15564 23992 15570
rect 23940 15506 23992 15512
rect 23848 15088 23900 15094
rect 23848 15030 23900 15036
rect 23846 14376 23902 14385
rect 23846 14311 23902 14320
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23756 13728 23808 13734
rect 23756 13670 23808 13676
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23768 12434 23796 13670
rect 23860 12481 23888 14311
rect 23952 13870 23980 15506
rect 23940 13864 23992 13870
rect 23940 13806 23992 13812
rect 23676 12406 23796 12434
rect 23846 12472 23902 12481
rect 23846 12407 23902 12416
rect 23112 11076 23164 11082
rect 23112 11018 23164 11024
rect 23308 11070 23520 11098
rect 23572 11144 23624 11150
rect 23572 11086 23624 11092
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 23124 10674 23152 11018
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 23112 10668 23164 10674
rect 23112 10610 23164 10616
rect 22744 10056 22796 10062
rect 22744 9998 22796 10004
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22756 8498 22784 9862
rect 22744 8492 22796 8498
rect 22744 8434 22796 8440
rect 22848 7478 22876 10610
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 23308 10062 23336 11070
rect 23572 11008 23624 11014
rect 23572 10950 23624 10956
rect 23386 10840 23442 10849
rect 23386 10775 23442 10784
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23400 9738 23428 10775
rect 23308 9710 23428 9738
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 23112 7880 23164 7886
rect 23112 7822 23164 7828
rect 23124 7546 23152 7822
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 22836 7472 22888 7478
rect 22836 7414 22888 7420
rect 22848 7002 22876 7414
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22836 6996 22888 7002
rect 22836 6938 22888 6944
rect 23308 6905 23336 9710
rect 23584 9654 23612 10950
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23388 8492 23440 8498
rect 23388 8434 23440 8440
rect 23400 8090 23428 8434
rect 23388 8084 23440 8090
rect 23388 8026 23440 8032
rect 23294 6896 23350 6905
rect 23294 6831 23350 6840
rect 23020 6724 23072 6730
rect 23020 6666 23072 6672
rect 23204 6724 23256 6730
rect 23204 6666 23256 6672
rect 23032 6458 23060 6666
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23216 6361 23244 6666
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23202 6352 23258 6361
rect 22836 6316 22888 6322
rect 23308 6322 23336 6394
rect 23202 6287 23258 6296
rect 23296 6316 23348 6322
rect 22836 6258 22888 6264
rect 23296 6258 23348 6264
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22572 4690 22600 4966
rect 22848 4826 22876 6258
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 23308 5234 23336 6054
rect 23676 5302 23704 12406
rect 23754 12200 23810 12209
rect 23754 12135 23810 12144
rect 23768 9602 23796 12135
rect 23952 12084 23980 13806
rect 24044 13734 24072 17870
rect 24122 17847 24178 17856
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 24136 16794 24164 17070
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 24228 16674 24256 26302
rect 24766 26200 24822 26302
rect 25410 26200 25466 27000
rect 25964 26648 26016 26654
rect 25964 26590 26016 26596
rect 24306 25392 24362 25401
rect 24306 25327 24362 25336
rect 24320 20369 24348 25327
rect 24584 25084 24636 25090
rect 24584 25026 24636 25032
rect 24596 24886 24624 25026
rect 24584 24880 24636 24886
rect 24584 24822 24636 24828
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24492 24064 24544 24070
rect 24492 24006 24544 24012
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24504 23202 24532 24006
rect 24596 23497 24624 24006
rect 24582 23488 24638 23497
rect 24582 23423 24638 23432
rect 24504 23174 24624 23202
rect 24400 21888 24452 21894
rect 24400 21830 24452 21836
rect 24412 21350 24440 21830
rect 24490 21720 24546 21729
rect 24490 21655 24546 21664
rect 24400 21344 24452 21350
rect 24400 21286 24452 21292
rect 24504 20505 24532 21655
rect 24490 20496 24546 20505
rect 24490 20431 24546 20440
rect 24306 20360 24362 20369
rect 24306 20295 24362 20304
rect 24308 19712 24360 19718
rect 24308 19654 24360 19660
rect 24320 18698 24348 19654
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 24308 18692 24360 18698
rect 24308 18634 24360 18640
rect 24308 17876 24360 17882
rect 24308 17818 24360 17824
rect 24320 17542 24348 17818
rect 24308 17536 24360 17542
rect 24308 17478 24360 17484
rect 24320 17270 24348 17478
rect 24308 17264 24360 17270
rect 24308 17206 24360 17212
rect 24320 17105 24348 17206
rect 24412 17134 24440 19246
rect 24492 19168 24544 19174
rect 24492 19110 24544 19116
rect 24504 18193 24532 19110
rect 24490 18184 24546 18193
rect 24490 18119 24546 18128
rect 24400 17128 24452 17134
rect 24306 17096 24362 17105
rect 24400 17070 24452 17076
rect 24306 17031 24362 17040
rect 24228 16646 24532 16674
rect 24122 16416 24178 16425
rect 24122 16351 24178 16360
rect 24032 13728 24084 13734
rect 24032 13670 24084 13676
rect 24136 13512 24164 16351
rect 24504 15910 24532 16646
rect 24596 15994 24624 23174
rect 24688 22438 24716 24822
rect 24766 24440 24822 24449
rect 24766 24375 24768 24384
rect 24820 24375 24822 24384
rect 24768 24346 24820 24352
rect 24860 24336 24912 24342
rect 24860 24278 24912 24284
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24780 23746 24808 24142
rect 24872 23866 24900 24278
rect 25136 24268 25188 24274
rect 25136 24210 25188 24216
rect 25148 23905 25176 24210
rect 25134 23896 25190 23905
rect 24860 23860 24912 23866
rect 25134 23831 25190 23840
rect 24860 23802 24912 23808
rect 25044 23792 25096 23798
rect 24780 23718 24992 23746
rect 25044 23734 25096 23740
rect 24860 23656 24912 23662
rect 24860 23598 24912 23604
rect 24872 23526 24900 23598
rect 24860 23520 24912 23526
rect 24860 23462 24912 23468
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24780 22642 24808 23190
rect 24768 22636 24820 22642
rect 24768 22578 24820 22584
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24676 22432 24728 22438
rect 24676 22374 24728 22380
rect 24676 21412 24728 21418
rect 24676 21354 24728 21360
rect 24688 21185 24716 21354
rect 24674 21176 24730 21185
rect 24674 21111 24730 21120
rect 24780 21026 24808 22471
rect 24872 21185 24900 23258
rect 24964 23050 24992 23718
rect 24952 23044 25004 23050
rect 24952 22986 25004 22992
rect 24964 21706 24992 22986
rect 25056 22273 25084 23734
rect 25320 23248 25372 23254
rect 25320 23190 25372 23196
rect 25228 22704 25280 22710
rect 25228 22646 25280 22652
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25042 22264 25098 22273
rect 25042 22199 25098 22208
rect 25148 22137 25176 22578
rect 25134 22128 25190 22137
rect 25134 22063 25136 22072
rect 25188 22063 25190 22072
rect 25136 22034 25188 22040
rect 24964 21690 25084 21706
rect 24964 21684 25096 21690
rect 24964 21678 25044 21684
rect 25044 21626 25096 21632
rect 25134 21448 25190 21457
rect 25134 21383 25136 21392
rect 25188 21383 25190 21392
rect 25136 21354 25188 21360
rect 24858 21176 24914 21185
rect 24858 21111 24914 21120
rect 24780 20998 24900 21026
rect 25240 21010 25268 22646
rect 25332 22409 25360 23190
rect 25424 23089 25452 26200
rect 25976 24818 26004 26590
rect 26054 26330 26110 27000
rect 26698 26330 26754 27000
rect 26054 26302 26188 26330
rect 26054 26200 26110 26302
rect 26054 24848 26110 24857
rect 25964 24812 26016 24818
rect 26054 24783 26110 24792
rect 25964 24754 26016 24760
rect 25780 24676 25832 24682
rect 25780 24618 25832 24624
rect 25792 24410 25820 24618
rect 26068 24614 26096 24783
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25780 24404 25832 24410
rect 25780 24346 25832 24352
rect 25964 24404 26016 24410
rect 25964 24346 26016 24352
rect 25872 24064 25924 24070
rect 25872 24006 25924 24012
rect 25780 23180 25832 23186
rect 25780 23122 25832 23128
rect 25410 23080 25466 23089
rect 25410 23015 25466 23024
rect 25504 22976 25556 22982
rect 25504 22918 25556 22924
rect 25596 22976 25648 22982
rect 25792 22953 25820 23122
rect 25884 22982 25912 24006
rect 25976 23186 26004 24346
rect 26068 24274 26096 24550
rect 26056 24268 26108 24274
rect 26056 24210 26108 24216
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26068 23225 26096 23258
rect 26054 23216 26110 23225
rect 25964 23180 26016 23186
rect 26160 23202 26188 26302
rect 26698 26314 27016 26330
rect 26698 26308 27028 26314
rect 26698 26302 26976 26308
rect 26698 26200 26754 26302
rect 26976 26250 27028 26256
rect 26884 26240 26936 26246
rect 27342 26200 27398 27000
rect 27986 26330 28042 27000
rect 28264 26376 28316 26382
rect 27986 26324 28264 26330
rect 27986 26318 28316 26324
rect 27986 26302 28304 26318
rect 27986 26200 28042 26302
rect 28630 26200 28686 27000
rect 29274 26200 29330 27000
rect 29828 26784 29880 26790
rect 29828 26726 29880 26732
rect 26884 26182 26936 26188
rect 26240 25084 26292 25090
rect 26240 25026 26292 25032
rect 26252 24818 26280 25026
rect 26896 24993 26924 26182
rect 26882 24984 26938 24993
rect 26882 24919 26938 24928
rect 26976 24948 27028 24954
rect 26976 24890 27028 24896
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 26608 24676 26660 24682
rect 26608 24618 26660 24624
rect 26252 24274 26464 24290
rect 26252 24268 26476 24274
rect 26252 24262 26424 24268
rect 26252 24177 26280 24262
rect 26424 24210 26476 24216
rect 26238 24168 26294 24177
rect 26238 24103 26294 24112
rect 26422 24168 26478 24177
rect 26422 24103 26478 24112
rect 26332 24064 26384 24070
rect 26332 24006 26384 24012
rect 26344 23225 26372 24006
rect 26436 23662 26464 24103
rect 26516 24064 26568 24070
rect 26516 24006 26568 24012
rect 26424 23656 26476 23662
rect 26424 23598 26476 23604
rect 26330 23216 26386 23225
rect 26160 23174 26280 23202
rect 26054 23151 26110 23160
rect 25964 23122 26016 23128
rect 26148 23112 26200 23118
rect 26146 23080 26148 23089
rect 26200 23080 26202 23089
rect 26146 23015 26202 23024
rect 25872 22976 25924 22982
rect 25596 22918 25648 22924
rect 25778 22944 25834 22953
rect 25318 22400 25374 22409
rect 25318 22335 25374 22344
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25412 21888 25464 21894
rect 25412 21830 25464 21836
rect 25332 21554 25360 21830
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25424 21078 25452 21830
rect 25412 21072 25464 21078
rect 25412 21014 25464 21020
rect 24676 20800 24728 20806
rect 24674 20768 24676 20777
rect 24728 20768 24730 20777
rect 24674 20703 24730 20712
rect 24872 20262 24900 20998
rect 25136 21004 25188 21010
rect 25136 20946 25188 20952
rect 25228 21004 25280 21010
rect 25228 20946 25280 20952
rect 25320 21004 25372 21010
rect 25320 20946 25372 20952
rect 25148 20534 25176 20946
rect 25136 20528 25188 20534
rect 25136 20470 25188 20476
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24952 20052 25004 20058
rect 24952 19994 25004 20000
rect 24676 19712 24728 19718
rect 24676 19654 24728 19660
rect 24688 19446 24716 19654
rect 24860 19508 24912 19514
rect 24860 19450 24912 19456
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24676 18828 24728 18834
rect 24676 18770 24728 18776
rect 24688 18358 24716 18770
rect 24676 18352 24728 18358
rect 24676 18294 24728 18300
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17202 24716 17682
rect 24676 17196 24728 17202
rect 24676 17138 24728 17144
rect 24688 16114 24716 17138
rect 24780 16572 24808 18906
rect 24872 16726 24900 19450
rect 24964 19446 24992 19994
rect 25228 19916 25280 19922
rect 25228 19858 25280 19864
rect 25044 19712 25096 19718
rect 25044 19654 25096 19660
rect 24952 19440 25004 19446
rect 24952 19382 25004 19388
rect 24952 18692 25004 18698
rect 24952 18634 25004 18640
rect 24964 18465 24992 18634
rect 24950 18456 25006 18465
rect 24950 18391 25006 18400
rect 25056 16794 25084 19654
rect 25240 18714 25268 19858
rect 25332 19854 25360 20946
rect 25412 20256 25464 20262
rect 25412 20198 25464 20204
rect 25320 19848 25372 19854
rect 25320 19790 25372 19796
rect 25320 18964 25372 18970
rect 25320 18906 25372 18912
rect 25148 18686 25268 18714
rect 25148 18222 25176 18686
rect 25228 18624 25280 18630
rect 25332 18601 25360 18906
rect 25228 18566 25280 18572
rect 25318 18592 25374 18601
rect 25240 18290 25268 18566
rect 25318 18527 25374 18536
rect 25228 18284 25280 18290
rect 25228 18226 25280 18232
rect 25136 18216 25188 18222
rect 25136 18158 25188 18164
rect 25044 16788 25096 16794
rect 25044 16730 25096 16736
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 25136 16584 25188 16590
rect 24780 16544 24900 16572
rect 24768 16448 24820 16454
rect 24768 16390 24820 16396
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24780 16046 24808 16390
rect 24768 16040 24820 16046
rect 24596 15966 24716 15994
rect 24768 15982 24820 15988
rect 24400 15904 24452 15910
rect 24400 15846 24452 15852
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24216 15428 24268 15434
rect 24216 15370 24268 15376
rect 24228 15026 24256 15370
rect 24308 15088 24360 15094
rect 24308 15030 24360 15036
rect 24216 15020 24268 15026
rect 24216 14962 24268 14968
rect 24228 14793 24256 14962
rect 24214 14784 24270 14793
rect 24214 14719 24270 14728
rect 24216 14544 24268 14550
rect 24216 14486 24268 14492
rect 24228 14346 24256 14486
rect 24216 14340 24268 14346
rect 24216 14282 24268 14288
rect 24228 14074 24256 14282
rect 24320 14278 24348 15030
rect 24308 14272 24360 14278
rect 24308 14214 24360 14220
rect 24216 14068 24268 14074
rect 24216 14010 24268 14016
rect 24136 13484 24256 13512
rect 24228 13394 24256 13484
rect 24124 13388 24176 13394
rect 24124 13330 24176 13336
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24032 13184 24084 13190
rect 24032 13126 24084 13132
rect 24044 12186 24072 13126
rect 24136 12374 24164 13330
rect 24320 12850 24348 14214
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24320 12646 24348 12786
rect 24308 12640 24360 12646
rect 24308 12582 24360 12588
rect 24124 12368 24176 12374
rect 24124 12310 24176 12316
rect 24308 12300 24360 12306
rect 24308 12242 24360 12248
rect 24044 12158 24164 12186
rect 24032 12096 24084 12102
rect 23952 12056 24032 12084
rect 24032 12038 24084 12044
rect 23848 11552 23900 11558
rect 23846 11520 23848 11529
rect 23940 11552 23992 11558
rect 23900 11520 23902 11529
rect 23940 11494 23992 11500
rect 23846 11455 23902 11464
rect 23952 10674 23980 11494
rect 24044 10674 24072 12038
rect 24136 11014 24164 12158
rect 24216 11824 24268 11830
rect 24216 11766 24268 11772
rect 24228 11082 24256 11766
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24124 11008 24176 11014
rect 24124 10950 24176 10956
rect 24124 10736 24176 10742
rect 24124 10678 24176 10684
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23860 10198 23888 10406
rect 23848 10192 23900 10198
rect 23848 10134 23900 10140
rect 23768 9574 23888 9602
rect 23756 9444 23808 9450
rect 23756 9386 23808 9392
rect 23768 8634 23796 9386
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23756 7540 23808 7546
rect 23756 7482 23808 7488
rect 23768 6186 23796 7482
rect 23756 6180 23808 6186
rect 23756 6122 23808 6128
rect 23860 5914 23888 9574
rect 23952 8294 23980 10610
rect 24030 10296 24086 10305
rect 24030 10231 24086 10240
rect 24044 10062 24072 10231
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 24136 8634 24164 10678
rect 24216 10532 24268 10538
rect 24216 10474 24268 10480
rect 24228 10130 24256 10474
rect 24216 10124 24268 10130
rect 24216 10066 24268 10072
rect 24124 8628 24176 8634
rect 24124 8570 24176 8576
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24136 6662 24164 7686
rect 24124 6656 24176 6662
rect 24124 6598 24176 6604
rect 23848 5908 23900 5914
rect 23848 5850 23900 5856
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 23664 5296 23716 5302
rect 23664 5238 23716 5244
rect 23296 5228 23348 5234
rect 23296 5170 23348 5176
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22836 4820 22888 4826
rect 22836 4762 22888 4768
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22848 4214 22876 4762
rect 23768 4758 23796 5510
rect 24320 5166 24348 12242
rect 24412 12238 24440 15846
rect 24582 15192 24638 15201
rect 24582 15127 24638 15136
rect 24596 14929 24624 15127
rect 24582 14920 24638 14929
rect 24582 14855 24638 14864
rect 24490 14784 24546 14793
rect 24490 14719 24546 14728
rect 24504 14482 24532 14719
rect 24582 14648 24638 14657
rect 24582 14583 24638 14592
rect 24596 14550 24624 14583
rect 24584 14544 24636 14550
rect 24584 14486 24636 14492
rect 24492 14476 24544 14482
rect 24492 14418 24544 14424
rect 24400 12232 24452 12238
rect 24400 12174 24452 12180
rect 24504 8294 24532 14418
rect 24584 14408 24636 14414
rect 24584 14350 24636 14356
rect 24596 13938 24624 14350
rect 24584 13932 24636 13938
rect 24584 13874 24636 13880
rect 24584 13388 24636 13394
rect 24584 13330 24636 13336
rect 24596 12306 24624 13330
rect 24584 12300 24636 12306
rect 24584 12242 24636 12248
rect 24688 12170 24716 15966
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24780 15450 24808 15846
rect 24872 15570 24900 16544
rect 24950 16552 25006 16561
rect 25136 16526 25188 16532
rect 24950 16487 25006 16496
rect 24860 15564 24912 15570
rect 24860 15506 24912 15512
rect 24964 15484 24992 16487
rect 25148 16454 25176 16526
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 15706 25176 16390
rect 25136 15700 25188 15706
rect 25136 15642 25188 15648
rect 24964 15456 25176 15484
rect 24780 15422 24900 15450
rect 24872 15416 24900 15422
rect 24872 15388 25084 15416
rect 24768 15360 24820 15366
rect 24768 15302 24820 15308
rect 24780 15094 24808 15302
rect 24768 15088 24820 15094
rect 24768 15030 24820 15036
rect 24860 14816 24912 14822
rect 24860 14758 24912 14764
rect 24766 14376 24822 14385
rect 24766 14311 24822 14320
rect 24780 14278 24808 14311
rect 24768 14272 24820 14278
rect 24768 14214 24820 14220
rect 24780 13870 24808 14214
rect 24872 13870 24900 14758
rect 24952 14272 25004 14278
rect 24952 14214 25004 14220
rect 24964 14006 24992 14214
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 24768 13864 24820 13870
rect 24768 13806 24820 13812
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24952 13728 25004 13734
rect 24952 13670 25004 13676
rect 24964 13326 24992 13670
rect 24952 13320 25004 13326
rect 24952 13262 25004 13268
rect 24860 12708 24912 12714
rect 24860 12650 24912 12656
rect 24676 12164 24728 12170
rect 24676 12106 24728 12112
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24674 12064 24730 12073
rect 24596 11898 24624 12038
rect 24674 11999 24730 12008
rect 24584 11892 24636 11898
rect 24584 11834 24636 11840
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 11150 24624 11494
rect 24584 11144 24636 11150
rect 24584 11086 24636 11092
rect 24688 10198 24716 11999
rect 24872 11082 24900 12650
rect 24952 11824 25004 11830
rect 24952 11766 25004 11772
rect 24964 11626 24992 11766
rect 24952 11620 25004 11626
rect 24952 11562 25004 11568
rect 24860 11076 24912 11082
rect 24860 11018 24912 11024
rect 24766 10976 24822 10985
rect 24766 10911 24822 10920
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24412 8266 24532 8294
rect 24412 8090 24440 8266
rect 24400 8084 24452 8090
rect 24400 8026 24452 8032
rect 24780 7886 24808 10911
rect 25056 9110 25084 15388
rect 25148 13841 25176 15456
rect 25134 13832 25190 13841
rect 25240 13802 25268 18226
rect 25424 16833 25452 20198
rect 25516 19446 25544 22918
rect 25608 20641 25636 22918
rect 25872 22918 25924 22924
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 25778 22879 25834 22888
rect 25792 22681 25820 22879
rect 25778 22672 25834 22681
rect 25778 22607 25834 22616
rect 25780 22568 25832 22574
rect 25964 22568 26016 22574
rect 25780 22510 25832 22516
rect 25962 22536 25964 22545
rect 26016 22536 26018 22545
rect 25792 22409 25820 22510
rect 25962 22471 26018 22480
rect 25872 22432 25924 22438
rect 25778 22400 25834 22409
rect 25872 22374 25924 22380
rect 25778 22335 25834 22344
rect 25688 22160 25740 22166
rect 25688 22102 25740 22108
rect 25700 21434 25728 22102
rect 25778 21992 25834 22001
rect 25778 21927 25834 21936
rect 25792 21729 25820 21927
rect 25778 21720 25834 21729
rect 25778 21655 25834 21664
rect 25700 21406 25820 21434
rect 25688 21344 25740 21350
rect 25688 21286 25740 21292
rect 25700 20777 25728 21286
rect 25686 20768 25742 20777
rect 25686 20703 25742 20712
rect 25594 20632 25650 20641
rect 25792 20618 25820 21406
rect 25594 20567 25650 20576
rect 25700 20590 25820 20618
rect 25504 19440 25556 19446
rect 25504 19382 25556 19388
rect 25596 19372 25648 19378
rect 25596 19314 25648 19320
rect 25504 18964 25556 18970
rect 25504 18906 25556 18912
rect 25516 18442 25544 18906
rect 25608 18601 25636 19314
rect 25594 18592 25650 18601
rect 25594 18527 25650 18536
rect 25516 18414 25636 18442
rect 25504 18080 25556 18086
rect 25504 18022 25556 18028
rect 25410 16824 25466 16833
rect 25410 16759 25466 16768
rect 25320 16652 25372 16658
rect 25320 16594 25372 16600
rect 25332 14822 25360 16594
rect 25516 16454 25544 18022
rect 25412 16448 25464 16454
rect 25412 16390 25464 16396
rect 25504 16448 25556 16454
rect 25504 16390 25556 16396
rect 25424 15502 25452 16390
rect 25502 16008 25558 16017
rect 25502 15943 25558 15952
rect 25412 15496 25464 15502
rect 25412 15438 25464 15444
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25516 14634 25544 15943
rect 25608 15337 25636 18414
rect 25700 16640 25728 20590
rect 25780 19848 25832 19854
rect 25780 19790 25832 19796
rect 25792 19310 25820 19790
rect 25780 19304 25832 19310
rect 25780 19246 25832 19252
rect 25792 18834 25820 19246
rect 25884 18834 25912 22374
rect 26068 22098 26096 22918
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 26056 22092 26108 22098
rect 26056 22034 26108 22040
rect 26054 21992 26110 22001
rect 25964 21956 26016 21962
rect 26054 21927 26110 21936
rect 25964 21898 26016 21904
rect 25976 20942 26004 21898
rect 26068 21622 26096 21927
rect 26160 21622 26188 22170
rect 26252 22137 26280 23174
rect 26330 23151 26386 23160
rect 26332 22432 26384 22438
rect 26332 22374 26384 22380
rect 26238 22128 26294 22137
rect 26238 22063 26294 22072
rect 26344 21962 26372 22374
rect 26422 22128 26478 22137
rect 26422 22063 26478 22072
rect 26332 21956 26384 21962
rect 26332 21898 26384 21904
rect 26240 21888 26292 21894
rect 26240 21830 26292 21836
rect 26056 21616 26108 21622
rect 26056 21558 26108 21564
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 25964 20936 26016 20942
rect 25964 20878 26016 20884
rect 25780 18828 25832 18834
rect 25780 18770 25832 18776
rect 25872 18828 25924 18834
rect 25872 18770 25924 18776
rect 25792 17746 25820 18770
rect 25976 18358 26004 20878
rect 26252 20874 26280 21830
rect 26436 20913 26464 22063
rect 26528 21418 26556 24006
rect 26620 23594 26648 24618
rect 26790 24032 26846 24041
rect 26790 23967 26846 23976
rect 26608 23588 26660 23594
rect 26608 23530 26660 23536
rect 26620 23361 26648 23530
rect 26606 23352 26662 23361
rect 26606 23287 26662 23296
rect 26700 23248 26752 23254
rect 26700 23190 26752 23196
rect 26712 23050 26740 23190
rect 26700 23044 26752 23050
rect 26700 22986 26752 22992
rect 26606 22672 26662 22681
rect 26606 22607 26662 22616
rect 26620 22137 26648 22607
rect 26606 22128 26662 22137
rect 26606 22063 26662 22072
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26608 21412 26660 21418
rect 26608 21354 26660 21360
rect 26422 20904 26478 20913
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26240 20868 26292 20874
rect 26422 20839 26478 20848
rect 26240 20810 26292 20816
rect 26160 20754 26188 20810
rect 26160 20726 26280 20754
rect 26252 18834 26280 20726
rect 26528 20466 26556 21354
rect 26620 20534 26648 21354
rect 26804 20602 26832 23967
rect 26884 22976 26936 22982
rect 26988 22953 27016 24890
rect 27160 24336 27212 24342
rect 27158 24304 27160 24313
rect 27212 24304 27214 24313
rect 27158 24239 27214 24248
rect 27252 24132 27304 24138
rect 27252 24074 27304 24080
rect 27068 23792 27120 23798
rect 27068 23734 27120 23740
rect 26884 22918 26936 22924
rect 26974 22944 27030 22953
rect 26896 22681 26924 22918
rect 26974 22879 27030 22888
rect 26882 22672 26938 22681
rect 26882 22607 26938 22616
rect 26896 22438 26924 22607
rect 26884 22432 26936 22438
rect 26884 22374 26936 22380
rect 26792 20596 26844 20602
rect 26792 20538 26844 20544
rect 26608 20528 26660 20534
rect 26608 20470 26660 20476
rect 26516 20460 26568 20466
rect 26516 20402 26568 20408
rect 26620 19786 26648 20470
rect 26608 19780 26660 19786
rect 26608 19722 26660 19728
rect 26516 19168 26568 19174
rect 26514 19136 26516 19145
rect 26568 19136 26570 19145
rect 26514 19071 26570 19080
rect 26148 18828 26200 18834
rect 26148 18770 26200 18776
rect 26240 18828 26292 18834
rect 26240 18770 26292 18776
rect 26054 18728 26110 18737
rect 26054 18663 26110 18672
rect 25964 18352 26016 18358
rect 25964 18294 26016 18300
rect 25780 17740 25832 17746
rect 25780 17682 25832 17688
rect 26068 17660 26096 18663
rect 26160 18358 26188 18770
rect 26620 18714 26648 19722
rect 26698 19680 26754 19689
rect 26698 19615 26754 19624
rect 26252 18698 26648 18714
rect 26240 18692 26648 18698
rect 26292 18686 26648 18692
rect 26240 18634 26292 18640
rect 26148 18352 26200 18358
rect 26148 18294 26200 18300
rect 26148 18216 26200 18222
rect 26148 18158 26200 18164
rect 26160 17814 26188 18158
rect 26516 18148 26568 18154
rect 26516 18090 26568 18096
rect 26422 17912 26478 17921
rect 26422 17847 26478 17856
rect 26148 17808 26200 17814
rect 26148 17750 26200 17756
rect 26068 17632 26188 17660
rect 26160 17218 26188 17632
rect 26160 17190 26280 17218
rect 26148 17128 26200 17134
rect 26148 17070 26200 17076
rect 25700 16612 26004 16640
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25780 16448 25832 16454
rect 25780 16390 25832 16396
rect 25700 15570 25728 16390
rect 25688 15564 25740 15570
rect 25688 15506 25740 15512
rect 25594 15328 25650 15337
rect 25594 15263 25650 15272
rect 25332 14606 25544 14634
rect 25134 13767 25190 13776
rect 25228 13796 25280 13802
rect 25228 13738 25280 13744
rect 25136 13388 25188 13394
rect 25136 13330 25188 13336
rect 25148 11830 25176 13330
rect 25240 12918 25268 13738
rect 25228 12912 25280 12918
rect 25228 12854 25280 12860
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25240 11830 25268 12378
rect 25136 11824 25188 11830
rect 25136 11766 25188 11772
rect 25228 11824 25280 11830
rect 25228 11766 25280 11772
rect 25136 11348 25188 11354
rect 25136 11290 25188 11296
rect 25044 9104 25096 9110
rect 25044 9046 25096 9052
rect 24858 7984 24914 7993
rect 24858 7919 24860 7928
rect 24912 7919 24914 7928
rect 24860 7890 24912 7896
rect 24768 7880 24820 7886
rect 24768 7822 24820 7828
rect 24860 7812 24912 7818
rect 24860 7754 24912 7760
rect 24872 7342 24900 7754
rect 24860 7336 24912 7342
rect 24398 7304 24454 7313
rect 24860 7278 24912 7284
rect 24398 7239 24400 7248
rect 24452 7239 24454 7248
rect 24400 7210 24452 7216
rect 24952 5636 25004 5642
rect 24952 5578 25004 5584
rect 24964 5302 24992 5578
rect 24952 5296 25004 5302
rect 24952 5238 25004 5244
rect 24308 5160 24360 5166
rect 24308 5102 24360 5108
rect 23756 4752 23808 4758
rect 23756 4694 23808 4700
rect 23480 4616 23532 4622
rect 23480 4558 23532 4564
rect 22836 4208 22888 4214
rect 22836 4150 22888 4156
rect 23492 3942 23520 4558
rect 25148 4282 25176 11290
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25240 9586 25268 10610
rect 25332 10062 25360 14606
rect 25502 14512 25558 14521
rect 25502 14447 25558 14456
rect 25516 14414 25544 14447
rect 25504 14408 25556 14414
rect 25700 14362 25728 15506
rect 25504 14350 25556 14356
rect 25410 14104 25466 14113
rect 25516 14074 25544 14350
rect 25608 14334 25728 14362
rect 25410 14039 25466 14048
rect 25504 14068 25556 14074
rect 25424 13954 25452 14039
rect 25504 14010 25556 14016
rect 25608 13954 25636 14334
rect 25688 14272 25740 14278
rect 25686 14240 25688 14249
rect 25740 14240 25742 14249
rect 25686 14175 25742 14184
rect 25700 14074 25728 14175
rect 25688 14068 25740 14074
rect 25688 14010 25740 14016
rect 25424 13926 25544 13954
rect 25608 13926 25728 13954
rect 25410 13832 25466 13841
rect 25410 13767 25466 13776
rect 25424 11200 25452 13767
rect 25516 11354 25544 13926
rect 25596 13864 25648 13870
rect 25596 13806 25648 13812
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25424 11172 25544 11200
rect 25410 11112 25466 11121
rect 25410 11047 25466 11056
rect 25424 11014 25452 11047
rect 25412 11008 25464 11014
rect 25412 10950 25464 10956
rect 25320 10056 25372 10062
rect 25320 9998 25372 10004
rect 25228 9580 25280 9586
rect 25228 9522 25280 9528
rect 25320 9580 25372 9586
rect 25320 9522 25372 9528
rect 25228 8832 25280 8838
rect 25228 8774 25280 8780
rect 25240 6254 25268 8774
rect 25332 8022 25360 9522
rect 25516 8090 25544 11172
rect 25608 10742 25636 13806
rect 25596 10736 25648 10742
rect 25596 10678 25648 10684
rect 25700 9058 25728 13926
rect 25608 9030 25728 9058
rect 25504 8084 25556 8090
rect 25504 8026 25556 8032
rect 25320 8016 25372 8022
rect 25320 7958 25372 7964
rect 25608 7954 25636 9030
rect 25688 8968 25740 8974
rect 25688 8910 25740 8916
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25608 7818 25636 7890
rect 25596 7812 25648 7818
rect 25596 7754 25648 7760
rect 25700 7546 25728 8910
rect 25688 7540 25740 7546
rect 25688 7482 25740 7488
rect 25792 7206 25820 16390
rect 25872 14816 25924 14822
rect 25872 14758 25924 14764
rect 25884 14482 25912 14758
rect 25872 14476 25924 14482
rect 25872 14418 25924 14424
rect 25976 13802 26004 16612
rect 26160 15978 26188 17070
rect 26252 16561 26280 17190
rect 26238 16552 26294 16561
rect 26238 16487 26294 16496
rect 26436 16425 26464 17847
rect 26528 16658 26556 18090
rect 26608 16720 26660 16726
rect 26608 16662 26660 16668
rect 26516 16652 26568 16658
rect 26516 16594 26568 16600
rect 26620 16454 26648 16662
rect 26608 16448 26660 16454
rect 26422 16416 26478 16425
rect 26608 16390 26660 16396
rect 26422 16351 26478 16360
rect 26712 16182 26740 19615
rect 26804 19446 26832 20538
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26792 19236 26844 19242
rect 26792 19178 26844 19184
rect 26804 18902 26832 19178
rect 26792 18896 26844 18902
rect 26792 18838 26844 18844
rect 26790 18320 26846 18329
rect 26790 18255 26846 18264
rect 26804 17678 26832 18255
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26804 17202 26832 17614
rect 26896 17218 26924 22374
rect 27080 21962 27108 23734
rect 27264 23526 27292 24074
rect 27160 23520 27212 23526
rect 27160 23462 27212 23468
rect 27252 23520 27304 23526
rect 27356 23497 27384 26200
rect 28356 24744 28408 24750
rect 28356 24686 28408 24692
rect 27540 24274 27752 24290
rect 27540 24268 27764 24274
rect 27540 24262 27712 24268
rect 27436 24132 27488 24138
rect 27436 24074 27488 24080
rect 27448 23662 27476 24074
rect 27436 23656 27488 23662
rect 27436 23598 27488 23604
rect 27252 23462 27304 23468
rect 27342 23488 27398 23497
rect 27172 23186 27200 23462
rect 27342 23423 27398 23432
rect 27540 23361 27568 24262
rect 27712 24210 27764 24216
rect 27804 24268 27856 24274
rect 27804 24210 27856 24216
rect 27816 24041 27844 24210
rect 28368 24206 28396 24686
rect 28356 24200 28408 24206
rect 28356 24142 28408 24148
rect 27802 24032 27858 24041
rect 27802 23967 27858 23976
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27802 23896 27858 23905
rect 27950 23899 28258 23908
rect 27802 23831 27858 23840
rect 27712 23792 27764 23798
rect 27816 23780 27844 23831
rect 27816 23752 27936 23780
rect 27712 23734 27764 23740
rect 27724 23644 27752 23734
rect 27804 23656 27856 23662
rect 27724 23616 27804 23644
rect 27526 23352 27582 23361
rect 27526 23287 27582 23296
rect 27252 23248 27304 23254
rect 27540 23236 27568 23287
rect 27304 23208 27568 23236
rect 27252 23190 27304 23196
rect 27160 23180 27212 23186
rect 27160 23122 27212 23128
rect 27172 22710 27200 23122
rect 27724 23050 27752 23616
rect 27804 23598 27856 23604
rect 27802 23488 27858 23497
rect 27802 23423 27858 23432
rect 27712 23044 27764 23050
rect 27712 22986 27764 22992
rect 27434 22944 27490 22953
rect 27434 22879 27490 22888
rect 27250 22808 27306 22817
rect 27250 22743 27306 22752
rect 27160 22704 27212 22710
rect 27160 22646 27212 22652
rect 27160 22568 27212 22574
rect 27160 22510 27212 22516
rect 27172 21978 27200 22510
rect 27264 22234 27292 22743
rect 27252 22228 27304 22234
rect 27252 22170 27304 22176
rect 27344 22024 27396 22030
rect 27172 21972 27344 21978
rect 27172 21966 27396 21972
rect 27068 21956 27120 21962
rect 27068 21898 27120 21904
rect 27172 21950 27384 21966
rect 26974 21584 27030 21593
rect 26974 21519 27030 21528
rect 26988 21049 27016 21519
rect 27080 21418 27108 21898
rect 27068 21412 27120 21418
rect 27068 21354 27120 21360
rect 27066 21176 27122 21185
rect 27066 21111 27122 21120
rect 26974 21040 27030 21049
rect 26974 20975 27030 20984
rect 26976 20528 27028 20534
rect 26976 20470 27028 20476
rect 26988 17678 27016 20470
rect 27080 18329 27108 21111
rect 27172 20534 27200 21950
rect 27448 21842 27476 22879
rect 27618 22672 27674 22681
rect 27618 22607 27620 22616
rect 27672 22607 27674 22616
rect 27620 22578 27672 22584
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 27528 22500 27580 22506
rect 27528 22442 27580 22448
rect 27540 22098 27568 22442
rect 27724 22409 27752 22510
rect 27710 22400 27766 22409
rect 27710 22335 27766 22344
rect 27816 22250 27844 23423
rect 27908 22964 27936 23752
rect 27908 22936 28396 22964
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27724 22222 27844 22250
rect 27896 22228 27948 22234
rect 27528 22092 27580 22098
rect 27528 22034 27580 22040
rect 27356 21814 27476 21842
rect 27620 21888 27672 21894
rect 27620 21830 27672 21836
rect 27356 21593 27384 21814
rect 27528 21684 27580 21690
rect 27528 21626 27580 21632
rect 27342 21584 27398 21593
rect 27540 21554 27568 21626
rect 27342 21519 27398 21528
rect 27436 21548 27488 21554
rect 27436 21490 27488 21496
rect 27528 21548 27580 21554
rect 27528 21490 27580 21496
rect 27344 21412 27396 21418
rect 27344 21354 27396 21360
rect 27252 21344 27304 21350
rect 27252 21286 27304 21292
rect 27264 21146 27292 21286
rect 27252 21140 27304 21146
rect 27252 21082 27304 21088
rect 27356 20942 27384 21354
rect 27448 21078 27476 21490
rect 27528 21344 27580 21350
rect 27528 21286 27580 21292
rect 27436 21072 27488 21078
rect 27436 21014 27488 21020
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 27540 20806 27568 21286
rect 27528 20800 27580 20806
rect 27528 20742 27580 20748
rect 27436 20596 27488 20602
rect 27436 20538 27488 20544
rect 27160 20528 27212 20534
rect 27160 20470 27212 20476
rect 27448 20398 27476 20538
rect 27436 20392 27488 20398
rect 27436 20334 27488 20340
rect 27252 20324 27304 20330
rect 27252 20266 27304 20272
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27172 20058 27200 20198
rect 27160 20052 27212 20058
rect 27160 19994 27212 20000
rect 27160 19712 27212 19718
rect 27160 19654 27212 19660
rect 27172 18630 27200 19654
rect 27160 18624 27212 18630
rect 27160 18566 27212 18572
rect 27066 18320 27122 18329
rect 27066 18255 27122 18264
rect 27160 18216 27212 18222
rect 27160 18158 27212 18164
rect 27068 18080 27120 18086
rect 27068 18022 27120 18028
rect 26976 17672 27028 17678
rect 26976 17614 27028 17620
rect 27080 17610 27108 18022
rect 27068 17604 27120 17610
rect 27068 17546 27120 17552
rect 27080 17270 27108 17546
rect 27068 17264 27120 17270
rect 26792 17196 26844 17202
rect 26896 17190 27016 17218
rect 27068 17206 27120 17212
rect 26792 17138 26844 17144
rect 26804 16658 26832 17138
rect 26792 16652 26844 16658
rect 26792 16594 26844 16600
rect 26790 16552 26846 16561
rect 26790 16487 26846 16496
rect 26700 16176 26752 16182
rect 26700 16118 26752 16124
rect 26148 15972 26200 15978
rect 26148 15914 26200 15920
rect 26608 15564 26660 15570
rect 26608 15506 26660 15512
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 25964 13796 26016 13802
rect 25964 13738 26016 13744
rect 26056 13456 26108 13462
rect 26056 13398 26108 13404
rect 26068 12986 26096 13398
rect 26344 13274 26372 15302
rect 26422 15192 26478 15201
rect 26422 15127 26478 15136
rect 26436 14074 26464 15127
rect 26620 14822 26648 15506
rect 26608 14816 26660 14822
rect 26608 14758 26660 14764
rect 26516 14272 26568 14278
rect 26516 14214 26568 14220
rect 26424 14068 26476 14074
rect 26424 14010 26476 14016
rect 26160 13246 26372 13274
rect 26160 13190 26188 13246
rect 26528 13190 26556 14214
rect 26620 13938 26648 14758
rect 26804 14550 26832 16487
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26792 14544 26844 14550
rect 26792 14486 26844 14492
rect 26700 14476 26752 14482
rect 26700 14418 26752 14424
rect 26712 14278 26740 14418
rect 26700 14272 26752 14278
rect 26700 14214 26752 14220
rect 26608 13932 26660 13938
rect 26608 13874 26660 13880
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26148 13184 26200 13190
rect 26148 13126 26200 13132
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26056 12980 26108 12986
rect 26056 12922 26108 12928
rect 25964 12912 26016 12918
rect 25964 12854 26016 12860
rect 25872 11892 25924 11898
rect 25872 11834 25924 11840
rect 25884 11626 25912 11834
rect 25872 11620 25924 11626
rect 25872 11562 25924 11568
rect 25976 11218 26004 12854
rect 26252 11762 26280 13126
rect 26514 12472 26570 12481
rect 26514 12407 26570 12416
rect 26240 11756 26292 11762
rect 26240 11698 26292 11704
rect 25964 11212 26016 11218
rect 25964 11154 26016 11160
rect 26146 10160 26202 10169
rect 26146 10095 26202 10104
rect 26056 9920 26108 9926
rect 26056 9862 26108 9868
rect 25870 8800 25926 8809
rect 25870 8735 25926 8744
rect 25780 7200 25832 7206
rect 25780 7142 25832 7148
rect 25320 6996 25372 7002
rect 25320 6938 25372 6944
rect 25228 6248 25280 6254
rect 25228 6190 25280 6196
rect 25136 4276 25188 4282
rect 25136 4218 25188 4224
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 22744 3120 22796 3126
rect 22744 3062 22796 3068
rect 22388 2746 22508 2774
rect 22192 1352 22244 1358
rect 22098 1320 22154 1329
rect 22192 1294 22244 1300
rect 22098 1255 22154 1264
rect 22112 1222 22140 1255
rect 22480 1222 22508 2746
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 22572 2446 22600 2586
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 21456 1216 21508 1222
rect 21456 1158 21508 1164
rect 22100 1216 22152 1222
rect 22100 1158 22152 1164
rect 22468 1216 22520 1222
rect 22468 1158 22520 1164
rect 22756 800 22784 3062
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 23386 2680 23442 2689
rect 23386 2615 23388 2624
rect 23440 2615 23442 2624
rect 23388 2586 23440 2592
rect 25332 1290 25360 6938
rect 25504 5092 25556 5098
rect 25504 5034 25556 5040
rect 25516 2650 25544 5034
rect 25884 2774 25912 8735
rect 25962 8664 26018 8673
rect 25962 8599 25964 8608
rect 26016 8599 26018 8608
rect 25964 8570 26016 8576
rect 26068 6390 26096 9862
rect 26160 9518 26188 10095
rect 26238 9616 26294 9625
rect 26238 9551 26294 9560
rect 26332 9580 26384 9586
rect 26148 9512 26200 9518
rect 26148 9454 26200 9460
rect 26252 9450 26280 9551
rect 26332 9522 26384 9528
rect 26240 9444 26292 9450
rect 26240 9386 26292 9392
rect 26344 9178 26372 9522
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26240 8900 26292 8906
rect 26240 8842 26292 8848
rect 26252 6458 26280 8842
rect 26528 8566 26556 12407
rect 26712 11286 26740 13262
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26700 11280 26752 11286
rect 26700 11222 26752 11228
rect 26700 11076 26752 11082
rect 26700 11018 26752 11024
rect 26712 9994 26740 11018
rect 26700 9988 26752 9994
rect 26700 9930 26752 9936
rect 26608 9920 26660 9926
rect 26608 9862 26660 9868
rect 26516 8560 26568 8566
rect 26516 8502 26568 8508
rect 26240 6452 26292 6458
rect 26240 6394 26292 6400
rect 26056 6384 26108 6390
rect 26056 6326 26108 6332
rect 26148 6180 26200 6186
rect 26148 6122 26200 6128
rect 26160 4593 26188 6122
rect 26146 4584 26202 4593
rect 26146 4519 26202 4528
rect 25884 2746 26004 2774
rect 25504 2644 25556 2650
rect 25504 2586 25556 2592
rect 25412 2440 25464 2446
rect 25412 2382 25464 2388
rect 25320 1284 25372 1290
rect 25320 1226 25372 1232
rect 25424 800 25452 2382
rect 25976 1154 26004 2746
rect 25964 1148 26016 1154
rect 25964 1090 26016 1096
rect 26620 1057 26648 9862
rect 26804 9382 26832 12174
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26896 7002 26924 14826
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 26884 6860 26936 6866
rect 26884 6802 26936 6808
rect 26896 6458 26924 6802
rect 26884 6452 26936 6458
rect 26884 6394 26936 6400
rect 26988 4672 27016 17190
rect 27080 16454 27108 17206
rect 27172 16590 27200 18158
rect 27264 17218 27292 20266
rect 27436 19780 27488 19786
rect 27436 19722 27488 19728
rect 27344 19236 27396 19242
rect 27344 19178 27396 19184
rect 27356 17338 27384 19178
rect 27448 17610 27476 19722
rect 27632 19394 27660 21830
rect 27724 21729 27752 22222
rect 27896 22170 27948 22176
rect 27908 22094 27936 22170
rect 27816 22066 27936 22094
rect 27710 21720 27766 21729
rect 27710 21655 27766 21664
rect 27712 21480 27764 21486
rect 27712 21422 27764 21428
rect 27724 21146 27752 21422
rect 27712 21140 27764 21146
rect 27712 21082 27764 21088
rect 27816 21049 27844 22066
rect 28368 21865 28396 22936
rect 28448 22636 28500 22642
rect 28448 22578 28500 22584
rect 28460 22234 28488 22578
rect 28448 22228 28500 22234
rect 28448 22170 28500 22176
rect 28354 21856 28410 21865
rect 27950 21788 28258 21797
rect 28354 21791 28410 21800
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28354 21720 28410 21729
rect 28354 21655 28356 21664
rect 28408 21655 28410 21664
rect 28356 21626 28408 21632
rect 27896 21616 27948 21622
rect 27896 21558 27948 21564
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 27908 21486 27936 21558
rect 27896 21480 27948 21486
rect 27896 21422 27948 21428
rect 28000 21418 28028 21558
rect 28460 21554 28488 22170
rect 28080 21548 28132 21554
rect 28080 21490 28132 21496
rect 28448 21548 28500 21554
rect 28448 21490 28500 21496
rect 27988 21412 28040 21418
rect 27988 21354 28040 21360
rect 27802 21040 27858 21049
rect 27802 20975 27858 20984
rect 28000 20942 28028 21354
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27988 20936 28040 20942
rect 27988 20878 28040 20884
rect 27724 20058 27752 20878
rect 27804 20868 27856 20874
rect 27804 20810 27856 20816
rect 27816 20534 27844 20810
rect 28092 20806 28120 21490
rect 28460 21146 28488 21490
rect 28448 21140 28500 21146
rect 28448 21082 28500 21088
rect 28080 20800 28132 20806
rect 28080 20742 28132 20748
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27804 20528 27856 20534
rect 27804 20470 27856 20476
rect 27816 20398 27844 20470
rect 28460 20466 28488 21082
rect 28448 20460 28500 20466
rect 28448 20402 28500 20408
rect 27804 20392 27856 20398
rect 27804 20334 27856 20340
rect 28460 20058 28488 20402
rect 28538 20088 28594 20097
rect 27712 20052 27764 20058
rect 27712 19994 27764 20000
rect 28448 20052 28500 20058
rect 28538 20023 28594 20032
rect 28448 19994 28500 20000
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27540 19366 27660 19394
rect 27712 19440 27764 19446
rect 27712 19382 27764 19388
rect 27540 18970 27568 19366
rect 27620 19304 27672 19310
rect 27620 19246 27672 19252
rect 27632 18970 27660 19246
rect 27528 18964 27580 18970
rect 27528 18906 27580 18912
rect 27620 18964 27672 18970
rect 27620 18906 27672 18912
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27528 18284 27580 18290
rect 27528 18226 27580 18232
rect 27436 17604 27488 17610
rect 27436 17546 27488 17552
rect 27344 17332 27396 17338
rect 27344 17274 27396 17280
rect 27264 17190 27384 17218
rect 27540 17202 27568 18226
rect 27252 17128 27304 17134
rect 27252 17070 27304 17076
rect 27264 16590 27292 17070
rect 27160 16584 27212 16590
rect 27160 16526 27212 16532
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16114 27108 16390
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 27172 16114 27200 16186
rect 27068 16108 27120 16114
rect 27068 16050 27120 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 27080 14822 27108 16050
rect 27356 15638 27384 17190
rect 27528 17196 27580 17202
rect 27528 17138 27580 17144
rect 27632 16794 27660 18294
rect 27620 16788 27672 16794
rect 27620 16730 27672 16736
rect 27436 16652 27488 16658
rect 27436 16594 27488 16600
rect 27344 15632 27396 15638
rect 27344 15574 27396 15580
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27264 14890 27292 15370
rect 27342 15328 27398 15337
rect 27342 15263 27398 15272
rect 27252 14884 27304 14890
rect 27252 14826 27304 14832
rect 27068 14816 27120 14822
rect 27068 14758 27120 14764
rect 27080 12646 27108 14758
rect 27068 12640 27120 12646
rect 27068 12582 27120 12588
rect 27356 12434 27384 15263
rect 27264 12406 27384 12434
rect 27448 12434 27476 16594
rect 27618 16416 27674 16425
rect 27618 16351 27674 16360
rect 27528 16176 27580 16182
rect 27528 16118 27580 16124
rect 27540 15473 27568 16118
rect 27526 15464 27582 15473
rect 27526 15399 27582 15408
rect 27632 15348 27660 16351
rect 27724 16017 27752 19382
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28264 18828 28316 18834
rect 28264 18770 28316 18776
rect 28276 18630 28304 18770
rect 27804 18624 27856 18630
rect 27802 18592 27804 18601
rect 28264 18624 28316 18630
rect 27856 18592 27858 18601
rect 28264 18566 28316 18572
rect 27802 18527 27858 18536
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27802 18456 27858 18465
rect 27950 18459 28258 18468
rect 27858 18400 27936 18408
rect 27802 18391 27936 18400
rect 27816 18380 27936 18391
rect 27804 18080 27856 18086
rect 27802 18048 27804 18057
rect 27856 18048 27858 18057
rect 27802 17983 27858 17992
rect 27908 17921 27936 18380
rect 28368 18358 28396 19246
rect 28356 18352 28408 18358
rect 28356 18294 28408 18300
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27894 17912 27950 17921
rect 27894 17847 27950 17856
rect 28000 17746 28028 18226
rect 28262 18184 28318 18193
rect 28262 18119 28318 18128
rect 27988 17740 28040 17746
rect 27988 17682 28040 17688
rect 28276 17542 28304 18119
rect 28552 17864 28580 20023
rect 28644 19553 28672 26200
rect 28724 25084 28776 25090
rect 28724 25026 28776 25032
rect 28736 22710 28764 25026
rect 28816 24948 28868 24954
rect 28816 24890 28868 24896
rect 28828 23798 28856 24890
rect 29184 24880 29236 24886
rect 29184 24822 29236 24828
rect 28998 24712 29054 24721
rect 28998 24647 29054 24656
rect 28816 23792 28868 23798
rect 28816 23734 28868 23740
rect 28908 23792 28960 23798
rect 28908 23734 28960 23740
rect 28816 23656 28868 23662
rect 28816 23598 28868 23604
rect 28724 22704 28776 22710
rect 28724 22646 28776 22652
rect 28828 22556 28856 23598
rect 28920 23186 28948 23734
rect 29012 23730 29040 24647
rect 29092 24336 29144 24342
rect 29092 24278 29144 24284
rect 29000 23724 29052 23730
rect 29000 23666 29052 23672
rect 29000 23520 29052 23526
rect 29000 23462 29052 23468
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 29012 23050 29040 23462
rect 29104 23254 29132 24278
rect 29196 24274 29224 24822
rect 29288 24274 29316 26200
rect 29552 25696 29604 25702
rect 29552 25638 29604 25644
rect 29460 24608 29512 24614
rect 29460 24550 29512 24556
rect 29184 24268 29236 24274
rect 29184 24210 29236 24216
rect 29276 24268 29328 24274
rect 29276 24210 29328 24216
rect 29276 24064 29328 24070
rect 29276 24006 29328 24012
rect 29368 24064 29420 24070
rect 29368 24006 29420 24012
rect 29288 23526 29316 24006
rect 29380 23866 29408 24006
rect 29368 23860 29420 23866
rect 29368 23802 29420 23808
rect 29472 23594 29500 24550
rect 29460 23588 29512 23594
rect 29460 23530 29512 23536
rect 29276 23520 29328 23526
rect 29276 23462 29328 23468
rect 29092 23248 29144 23254
rect 29092 23190 29144 23196
rect 29288 23118 29316 23462
rect 29276 23112 29328 23118
rect 29276 23054 29328 23060
rect 29000 23044 29052 23050
rect 29000 22986 29052 22992
rect 28736 22528 28856 22556
rect 28736 21622 28764 22528
rect 28908 22432 28960 22438
rect 28908 22374 28960 22380
rect 28920 22273 28948 22374
rect 28906 22264 28962 22273
rect 29288 22234 29316 23054
rect 29472 22778 29500 23530
rect 29368 22772 29420 22778
rect 29368 22714 29420 22720
rect 29460 22772 29512 22778
rect 29460 22714 29512 22720
rect 28906 22199 28962 22208
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 28906 22128 28962 22137
rect 28906 22063 28962 22072
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28920 21978 28948 22063
rect 28724 21616 28776 21622
rect 28724 21558 28776 21564
rect 28828 21078 28856 21966
rect 28920 21950 29040 21978
rect 28908 21888 28960 21894
rect 28908 21830 28960 21836
rect 28920 21729 28948 21830
rect 28906 21720 28962 21729
rect 28906 21655 28962 21664
rect 29012 21570 29040 21950
rect 28920 21542 29040 21570
rect 29182 21584 29238 21593
rect 28724 21072 28776 21078
rect 28724 21014 28776 21020
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28630 19544 28686 19553
rect 28630 19479 28686 19488
rect 28552 17836 28672 17864
rect 28448 17808 28500 17814
rect 28448 17750 28500 17756
rect 28460 17678 28488 17750
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28264 17536 28316 17542
rect 27802 17504 27858 17513
rect 28264 17478 28316 17484
rect 27802 17439 27858 17448
rect 27816 16640 27844 17439
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 28460 17270 28488 17614
rect 28538 17504 28594 17513
rect 28538 17439 28594 17448
rect 28448 17264 28500 17270
rect 28448 17206 28500 17212
rect 27988 16652 28040 16658
rect 27816 16612 27988 16640
rect 27988 16594 28040 16600
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27802 16280 27858 16289
rect 27950 16283 28258 16292
rect 27858 16224 28028 16232
rect 27802 16215 28028 16224
rect 27816 16204 28028 16215
rect 28000 16153 28028 16204
rect 27802 16144 27858 16153
rect 27802 16079 27858 16088
rect 27986 16144 28042 16153
rect 27986 16079 28042 16088
rect 28264 16108 28316 16114
rect 27710 16008 27766 16017
rect 27710 15943 27766 15952
rect 27816 15706 27844 16079
rect 28264 16050 28316 16056
rect 27986 15736 28042 15745
rect 27804 15700 27856 15706
rect 27986 15671 27988 15680
rect 27804 15642 27856 15648
rect 28040 15671 28042 15680
rect 27988 15642 28040 15648
rect 28000 15502 28028 15642
rect 28276 15638 28304 16050
rect 28264 15632 28316 15638
rect 28264 15574 28316 15580
rect 27712 15496 27764 15502
rect 27710 15464 27712 15473
rect 27988 15496 28040 15502
rect 27764 15464 27766 15473
rect 27988 15438 28040 15444
rect 27710 15399 27766 15408
rect 27632 15320 27752 15348
rect 27724 15094 27752 15320
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27712 15088 27764 15094
rect 27712 15030 27764 15036
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 12442 27660 14962
rect 28368 14929 28396 16526
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28460 14958 28488 16390
rect 28552 15042 28580 17439
rect 28644 16402 28672 17836
rect 28736 16522 28764 21014
rect 28816 20800 28868 20806
rect 28816 20742 28868 20748
rect 28828 19334 28856 20742
rect 28920 19938 28948 21542
rect 29182 21519 29238 21528
rect 28920 19910 29132 19938
rect 28998 19816 29054 19825
rect 28998 19751 29054 19760
rect 28906 19544 28962 19553
rect 28906 19479 28962 19488
rect 28920 19446 28948 19479
rect 28908 19440 28960 19446
rect 28908 19382 28960 19388
rect 28828 19306 28948 19334
rect 28816 19168 28868 19174
rect 28816 19110 28868 19116
rect 28828 18766 28856 19110
rect 28816 18760 28868 18766
rect 28816 18702 28868 18708
rect 28828 16572 28856 18702
rect 28920 17490 28948 19306
rect 29012 18193 29040 19751
rect 29104 19145 29132 19910
rect 29090 19136 29146 19145
rect 29090 19071 29146 19080
rect 29092 18828 29144 18834
rect 29092 18770 29144 18776
rect 29104 18465 29132 18770
rect 29196 18601 29224 21519
rect 29276 21140 29328 21146
rect 29276 21082 29328 21088
rect 29288 20806 29316 21082
rect 29276 20800 29328 20806
rect 29276 20742 29328 20748
rect 29380 20262 29408 22714
rect 29564 22250 29592 25638
rect 29736 24268 29788 24274
rect 29736 24210 29788 24216
rect 29644 23656 29696 23662
rect 29644 23598 29696 23604
rect 29656 23322 29684 23598
rect 29748 23594 29776 24210
rect 29736 23588 29788 23594
rect 29736 23530 29788 23536
rect 29644 23316 29696 23322
rect 29644 23258 29696 23264
rect 29644 23044 29696 23050
rect 29644 22986 29696 22992
rect 29472 22222 29592 22250
rect 29656 22234 29684 22986
rect 29736 22976 29788 22982
rect 29736 22918 29788 22924
rect 29748 22506 29776 22918
rect 29736 22500 29788 22506
rect 29736 22442 29788 22448
rect 29644 22228 29696 22234
rect 29472 20777 29500 22222
rect 29644 22170 29696 22176
rect 29840 22094 29868 26726
rect 29918 26330 29974 27000
rect 30562 26330 30618 27000
rect 31206 26330 31262 27000
rect 31850 26330 31906 27000
rect 32494 26330 32550 27000
rect 33138 26330 33194 27000
rect 33692 26852 33744 26858
rect 33692 26794 33744 26800
rect 29918 26302 30236 26330
rect 29918 26200 29974 26302
rect 29920 24676 29972 24682
rect 29920 24618 29972 24624
rect 29932 24342 29960 24618
rect 29920 24336 29972 24342
rect 29920 24278 29972 24284
rect 30208 23322 30236 26302
rect 30562 26302 30880 26330
rect 30562 26200 30618 26302
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30196 23316 30248 23322
rect 30196 23258 30248 23264
rect 30104 23044 30156 23050
rect 30104 22986 30156 22992
rect 30012 22772 30064 22778
rect 30012 22714 30064 22720
rect 29920 22432 29972 22438
rect 29920 22374 29972 22380
rect 29564 22066 29868 22094
rect 29458 20768 29514 20777
rect 29458 20703 29514 20712
rect 29276 20256 29328 20262
rect 29276 20198 29328 20204
rect 29368 20256 29420 20262
rect 29368 20198 29420 20204
rect 29288 19310 29316 20198
rect 29564 20058 29592 22066
rect 29828 22024 29880 22030
rect 29828 21966 29880 21972
rect 29736 21548 29788 21554
rect 29736 21490 29788 21496
rect 29748 20534 29776 21490
rect 29736 20528 29788 20534
rect 29736 20470 29788 20476
rect 29552 20052 29604 20058
rect 29552 19994 29604 20000
rect 29368 19712 29420 19718
rect 29368 19654 29420 19660
rect 29380 19334 29408 19654
rect 29644 19508 29696 19514
rect 29644 19450 29696 19456
rect 29276 19304 29328 19310
rect 29380 19306 29592 19334
rect 29276 19246 29328 19252
rect 29460 18828 29512 18834
rect 29460 18770 29512 18776
rect 29368 18624 29420 18630
rect 29182 18592 29238 18601
rect 29472 18601 29500 18770
rect 29368 18566 29420 18572
rect 29458 18592 29514 18601
rect 29182 18527 29238 18536
rect 29090 18456 29146 18465
rect 29380 18426 29408 18566
rect 29458 18527 29514 18536
rect 29090 18391 29146 18400
rect 29368 18420 29420 18426
rect 29368 18362 29420 18368
rect 29460 18284 29512 18290
rect 29460 18226 29512 18232
rect 28998 18184 29054 18193
rect 28998 18119 29054 18128
rect 29472 17746 29500 18226
rect 29564 17785 29592 19306
rect 29550 17776 29606 17785
rect 29460 17740 29512 17746
rect 29550 17711 29606 17720
rect 29460 17682 29512 17688
rect 29276 17604 29328 17610
rect 29276 17546 29328 17552
rect 29288 17513 29316 17546
rect 29274 17504 29330 17513
rect 28920 17462 29132 17490
rect 28906 17368 28962 17377
rect 28906 17303 28962 17312
rect 28920 17134 28948 17303
rect 28908 17128 28960 17134
rect 28908 17070 28960 17076
rect 28908 16788 28960 16794
rect 28908 16730 28960 16736
rect 28920 16674 28948 16730
rect 28920 16646 29040 16674
rect 28908 16584 28960 16590
rect 28828 16544 28908 16572
rect 28908 16526 28960 16532
rect 28724 16516 28776 16522
rect 28724 16458 28776 16464
rect 28816 16448 28868 16454
rect 28644 16374 28764 16402
rect 29012 16436 29040 16646
rect 29104 16538 29132 17462
rect 29274 17439 29330 17448
rect 29472 17270 29500 17682
rect 29656 17542 29684 19450
rect 29748 19378 29776 20470
rect 29840 19922 29868 21966
rect 29932 21486 29960 22374
rect 30024 22234 30052 22714
rect 30116 22710 30144 22986
rect 30196 22976 30248 22982
rect 30196 22918 30248 22924
rect 30104 22704 30156 22710
rect 30104 22646 30156 22652
rect 30012 22228 30064 22234
rect 30012 22170 30064 22176
rect 30010 22128 30066 22137
rect 30010 22063 30066 22072
rect 30024 21894 30052 22063
rect 30012 21888 30064 21894
rect 30012 21830 30064 21836
rect 29920 21480 29972 21486
rect 29920 21422 29972 21428
rect 30116 21418 30144 22646
rect 30208 22438 30236 22918
rect 30196 22432 30248 22438
rect 30196 22374 30248 22380
rect 30288 22432 30340 22438
rect 30288 22374 30340 22380
rect 30300 22166 30328 22374
rect 30288 22160 30340 22166
rect 30392 22137 30420 25230
rect 30656 24880 30708 24886
rect 30656 24822 30708 24828
rect 30562 22264 30618 22273
rect 30562 22199 30564 22208
rect 30616 22199 30618 22208
rect 30564 22170 30616 22176
rect 30288 22102 30340 22108
rect 30378 22128 30434 22137
rect 30668 22094 30696 24822
rect 30748 23724 30800 23730
rect 30748 23666 30800 23672
rect 30378 22063 30434 22072
rect 30576 22066 30696 22094
rect 30288 21888 30340 21894
rect 30288 21830 30340 21836
rect 30104 21412 30156 21418
rect 30104 21354 30156 21360
rect 30010 21176 30066 21185
rect 30010 21111 30066 21120
rect 29918 20904 29974 20913
rect 29918 20839 29974 20848
rect 29828 19916 29880 19922
rect 29828 19858 29880 19864
rect 29840 19718 29868 19858
rect 29828 19712 29880 19718
rect 29828 19654 29880 19660
rect 29736 19372 29788 19378
rect 29736 19314 29788 19320
rect 29748 18426 29776 19314
rect 29828 18964 29880 18970
rect 29828 18906 29880 18912
rect 29736 18420 29788 18426
rect 29736 18362 29788 18368
rect 29840 18034 29868 18906
rect 29748 18006 29868 18034
rect 29644 17536 29696 17542
rect 29644 17478 29696 17484
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29184 17128 29236 17134
rect 29184 17070 29236 17076
rect 29196 16658 29224 17070
rect 29472 16794 29500 17206
rect 29642 16824 29698 16833
rect 29460 16788 29512 16794
rect 29642 16759 29644 16768
rect 29460 16730 29512 16736
rect 29696 16759 29698 16768
rect 29644 16730 29696 16736
rect 29656 16658 29684 16730
rect 29184 16652 29236 16658
rect 29184 16594 29236 16600
rect 29644 16652 29696 16658
rect 29644 16594 29696 16600
rect 29748 16590 29776 18006
rect 29826 17912 29882 17921
rect 29826 17847 29882 17856
rect 29840 16708 29868 17847
rect 29932 16833 29960 20839
rect 29918 16824 29974 16833
rect 29918 16759 29974 16768
rect 29840 16680 29960 16708
rect 29736 16584 29788 16590
rect 29104 16510 29316 16538
rect 29736 16526 29788 16532
rect 28816 16390 28868 16396
rect 28920 16408 29040 16436
rect 29092 16448 29144 16454
rect 28632 15496 28684 15502
rect 28632 15438 28684 15444
rect 28644 15162 28672 15438
rect 28736 15366 28764 16374
rect 28724 15360 28776 15366
rect 28724 15302 28776 15308
rect 28632 15156 28684 15162
rect 28632 15098 28684 15104
rect 28722 15056 28778 15065
rect 28552 15014 28672 15042
rect 28448 14952 28500 14958
rect 28354 14920 28410 14929
rect 28448 14894 28500 14900
rect 28354 14855 28410 14864
rect 28448 14544 28500 14550
rect 28448 14486 28500 14492
rect 27712 14272 27764 14278
rect 27712 14214 27764 14220
rect 27724 13274 27752 14214
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27804 13728 27856 13734
rect 27804 13670 27856 13676
rect 27894 13696 27950 13705
rect 27816 13394 27844 13670
rect 27894 13631 27950 13640
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27724 13246 27844 13274
rect 27712 13184 27764 13190
rect 27712 13126 27764 13132
rect 27620 12436 27672 12442
rect 27448 12406 27568 12434
rect 27160 11756 27212 11762
rect 27160 11698 27212 11704
rect 27172 11354 27200 11698
rect 27160 11348 27212 11354
rect 27160 11290 27212 11296
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 27080 5574 27108 11086
rect 27172 10577 27200 11086
rect 27158 10568 27214 10577
rect 27158 10503 27214 10512
rect 27068 5568 27120 5574
rect 27068 5510 27120 5516
rect 27068 5024 27120 5030
rect 27120 4972 27200 4978
rect 27068 4966 27200 4972
rect 27080 4950 27200 4966
rect 27172 4690 27200 4950
rect 27068 4684 27120 4690
rect 26988 4644 27068 4672
rect 27068 4626 27120 4632
rect 27160 4684 27212 4690
rect 27160 4626 27212 4632
rect 27080 3466 27108 4626
rect 27068 3460 27120 3466
rect 27068 3402 27120 3408
rect 26606 1048 26662 1057
rect 26606 983 26662 992
rect 27264 921 27292 12406
rect 27344 12300 27396 12306
rect 27344 12242 27396 12248
rect 27356 11529 27384 12242
rect 27342 11520 27398 11529
rect 27342 11455 27398 11464
rect 27436 11280 27488 11286
rect 27434 11248 27436 11257
rect 27488 11248 27490 11257
rect 27434 11183 27490 11192
rect 27434 10840 27490 10849
rect 27434 10775 27490 10784
rect 27448 10674 27476 10775
rect 27436 10668 27488 10674
rect 27436 10610 27488 10616
rect 27540 5302 27568 12406
rect 27620 12378 27672 12384
rect 27724 12374 27752 13126
rect 27712 12368 27764 12374
rect 27712 12310 27764 12316
rect 27620 12096 27672 12102
rect 27816 12050 27844 13246
rect 27908 13190 27936 13631
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 28356 12640 28408 12646
rect 28356 12582 28408 12588
rect 27620 12038 27672 12044
rect 27632 9654 27660 12038
rect 27724 12022 27844 12050
rect 27724 11558 27752 12022
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27802 11928 27858 11937
rect 27950 11931 28258 11940
rect 27802 11863 27804 11872
rect 27856 11863 27858 11872
rect 27804 11834 27856 11840
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27804 11552 27856 11558
rect 27804 11494 27856 11500
rect 27816 11082 27844 11494
rect 27804 11076 27856 11082
rect 27804 11018 27856 11024
rect 27712 11008 27764 11014
rect 27712 10950 27764 10956
rect 27724 10470 27752 10950
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27724 9897 27752 10406
rect 27710 9888 27766 9897
rect 27710 9823 27766 9832
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27620 9648 27672 9654
rect 27620 9590 27672 9596
rect 27712 9648 27764 9654
rect 27712 9590 27764 9596
rect 27724 9110 27752 9590
rect 27712 9104 27764 9110
rect 28368 9081 28396 12582
rect 28460 12442 28488 14486
rect 28540 13932 28592 13938
rect 28540 13874 28592 13880
rect 28448 12436 28500 12442
rect 28448 12378 28500 12384
rect 28552 10538 28580 13874
rect 28644 13394 28672 15014
rect 28722 14991 28724 15000
rect 28776 14991 28778 15000
rect 28724 14962 28776 14968
rect 28722 14920 28778 14929
rect 28722 14855 28778 14864
rect 28736 14657 28764 14855
rect 28722 14648 28778 14657
rect 28722 14583 28778 14592
rect 28632 13388 28684 13394
rect 28632 13330 28684 13336
rect 28736 11286 28764 14583
rect 28828 14550 28856 16390
rect 28816 14544 28868 14550
rect 28816 14486 28868 14492
rect 28816 14272 28868 14278
rect 28816 14214 28868 14220
rect 28828 12434 28856 14214
rect 28920 13802 28948 16408
rect 29092 16390 29144 16396
rect 29000 15904 29052 15910
rect 29000 15846 29052 15852
rect 29012 14618 29040 15846
rect 29000 14612 29052 14618
rect 29000 14554 29052 14560
rect 28908 13796 28960 13802
rect 28908 13738 28960 13744
rect 28906 13288 28962 13297
rect 28906 13223 28908 13232
rect 28960 13223 28962 13232
rect 28908 13194 28960 13200
rect 28908 12776 28960 12782
rect 28906 12744 28908 12753
rect 28960 12744 28962 12753
rect 28906 12679 28962 12688
rect 28828 12406 28948 12434
rect 28724 11280 28776 11286
rect 28724 11222 28776 11228
rect 28632 11076 28684 11082
rect 28632 11018 28684 11024
rect 28724 11076 28776 11082
rect 28724 11018 28776 11024
rect 28540 10532 28592 10538
rect 28540 10474 28592 10480
rect 28448 9920 28500 9926
rect 28448 9862 28500 9868
rect 27712 9046 27764 9052
rect 28354 9072 28410 9081
rect 28354 9007 28410 9016
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27632 7857 27660 8910
rect 27712 8832 27764 8838
rect 27712 8774 27764 8780
rect 28356 8832 28408 8838
rect 28356 8774 28408 8780
rect 27618 7848 27674 7857
rect 27618 7783 27674 7792
rect 27620 6248 27672 6254
rect 27620 6190 27672 6196
rect 27528 5296 27580 5302
rect 27528 5238 27580 5244
rect 27344 5160 27396 5166
rect 27344 5102 27396 5108
rect 27356 4826 27384 5102
rect 27344 4820 27396 4826
rect 27344 4762 27396 4768
rect 27632 3505 27660 6190
rect 27724 5778 27752 8774
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 28368 8634 28396 8774
rect 28356 8628 28408 8634
rect 28356 8570 28408 8576
rect 27804 8424 27856 8430
rect 27804 8366 27856 8372
rect 27816 7750 27844 8366
rect 27804 7744 27856 7750
rect 27804 7686 27856 7692
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27712 5772 27764 5778
rect 27712 5714 27764 5720
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27804 4480 27856 4486
rect 27804 4422 27856 4428
rect 27618 3496 27674 3505
rect 27618 3431 27674 3440
rect 27816 2650 27844 4422
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28356 2440 28408 2446
rect 28356 2382 28408 2388
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 27250 912 27306 921
rect 27250 847 27306 856
rect 28092 870 28212 898
rect 28092 800 28120 870
rect 21272 604 21324 610
rect 21272 546 21324 552
rect 20812 196 20864 202
rect 20812 138 20864 144
rect 22742 0 22798 800
rect 25410 0 25466 800
rect 28078 0 28134 800
rect 28184 762 28212 870
rect 28368 762 28396 2382
rect 28460 1873 28488 9862
rect 28644 2774 28672 11018
rect 28736 3670 28764 11018
rect 28816 10668 28868 10674
rect 28816 10610 28868 10616
rect 28828 9722 28856 10610
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28920 5166 28948 12406
rect 29000 9036 29052 9042
rect 29000 8978 29052 8984
rect 29012 7478 29040 8978
rect 29000 7472 29052 7478
rect 29000 7414 29052 7420
rect 28908 5160 28960 5166
rect 28908 5102 28960 5108
rect 28724 3664 28776 3670
rect 28724 3606 28776 3612
rect 28920 3534 28948 5102
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28644 2746 28764 2774
rect 28736 2378 28764 2746
rect 28724 2372 28776 2378
rect 28724 2314 28776 2320
rect 28446 1864 28502 1873
rect 28446 1799 28502 1808
rect 28184 734 28396 762
rect 29104 649 29132 16390
rect 29182 16144 29238 16153
rect 29182 16079 29238 16088
rect 29196 15162 29224 16079
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 29288 14278 29316 16510
rect 29552 15904 29604 15910
rect 29552 15846 29604 15852
rect 29460 15020 29512 15026
rect 29460 14962 29512 14968
rect 29368 14816 29420 14822
rect 29368 14758 29420 14764
rect 29380 14414 29408 14758
rect 29368 14408 29420 14414
rect 29368 14350 29420 14356
rect 29276 14272 29328 14278
rect 29276 14214 29328 14220
rect 29368 14272 29420 14278
rect 29472 14226 29500 14962
rect 29420 14220 29500 14226
rect 29368 14214 29500 14220
rect 29380 14198 29500 14214
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 29288 12442 29316 14010
rect 29276 12436 29328 12442
rect 29276 12378 29328 12384
rect 29380 11098 29408 14198
rect 29196 11070 29408 11098
rect 29196 8945 29224 11070
rect 29564 10826 29592 15846
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29656 12306 29684 15438
rect 29736 14612 29788 14618
rect 29736 14554 29788 14560
rect 29748 14414 29776 14554
rect 29736 14408 29788 14414
rect 29736 14350 29788 14356
rect 29748 13462 29776 14350
rect 29828 13932 29880 13938
rect 29828 13874 29880 13880
rect 29736 13456 29788 13462
rect 29736 13398 29788 13404
rect 29840 12617 29868 13874
rect 29932 13734 29960 16680
rect 30024 15994 30052 21111
rect 30116 20874 30144 21354
rect 30104 20868 30156 20874
rect 30104 20810 30156 20816
rect 30300 20040 30328 21830
rect 30300 20012 30420 20040
rect 30288 19916 30340 19922
rect 30288 19858 30340 19864
rect 30104 19848 30156 19854
rect 30104 19790 30156 19796
rect 30116 18358 30144 19790
rect 30196 19712 30248 19718
rect 30194 19680 30196 19689
rect 30248 19680 30250 19689
rect 30194 19615 30250 19624
rect 30196 18624 30248 18630
rect 30194 18592 30196 18601
rect 30248 18592 30250 18601
rect 30194 18527 30250 18536
rect 30104 18352 30156 18358
rect 30104 18294 30156 18300
rect 30196 17808 30248 17814
rect 30300 17796 30328 19858
rect 30392 19825 30420 20012
rect 30378 19816 30434 19825
rect 30576 19786 30604 22066
rect 30760 22012 30788 23666
rect 30668 21984 30788 22012
rect 30668 21554 30696 21984
rect 30748 21888 30800 21894
rect 30748 21830 30800 21836
rect 30760 21554 30788 21830
rect 30656 21548 30708 21554
rect 30656 21490 30708 21496
rect 30748 21548 30800 21554
rect 30748 21490 30800 21496
rect 30668 20874 30696 21490
rect 30760 21146 30788 21490
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30656 20868 30708 20874
rect 30656 20810 30708 20816
rect 30746 20768 30802 20777
rect 30746 20703 30802 20712
rect 30656 20324 30708 20330
rect 30656 20266 30708 20272
rect 30378 19751 30434 19760
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30564 19780 30616 19786
rect 30564 19722 30616 19728
rect 30484 19378 30512 19722
rect 30472 19372 30524 19378
rect 30472 19314 30524 19320
rect 30380 18624 30432 18630
rect 30380 18566 30432 18572
rect 30564 18624 30616 18630
rect 30564 18566 30616 18572
rect 30392 17882 30420 18566
rect 30470 18320 30526 18329
rect 30576 18290 30604 18566
rect 30470 18255 30526 18264
rect 30564 18284 30616 18290
rect 30380 17876 30432 17882
rect 30380 17818 30432 17824
rect 30248 17768 30328 17796
rect 30196 17750 30248 17756
rect 30102 17640 30158 17649
rect 30102 17575 30158 17584
rect 30116 17542 30144 17575
rect 30104 17536 30156 17542
rect 30104 17478 30156 17484
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17105 30236 17478
rect 30300 17202 30328 17768
rect 30484 17490 30512 18255
rect 30564 18226 30616 18232
rect 30564 18148 30616 18154
rect 30564 18090 30616 18096
rect 30576 17542 30604 18090
rect 30392 17462 30512 17490
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30288 17196 30340 17202
rect 30288 17138 30340 17144
rect 30194 17096 30250 17105
rect 30194 17031 30250 17040
rect 30392 16572 30420 17462
rect 30668 17320 30696 20266
rect 30484 17292 30696 17320
rect 30484 16726 30512 17292
rect 30654 17232 30710 17241
rect 30654 17167 30710 17176
rect 30564 16992 30616 16998
rect 30564 16934 30616 16940
rect 30472 16720 30524 16726
rect 30472 16662 30524 16668
rect 30392 16544 30512 16572
rect 30104 16448 30156 16454
rect 30104 16390 30156 16396
rect 30116 16114 30144 16390
rect 30104 16108 30156 16114
rect 30104 16050 30156 16056
rect 30024 15966 30144 15994
rect 30116 15502 30144 15966
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30104 15496 30156 15502
rect 30104 15438 30156 15444
rect 29920 13728 29972 13734
rect 29920 13670 29972 13676
rect 29826 12608 29882 12617
rect 29826 12543 29882 12552
rect 29736 12436 29788 12442
rect 29736 12378 29788 12384
rect 29644 12300 29696 12306
rect 29644 12242 29696 12248
rect 29644 11280 29696 11286
rect 29644 11222 29696 11228
rect 29380 10810 29592 10826
rect 29368 10804 29592 10810
rect 29420 10798 29592 10804
rect 29368 10746 29420 10752
rect 29182 8936 29238 8945
rect 29182 8871 29238 8880
rect 29656 7449 29684 11222
rect 29748 8498 29776 12378
rect 30024 12345 30052 15438
rect 30380 14816 30432 14822
rect 30380 14758 30432 14764
rect 30288 14476 30340 14482
rect 30288 14418 30340 14424
rect 30300 14278 30328 14418
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30392 12434 30420 14758
rect 30484 13938 30512 16544
rect 30576 16114 30604 16934
rect 30668 16658 30696 17167
rect 30656 16652 30708 16658
rect 30656 16594 30708 16600
rect 30564 16108 30616 16114
rect 30564 16050 30616 16056
rect 30472 13932 30524 13938
rect 30472 13874 30524 13880
rect 30392 12406 30512 12434
rect 30010 12336 30066 12345
rect 30010 12271 30066 12280
rect 30380 11892 30432 11898
rect 30380 11834 30432 11840
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30024 10810 30052 11018
rect 30012 10804 30064 10810
rect 30012 10746 30064 10752
rect 30392 10130 30420 11834
rect 30380 10124 30432 10130
rect 30380 10066 30432 10072
rect 29736 8492 29788 8498
rect 29736 8434 29788 8440
rect 29642 7440 29698 7449
rect 29642 7375 29698 7384
rect 30484 6662 30512 12406
rect 30576 11801 30604 16050
rect 30654 15600 30710 15609
rect 30654 15535 30710 15544
rect 30562 11792 30618 11801
rect 30562 11727 30618 11736
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30668 5846 30696 15535
rect 30760 14482 30788 20703
rect 30852 19122 30880 26302
rect 31206 26302 31340 26330
rect 31206 26200 31262 26302
rect 31116 24948 31168 24954
rect 31116 24890 31168 24896
rect 31024 24200 31076 24206
rect 31024 24142 31076 24148
rect 31036 23866 31064 24142
rect 31024 23860 31076 23866
rect 31024 23802 31076 23808
rect 31128 23662 31156 24890
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31312 22710 31340 26302
rect 31850 26302 32168 26330
rect 31850 26200 31906 26302
rect 31944 25628 31996 25634
rect 31944 25570 31996 25576
rect 31392 23792 31444 23798
rect 31444 23752 31708 23780
rect 31392 23734 31444 23740
rect 31680 23662 31708 23752
rect 31668 23656 31720 23662
rect 31668 23598 31720 23604
rect 31760 23520 31812 23526
rect 31760 23462 31812 23468
rect 31850 23488 31906 23497
rect 31772 23254 31800 23462
rect 31956 23474 31984 25570
rect 32036 24064 32088 24070
rect 32036 24006 32088 24012
rect 32048 23798 32076 24006
rect 32036 23792 32088 23798
rect 32036 23734 32088 23740
rect 31956 23446 32076 23474
rect 31850 23423 31906 23432
rect 31760 23248 31812 23254
rect 31760 23190 31812 23196
rect 31392 23112 31444 23118
rect 31392 23054 31444 23060
rect 31404 22778 31432 23054
rect 31576 22976 31628 22982
rect 31576 22918 31628 22924
rect 31482 22808 31538 22817
rect 31392 22772 31444 22778
rect 31482 22743 31538 22752
rect 31392 22714 31444 22720
rect 31208 22704 31260 22710
rect 31022 22672 31078 22681
rect 31208 22646 31260 22652
rect 31300 22704 31352 22710
rect 31300 22646 31352 22652
rect 31022 22607 31078 22616
rect 30932 22024 30984 22030
rect 30932 21966 30984 21972
rect 30944 21690 30972 21966
rect 30932 21684 30984 21690
rect 30932 21626 30984 21632
rect 31036 20466 31064 22607
rect 31114 21584 31170 21593
rect 31114 21519 31116 21528
rect 31168 21519 31170 21528
rect 31116 21490 31168 21496
rect 31116 20800 31168 20806
rect 31114 20768 31116 20777
rect 31168 20768 31170 20777
rect 31114 20703 31170 20712
rect 31024 20460 31076 20466
rect 31024 20402 31076 20408
rect 31036 19922 31064 20402
rect 31116 20392 31168 20398
rect 31116 20334 31168 20340
rect 31024 19916 31076 19922
rect 31024 19858 31076 19864
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19242 30972 19654
rect 30932 19236 30984 19242
rect 30932 19178 30984 19184
rect 30852 19094 30972 19122
rect 30840 18760 30892 18766
rect 30840 18702 30892 18708
rect 30852 18086 30880 18702
rect 30840 18080 30892 18086
rect 30840 18022 30892 18028
rect 30840 17672 30892 17678
rect 30840 17614 30892 17620
rect 30852 17270 30880 17614
rect 30840 17264 30892 17270
rect 30840 17206 30892 17212
rect 30944 16114 30972 19094
rect 31022 18320 31078 18329
rect 31022 18255 31078 18264
rect 31036 17746 31064 18255
rect 31024 17740 31076 17746
rect 31024 17682 31076 17688
rect 31128 17202 31156 20334
rect 31220 18834 31248 22646
rect 31496 22642 31524 22743
rect 31484 22636 31536 22642
rect 31484 22578 31536 22584
rect 31496 21146 31524 22578
rect 31588 22574 31616 22918
rect 31772 22778 31800 23190
rect 31760 22772 31812 22778
rect 31760 22714 31812 22720
rect 31576 22568 31628 22574
rect 31576 22510 31628 22516
rect 31760 22432 31812 22438
rect 31758 22400 31760 22409
rect 31812 22400 31814 22409
rect 31758 22335 31814 22344
rect 31864 22094 31892 23423
rect 31942 23352 31998 23361
rect 31942 23287 31998 23296
rect 31956 22982 31984 23287
rect 31944 22976 31996 22982
rect 31944 22918 31996 22924
rect 31864 22066 31984 22094
rect 31760 21616 31812 21622
rect 31760 21558 31812 21564
rect 31574 21312 31630 21321
rect 31574 21247 31630 21256
rect 31484 21140 31536 21146
rect 31484 21082 31536 21088
rect 31390 20632 31446 20641
rect 31390 20567 31446 20576
rect 31300 20392 31352 20398
rect 31300 20334 31352 20340
rect 31312 19446 31340 20334
rect 31404 20262 31432 20567
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31392 20052 31444 20058
rect 31392 19994 31444 20000
rect 31300 19440 31352 19446
rect 31300 19382 31352 19388
rect 31300 19236 31352 19242
rect 31300 19178 31352 19184
rect 31208 18828 31260 18834
rect 31208 18770 31260 18776
rect 31208 17536 31260 17542
rect 31208 17478 31260 17484
rect 31116 17196 31168 17202
rect 31116 17138 31168 17144
rect 31220 16250 31248 17478
rect 31312 17134 31340 19178
rect 31404 17660 31432 19994
rect 31496 19242 31524 21082
rect 31484 19236 31536 19242
rect 31484 19178 31536 19184
rect 31496 19009 31524 19178
rect 31482 19000 31538 19009
rect 31482 18935 31538 18944
rect 31588 17814 31616 21247
rect 31668 20936 31720 20942
rect 31666 20904 31668 20913
rect 31720 20904 31722 20913
rect 31666 20839 31722 20848
rect 31772 20806 31800 21558
rect 31956 21418 31984 22066
rect 31944 21412 31996 21418
rect 31944 21354 31996 21360
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31864 21146 31892 21286
rect 31852 21140 31904 21146
rect 31852 21082 31904 21088
rect 31760 20800 31812 20806
rect 31760 20742 31812 20748
rect 31772 20534 31800 20742
rect 31760 20528 31812 20534
rect 31760 20470 31812 20476
rect 31772 19378 31800 20470
rect 31864 20346 31892 21082
rect 31944 20936 31996 20942
rect 31944 20878 31996 20884
rect 31956 20777 31984 20878
rect 31942 20768 31998 20777
rect 31942 20703 31998 20712
rect 31864 20318 31984 20346
rect 31956 20262 31984 20318
rect 31944 20256 31996 20262
rect 31944 20198 31996 20204
rect 31956 20058 31984 20198
rect 31944 20052 31996 20058
rect 31944 19994 31996 20000
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31944 19304 31996 19310
rect 31944 19246 31996 19252
rect 31760 19168 31812 19174
rect 31758 19136 31760 19145
rect 31812 19136 31814 19145
rect 31758 19071 31814 19080
rect 31760 18692 31812 18698
rect 31956 18680 31984 19246
rect 31812 18652 31984 18680
rect 31760 18634 31812 18640
rect 31668 18080 31720 18086
rect 31666 18048 31668 18057
rect 31720 18048 31722 18057
rect 31666 17983 31722 17992
rect 31576 17808 31628 17814
rect 31576 17750 31628 17756
rect 31404 17632 31524 17660
rect 31300 17128 31352 17134
rect 31300 17070 31352 17076
rect 31300 16788 31352 16794
rect 31300 16730 31352 16736
rect 31208 16244 31260 16250
rect 31208 16186 31260 16192
rect 30932 16108 30984 16114
rect 30932 16050 30984 16056
rect 31116 15428 31168 15434
rect 31116 15370 31168 15376
rect 31024 15360 31076 15366
rect 31024 15302 31076 15308
rect 30932 15020 30984 15026
rect 30932 14962 30984 14968
rect 30944 14618 30972 14962
rect 30932 14612 30984 14618
rect 30932 14554 30984 14560
rect 30748 14476 30800 14482
rect 30748 14418 30800 14424
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30852 13530 30880 14350
rect 30840 13524 30892 13530
rect 30840 13466 30892 13472
rect 30838 13152 30894 13161
rect 30838 13087 30894 13096
rect 30852 12434 30880 13087
rect 30760 12406 30880 12434
rect 30656 5840 30708 5846
rect 30656 5782 30708 5788
rect 29736 5364 29788 5370
rect 29736 5306 29788 5312
rect 29644 5160 29696 5166
rect 29644 5102 29696 5108
rect 29656 4758 29684 5102
rect 29748 4758 29776 5306
rect 29644 4752 29696 4758
rect 29644 4694 29696 4700
rect 29736 4752 29788 4758
rect 29736 4694 29788 4700
rect 30760 4690 30788 12406
rect 31036 8430 31064 15302
rect 31128 15094 31156 15370
rect 31116 15088 31168 15094
rect 31116 15030 31168 15036
rect 31206 15056 31262 15065
rect 31206 14991 31262 15000
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 30840 5024 30892 5030
rect 30840 4966 30892 4972
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 30852 2650 30880 4966
rect 31220 4010 31248 14991
rect 31312 14958 31340 16730
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31300 14952 31352 14958
rect 31300 14894 31352 14900
rect 31300 11076 31352 11082
rect 31300 11018 31352 11024
rect 31312 9178 31340 11018
rect 31404 10305 31432 16594
rect 31496 16046 31524 17632
rect 31680 17270 31708 17983
rect 31772 17649 31800 18634
rect 32048 18358 32076 23446
rect 32140 21350 32168 26302
rect 32494 26302 32904 26330
rect 32494 26200 32550 26302
rect 32680 24948 32732 24954
rect 32680 24890 32732 24896
rect 32586 24440 32642 24449
rect 32586 24375 32642 24384
rect 32220 24268 32272 24274
rect 32220 24210 32272 24216
rect 32232 23798 32260 24210
rect 32220 23792 32272 23798
rect 32220 23734 32272 23740
rect 32312 23724 32364 23730
rect 32312 23666 32364 23672
rect 32324 23322 32352 23666
rect 32220 23316 32272 23322
rect 32220 23258 32272 23264
rect 32312 23316 32364 23322
rect 32312 23258 32364 23264
rect 32128 21344 32180 21350
rect 32128 21286 32180 21292
rect 32128 21004 32180 21010
rect 32128 20946 32180 20952
rect 32140 19718 32168 20946
rect 32232 20806 32260 23258
rect 32402 23216 32458 23225
rect 32402 23151 32458 23160
rect 32496 23180 32548 23186
rect 32220 20800 32272 20806
rect 32220 20742 32272 20748
rect 32312 20460 32364 20466
rect 32312 20402 32364 20408
rect 32220 20256 32272 20262
rect 32220 20198 32272 20204
rect 32232 19854 32260 20198
rect 32220 19848 32272 19854
rect 32220 19790 32272 19796
rect 32128 19712 32180 19718
rect 32128 19654 32180 19660
rect 32220 19712 32272 19718
rect 32220 19654 32272 19660
rect 32128 19372 32180 19378
rect 32128 19314 32180 19320
rect 32140 18426 32168 19314
rect 32232 18766 32260 19654
rect 32324 19514 32352 20402
rect 32312 19508 32364 19514
rect 32312 19450 32364 19456
rect 32312 19168 32364 19174
rect 32312 19110 32364 19116
rect 32324 18766 32352 19110
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32312 18760 32364 18766
rect 32312 18702 32364 18708
rect 32128 18420 32180 18426
rect 32128 18362 32180 18368
rect 32036 18352 32088 18358
rect 32036 18294 32088 18300
rect 32416 18272 32444 23151
rect 32496 23122 32548 23128
rect 32508 22778 32536 23122
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32508 21078 32536 22374
rect 32600 21622 32628 24375
rect 32588 21616 32640 21622
rect 32588 21558 32640 21564
rect 32588 21344 32640 21350
rect 32588 21286 32640 21292
rect 32496 21072 32548 21078
rect 32496 21014 32548 21020
rect 32600 21010 32628 21286
rect 32588 21004 32640 21010
rect 32588 20946 32640 20952
rect 32588 20052 32640 20058
rect 32588 19994 32640 20000
rect 32496 18760 32548 18766
rect 32496 18702 32548 18708
rect 32508 18601 32536 18702
rect 32494 18592 32550 18601
rect 32494 18527 32550 18536
rect 32232 18244 32444 18272
rect 32036 17672 32088 17678
rect 31758 17640 31814 17649
rect 32036 17614 32088 17620
rect 31758 17575 31814 17584
rect 32048 17338 32076 17614
rect 32036 17332 32088 17338
rect 32036 17274 32088 17280
rect 31668 17264 31720 17270
rect 31668 17206 31720 17212
rect 31944 17060 31996 17066
rect 31944 17002 31996 17008
rect 31666 16824 31722 16833
rect 31666 16759 31722 16768
rect 31680 16114 31708 16759
rect 31852 16244 31904 16250
rect 31852 16186 31904 16192
rect 31668 16108 31720 16114
rect 31668 16050 31720 16056
rect 31760 16108 31812 16114
rect 31760 16050 31812 16056
rect 31484 16040 31536 16046
rect 31484 15982 31536 15988
rect 31574 16008 31630 16017
rect 31574 15943 31630 15952
rect 31588 15910 31616 15943
rect 31576 15904 31628 15910
rect 31576 15846 31628 15852
rect 31668 15904 31720 15910
rect 31668 15846 31720 15852
rect 31680 15706 31708 15846
rect 31772 15706 31800 16050
rect 31668 15700 31720 15706
rect 31668 15642 31720 15648
rect 31760 15700 31812 15706
rect 31760 15642 31812 15648
rect 31864 15638 31892 16186
rect 31852 15632 31904 15638
rect 31758 15600 31814 15609
rect 31852 15574 31904 15580
rect 31758 15535 31814 15544
rect 31668 15496 31720 15502
rect 31668 15438 31720 15444
rect 31680 14822 31708 15438
rect 31576 14816 31628 14822
rect 31576 14758 31628 14764
rect 31668 14816 31720 14822
rect 31668 14758 31720 14764
rect 31588 12850 31616 14758
rect 31576 12844 31628 12850
rect 31576 12786 31628 12792
rect 31680 12238 31708 14758
rect 31668 12232 31720 12238
rect 31668 12174 31720 12180
rect 31390 10296 31446 10305
rect 31390 10231 31446 10240
rect 31300 9172 31352 9178
rect 31300 9114 31352 9120
rect 31772 5302 31800 15535
rect 31852 14544 31904 14550
rect 31852 14486 31904 14492
rect 31864 9518 31892 14486
rect 31956 13569 31984 17002
rect 32232 15638 32260 18244
rect 32600 17490 32628 19994
rect 32692 19961 32720 24890
rect 32876 21622 32904 26302
rect 33138 26302 33640 26330
rect 33138 26200 33194 26302
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 33416 23248 33468 23254
rect 33416 23190 33468 23196
rect 33140 23112 33192 23118
rect 33140 23054 33192 23060
rect 33048 22976 33100 22982
rect 33048 22918 33100 22924
rect 33060 22506 33088 22918
rect 33152 22545 33180 23054
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 33138 22536 33194 22545
rect 33048 22500 33100 22506
rect 33138 22471 33194 22480
rect 33048 22442 33100 22448
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33336 22098 33364 22578
rect 33324 22092 33376 22098
rect 33324 22034 33376 22040
rect 33428 22030 33456 23190
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33048 22024 33100 22030
rect 32968 21972 33048 21978
rect 32968 21966 33100 21972
rect 33416 22024 33468 22030
rect 33416 21966 33468 21972
rect 32968 21950 33088 21966
rect 32772 21616 32824 21622
rect 32772 21558 32824 21564
rect 32864 21616 32916 21622
rect 32864 21558 32916 21564
rect 32784 21026 32812 21558
rect 32968 21434 32996 21950
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33060 21690 33088 21830
rect 33048 21684 33100 21690
rect 33048 21626 33100 21632
rect 33324 21548 33376 21554
rect 33520 21536 33548 22918
rect 33376 21508 33548 21536
rect 33324 21490 33376 21496
rect 32876 21406 32996 21434
rect 32876 21146 32904 21406
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32864 21140 32916 21146
rect 32864 21082 32916 21088
rect 32784 20998 33088 21026
rect 33060 20262 33088 20998
rect 33520 20942 33548 21286
rect 33508 20936 33560 20942
rect 33508 20878 33560 20884
rect 33414 20632 33470 20641
rect 33414 20567 33470 20576
rect 33428 20466 33456 20567
rect 33416 20460 33468 20466
rect 33416 20402 33468 20408
rect 33048 20256 33100 20262
rect 33048 20198 33100 20204
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33140 19984 33192 19990
rect 32678 19952 32734 19961
rect 33140 19926 33192 19932
rect 32678 19887 32734 19896
rect 33048 19780 33100 19786
rect 33048 19722 33100 19728
rect 32770 19408 32826 19417
rect 32770 19343 32826 19352
rect 32508 17462 32628 17490
rect 32680 17536 32732 17542
rect 32680 17478 32732 17484
rect 32404 16992 32456 16998
rect 32404 16934 32456 16940
rect 32312 16652 32364 16658
rect 32312 16594 32364 16600
rect 32220 15632 32272 15638
rect 32220 15574 32272 15580
rect 32036 15496 32088 15502
rect 32036 15438 32088 15444
rect 31942 13560 31998 13569
rect 31942 13495 31998 13504
rect 32048 9654 32076 15438
rect 32220 15360 32272 15366
rect 32220 15302 32272 15308
rect 32232 11626 32260 15302
rect 32220 11620 32272 11626
rect 32220 11562 32272 11568
rect 32232 11354 32260 11562
rect 32220 11348 32272 11354
rect 32220 11290 32272 11296
rect 32036 9648 32088 9654
rect 32036 9590 32088 9596
rect 31852 9512 31904 9518
rect 31852 9454 31904 9460
rect 32324 8362 32352 16594
rect 32416 15978 32444 16934
rect 32404 15972 32456 15978
rect 32404 15914 32456 15920
rect 32508 15366 32536 17462
rect 32588 16584 32640 16590
rect 32588 16526 32640 16532
rect 32600 15366 32628 16526
rect 32692 16250 32720 17478
rect 32784 17134 32812 19343
rect 33060 19242 33088 19722
rect 33152 19310 33180 19926
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33048 19236 33100 19242
rect 33048 19178 33100 19184
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 33414 19000 33470 19009
rect 33324 18964 33376 18970
rect 33376 18944 33414 18952
rect 33376 18935 33470 18944
rect 33376 18924 33456 18935
rect 33324 18906 33376 18912
rect 32862 18728 32918 18737
rect 32862 18663 32918 18672
rect 32876 17814 32904 18663
rect 32956 18624 33008 18630
rect 32956 18566 33008 18572
rect 33508 18624 33560 18630
rect 33508 18566 33560 18572
rect 32968 18222 32996 18566
rect 32956 18216 33008 18222
rect 32956 18158 33008 18164
rect 33416 18216 33468 18222
rect 33416 18158 33468 18164
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 32864 17808 32916 17814
rect 32864 17750 32916 17756
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 32772 17128 32824 17134
rect 32772 17070 32824 17076
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33336 16674 33364 17614
rect 33244 16646 33364 16674
rect 33244 16454 33272 16646
rect 33324 16584 33376 16590
rect 33324 16526 33376 16532
rect 33232 16448 33284 16454
rect 33232 16390 33284 16396
rect 32680 16244 32732 16250
rect 32680 16186 32732 16192
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32404 11756 32456 11762
rect 32404 11698 32456 11704
rect 32312 8356 32364 8362
rect 32312 8298 32364 8304
rect 31760 5296 31812 5302
rect 31760 5238 31812 5244
rect 31772 4826 31800 5238
rect 31760 4820 31812 4826
rect 31760 4762 31812 4768
rect 31208 4004 31260 4010
rect 31208 3946 31260 3952
rect 30840 2644 30892 2650
rect 30840 2586 30892 2592
rect 32416 2582 32444 11698
rect 32600 10606 32628 15302
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32588 10600 32640 10606
rect 32588 10542 32640 10548
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 33336 9994 33364 16526
rect 33428 11830 33456 18158
rect 33520 15162 33548 18566
rect 33612 18426 33640 26302
rect 33704 23866 33732 26794
rect 33782 26330 33838 27000
rect 34426 26330 34482 27000
rect 34612 26648 34664 26654
rect 34612 26590 34664 26596
rect 33782 26302 34192 26330
rect 33782 26200 33838 26302
rect 33876 26172 33928 26178
rect 33876 26114 33928 26120
rect 33784 25560 33836 25566
rect 33784 25502 33836 25508
rect 33692 23860 33744 23866
rect 33692 23802 33744 23808
rect 33796 22094 33824 25502
rect 33704 22066 33824 22094
rect 33704 18970 33732 22066
rect 33692 18964 33744 18970
rect 33692 18906 33744 18912
rect 33784 18760 33836 18766
rect 33784 18702 33836 18708
rect 33692 18692 33744 18698
rect 33692 18634 33744 18640
rect 33600 18420 33652 18426
rect 33600 18362 33652 18368
rect 33508 15156 33560 15162
rect 33508 15098 33560 15104
rect 33600 15020 33652 15026
rect 33600 14962 33652 14968
rect 33612 14822 33640 14962
rect 33600 14816 33652 14822
rect 33600 14758 33652 14764
rect 33416 11824 33468 11830
rect 33416 11766 33468 11772
rect 33324 9988 33376 9994
rect 33324 9930 33376 9936
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32772 9104 32824 9110
rect 32772 9046 32824 9052
rect 32784 2961 32812 9046
rect 33704 8537 33732 18634
rect 33690 8528 33746 8537
rect 33690 8463 33746 8472
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 33508 5092 33560 5098
rect 33508 5034 33560 5040
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32770 2952 32826 2961
rect 32770 2887 32826 2896
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33520 2650 33548 5034
rect 33508 2644 33560 2650
rect 33508 2586 33560 2592
rect 32404 2576 32456 2582
rect 32404 2518 32456 2524
rect 30748 2440 30800 2446
rect 30748 2382 30800 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 30760 800 30788 2382
rect 33428 800 33456 2382
rect 33796 2009 33824 18702
rect 33888 16658 33916 26114
rect 33968 23044 34020 23050
rect 33968 22986 34020 22992
rect 33980 22642 34008 22986
rect 34164 22681 34192 26302
rect 34256 26302 34482 26330
rect 34150 22672 34206 22681
rect 33968 22636 34020 22642
rect 34150 22607 34206 22616
rect 33968 22578 34020 22584
rect 34152 20800 34204 20806
rect 34152 20742 34204 20748
rect 34164 20602 34192 20742
rect 34152 20596 34204 20602
rect 34152 20538 34204 20544
rect 34060 20392 34112 20398
rect 34060 20334 34112 20340
rect 34072 19922 34100 20334
rect 34060 19916 34112 19922
rect 34060 19858 34112 19864
rect 34060 19712 34112 19718
rect 34060 19654 34112 19660
rect 34072 19553 34100 19654
rect 34058 19544 34114 19553
rect 34058 19479 34114 19488
rect 34256 18970 34284 26302
rect 34426 26200 34482 26302
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 34348 22817 34376 24142
rect 34334 22808 34390 22817
rect 34334 22743 34336 22752
rect 34388 22743 34390 22752
rect 34336 22714 34388 22720
rect 34520 22024 34572 22030
rect 34520 21966 34572 21972
rect 34336 21888 34388 21894
rect 34336 21830 34388 21836
rect 34428 21888 34480 21894
rect 34428 21830 34480 21836
rect 34348 21729 34376 21830
rect 34334 21720 34390 21729
rect 34334 21655 34390 21664
rect 34440 21554 34468 21830
rect 34428 21548 34480 21554
rect 34428 21490 34480 21496
rect 34532 21457 34560 21966
rect 34518 21448 34574 21457
rect 34518 21383 34574 21392
rect 34624 20602 34652 26590
rect 35070 26200 35126 27000
rect 35714 26200 35770 27000
rect 36358 26200 36414 27000
rect 36544 26716 36596 26722
rect 36544 26658 36596 26664
rect 34704 25968 34756 25974
rect 34704 25910 34756 25916
rect 34716 21146 34744 25910
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34808 22506 34836 22918
rect 34796 22500 34848 22506
rect 34796 22442 34848 22448
rect 34808 21962 34836 22442
rect 35084 22166 35112 26200
rect 35624 24132 35676 24138
rect 35624 24074 35676 24080
rect 35440 24064 35492 24070
rect 35440 24006 35492 24012
rect 35452 22778 35480 24006
rect 35636 23730 35664 24074
rect 35624 23724 35676 23730
rect 35624 23666 35676 23672
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35072 22160 35124 22166
rect 35072 22102 35124 22108
rect 34980 22024 35032 22030
rect 34980 21966 35032 21972
rect 34796 21956 34848 21962
rect 34796 21898 34848 21904
rect 34992 21486 35020 21966
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 35636 21554 35664 21830
rect 35624 21548 35676 21554
rect 35624 21490 35676 21496
rect 34980 21480 35032 21486
rect 34980 21422 35032 21428
rect 35256 21344 35308 21350
rect 35256 21286 35308 21292
rect 34704 21140 34756 21146
rect 34704 21082 34756 21088
rect 34612 20596 34664 20602
rect 34612 20538 34664 20544
rect 34336 20392 34388 20398
rect 34334 20360 34336 20369
rect 34388 20360 34390 20369
rect 34334 20295 34390 20304
rect 34428 19848 34480 19854
rect 34428 19790 34480 19796
rect 34336 19168 34388 19174
rect 34336 19110 34388 19116
rect 34244 18964 34296 18970
rect 34244 18906 34296 18912
rect 34348 18698 34376 19110
rect 34336 18692 34388 18698
rect 34336 18634 34388 18640
rect 34244 18284 34296 18290
rect 34244 18226 34296 18232
rect 34060 17536 34112 17542
rect 34060 17478 34112 17484
rect 34072 17202 34100 17478
rect 34060 17196 34112 17202
rect 34060 17138 34112 17144
rect 33876 16652 33928 16658
rect 33876 16594 33928 16600
rect 33876 15496 33928 15502
rect 33876 15438 33928 15444
rect 33888 6458 33916 15438
rect 34072 6769 34100 17138
rect 34256 10713 34284 18226
rect 34440 17105 34468 19790
rect 35164 19712 35216 19718
rect 35164 19654 35216 19660
rect 34612 19236 34664 19242
rect 34612 19178 34664 19184
rect 34624 19009 34652 19178
rect 34610 19000 34666 19009
rect 34610 18935 34666 18944
rect 34888 18760 34940 18766
rect 34888 18702 34940 18708
rect 34900 18630 34928 18702
rect 34888 18624 34940 18630
rect 34888 18566 34940 18572
rect 34520 18216 34572 18222
rect 34520 18158 34572 18164
rect 34532 17338 34560 18158
rect 34612 17672 34664 17678
rect 34612 17614 34664 17620
rect 34624 17542 34652 17614
rect 34612 17536 34664 17542
rect 34612 17478 34664 17484
rect 34520 17332 34572 17338
rect 34520 17274 34572 17280
rect 34520 17196 34572 17202
rect 34520 17138 34572 17144
rect 34426 17096 34482 17105
rect 34426 17031 34482 17040
rect 34532 11898 34560 17138
rect 34624 16590 34652 17478
rect 34796 17128 34848 17134
rect 34796 17070 34848 17076
rect 34704 16992 34756 16998
rect 34704 16934 34756 16940
rect 34612 16584 34664 16590
rect 34612 16526 34664 16532
rect 34520 11892 34572 11898
rect 34520 11834 34572 11840
rect 34242 10704 34298 10713
rect 34242 10639 34298 10648
rect 34058 6760 34114 6769
rect 34058 6695 34114 6704
rect 33876 6452 33928 6458
rect 33876 6394 33928 6400
rect 34716 4758 34744 16934
rect 34808 14929 34836 17070
rect 34900 16153 34928 18566
rect 35176 16794 35204 19654
rect 35164 16788 35216 16794
rect 35164 16730 35216 16736
rect 34980 16516 35032 16522
rect 34980 16458 35032 16464
rect 34886 16144 34942 16153
rect 34886 16079 34942 16088
rect 34794 14920 34850 14929
rect 34794 14855 34850 14864
rect 34704 4752 34756 4758
rect 34704 4694 34756 4700
rect 33782 2000 33838 2009
rect 33782 1935 33838 1944
rect 29090 640 29146 649
rect 29090 575 29146 584
rect 30746 0 30802 800
rect 33414 0 33470 800
rect 34992 746 35020 16458
rect 35072 16448 35124 16454
rect 35072 16390 35124 16396
rect 35084 15201 35112 16390
rect 35070 15192 35126 15201
rect 35070 15127 35126 15136
rect 35268 13161 35296 21286
rect 35440 20936 35492 20942
rect 35440 20878 35492 20884
rect 35254 13152 35310 13161
rect 35254 13087 35310 13096
rect 35452 1222 35480 20878
rect 35532 20460 35584 20466
rect 35532 20402 35584 20408
rect 35544 20058 35572 20402
rect 35532 20052 35584 20058
rect 35532 19994 35584 20000
rect 35532 19372 35584 19378
rect 35532 19314 35584 19320
rect 35544 17377 35572 19314
rect 35728 18970 35756 26200
rect 36176 25152 36228 25158
rect 36176 25094 36228 25100
rect 35808 25016 35860 25022
rect 35808 24958 35860 24964
rect 35820 23474 35848 24958
rect 35992 23520 36044 23526
rect 35820 23446 35940 23474
rect 35992 23462 36044 23468
rect 35912 22778 35940 23446
rect 36004 23118 36032 23462
rect 35992 23112 36044 23118
rect 35992 23054 36044 23060
rect 35900 22772 35952 22778
rect 35900 22714 35952 22720
rect 36084 21956 36136 21962
rect 36084 21898 36136 21904
rect 35900 21548 35952 21554
rect 35900 21490 35952 21496
rect 35912 20602 35940 21490
rect 35992 21344 36044 21350
rect 35992 21286 36044 21292
rect 35900 20596 35952 20602
rect 35900 20538 35952 20544
rect 36004 20466 36032 21286
rect 36096 21049 36124 21898
rect 36082 21040 36138 21049
rect 36188 21010 36216 25094
rect 36372 23254 36400 26200
rect 36360 23248 36412 23254
rect 36360 23190 36412 23196
rect 36556 21690 36584 26658
rect 37002 26330 37058 27000
rect 36820 26308 36872 26314
rect 36820 26250 36872 26256
rect 36924 26302 37058 26330
rect 36636 25220 36688 25226
rect 36636 25162 36688 25168
rect 36648 24342 36676 25162
rect 36636 24336 36688 24342
rect 36636 24278 36688 24284
rect 36832 23118 36860 26250
rect 36820 23112 36872 23118
rect 36820 23054 36872 23060
rect 36832 22778 36860 23054
rect 36820 22772 36872 22778
rect 36820 22714 36872 22720
rect 36544 21684 36596 21690
rect 36544 21626 36596 21632
rect 36544 21344 36596 21350
rect 36544 21286 36596 21292
rect 36082 20975 36138 20984
rect 36176 21004 36228 21010
rect 36176 20946 36228 20952
rect 36268 20936 36320 20942
rect 36268 20878 36320 20884
rect 35992 20460 36044 20466
rect 35992 20402 36044 20408
rect 35992 19712 36044 19718
rect 35992 19654 36044 19660
rect 36004 19378 36032 19654
rect 35992 19372 36044 19378
rect 35992 19314 36044 19320
rect 35624 18964 35676 18970
rect 35624 18906 35676 18912
rect 35716 18964 35768 18970
rect 35716 18906 35768 18912
rect 35636 18630 35664 18906
rect 35806 18864 35862 18873
rect 35806 18799 35862 18808
rect 35624 18624 35676 18630
rect 35624 18566 35676 18572
rect 35820 18290 35848 18799
rect 35808 18284 35860 18290
rect 35808 18226 35860 18232
rect 35898 17912 35954 17921
rect 35898 17847 35954 17856
rect 35912 17678 35940 17847
rect 36280 17746 36308 20878
rect 36452 18080 36504 18086
rect 36452 18022 36504 18028
rect 36268 17740 36320 17746
rect 36268 17682 36320 17688
rect 35900 17672 35952 17678
rect 35900 17614 35952 17620
rect 35530 17368 35586 17377
rect 35912 17338 35940 17614
rect 36084 17536 36136 17542
rect 36084 17478 36136 17484
rect 35530 17303 35586 17312
rect 35900 17332 35952 17338
rect 35900 17274 35952 17280
rect 35992 17128 36044 17134
rect 35992 17070 36044 17076
rect 36004 12374 36032 17070
rect 35992 12368 36044 12374
rect 35992 12310 36044 12316
rect 36096 10674 36124 17478
rect 36464 16046 36492 18022
rect 36452 16040 36504 16046
rect 36452 15982 36504 15988
rect 36556 13802 36584 21286
rect 36728 20596 36780 20602
rect 36728 20538 36780 20544
rect 36636 20392 36688 20398
rect 36636 20334 36688 20340
rect 36648 19514 36676 20334
rect 36740 19689 36768 20538
rect 36726 19680 36782 19689
rect 36726 19615 36782 19624
rect 36636 19508 36688 19514
rect 36636 19450 36688 19456
rect 36636 19304 36688 19310
rect 36636 19246 36688 19252
rect 36648 19174 36676 19246
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36648 17814 36676 19110
rect 36924 18426 36952 26302
rect 37002 26200 37058 26302
rect 37280 26240 37332 26246
rect 37646 26200 37702 27000
rect 38290 26330 38346 27000
rect 38290 26302 38424 26330
rect 38290 26200 38346 26302
rect 37280 26182 37332 26188
rect 37004 25832 37056 25838
rect 37004 25774 37056 25780
rect 37016 24342 37044 25774
rect 37004 24336 37056 24342
rect 37004 24278 37056 24284
rect 37096 23520 37148 23526
rect 37096 23462 37148 23468
rect 37108 23186 37136 23462
rect 37096 23180 37148 23186
rect 37096 23122 37148 23128
rect 37094 23080 37150 23089
rect 37094 23015 37150 23024
rect 37108 22982 37136 23015
rect 37096 22976 37148 22982
rect 37096 22918 37148 22924
rect 37188 22636 37240 22642
rect 37188 22578 37240 22584
rect 37004 22500 37056 22506
rect 37004 22442 37056 22448
rect 37016 22098 37044 22442
rect 37200 22098 37228 22578
rect 37004 22092 37056 22098
rect 37004 22034 37056 22040
rect 37188 22092 37240 22098
rect 37292 22094 37320 26182
rect 37464 24608 37516 24614
rect 37464 24550 37516 24556
rect 37476 24206 37504 24550
rect 37372 24200 37424 24206
rect 37372 24142 37424 24148
rect 37464 24200 37516 24206
rect 37464 24142 37516 24148
rect 37384 22778 37412 24142
rect 37464 24064 37516 24070
rect 37464 24006 37516 24012
rect 37372 22772 37424 22778
rect 37372 22714 37424 22720
rect 37476 22642 37504 24006
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37292 22066 37412 22094
rect 37188 22034 37240 22040
rect 37096 21956 37148 21962
rect 37096 21898 37148 21904
rect 37108 21690 37136 21898
rect 37188 21888 37240 21894
rect 37188 21830 37240 21836
rect 37096 21684 37148 21690
rect 37096 21626 37148 21632
rect 37004 21480 37056 21486
rect 37004 21422 37056 21428
rect 37016 21350 37044 21422
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 37200 21078 37228 21830
rect 37188 21072 37240 21078
rect 37188 21014 37240 21020
rect 37384 20466 37412 22066
rect 37372 20460 37424 20466
rect 37372 20402 37424 20408
rect 37004 20256 37056 20262
rect 37004 20198 37056 20204
rect 37016 19786 37044 20198
rect 37096 19848 37148 19854
rect 37096 19790 37148 19796
rect 37004 19780 37056 19786
rect 37004 19722 37056 19728
rect 36912 18420 36964 18426
rect 36912 18362 36964 18368
rect 36818 18320 36874 18329
rect 36818 18255 36874 18264
rect 36832 18222 36860 18255
rect 36820 18216 36872 18222
rect 36820 18158 36872 18164
rect 36728 18080 36780 18086
rect 36728 18022 36780 18028
rect 36636 17808 36688 17814
rect 36636 17750 36688 17756
rect 36544 13796 36596 13802
rect 36544 13738 36596 13744
rect 36740 12986 36768 18022
rect 36912 17808 36964 17814
rect 36910 17776 36912 17785
rect 36964 17776 36966 17785
rect 36910 17711 36966 17720
rect 37016 17678 37044 19722
rect 37108 18970 37136 19790
rect 37660 19786 37688 26200
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 37738 23624 37794 23633
rect 37738 23559 37794 23568
rect 37752 21554 37780 23559
rect 38292 23044 38344 23050
rect 38292 22986 38344 22992
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37832 22024 37884 22030
rect 37832 21966 37884 21972
rect 37844 21690 37872 21966
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 38304 21690 38332 22986
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 38292 21684 38344 21690
rect 38292 21626 38344 21632
rect 37740 21548 37792 21554
rect 37740 21490 37792 21496
rect 38200 21344 38252 21350
rect 38200 21286 38252 21292
rect 38212 20942 38240 21286
rect 38200 20936 38252 20942
rect 38200 20878 38252 20884
rect 37740 20800 37792 20806
rect 37740 20742 37792 20748
rect 37648 19780 37700 19786
rect 37648 19722 37700 19728
rect 37556 19712 37608 19718
rect 37556 19654 37608 19660
rect 37096 18964 37148 18970
rect 37096 18906 37148 18912
rect 37464 18760 37516 18766
rect 37464 18702 37516 18708
rect 37188 18284 37240 18290
rect 37188 18226 37240 18232
rect 37200 18086 37228 18226
rect 37188 18080 37240 18086
rect 37188 18022 37240 18028
rect 37476 17882 37504 18702
rect 37464 17876 37516 17882
rect 37464 17818 37516 17824
rect 37004 17672 37056 17678
rect 37004 17614 37056 17620
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 37372 17536 37424 17542
rect 37370 17504 37372 17513
rect 37424 17504 37426 17513
rect 37370 17439 37426 17448
rect 37280 17196 37332 17202
rect 37280 17138 37332 17144
rect 37292 15570 37320 17138
rect 37280 15564 37332 15570
rect 37280 15506 37332 15512
rect 36728 12980 36780 12986
rect 36728 12922 36780 12928
rect 37476 12209 37504 17614
rect 37568 13326 37596 19654
rect 37752 18358 37780 20742
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 38396 19446 38424 26302
rect 38934 26200 38990 27000
rect 39578 26200 39634 27000
rect 40222 26200 40278 27000
rect 40866 26200 40922 27000
rect 40960 26444 41012 26450
rect 40960 26386 41012 26392
rect 38568 23520 38620 23526
rect 38568 23462 38620 23468
rect 38580 22642 38608 23462
rect 38948 22778 38976 26200
rect 39120 26104 39172 26110
rect 39120 26046 39172 26052
rect 38936 22772 38988 22778
rect 38936 22714 38988 22720
rect 38568 22636 38620 22642
rect 38568 22578 38620 22584
rect 38844 22024 38896 22030
rect 38750 21992 38806 22001
rect 38844 21966 38896 21972
rect 38750 21927 38806 21936
rect 38764 21894 38792 21927
rect 38752 21888 38804 21894
rect 38752 21830 38804 21836
rect 38764 21554 38792 21830
rect 38752 21548 38804 21554
rect 38752 21490 38804 21496
rect 38856 21146 38884 21966
rect 38844 21140 38896 21146
rect 38844 21082 38896 21088
rect 39026 20496 39082 20505
rect 39026 20431 39028 20440
rect 39080 20431 39082 20440
rect 39028 20402 39080 20408
rect 38568 19780 38620 19786
rect 38568 19722 38620 19728
rect 38384 19440 38436 19446
rect 38384 19382 38436 19388
rect 38580 19378 38608 19722
rect 38660 19712 38712 19718
rect 38660 19654 38712 19660
rect 38476 19372 38528 19378
rect 38476 19314 38528 19320
rect 38568 19372 38620 19378
rect 38568 19314 38620 19320
rect 37832 18624 37884 18630
rect 37832 18566 37884 18572
rect 37740 18352 37792 18358
rect 37740 18294 37792 18300
rect 37648 18080 37700 18086
rect 37648 18022 37700 18028
rect 37660 14550 37688 18022
rect 37844 16726 37872 18566
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 38384 18080 38436 18086
rect 38384 18022 38436 18028
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 37832 16720 37884 16726
rect 37832 16662 37884 16668
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 37648 14544 37700 14550
rect 37648 14486 37700 14492
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 37556 13320 37608 13326
rect 37556 13262 37608 13268
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37462 12200 37518 12209
rect 37462 12135 37518 12144
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 36084 10668 36136 10674
rect 36084 10610 36136 10616
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 36360 8628 36412 8634
rect 36360 8570 36412 8576
rect 36372 2514 36400 8570
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 38396 6905 38424 18022
rect 38488 9042 38516 19314
rect 38672 18290 38700 19654
rect 39132 19310 39160 26046
rect 39212 25084 39264 25090
rect 39212 25026 39264 25032
rect 39224 22642 39252 25026
rect 39396 24336 39448 24342
rect 39396 24278 39448 24284
rect 39212 22636 39264 22642
rect 39212 22578 39264 22584
rect 39212 20936 39264 20942
rect 39212 20878 39264 20884
rect 39120 19304 39172 19310
rect 39120 19246 39172 19252
rect 38752 18624 38804 18630
rect 38752 18566 38804 18572
rect 38660 18284 38712 18290
rect 38660 18226 38712 18232
rect 38660 17876 38712 17882
rect 38660 17818 38712 17824
rect 38672 15473 38700 17818
rect 38764 15502 38792 18566
rect 38936 18080 38988 18086
rect 38936 18022 38988 18028
rect 38948 17066 38976 18022
rect 39224 17134 39252 20878
rect 39304 20800 39356 20806
rect 39304 20742 39356 20748
rect 39316 17610 39344 20742
rect 39408 20482 39436 24278
rect 39488 24064 39540 24070
rect 39488 24006 39540 24012
rect 39500 23066 39528 24006
rect 39592 23254 39620 26200
rect 39764 26036 39816 26042
rect 39764 25978 39816 25984
rect 39672 24064 39724 24070
rect 39672 24006 39724 24012
rect 39684 23730 39712 24006
rect 39672 23724 39724 23730
rect 39672 23666 39724 23672
rect 39580 23248 39632 23254
rect 39580 23190 39632 23196
rect 39500 23038 39620 23066
rect 39488 22976 39540 22982
rect 39488 22918 39540 22924
rect 39500 21554 39528 22918
rect 39592 22624 39620 23038
rect 39776 22982 39804 25978
rect 39948 23588 40000 23594
rect 39948 23530 40000 23536
rect 39764 22976 39816 22982
rect 39764 22918 39816 22924
rect 39672 22636 39724 22642
rect 39592 22596 39672 22624
rect 39672 22578 39724 22584
rect 39684 22234 39712 22578
rect 39672 22228 39724 22234
rect 39672 22170 39724 22176
rect 39488 21548 39540 21554
rect 39488 21490 39540 21496
rect 39856 21548 39908 21554
rect 39856 21490 39908 21496
rect 39488 21344 39540 21350
rect 39488 21286 39540 21292
rect 39500 20942 39528 21286
rect 39488 20936 39540 20942
rect 39488 20878 39540 20884
rect 39408 20454 39712 20482
rect 39488 20392 39540 20398
rect 39488 20334 39540 20340
rect 39396 19848 39448 19854
rect 39396 19790 39448 19796
rect 39408 19242 39436 19790
rect 39396 19236 39448 19242
rect 39396 19178 39448 19184
rect 39304 17604 39356 17610
rect 39304 17546 39356 17552
rect 39212 17128 39264 17134
rect 39212 17070 39264 17076
rect 38936 17060 38988 17066
rect 38936 17002 38988 17008
rect 38752 15496 38804 15502
rect 38658 15464 38714 15473
rect 38752 15438 38804 15444
rect 38658 15399 38714 15408
rect 38476 9036 38528 9042
rect 38476 8978 38528 8984
rect 39408 8090 39436 19178
rect 39500 19174 39528 20334
rect 39488 19168 39540 19174
rect 39488 19110 39540 19116
rect 39580 18964 39632 18970
rect 39580 18906 39632 18912
rect 39592 8401 39620 18906
rect 39684 13734 39712 20454
rect 39868 18222 39896 21490
rect 39856 18216 39908 18222
rect 39856 18158 39908 18164
rect 39672 13728 39724 13734
rect 39672 13670 39724 13676
rect 39960 12889 39988 23530
rect 40040 23112 40092 23118
rect 40040 23054 40092 23060
rect 40052 22574 40080 23054
rect 40040 22568 40092 22574
rect 40040 22510 40092 22516
rect 40132 22432 40184 22438
rect 40132 22374 40184 22380
rect 40144 21962 40172 22374
rect 40236 22234 40264 26200
rect 40316 25492 40368 25498
rect 40316 25434 40368 25440
rect 40328 23866 40356 25434
rect 40408 25424 40460 25430
rect 40408 25366 40460 25372
rect 40316 23860 40368 23866
rect 40316 23802 40368 23808
rect 40316 23044 40368 23050
rect 40316 22986 40368 22992
rect 40224 22228 40276 22234
rect 40224 22170 40276 22176
rect 40132 21956 40184 21962
rect 40132 21898 40184 21904
rect 40224 21344 40276 21350
rect 40224 21286 40276 21292
rect 40040 20936 40092 20942
rect 40040 20878 40092 20884
rect 40052 20058 40080 20878
rect 40040 20052 40092 20058
rect 40040 19994 40092 20000
rect 40236 19514 40264 21286
rect 40328 20466 40356 22986
rect 40420 22098 40448 25366
rect 40500 23656 40552 23662
rect 40500 23598 40552 23604
rect 40512 23322 40540 23598
rect 40500 23316 40552 23322
rect 40500 23258 40552 23264
rect 40500 22772 40552 22778
rect 40500 22714 40552 22720
rect 40408 22092 40460 22098
rect 40408 22034 40460 22040
rect 40408 21956 40460 21962
rect 40408 21898 40460 21904
rect 40316 20460 40368 20466
rect 40316 20402 40368 20408
rect 40224 19508 40276 19514
rect 40224 19450 40276 19456
rect 40224 19372 40276 19378
rect 40224 19314 40276 19320
rect 40236 18902 40264 19314
rect 40224 18896 40276 18902
rect 40224 18838 40276 18844
rect 40420 14822 40448 21898
rect 40512 19446 40540 22714
rect 40880 22438 40908 26200
rect 40868 22432 40920 22438
rect 40868 22374 40920 22380
rect 40684 22024 40736 22030
rect 40684 21966 40736 21972
rect 40696 21146 40724 21966
rect 40684 21140 40736 21146
rect 40684 21082 40736 21088
rect 40592 20256 40644 20262
rect 40592 20198 40644 20204
rect 40868 20256 40920 20262
rect 40868 20198 40920 20204
rect 40604 19786 40632 20198
rect 40880 19854 40908 20198
rect 40972 19990 41000 26386
rect 41510 26330 41566 27000
rect 41604 26512 41656 26518
rect 41604 26454 41656 26460
rect 41432 26302 41566 26330
rect 41144 25764 41196 25770
rect 41144 25706 41196 25712
rect 41156 23225 41184 25706
rect 41432 24206 41460 26302
rect 41510 26200 41566 26302
rect 41420 24200 41472 24206
rect 41420 24142 41472 24148
rect 41512 24200 41564 24206
rect 41512 24142 41564 24148
rect 41432 23866 41460 24142
rect 41420 23860 41472 23866
rect 41420 23802 41472 23808
rect 41236 23248 41288 23254
rect 41142 23216 41198 23225
rect 41236 23190 41288 23196
rect 41142 23151 41198 23160
rect 41156 23118 41184 23151
rect 41144 23112 41196 23118
rect 41144 23054 41196 23060
rect 41052 22976 41104 22982
rect 41052 22918 41104 22924
rect 41064 22642 41092 22918
rect 41052 22636 41104 22642
rect 41052 22578 41104 22584
rect 41248 20466 41276 23190
rect 41328 21412 41380 21418
rect 41328 21354 41380 21360
rect 41340 20874 41368 21354
rect 41328 20868 41380 20874
rect 41328 20810 41380 20816
rect 41236 20460 41288 20466
rect 41236 20402 41288 20408
rect 41248 20058 41276 20402
rect 41236 20052 41288 20058
rect 41236 19994 41288 20000
rect 40960 19984 41012 19990
rect 40960 19926 41012 19932
rect 40868 19848 40920 19854
rect 40868 19790 40920 19796
rect 40592 19780 40644 19786
rect 40592 19722 40644 19728
rect 40500 19440 40552 19446
rect 40500 19382 40552 19388
rect 40408 14816 40460 14822
rect 40408 14758 40460 14764
rect 40040 14000 40092 14006
rect 40040 13942 40092 13948
rect 39946 12880 40002 12889
rect 39946 12815 40002 12824
rect 40052 11762 40080 13942
rect 40040 11756 40092 11762
rect 40040 11698 40092 11704
rect 40604 9110 40632 19722
rect 40960 19712 41012 19718
rect 40960 19654 41012 19660
rect 40774 19272 40830 19281
rect 40774 19207 40830 19216
rect 40788 19174 40816 19207
rect 40776 19168 40828 19174
rect 40776 19110 40828 19116
rect 40972 11665 41000 19654
rect 41236 19508 41288 19514
rect 41236 19450 41288 19456
rect 41248 15434 41276 19450
rect 41236 15428 41288 15434
rect 41236 15370 41288 15376
rect 40958 11656 41014 11665
rect 40958 11591 41014 11600
rect 40592 9104 40644 9110
rect 40592 9046 40644 9052
rect 41340 8974 41368 20810
rect 41524 20534 41552 24142
rect 41616 22098 41644 26454
rect 42154 26200 42210 27000
rect 42798 26200 42854 27000
rect 42892 26580 42944 26586
rect 42892 26522 42944 26528
rect 42904 26058 42932 26522
rect 43442 26200 43498 27000
rect 44086 26200 44142 27000
rect 44730 26330 44786 27000
rect 44730 26302 45140 26330
rect 44730 26200 44786 26302
rect 42812 26030 42932 26058
rect 41880 25900 41932 25906
rect 41880 25842 41932 25848
rect 41788 23724 41840 23730
rect 41788 23666 41840 23672
rect 41800 23322 41828 23666
rect 41892 23594 41920 25842
rect 41970 25800 42026 25809
rect 41970 25735 42026 25744
rect 41880 23588 41932 23594
rect 41880 23530 41932 23536
rect 41788 23316 41840 23322
rect 41788 23258 41840 23264
rect 41880 22568 41932 22574
rect 41880 22510 41932 22516
rect 41696 22228 41748 22234
rect 41696 22170 41748 22176
rect 41604 22092 41656 22098
rect 41604 22034 41656 22040
rect 41512 20528 41564 20534
rect 41512 20470 41564 20476
rect 41420 20392 41472 20398
rect 41420 20334 41472 20340
rect 41432 15094 41460 20334
rect 41524 19514 41552 20470
rect 41708 19854 41736 22170
rect 41788 21548 41840 21554
rect 41788 21490 41840 21496
rect 41696 19848 41748 19854
rect 41696 19790 41748 19796
rect 41604 19712 41656 19718
rect 41604 19654 41656 19660
rect 41512 19508 41564 19514
rect 41512 19450 41564 19456
rect 41616 17338 41644 19654
rect 41800 19310 41828 21490
rect 41788 19304 41840 19310
rect 41788 19246 41840 19252
rect 41604 17332 41656 17338
rect 41604 17274 41656 17280
rect 41420 15088 41472 15094
rect 41420 15030 41472 15036
rect 41892 10577 41920 22510
rect 41984 21146 42012 25735
rect 42064 24948 42116 24954
rect 42064 24890 42116 24896
rect 41972 21140 42024 21146
rect 41972 21082 42024 21088
rect 42076 20942 42104 24890
rect 42812 24206 42840 26030
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 42800 24200 42852 24206
rect 42800 24142 42852 24148
rect 42708 24132 42760 24138
rect 42708 24074 42760 24080
rect 42720 23798 42748 24074
rect 42892 24064 42944 24070
rect 42892 24006 42944 24012
rect 42904 23798 42932 24006
rect 42708 23792 42760 23798
rect 42706 23760 42708 23769
rect 42892 23792 42944 23798
rect 42760 23760 42762 23769
rect 42892 23734 42944 23740
rect 43456 23746 43484 26200
rect 43628 25356 43680 25362
rect 43628 25298 43680 25304
rect 42706 23695 42762 23704
rect 42800 23724 42852 23730
rect 42800 23666 42852 23672
rect 43352 23724 43404 23730
rect 43456 23718 43576 23746
rect 43352 23666 43404 23672
rect 42812 23050 42840 23666
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 43168 23316 43220 23322
rect 43168 23258 43220 23264
rect 42800 23044 42852 23050
rect 42800 22986 42852 22992
rect 43180 22574 43208 23258
rect 43168 22568 43220 22574
rect 43168 22510 43220 22516
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43260 21888 43312 21894
rect 43260 21830 43312 21836
rect 43272 21690 43300 21830
rect 43260 21684 43312 21690
rect 43260 21626 43312 21632
rect 42524 21548 42576 21554
rect 42524 21490 42576 21496
rect 42064 20936 42116 20942
rect 42116 20896 42196 20924
rect 42064 20878 42116 20884
rect 42064 20800 42116 20806
rect 42064 20742 42116 20748
rect 41878 10568 41934 10577
rect 41878 10503 41934 10512
rect 41328 8968 41380 8974
rect 41328 8910 41380 8916
rect 39578 8392 39634 8401
rect 39578 8327 39634 8336
rect 39396 8084 39448 8090
rect 39396 8026 39448 8032
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 38382 6896 38438 6905
rect 38382 6831 38438 6840
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 36360 2508 36412 2514
rect 36360 2450 36412 2456
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 35440 1216 35492 1222
rect 35440 1158 35492 1164
rect 36096 800 36124 2382
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38764 800 38792 7686
rect 42076 6186 42104 20742
rect 42168 20058 42196 20896
rect 42156 20052 42208 20058
rect 42156 19994 42208 20000
rect 42536 19718 42564 21490
rect 42800 21344 42852 21350
rect 42800 21286 42852 21292
rect 42708 20868 42760 20874
rect 42708 20810 42760 20816
rect 42720 20330 42748 20810
rect 42708 20324 42760 20330
rect 42708 20266 42760 20272
rect 42524 19712 42576 19718
rect 42524 19654 42576 19660
rect 42536 14618 42564 19654
rect 42524 14612 42576 14618
rect 42524 14554 42576 14560
rect 42720 13530 42748 20266
rect 42812 14006 42840 21286
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43364 21026 43392 23666
rect 43444 23656 43496 23662
rect 43444 23598 43496 23604
rect 43456 23322 43484 23598
rect 43444 23316 43496 23322
rect 43444 23258 43496 23264
rect 43444 22432 43496 22438
rect 43444 22374 43496 22380
rect 43272 20998 43392 21026
rect 43272 20618 43300 20998
rect 43456 20942 43484 22374
rect 43548 22234 43576 23718
rect 43640 23254 43668 25298
rect 43718 24848 43774 24857
rect 43718 24783 43774 24792
rect 43628 23248 43680 23254
rect 43628 23190 43680 23196
rect 43732 22642 43760 24783
rect 43904 24200 43956 24206
rect 43904 24142 43956 24148
rect 43812 24064 43864 24070
rect 43812 24006 43864 24012
rect 43720 22636 43772 22642
rect 43720 22578 43772 22584
rect 43536 22228 43588 22234
rect 43536 22170 43588 22176
rect 43628 21548 43680 21554
rect 43628 21490 43680 21496
rect 43536 21344 43588 21350
rect 43536 21286 43588 21292
rect 43444 20936 43496 20942
rect 43350 20904 43406 20913
rect 43444 20878 43496 20884
rect 43350 20839 43406 20848
rect 43364 20806 43392 20839
rect 43352 20800 43404 20806
rect 43352 20742 43404 20748
rect 43272 20590 43392 20618
rect 43456 20602 43484 20878
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 42800 14000 42852 14006
rect 42800 13942 42852 13948
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 42708 13524 42760 13530
rect 42708 13466 42760 13472
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 42064 6180 42116 6186
rect 42064 6122 42116 6128
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 43364 5137 43392 20590
rect 43444 20596 43496 20602
rect 43444 20538 43496 20544
rect 43548 18970 43576 21286
rect 43640 20262 43668 21490
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43536 18964 43588 18970
rect 43536 18906 43588 18912
rect 43640 6254 43668 20198
rect 43628 6248 43680 6254
rect 43628 6190 43680 6196
rect 43350 5128 43406 5137
rect 43350 5063 43406 5072
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 41420 4820 41472 4826
rect 41420 4762 41472 4768
rect 41432 800 41460 4762
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 43824 2417 43852 24006
rect 43916 22778 43944 24142
rect 43904 22772 43956 22778
rect 43904 22714 43956 22720
rect 43996 22568 44048 22574
rect 43996 22510 44048 22516
rect 44008 21554 44036 22510
rect 44100 22114 44128 26200
rect 44364 25288 44416 25294
rect 44364 25230 44416 25236
rect 44180 23520 44232 23526
rect 44180 23462 44232 23468
rect 44192 23118 44220 23462
rect 44376 23322 44404 25230
rect 44916 24336 44968 24342
rect 44916 24278 44968 24284
rect 44456 24200 44508 24206
rect 44456 24142 44508 24148
rect 44822 24168 44878 24177
rect 44364 23316 44416 23322
rect 44364 23258 44416 23264
rect 44180 23112 44232 23118
rect 44180 23054 44232 23060
rect 44364 22500 44416 22506
rect 44364 22442 44416 22448
rect 44100 22086 44220 22114
rect 44192 21962 44220 22086
rect 44376 22030 44404 22442
rect 44364 22024 44416 22030
rect 44364 21966 44416 21972
rect 44180 21956 44232 21962
rect 44180 21898 44232 21904
rect 44088 21684 44140 21690
rect 44088 21626 44140 21632
rect 44100 21593 44128 21626
rect 44086 21584 44142 21593
rect 43996 21548 44048 21554
rect 44086 21519 44142 21528
rect 43996 21490 44048 21496
rect 44008 21162 44036 21490
rect 44468 21486 44496 24142
rect 44822 24103 44878 24112
rect 44548 24064 44600 24070
rect 44548 24006 44600 24012
rect 44560 23186 44588 24006
rect 44836 23730 44864 24103
rect 44824 23724 44876 23730
rect 44824 23666 44876 23672
rect 44928 23662 44956 24278
rect 44916 23656 44968 23662
rect 44916 23598 44968 23604
rect 44548 23180 44600 23186
rect 44548 23122 44600 23128
rect 44640 23112 44692 23118
rect 44640 23054 44692 23060
rect 44652 22710 44680 23054
rect 44640 22704 44692 22710
rect 44640 22646 44692 22652
rect 45112 22642 45140 26302
rect 45374 26200 45430 27000
rect 45928 26376 45980 26382
rect 45928 26318 45980 26324
rect 45388 22710 45416 26200
rect 45940 24410 45968 26318
rect 46018 26200 46074 27000
rect 46662 26200 46718 27000
rect 47306 26200 47362 27000
rect 47950 26200 48006 27000
rect 48594 26200 48650 27000
rect 45928 24404 45980 24410
rect 45928 24346 45980 24352
rect 45940 23662 45968 24346
rect 45928 23656 45980 23662
rect 45928 23598 45980 23604
rect 45836 22976 45888 22982
rect 45836 22918 45888 22924
rect 45376 22704 45428 22710
rect 45376 22646 45428 22652
rect 44916 22636 44968 22642
rect 44916 22578 44968 22584
rect 45008 22636 45060 22642
rect 45008 22578 45060 22584
rect 45100 22636 45152 22642
rect 45100 22578 45152 22584
rect 44824 22500 44876 22506
rect 44824 22442 44876 22448
rect 44548 22432 44600 22438
rect 44548 22374 44600 22380
rect 44456 21480 44508 21486
rect 44456 21422 44508 21428
rect 44008 21146 44128 21162
rect 44008 21140 44140 21146
rect 44008 21134 44088 21140
rect 44088 21082 44140 21088
rect 43904 20868 43956 20874
rect 43904 20810 43956 20816
rect 43916 16561 43944 20810
rect 44560 20534 44588 22374
rect 44732 21344 44784 21350
rect 44732 21286 44784 21292
rect 44548 20528 44600 20534
rect 44548 20470 44600 20476
rect 44744 19825 44772 21286
rect 44730 19816 44786 19825
rect 44730 19751 44786 19760
rect 43902 16552 43958 16561
rect 43902 16487 43958 16496
rect 44836 14890 44864 22442
rect 44928 21690 44956 22578
rect 45020 22166 45048 22578
rect 45652 22568 45704 22574
rect 45652 22510 45704 22516
rect 45192 22432 45244 22438
rect 45192 22374 45244 22380
rect 45008 22160 45060 22166
rect 45008 22102 45060 22108
rect 44916 21684 44968 21690
rect 44916 21626 44968 21632
rect 44824 14884 44876 14890
rect 44824 14826 44876 14832
rect 45204 9489 45232 22374
rect 45284 21956 45336 21962
rect 45284 21898 45336 21904
rect 45468 21956 45520 21962
rect 45468 21898 45520 21904
rect 45296 21690 45324 21898
rect 45376 21888 45428 21894
rect 45376 21830 45428 21836
rect 45284 21684 45336 21690
rect 45284 21626 45336 21632
rect 45388 17882 45416 21830
rect 45480 19242 45508 21898
rect 45664 21690 45692 22510
rect 45848 22098 45876 22918
rect 46032 22166 46060 26200
rect 46202 24848 46258 24857
rect 46202 24783 46258 24792
rect 46112 23248 46164 23254
rect 46110 23216 46112 23225
rect 46164 23216 46166 23225
rect 46110 23151 46166 23160
rect 46020 22160 46072 22166
rect 46020 22102 46072 22108
rect 45836 22092 45888 22098
rect 45836 22034 45888 22040
rect 45652 21684 45704 21690
rect 45652 21626 45704 21632
rect 45468 19236 45520 19242
rect 45468 19178 45520 19184
rect 45376 17876 45428 17882
rect 45376 17818 45428 17824
rect 46216 14346 46244 24783
rect 46386 23760 46442 23769
rect 46386 23695 46442 23704
rect 46400 14521 46428 23695
rect 46676 23322 46704 26200
rect 47320 23798 47348 26200
rect 47964 24154 47992 26200
rect 47872 24126 47992 24154
rect 48412 24200 48464 24206
rect 48412 24142 48464 24148
rect 47308 23792 47360 23798
rect 47308 23734 47360 23740
rect 47032 23724 47084 23730
rect 47032 23666 47084 23672
rect 46940 23588 46992 23594
rect 46940 23530 46992 23536
rect 46664 23316 46716 23322
rect 46664 23258 46716 23264
rect 46952 22710 46980 23530
rect 46940 22704 46992 22710
rect 46754 22672 46810 22681
rect 46480 22636 46532 22642
rect 46940 22646 46992 22652
rect 46754 22607 46810 22616
rect 46480 22578 46532 22584
rect 46492 22234 46520 22578
rect 46664 22432 46716 22438
rect 46664 22374 46716 22380
rect 46480 22228 46532 22234
rect 46480 22170 46532 22176
rect 46570 21992 46626 22001
rect 46570 21927 46626 21936
rect 46386 14512 46442 14521
rect 46386 14447 46442 14456
rect 46584 14385 46612 21927
rect 46676 19922 46704 22374
rect 46768 19990 46796 22607
rect 46940 22432 46992 22438
rect 46940 22374 46992 22380
rect 46952 20754 46980 22374
rect 47044 21690 47072 23666
rect 47216 22976 47268 22982
rect 47216 22918 47268 22924
rect 47032 21684 47084 21690
rect 47032 21626 47084 21632
rect 47228 21554 47256 22918
rect 47320 22710 47348 23734
rect 47308 22704 47360 22710
rect 47308 22646 47360 22652
rect 47872 22030 47900 24126
rect 48320 24064 48372 24070
rect 48320 24006 48372 24012
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 48332 22642 48360 24006
rect 48424 23866 48452 24142
rect 48504 24064 48556 24070
rect 48504 24006 48556 24012
rect 48412 23860 48464 23866
rect 48412 23802 48464 23808
rect 48516 23254 48544 24006
rect 48504 23248 48556 23254
rect 48504 23190 48556 23196
rect 48504 23112 48556 23118
rect 48504 23054 48556 23060
rect 48320 22636 48372 22642
rect 48320 22578 48372 22584
rect 48516 22098 48544 23054
rect 48504 22092 48556 22098
rect 48504 22034 48556 22040
rect 47860 22024 47912 22030
rect 47780 21972 47860 21978
rect 47780 21966 47912 21972
rect 47780 21950 47900 21966
rect 47400 21888 47452 21894
rect 47400 21830 47452 21836
rect 47216 21548 47268 21554
rect 47216 21490 47268 21496
rect 46860 20726 46980 20754
rect 46756 19984 46808 19990
rect 46756 19926 46808 19932
rect 46664 19916 46716 19922
rect 46664 19858 46716 19864
rect 46860 18154 46888 20726
rect 46848 18148 46900 18154
rect 46848 18090 46900 18096
rect 47412 17270 47440 21830
rect 47780 21690 47808 21950
rect 47860 21888 47912 21894
rect 47860 21830 47912 21836
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47768 21548 47820 21554
rect 47768 21490 47820 21496
rect 47780 20806 47808 21490
rect 47768 20800 47820 20806
rect 47768 20742 47820 20748
rect 47400 17264 47452 17270
rect 47400 17206 47452 17212
rect 46570 14376 46626 14385
rect 46204 14340 46256 14346
rect 46570 14311 46626 14320
rect 46204 14282 46256 14288
rect 47780 11082 47808 20742
rect 47872 14278 47900 21830
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 48608 21146 48636 26200
rect 49240 24200 49292 24206
rect 49240 24142 49292 24148
rect 48964 24064 49016 24070
rect 48964 24006 49016 24012
rect 48872 23724 48924 23730
rect 48872 23666 48924 23672
rect 48884 23322 48912 23666
rect 48872 23316 48924 23322
rect 48872 23258 48924 23264
rect 48688 22432 48740 22438
rect 48688 22374 48740 22380
rect 48700 22030 48728 22374
rect 48688 22024 48740 22030
rect 48688 21966 48740 21972
rect 48596 21140 48648 21146
rect 48596 21082 48648 21088
rect 48608 20942 48636 21082
rect 48596 20936 48648 20942
rect 48596 20878 48648 20884
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 48884 20602 48912 23258
rect 48872 20596 48924 20602
rect 48872 20538 48924 20544
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47860 14272 47912 14278
rect 47860 14214 47912 14220
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47768 11076 47820 11082
rect 47768 11018 47820 11024
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 48976 10033 49004 24006
rect 49056 23520 49108 23526
rect 49056 23462 49108 23468
rect 48962 10024 49018 10033
rect 48962 9959 49018 9968
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 45190 9480 45246 9489
rect 45190 9415 45246 9424
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 49068 8022 49096 23462
rect 49252 22545 49280 24142
rect 49332 24132 49384 24138
rect 49332 24074 49384 24080
rect 49344 23322 49372 24074
rect 49332 23316 49384 23322
rect 49332 23258 49384 23264
rect 49332 23112 49384 23118
rect 49332 23054 49384 23060
rect 49238 22536 49294 22545
rect 49238 22471 49294 22480
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21049 49188 21422
rect 49146 21040 49202 21049
rect 49146 20975 49202 20984
rect 49252 20534 49280 22471
rect 49344 21146 49372 23054
rect 49332 21140 49384 21146
rect 49332 21082 49384 21088
rect 49240 20528 49292 20534
rect 49240 20470 49292 20476
rect 49056 8016 49108 8022
rect 49056 7958 49108 7964
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 49424 5024 49476 5030
rect 49424 4966 49476 4972
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 44088 3528 44140 3534
rect 44088 3470 44140 3476
rect 43810 2408 43866 2417
rect 43810 2343 43866 2352
rect 44100 800 44128 3470
rect 46756 3460 46808 3466
rect 46756 3402 46808 3408
rect 46768 800 46796 3402
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 49436 800 49464 4966
rect 34980 740 35032 746
rect 34980 682 35032 688
rect 36082 0 36138 800
rect 38750 0 38806 800
rect 41418 0 41474 800
rect 44086 0 44142 800
rect 46754 0 46810 800
rect 49422 0 49478 800
<< via2 >>
rect 938 9424 994 9480
rect 1490 20304 1546 20360
rect 1398 19080 1454 19136
rect 1490 18672 1546 18728
rect 1674 20848 1730 20904
rect 1398 17856 1454 17912
rect 1214 17040 1270 17096
rect 1306 16632 1362 16688
rect 1306 16224 1362 16280
rect 1122 13368 1178 13424
rect 1306 15816 1362 15872
rect 1306 15408 1362 15464
rect 1306 15000 1362 15056
rect 1306 14592 1362 14648
rect 1306 14184 1362 14240
rect 1582 13932 1638 13968
rect 1582 13912 1584 13932
rect 1584 13912 1636 13932
rect 1636 13912 1638 13932
rect 1398 12144 1454 12200
rect 1582 13268 1584 13288
rect 1584 13268 1636 13288
rect 1636 13268 1638 13288
rect 1582 13232 1638 13268
rect 2042 19488 2098 19544
rect 2226 24248 2282 24304
rect 2226 21120 2282 21176
rect 2042 18264 2098 18320
rect 2042 17448 2098 17504
rect 2042 13776 2098 13832
rect 1766 11056 1822 11112
rect 1766 10784 1822 10840
rect 1398 9288 1454 9344
rect 1214 7520 1270 7576
rect 1306 6024 1362 6080
rect 1306 5652 1308 5672
rect 1308 5652 1360 5672
rect 1360 5652 1362 5672
rect 1306 5616 1362 5652
rect 1306 5208 1362 5264
rect 1674 9560 1730 9616
rect 1582 8744 1638 8800
rect 1950 10784 2006 10840
rect 1950 10512 2006 10568
rect 1950 9832 2006 9888
rect 1490 8200 1546 8256
rect 1490 4800 1546 4856
rect 1766 6704 1822 6760
rect 1306 2388 1308 2408
rect 1308 2388 1360 2408
rect 1360 2388 1362 2408
rect 1306 2352 1362 2388
rect 938 1808 994 1864
rect 1582 2760 1638 2816
rect 2778 24384 2834 24440
rect 3330 25200 3386 25256
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 3330 22480 3386 22536
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 3330 21936 3386 21992
rect 2686 21528 2742 21584
rect 3330 21256 3386 21312
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 2778 19896 2834 19952
rect 2594 19760 2650 19816
rect 2318 10104 2374 10160
rect 2318 8084 2374 8120
rect 2318 8064 2320 8084
rect 2320 8064 2372 8084
rect 2372 8064 2374 8084
rect 2134 6740 2136 6760
rect 2136 6740 2188 6760
rect 2188 6740 2190 6760
rect 2134 6704 2190 6740
rect 2410 7928 2466 7984
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 3698 23976 3754 24032
rect 3606 23196 3608 23216
rect 3608 23196 3660 23216
rect 3660 23196 3662 23216
rect 3606 23160 3662 23196
rect 3606 22072 3662 22128
rect 4066 25608 4122 25664
rect 3974 24792 4030 24848
rect 4802 25064 4858 25120
rect 4066 23568 4122 23624
rect 3882 23024 3938 23080
rect 3790 22752 3846 22808
rect 3790 20712 3846 20768
rect 3606 18264 3662 18320
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 3606 17740 3662 17776
rect 3606 17720 3608 17740
rect 3608 17720 3660 17740
rect 3660 17720 3662 17740
rect 3422 16668 3424 16688
rect 3424 16668 3476 16688
rect 3476 16668 3478 16688
rect 3422 16632 3478 16668
rect 3422 15428 3478 15464
rect 3422 15408 3424 15428
rect 3424 15408 3476 15428
rect 3476 15408 3478 15428
rect 3606 15580 3608 15600
rect 3608 15580 3660 15600
rect 3660 15580 3662 15600
rect 3606 15544 3662 15580
rect 3974 21528 4030 21584
rect 4066 20984 4122 21040
rect 3974 20168 4030 20224
rect 4066 18128 4122 18184
rect 4710 23432 4766 23488
rect 4342 17620 4344 17640
rect 4344 17620 4396 17640
rect 4396 17620 4398 17640
rect 4342 17584 4398 17620
rect 3882 16904 3938 16960
rect 3698 15136 3754 15192
rect 3606 14220 3608 14240
rect 3608 14220 3660 14240
rect 3660 14220 3662 14240
rect 3606 14184 3662 14220
rect 3514 13812 3516 13832
rect 3516 13812 3568 13832
rect 3568 13812 3570 13832
rect 3514 13776 3570 13812
rect 2870 13096 2926 13152
rect 2870 12960 2926 13016
rect 3238 12960 3294 13016
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 3330 12280 3386 12336
rect 3238 11736 3294 11792
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 2962 10784 3018 10840
rect 3054 10512 3110 10568
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 3146 10104 3202 10160
rect 2962 9424 3018 9480
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 2962 8336 3018 8392
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 2594 5480 2650 5536
rect 3238 6432 3294 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 3514 13232 3570 13288
rect 3974 15000 4030 15056
rect 3882 14864 3938 14920
rect 3790 13640 3846 13696
rect 3790 13368 3846 13424
rect 3698 12008 3754 12064
rect 3882 12416 3938 12472
rect 3514 7656 3570 7712
rect 3514 6568 3570 6624
rect 2962 5208 3018 5264
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 2686 4664 2742 4720
rect 3146 4664 3202 4720
rect 2962 4564 2964 4584
rect 2964 4564 3016 4584
rect 3016 4564 3018 4584
rect 2962 4528 3018 4564
rect 1858 1400 1914 1456
rect 2778 2488 2834 2544
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 3054 3440 3110 3496
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 3330 2624 3386 2680
rect 3790 11192 3846 11248
rect 3790 9560 3846 9616
rect 3790 6024 3846 6080
rect 4250 14728 4306 14784
rect 4250 13524 4306 13560
rect 4250 13504 4252 13524
rect 4252 13504 4304 13524
rect 4304 13504 4306 13524
rect 4894 19080 4950 19136
rect 5538 22616 5594 22672
rect 6182 25472 6238 25528
rect 5814 21528 5870 21584
rect 5630 20712 5686 20768
rect 5538 20440 5594 20496
rect 5906 20304 5962 20360
rect 6090 18536 6146 18592
rect 5538 15136 5594 15192
rect 4710 14048 4766 14104
rect 4066 10376 4122 10432
rect 4342 9968 4398 10024
rect 4250 9580 4306 9616
rect 4250 9560 4252 9580
rect 4252 9560 4304 9580
rect 4304 9560 4306 9580
rect 4250 8472 4306 8528
rect 4526 8064 4582 8120
rect 4802 11056 4858 11112
rect 4986 14068 5042 14104
rect 4986 14048 4988 14068
rect 4988 14048 5040 14068
rect 5040 14048 5042 14068
rect 5078 12824 5134 12880
rect 5078 12552 5134 12608
rect 5078 12280 5134 12336
rect 4986 12144 5042 12200
rect 5170 11872 5226 11928
rect 5078 9444 5134 9480
rect 5078 9424 5080 9444
rect 5080 9424 5132 9444
rect 5132 9424 5134 9444
rect 4986 8200 5042 8256
rect 4802 7928 4858 7984
rect 4434 6976 4490 7032
rect 4158 6296 4214 6352
rect 3698 4392 3754 4448
rect 3606 3576 3662 3632
rect 3514 1944 3570 2000
rect 3422 1536 3478 1592
rect 3790 3984 3846 4040
rect 3882 856 3938 912
rect 4618 6296 4674 6352
rect 4066 3168 4122 3224
rect 5078 7928 5134 7984
rect 5354 7384 5410 7440
rect 5630 9596 5632 9616
rect 5632 9596 5684 9616
rect 5684 9596 5686 9616
rect 5630 9560 5686 9596
rect 6918 21120 6974 21176
rect 6550 20712 6606 20768
rect 6458 20576 6514 20632
rect 5998 16088 6054 16144
rect 6826 19624 6882 19680
rect 6458 17040 6514 17096
rect 5998 12416 6054 12472
rect 5998 11872 6054 11928
rect 5814 8336 5870 8392
rect 5722 6296 5778 6352
rect 5170 5344 5226 5400
rect 5538 6160 5594 6216
rect 5446 5908 5502 5944
rect 5446 5888 5448 5908
rect 5448 5888 5500 5908
rect 5500 5888 5502 5908
rect 5354 4140 5410 4176
rect 5354 4120 5356 4140
rect 5356 4120 5408 4140
rect 5408 4120 5410 4140
rect 5262 3032 5318 3088
rect 5538 4664 5594 4720
rect 6366 12416 6422 12472
rect 6274 12280 6330 12336
rect 6274 11872 6330 11928
rect 6090 6024 6146 6080
rect 6090 5616 6146 5672
rect 6642 16108 6698 16144
rect 6642 16088 6644 16108
rect 6644 16088 6696 16108
rect 6696 16088 6698 16108
rect 6826 17992 6882 18048
rect 6918 16768 6974 16824
rect 7562 19624 7618 19680
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 8022 20848 8078 20904
rect 7194 17584 7250 17640
rect 6642 14320 6698 14376
rect 6550 14048 6606 14104
rect 6734 12960 6790 13016
rect 7010 15000 7066 15056
rect 7470 17720 7526 17776
rect 7378 15000 7434 15056
rect 7102 14728 7158 14784
rect 6550 12844 6606 12880
rect 6550 12824 6552 12844
rect 6552 12824 6604 12844
rect 6604 12824 6606 12844
rect 6642 12552 6698 12608
rect 6734 12008 6790 12064
rect 6550 10784 6606 10840
rect 6734 10240 6790 10296
rect 6642 9560 6698 9616
rect 6550 9288 6606 9344
rect 6826 9460 6828 9480
rect 6828 9460 6880 9480
rect 6880 9460 6882 9480
rect 6826 9424 6882 9460
rect 6642 9152 6698 9208
rect 6642 8336 6698 8392
rect 6366 6060 6368 6080
rect 6368 6060 6420 6080
rect 6420 6060 6422 6080
rect 6366 6024 6422 6060
rect 5814 3576 5870 3632
rect 5814 2352 5870 2408
rect 5446 720 5502 776
rect 6274 5072 6330 5128
rect 5998 3848 6054 3904
rect 6090 1264 6146 1320
rect 6550 5480 6606 5536
rect 6458 4800 6514 4856
rect 6550 3984 6606 4040
rect 6826 7656 6882 7712
rect 6734 7148 6736 7168
rect 6736 7148 6788 7168
rect 6788 7148 6790 7168
rect 6734 7112 6790 7148
rect 6734 6704 6790 6760
rect 7286 14320 7342 14376
rect 7286 14184 7342 14240
rect 7194 13232 7250 13288
rect 7654 16632 7710 16688
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 8482 23432 8538 23488
rect 8390 19896 8446 19952
rect 8022 18692 8078 18728
rect 8022 18672 8024 18692
rect 8024 18672 8076 18692
rect 8076 18672 8078 18692
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 8114 18128 8170 18184
rect 7838 17856 7894 17912
rect 8298 17856 8354 17912
rect 8206 17720 8262 17776
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 8206 17076 8208 17096
rect 8208 17076 8260 17096
rect 8260 17076 8262 17096
rect 8206 17040 8262 17076
rect 8022 16768 8078 16824
rect 7838 16632 7894 16688
rect 8114 16496 8170 16552
rect 8298 16496 8354 16552
rect 7654 15680 7710 15736
rect 7654 15564 7710 15600
rect 7654 15544 7656 15564
rect 7656 15544 7708 15564
rect 7708 15544 7710 15564
rect 7654 15156 7710 15192
rect 7654 15136 7656 15156
rect 7656 15136 7708 15156
rect 7708 15136 7710 15156
rect 7562 14048 7618 14104
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7930 15544 7986 15600
rect 7930 15428 7986 15464
rect 7930 15408 7932 15428
rect 7932 15408 7984 15428
rect 7984 15408 7986 15428
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 8022 14884 8078 14920
rect 8022 14864 8024 14884
rect 8024 14864 8076 14884
rect 8076 14864 8078 14884
rect 7654 13912 7710 13968
rect 7470 13776 7526 13832
rect 7930 14340 7986 14376
rect 7930 14320 7932 14340
rect 7932 14320 7984 14340
rect 7984 14320 7986 14340
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 7378 13504 7434 13560
rect 7378 13096 7434 13152
rect 7286 12960 7342 13016
rect 7102 10920 7158 10976
rect 7102 9560 7158 9616
rect 7470 12180 7472 12200
rect 7472 12180 7524 12200
rect 7524 12180 7526 12200
rect 7470 12144 7526 12180
rect 7378 9868 7380 9888
rect 7380 9868 7432 9888
rect 7432 9868 7434 9888
rect 7378 9832 7434 9868
rect 7838 13640 7894 13696
rect 8758 21836 8760 21856
rect 8760 21836 8812 21856
rect 8812 21836 8814 21856
rect 8758 21800 8814 21836
rect 9034 22208 9090 22264
rect 9034 21956 9090 21992
rect 9034 21936 9036 21956
rect 9036 21936 9088 21956
rect 9088 21936 9090 21956
rect 9034 20576 9090 20632
rect 9862 25200 9918 25256
rect 9678 23704 9734 23760
rect 9770 23432 9826 23488
rect 9310 21664 9366 21720
rect 9770 22072 9826 22128
rect 9586 21412 9642 21448
rect 9586 21392 9588 21412
rect 9588 21392 9640 21412
rect 9640 21392 9642 21412
rect 9678 20712 9734 20768
rect 8574 18128 8630 18184
rect 8942 19116 8944 19136
rect 8944 19116 8996 19136
rect 8996 19116 8998 19136
rect 8942 19080 8998 19116
rect 8574 16768 8630 16824
rect 8850 17176 8906 17232
rect 8574 16360 8630 16416
rect 8666 16244 8722 16280
rect 8666 16224 8668 16244
rect 8668 16224 8720 16244
rect 8720 16224 8722 16244
rect 8758 15952 8814 16008
rect 8574 15136 8630 15192
rect 8482 14356 8484 14376
rect 8484 14356 8536 14376
rect 8536 14356 8538 14376
rect 8482 14320 8538 14356
rect 8482 14048 8538 14104
rect 8206 13368 8262 13424
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 8206 12552 8262 12608
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 7562 9424 7618 9480
rect 7378 7792 7434 7848
rect 7286 7656 7342 7712
rect 7930 11056 7986 11112
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 8574 11328 8630 11384
rect 8298 10648 8354 10704
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 8574 10784 8630 10840
rect 8390 10376 8446 10432
rect 8390 9152 8446 9208
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 7746 6568 7802 6624
rect 7746 6432 7802 6488
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7930 6296 7986 6352
rect 8390 6432 8446 6488
rect 7838 5752 7894 5808
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7746 5364 7802 5400
rect 7746 5344 7748 5364
rect 7748 5344 7800 5364
rect 7800 5344 7802 5364
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 9218 17992 9274 18048
rect 9034 15680 9090 15736
rect 9034 14320 9090 14376
rect 8942 13912 8998 13968
rect 8942 13368 8998 13424
rect 8850 10376 8906 10432
rect 8850 9596 8852 9616
rect 8852 9596 8904 9616
rect 8904 9596 8906 9616
rect 8850 9560 8906 9596
rect 8850 8744 8906 8800
rect 9494 19352 9550 19408
rect 9494 18536 9550 18592
rect 9678 19216 9734 19272
rect 9862 18400 9918 18456
rect 9770 17992 9826 18048
rect 9402 17720 9458 17776
rect 9310 17176 9366 17232
rect 9218 16632 9274 16688
rect 9586 16632 9642 16688
rect 9954 16652 10010 16688
rect 9954 16632 9956 16652
rect 9956 16632 10008 16652
rect 10008 16632 10010 16652
rect 9402 16224 9458 16280
rect 9402 15136 9458 15192
rect 9494 13368 9550 13424
rect 9862 15136 9918 15192
rect 9678 13912 9734 13968
rect 9586 12960 9642 13016
rect 9770 13368 9826 13424
rect 9770 13096 9826 13152
rect 9954 14320 10010 14376
rect 11058 24828 11060 24848
rect 11060 24828 11112 24848
rect 11112 24828 11114 24848
rect 11058 24792 11114 24828
rect 10874 23976 10930 24032
rect 10598 23840 10654 23896
rect 10506 22072 10562 22128
rect 10322 19780 10378 19816
rect 10322 19760 10324 19780
rect 10324 19760 10376 19780
rect 10376 19760 10378 19780
rect 10690 23568 10746 23624
rect 11426 22616 11482 22672
rect 10782 19252 10784 19272
rect 10784 19252 10836 19272
rect 10836 19252 10838 19272
rect 10782 19216 10838 19252
rect 10782 18944 10838 19000
rect 10598 18692 10654 18728
rect 10598 18672 10600 18692
rect 10600 18672 10652 18692
rect 10652 18672 10654 18692
rect 11334 21664 11390 21720
rect 11334 20748 11336 20768
rect 11336 20748 11388 20768
rect 11388 20748 11390 20768
rect 10690 18284 10746 18320
rect 10690 18264 10692 18284
rect 10692 18264 10744 18284
rect 10744 18264 10746 18284
rect 10506 17448 10562 17504
rect 10322 16940 10324 16960
rect 10324 16940 10376 16960
rect 10376 16940 10378 16960
rect 10322 16904 10378 16940
rect 10322 15952 10378 16008
rect 10230 15680 10286 15736
rect 10690 16224 10746 16280
rect 10506 15136 10562 15192
rect 9586 12280 9642 12336
rect 9034 9968 9090 10024
rect 9126 8744 9182 8800
rect 9034 8472 9090 8528
rect 9126 8200 9182 8256
rect 9034 6740 9036 6760
rect 9036 6740 9088 6760
rect 9088 6740 9090 6760
rect 9034 6704 9090 6740
rect 8850 6160 8906 6216
rect 9034 6160 9090 6216
rect 9862 12008 9918 12064
rect 9402 9968 9458 10024
rect 9862 10920 9918 10976
rect 10046 10920 10102 10976
rect 9770 9968 9826 10024
rect 9678 8608 9734 8664
rect 9678 6296 9734 6352
rect 9954 10240 10010 10296
rect 9862 8608 9918 8664
rect 9862 8472 9918 8528
rect 9034 4528 9090 4584
rect 8574 3460 8630 3496
rect 8574 3440 8576 3460
rect 8576 3440 8628 3460
rect 8628 3440 8630 3460
rect 8758 2896 8814 2952
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 9402 4800 9458 4856
rect 9678 4392 9734 4448
rect 9310 4020 9312 4040
rect 9312 4020 9364 4040
rect 9364 4020 9366 4040
rect 9310 3984 9366 4020
rect 10230 9152 10286 9208
rect 10046 8608 10102 8664
rect 10046 8372 10048 8392
rect 10048 8372 10100 8392
rect 10100 8372 10102 8392
rect 10046 8336 10102 8372
rect 10046 7112 10102 7168
rect 9954 5072 10010 5128
rect 10414 10512 10470 10568
rect 10414 9696 10470 9752
rect 10414 9560 10470 9616
rect 10690 14592 10746 14648
rect 11058 16652 11114 16688
rect 11058 16632 11060 16652
rect 11060 16632 11112 16652
rect 11112 16632 11114 16652
rect 11058 16124 11060 16144
rect 11060 16124 11112 16144
rect 11112 16124 11114 16144
rect 11058 16088 11114 16124
rect 10966 14728 11022 14784
rect 10874 14320 10930 14376
rect 11150 15408 11206 15464
rect 11058 14048 11114 14104
rect 11334 20712 11390 20748
rect 11334 18264 11390 18320
rect 11334 17720 11390 17776
rect 11702 23432 11758 23488
rect 11978 25336 12034 25392
rect 11794 23024 11850 23080
rect 11978 22888 12034 22944
rect 11794 20460 11850 20496
rect 11794 20440 11796 20460
rect 11796 20440 11848 20460
rect 11848 20440 11850 20460
rect 11610 19488 11666 19544
rect 11610 18300 11612 18320
rect 11612 18300 11664 18320
rect 11664 18300 11666 18320
rect 11610 18264 11666 18300
rect 11518 17604 11574 17640
rect 11518 17584 11520 17604
rect 11520 17584 11572 17604
rect 11572 17584 11574 17604
rect 11426 16244 11482 16280
rect 11426 16224 11428 16244
rect 11428 16224 11480 16244
rect 11480 16224 11482 16244
rect 11518 16088 11574 16144
rect 11242 14864 11298 14920
rect 10782 13096 10838 13152
rect 10598 11192 10654 11248
rect 10598 9968 10654 10024
rect 11150 13504 11206 13560
rect 10966 11328 11022 11384
rect 11426 15272 11482 15328
rect 11426 13640 11482 13696
rect 11242 12280 11298 12336
rect 11242 11756 11298 11792
rect 11242 11736 11244 11756
rect 11244 11736 11296 11756
rect 11296 11736 11298 11756
rect 11242 11328 11298 11384
rect 11150 10512 11206 10568
rect 11242 10260 11298 10296
rect 12254 24656 12310 24712
rect 12530 24148 12532 24168
rect 12532 24148 12584 24168
rect 12584 24148 12586 24168
rect 12530 24112 12586 24148
rect 11794 17312 11850 17368
rect 11794 14764 11796 14784
rect 11796 14764 11848 14784
rect 11848 14764 11850 14784
rect 11794 14728 11850 14764
rect 11702 14592 11758 14648
rect 11978 15272 12034 15328
rect 11886 14320 11942 14376
rect 11886 13368 11942 13424
rect 11702 12860 11704 12880
rect 11704 12860 11756 12880
rect 11756 12860 11758 12880
rect 11702 12824 11758 12860
rect 11426 12008 11482 12064
rect 11426 11736 11482 11792
rect 11518 11464 11574 11520
rect 11518 11192 11574 11248
rect 11242 10240 11244 10260
rect 11244 10240 11296 10260
rect 11296 10240 11298 10260
rect 10782 8880 10838 8936
rect 10782 8336 10838 8392
rect 10230 6704 10286 6760
rect 10230 6604 10232 6624
rect 10232 6604 10284 6624
rect 10284 6604 10286 6624
rect 10230 6568 10286 6604
rect 10230 5908 10286 5944
rect 10230 5888 10232 5908
rect 10232 5888 10284 5908
rect 10284 5888 10286 5908
rect 9494 2624 9550 2680
rect 9126 856 9182 912
rect 10598 8200 10654 8256
rect 11150 9696 11206 9752
rect 10966 8472 11022 8528
rect 11150 8744 11206 8800
rect 11334 9152 11390 9208
rect 11242 8472 11298 8528
rect 11150 7656 11206 7712
rect 11334 7792 11390 7848
rect 11242 7520 11298 7576
rect 10874 6704 10930 6760
rect 10782 6432 10838 6488
rect 11058 5480 11114 5536
rect 10966 5072 11022 5128
rect 11150 4020 11152 4040
rect 11152 4020 11204 4040
rect 11204 4020 11206 4040
rect 11150 3984 11206 4020
rect 10874 3168 10930 3224
rect 11334 6160 11390 6216
rect 11334 5616 11390 5672
rect 11518 9152 11574 9208
rect 11518 8880 11574 8936
rect 11794 12552 11850 12608
rect 11702 10512 11758 10568
rect 11702 9288 11758 9344
rect 11610 5908 11666 5944
rect 11610 5888 11612 5908
rect 11612 5888 11664 5908
rect 11664 5888 11666 5908
rect 11702 5616 11758 5672
rect 12254 21428 12256 21448
rect 12256 21428 12308 21448
rect 12308 21428 12310 21448
rect 12254 21392 12310 21428
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 13358 23296 13414 23352
rect 12530 22752 12586 22808
rect 12438 22344 12494 22400
rect 12530 21256 12586 21312
rect 12714 22208 12770 22264
rect 12898 22752 12954 22808
rect 12898 22480 12954 22536
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12990 20340 12992 20360
rect 12992 20340 13044 20360
rect 13044 20340 13046 20360
rect 12990 20304 13046 20340
rect 12714 20168 12770 20224
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12714 19760 12770 19816
rect 12622 19216 12678 19272
rect 12714 18808 12770 18864
rect 12530 17856 12586 17912
rect 12530 16360 12586 16416
rect 12530 15544 12586 15600
rect 12346 15136 12402 15192
rect 12530 15136 12586 15192
rect 12530 13912 12586 13968
rect 13174 19216 13230 19272
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 13542 24248 13598 24304
rect 13910 24248 13966 24304
rect 14278 24112 14334 24168
rect 14094 22888 14150 22944
rect 13726 22072 13782 22128
rect 13818 20304 13874 20360
rect 14002 20168 14058 20224
rect 13726 19896 13782 19952
rect 13818 19796 13820 19816
rect 13820 19796 13872 19816
rect 13872 19796 13874 19816
rect 13818 19760 13874 19796
rect 13358 18400 13414 18456
rect 13358 17992 13414 18048
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 13358 16532 13360 16552
rect 13360 16532 13412 16552
rect 13412 16532 13414 16552
rect 12898 16124 12900 16144
rect 12900 16124 12952 16144
rect 12952 16124 12954 16144
rect 12898 16088 12954 16124
rect 13358 16496 13414 16532
rect 13358 16108 13414 16144
rect 13358 16088 13360 16108
rect 13360 16088 13412 16108
rect 13412 16088 13414 16108
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12806 14592 12862 14648
rect 12438 11892 12494 11928
rect 12438 11872 12440 11892
rect 12440 11872 12492 11892
rect 12492 11872 12494 11892
rect 11978 10104 12034 10160
rect 12162 10240 12218 10296
rect 12070 9968 12126 10024
rect 11886 9596 11888 9616
rect 11888 9596 11940 9616
rect 11940 9596 11942 9616
rect 11886 9560 11942 9596
rect 11978 9016 12034 9072
rect 11702 5208 11758 5264
rect 12346 9696 12402 9752
rect 12162 8064 12218 8120
rect 12162 7656 12218 7712
rect 12530 9560 12586 9616
rect 12438 9424 12494 9480
rect 12162 7248 12218 7304
rect 12162 7112 12218 7168
rect 12070 6740 12072 6760
rect 12072 6740 12124 6760
rect 12124 6740 12126 6760
rect 12070 6704 12126 6740
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 13174 12708 13230 12744
rect 13174 12688 13176 12708
rect 13176 12688 13228 12708
rect 13228 12688 13230 12708
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 13266 11056 13322 11112
rect 12806 10376 12862 10432
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 13910 18672 13966 18728
rect 14370 23160 14426 23216
rect 14370 22888 14426 22944
rect 14646 23160 14702 23216
rect 14278 22480 14334 22536
rect 14370 20440 14426 20496
rect 14278 19760 14334 19816
rect 14186 18128 14242 18184
rect 14462 18828 14518 18864
rect 14462 18808 14464 18828
rect 14464 18808 14516 18828
rect 14516 18808 14518 18828
rect 14370 17856 14426 17912
rect 15014 23976 15070 24032
rect 14922 23432 14978 23488
rect 14830 22380 14832 22400
rect 14832 22380 14884 22400
rect 14884 22380 14886 22400
rect 14830 22344 14886 22380
rect 14646 20032 14702 20088
rect 14646 19624 14702 19680
rect 14646 18672 14702 18728
rect 14278 17448 14334 17504
rect 14002 16904 14058 16960
rect 13726 16224 13782 16280
rect 13634 15036 13636 15056
rect 13636 15036 13688 15056
rect 13688 15036 13690 15056
rect 13634 15000 13690 15036
rect 14002 15680 14058 15736
rect 14646 17448 14702 17504
rect 14922 22072 14978 22128
rect 15658 24384 15714 24440
rect 15290 23704 15346 23760
rect 15474 23432 15530 23488
rect 14922 21936 14978 21992
rect 15198 21972 15200 21992
rect 15200 21972 15252 21992
rect 15252 21972 15254 21992
rect 15198 21936 15254 21972
rect 15566 22888 15622 22944
rect 15382 21800 15438 21856
rect 15106 21564 15108 21584
rect 15108 21564 15160 21584
rect 15160 21564 15162 21584
rect 15106 21528 15162 21564
rect 14830 20576 14886 20632
rect 14830 20168 14886 20224
rect 15106 20984 15162 21040
rect 15198 19896 15254 19952
rect 14830 17720 14886 17776
rect 14830 17448 14886 17504
rect 14738 17176 14794 17232
rect 14738 16632 14794 16688
rect 14094 15544 14150 15600
rect 13818 14728 13874 14784
rect 13726 14456 13782 14512
rect 13542 12008 13598 12064
rect 13542 11192 13598 11248
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 13266 8880 13322 8936
rect 12438 6704 12494 6760
rect 12438 4256 12494 4312
rect 10966 1808 11022 1864
rect 12714 6060 12716 6080
rect 12716 6060 12768 6080
rect 12768 6060 12770 6080
rect 12714 6024 12770 6060
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12898 7520 12954 7576
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12714 5752 12770 5808
rect 13542 8880 13598 8936
rect 13542 8472 13598 8528
rect 13450 6704 13506 6760
rect 14278 15408 14334 15464
rect 13910 12824 13966 12880
rect 13910 11872 13966 11928
rect 13818 11736 13874 11792
rect 13818 11212 13874 11248
rect 13818 11192 13820 11212
rect 13820 11192 13872 11212
rect 13872 11192 13874 11212
rect 13818 10956 13820 10976
rect 13820 10956 13872 10976
rect 13872 10956 13874 10976
rect 13818 10920 13874 10956
rect 13818 10784 13874 10840
rect 13818 10140 13820 10160
rect 13820 10140 13872 10160
rect 13872 10140 13874 10160
rect 13818 10104 13874 10140
rect 13818 9968 13874 10024
rect 13726 7248 13782 7304
rect 13634 6568 13690 6624
rect 13910 8064 13966 8120
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 13818 4528 13874 4584
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 13082 3168 13138 3224
rect 13358 3168 13414 3224
rect 13358 2796 13360 2816
rect 13360 2796 13412 2816
rect 13412 2796 13414 2816
rect 12438 2624 12494 2680
rect 13358 2760 13414 2796
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 13450 2624 13506 2680
rect 13726 1808 13782 1864
rect 14186 11464 14242 11520
rect 14094 9868 14096 9888
rect 14096 9868 14148 9888
rect 14148 9868 14150 9888
rect 14094 9832 14150 9868
rect 14186 9324 14188 9344
rect 14188 9324 14240 9344
rect 14240 9324 14242 9344
rect 14186 9288 14242 9324
rect 14094 8472 14150 8528
rect 14186 8336 14242 8392
rect 14094 6568 14150 6624
rect 14462 15972 14518 16008
rect 14462 15952 14464 15972
rect 14464 15952 14516 15972
rect 14516 15952 14518 15972
rect 14462 15680 14518 15736
rect 14370 11736 14426 11792
rect 14554 11736 14610 11792
rect 14554 10920 14610 10976
rect 14370 10648 14426 10704
rect 14278 7384 14334 7440
rect 14554 9968 14610 10024
rect 15290 19624 15346 19680
rect 15842 23296 15898 23352
rect 15934 21664 15990 21720
rect 16486 24792 16542 24848
rect 16394 23568 16450 23624
rect 15566 20304 15622 20360
rect 15106 17720 15162 17776
rect 15382 18164 15384 18184
rect 15384 18164 15436 18184
rect 15436 18164 15438 18184
rect 15382 18128 15438 18164
rect 15198 17312 15254 17368
rect 15382 16768 15438 16824
rect 14738 12552 14794 12608
rect 14922 11192 14978 11248
rect 14738 9596 14740 9616
rect 14740 9596 14792 9616
rect 14792 9596 14794 9616
rect 14738 9560 14794 9596
rect 14646 8492 14702 8528
rect 14646 8472 14648 8492
rect 14648 8472 14700 8492
rect 14700 8472 14702 8492
rect 14922 9152 14978 9208
rect 15658 19080 15714 19136
rect 16118 20440 16174 20496
rect 16302 21664 16358 21720
rect 16302 21292 16304 21312
rect 16304 21292 16356 21312
rect 16356 21292 16358 21312
rect 16302 21256 16358 21292
rect 16486 23432 16542 23488
rect 16670 23840 16726 23896
rect 16670 22208 16726 22264
rect 16578 21936 16634 21992
rect 17038 23840 17094 23896
rect 17038 23704 17094 23760
rect 16762 22108 16764 22128
rect 16764 22108 16816 22128
rect 16816 22108 16818 22128
rect 16762 22072 16818 22108
rect 16762 20848 16818 20904
rect 16578 20576 16634 20632
rect 16118 20168 16174 20224
rect 16302 19488 16358 19544
rect 15750 17992 15806 18048
rect 16118 18944 16174 19000
rect 16118 18536 16174 18592
rect 16026 18264 16082 18320
rect 16210 17992 16266 18048
rect 16486 20032 16542 20088
rect 16486 19352 16542 19408
rect 16394 18536 16450 18592
rect 15566 15816 15622 15872
rect 15474 14592 15530 14648
rect 15290 14320 15346 14376
rect 15290 11872 15346 11928
rect 15658 15428 15714 15464
rect 15658 15408 15660 15428
rect 15660 15408 15712 15428
rect 15712 15408 15714 15428
rect 15750 15000 15806 15056
rect 15474 12008 15530 12064
rect 14554 3712 14610 3768
rect 14186 1400 14242 1456
rect 13910 1128 13966 1184
rect 14830 3068 14832 3088
rect 14832 3068 14884 3088
rect 14884 3068 14886 3088
rect 14830 3032 14886 3068
rect 15842 13368 15898 13424
rect 16118 16632 16174 16688
rect 15842 11872 15898 11928
rect 16210 16496 16266 16552
rect 16854 20168 16910 20224
rect 16854 19624 16910 19680
rect 16946 19488 17002 19544
rect 17130 21392 17186 21448
rect 17130 21120 17186 21176
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17958 23024 18014 23080
rect 18602 24656 18658 24712
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 17406 21800 17462 21856
rect 17222 20848 17278 20904
rect 17406 20748 17408 20768
rect 17408 20748 17460 20768
rect 17460 20748 17462 20768
rect 17406 20712 17462 20748
rect 17130 20168 17186 20224
rect 17222 20032 17278 20088
rect 17682 20576 17738 20632
rect 17682 20032 17738 20088
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17958 21412 18014 21448
rect 17958 21392 17960 21412
rect 17960 21392 18012 21412
rect 18012 21392 18014 21412
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 18786 24248 18842 24304
rect 18786 24012 18788 24032
rect 18788 24012 18840 24032
rect 18840 24012 18842 24032
rect 18786 23976 18842 24012
rect 19062 23296 19118 23352
rect 18418 20712 18474 20768
rect 16578 18264 16634 18320
rect 16302 15000 16358 15056
rect 16762 18808 16818 18864
rect 17038 19080 17094 19136
rect 17130 18808 17186 18864
rect 16854 18400 16910 18456
rect 17038 17992 17094 18048
rect 16670 15544 16726 15600
rect 16854 15544 16910 15600
rect 16854 15272 16910 15328
rect 16486 14864 16542 14920
rect 16302 14456 16358 14512
rect 16486 14184 16542 14240
rect 16302 13524 16358 13560
rect 16302 13504 16304 13524
rect 16304 13504 16356 13524
rect 16356 13504 16358 13524
rect 16210 13096 16266 13152
rect 16302 12552 16358 12608
rect 16670 14864 16726 14920
rect 16670 14068 16726 14104
rect 16670 14048 16672 14068
rect 16672 14048 16724 14068
rect 16724 14048 16726 14068
rect 16670 13640 16726 13696
rect 16578 13504 16634 13560
rect 16854 13504 16910 13560
rect 16486 13096 16542 13152
rect 16486 12280 16542 12336
rect 16118 11736 16174 11792
rect 15198 6740 15200 6760
rect 15200 6740 15252 6760
rect 15252 6740 15254 6760
rect 15198 6704 15254 6740
rect 15014 3984 15070 4040
rect 15474 6740 15476 6760
rect 15476 6740 15528 6760
rect 15528 6740 15530 6760
rect 15474 6704 15530 6740
rect 15750 6568 15806 6624
rect 15290 3576 15346 3632
rect 15198 1128 15254 1184
rect 16118 8200 16174 8256
rect 15934 5752 15990 5808
rect 16394 11328 16450 11384
rect 17130 16224 17186 16280
rect 17130 15408 17186 15464
rect 17498 19488 17554 19544
rect 18694 22072 18750 22128
rect 18694 21664 18750 21720
rect 18878 21564 18880 21584
rect 18880 21564 18932 21584
rect 18932 21564 18934 21584
rect 18878 21528 18934 21564
rect 19154 21392 19210 21448
rect 19154 21120 19210 21176
rect 18510 19660 18512 19680
rect 18512 19660 18564 19680
rect 18564 19660 18566 19680
rect 18510 19624 18566 19660
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17774 19488 17830 19544
rect 18602 19488 18658 19544
rect 17774 19388 17776 19408
rect 17776 19388 17828 19408
rect 17828 19388 17830 19408
rect 17774 19352 17830 19388
rect 18602 19080 18658 19136
rect 17590 18536 17646 18592
rect 18050 18808 18106 18864
rect 18234 18808 18290 18864
rect 17682 18400 17738 18456
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17498 18264 17554 18320
rect 17958 18264 18014 18320
rect 18510 18400 18566 18456
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 18786 18808 18842 18864
rect 18786 17992 18842 18048
rect 18602 17448 18658 17504
rect 17774 16632 17830 16688
rect 18510 16904 18566 16960
rect 18418 16768 18474 16824
rect 17406 16360 17462 16416
rect 17590 16224 17646 16280
rect 17130 14884 17186 14920
rect 17130 14864 17132 14884
rect 17132 14864 17184 14884
rect 17184 14864 17186 14884
rect 17406 14864 17462 14920
rect 16486 9152 16542 9208
rect 16394 8608 16450 8664
rect 16946 11056 17002 11112
rect 16762 7540 16818 7576
rect 16762 7520 16764 7540
rect 16764 7520 16816 7540
rect 16816 7520 16818 7540
rect 16670 6432 16726 6488
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17590 15544 17646 15600
rect 17682 15272 17738 15328
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 18694 16496 18750 16552
rect 18602 16360 18658 16416
rect 18602 16088 18658 16144
rect 18970 20460 19026 20496
rect 18970 20440 18972 20460
rect 18972 20440 19024 20460
rect 19024 20440 19026 20460
rect 19706 23840 19762 23896
rect 19614 22752 19670 22808
rect 19430 22072 19486 22128
rect 19338 21800 19394 21856
rect 19062 19352 19118 19408
rect 18970 18400 19026 18456
rect 18970 16768 19026 16824
rect 18786 15680 18842 15736
rect 18510 15308 18512 15328
rect 18512 15308 18564 15328
rect 18564 15308 18566 15328
rect 18510 15272 18566 15308
rect 18694 15308 18696 15328
rect 18696 15308 18748 15328
rect 18748 15308 18750 15328
rect 18694 15272 18750 15308
rect 18418 15136 18474 15192
rect 18602 14456 18658 14512
rect 18510 14184 18566 14240
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 18694 13776 18750 13832
rect 18694 13252 18750 13288
rect 18694 13232 18696 13252
rect 18696 13232 18748 13252
rect 18748 13232 18750 13252
rect 17774 13096 17830 13152
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 18694 12960 18750 13016
rect 17774 12008 17830 12064
rect 17958 12416 18014 12472
rect 18142 12416 18198 12472
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17406 9832 17462 9888
rect 17406 9424 17462 9480
rect 17498 9288 17554 9344
rect 17590 9152 17646 9208
rect 17590 8880 17646 8936
rect 17590 7656 17646 7712
rect 17314 4664 17370 4720
rect 17314 4392 17370 4448
rect 17774 9832 17830 9888
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 18234 10240 18290 10296
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17866 9288 17922 9344
rect 17866 8900 17922 8936
rect 17866 8880 17868 8900
rect 17868 8880 17920 8900
rect 17920 8880 17922 8900
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 18050 8372 18052 8392
rect 18052 8372 18104 8392
rect 18104 8372 18106 8392
rect 18050 8336 18106 8372
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 18602 12008 18658 12064
rect 18970 16396 18972 16416
rect 18972 16396 19024 16416
rect 19024 16396 19026 16416
rect 18970 16360 19026 16396
rect 19154 18672 19210 18728
rect 19246 17992 19302 18048
rect 19154 17176 19210 17232
rect 18878 13232 18934 13288
rect 18878 12436 18934 12472
rect 18878 12416 18880 12436
rect 18880 12416 18932 12436
rect 18932 12416 18934 12436
rect 18878 11328 18934 11384
rect 18878 10920 18934 10976
rect 18786 9968 18842 10024
rect 18326 7248 18382 7304
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 18326 6296 18382 6352
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 18326 5072 18382 5128
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 18326 3848 18382 3904
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 17590 2488 17646 2544
rect 19890 22072 19946 22128
rect 19522 20848 19578 20904
rect 20074 22752 20130 22808
rect 20074 22344 20130 22400
rect 19614 20712 19670 20768
rect 20258 22480 20314 22536
rect 20350 21972 20352 21992
rect 20352 21972 20404 21992
rect 20404 21972 20406 21992
rect 20350 21936 20406 21972
rect 19522 18284 19578 18320
rect 19522 18264 19524 18284
rect 19524 18264 19576 18284
rect 19576 18264 19578 18284
rect 19430 16360 19486 16416
rect 19614 17992 19670 18048
rect 19614 17720 19670 17776
rect 19522 15272 19578 15328
rect 19246 13232 19302 13288
rect 19338 13096 19394 13152
rect 19062 9696 19118 9752
rect 19246 11872 19302 11928
rect 19798 17720 19854 17776
rect 20258 18672 20314 18728
rect 19982 17992 20038 18048
rect 19982 17720 20038 17776
rect 20442 18536 20498 18592
rect 20442 18264 20498 18320
rect 19890 15544 19946 15600
rect 20166 15564 20222 15600
rect 20166 15544 20168 15564
rect 20168 15544 20220 15564
rect 20220 15544 20222 15564
rect 20258 14728 20314 14784
rect 19798 14068 19854 14104
rect 19798 14048 19800 14068
rect 19800 14048 19852 14068
rect 19852 14048 19854 14068
rect 19798 13640 19854 13696
rect 19798 12960 19854 13016
rect 19338 6160 19394 6216
rect 19246 5752 19302 5808
rect 18878 4936 18934 4992
rect 19614 9288 19670 9344
rect 20074 14320 20130 14376
rect 20626 19624 20682 19680
rect 20534 17992 20590 18048
rect 20718 17584 20774 17640
rect 20534 16904 20590 16960
rect 20994 22888 21050 22944
rect 21086 21564 21088 21584
rect 21088 21564 21140 21584
rect 21140 21564 21142 21584
rect 21086 21528 21142 21564
rect 21086 21120 21142 21176
rect 21086 20304 21142 20360
rect 20994 19080 21050 19136
rect 21270 22752 21326 22808
rect 21362 22072 21418 22128
rect 21730 22344 21786 22400
rect 21730 22208 21786 22264
rect 21638 22072 21694 22128
rect 21454 21800 21510 21856
rect 21454 21256 21510 21312
rect 21546 20576 21602 20632
rect 21454 20032 21510 20088
rect 21086 18672 21142 18728
rect 20994 18264 21050 18320
rect 20534 15580 20536 15600
rect 20536 15580 20588 15600
rect 20588 15580 20590 15600
rect 20534 15544 20590 15580
rect 20166 11872 20222 11928
rect 19982 10240 20038 10296
rect 19982 9968 20038 10024
rect 19706 7112 19762 7168
rect 19706 6704 19762 6760
rect 19982 5228 20038 5264
rect 19982 5208 19984 5228
rect 19984 5208 20036 5228
rect 20036 5208 20038 5228
rect 19338 3984 19394 4040
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 20350 10240 20406 10296
rect 20534 14456 20590 14512
rect 20902 13912 20958 13968
rect 20718 13640 20774 13696
rect 20626 12008 20682 12064
rect 21086 13776 21142 13832
rect 20902 12552 20958 12608
rect 21638 18944 21694 19000
rect 21822 20848 21878 20904
rect 21822 20576 21878 20632
rect 22006 23432 22062 23488
rect 22006 22480 22062 22536
rect 22466 24928 22522 24984
rect 22466 23296 22522 23352
rect 22466 22752 22522 22808
rect 22282 22208 22338 22264
rect 22466 22072 22522 22128
rect 22190 20712 22246 20768
rect 22926 24792 22982 24848
rect 23386 24520 23442 24576
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 21822 17992 21878 18048
rect 20902 11464 20958 11520
rect 20166 2488 20222 2544
rect 21454 13932 21510 13968
rect 21454 13912 21456 13932
rect 21456 13912 21508 13932
rect 21508 13912 21510 13932
rect 21086 9152 21142 9208
rect 20810 3576 20866 3632
rect 21730 14764 21732 14784
rect 21732 14764 21784 14784
rect 21784 14764 21786 14784
rect 21730 14728 21786 14764
rect 22190 17448 22246 17504
rect 22098 17060 22154 17096
rect 22098 17040 22100 17060
rect 22100 17040 22152 17060
rect 22152 17040 22154 17060
rect 21914 12552 21970 12608
rect 21914 11872 21970 11928
rect 22374 19488 22430 19544
rect 22742 21256 22798 21312
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 23754 23296 23810 23352
rect 23662 22344 23718 22400
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 22742 20168 22798 20224
rect 22742 19488 22798 19544
rect 22650 19352 22706 19408
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 24122 22752 24178 22808
rect 23478 21140 23534 21176
rect 23478 21120 23480 21140
rect 23480 21120 23532 21140
rect 23532 21120 23534 21140
rect 23754 20848 23810 20904
rect 23570 20596 23626 20632
rect 23570 20576 23572 20596
rect 23572 20576 23624 20596
rect 23624 20576 23626 20596
rect 22926 19372 22982 19408
rect 22926 19352 22928 19372
rect 22928 19352 22980 19372
rect 22980 19352 22982 19372
rect 23110 19352 23166 19408
rect 22558 18536 22614 18592
rect 22558 18400 22614 18456
rect 22742 17040 22798 17096
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 23202 17720 23258 17776
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22650 16224 22706 16280
rect 22466 13912 22522 13968
rect 22650 13912 22706 13968
rect 22558 13776 22614 13832
rect 21454 7540 21510 7576
rect 21454 7520 21456 7540
rect 21456 7520 21508 7540
rect 21508 7520 21510 7540
rect 22098 11620 22154 11656
rect 22098 11600 22100 11620
rect 22100 11600 22152 11620
rect 22152 11600 22154 11620
rect 22006 9016 22062 9072
rect 21914 4684 21970 4720
rect 21914 4664 21916 4684
rect 21916 4664 21968 4684
rect 21968 4664 21970 4684
rect 22282 12552 22338 12608
rect 22282 10104 22338 10160
rect 22282 9696 22338 9752
rect 22190 6840 22246 6896
rect 22098 3712 22154 3768
rect 22006 2644 22062 2680
rect 22006 2624 22008 2644
rect 22008 2624 22060 2644
rect 22060 2624 22062 2644
rect 23570 19352 23626 19408
rect 23754 20032 23810 20088
rect 23662 19080 23718 19136
rect 23846 18400 23902 18456
rect 24122 18264 24178 18320
rect 24030 17992 24086 18048
rect 23754 17620 23756 17640
rect 23756 17620 23808 17640
rect 23808 17620 23810 17640
rect 23202 16360 23258 16416
rect 23754 17584 23810 17620
rect 23846 17484 23848 17504
rect 23848 17484 23900 17504
rect 23900 17484 23902 17504
rect 23846 17448 23902 17484
rect 23570 16788 23626 16824
rect 23570 16768 23572 16788
rect 23572 16768 23624 16788
rect 23624 16768 23626 16788
rect 23570 16224 23626 16280
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 23202 14864 23258 14920
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22834 11736 22890 11792
rect 23294 12280 23350 12336
rect 23294 11736 23350 11792
rect 23202 11600 23258 11656
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 23846 14320 23902 14376
rect 23846 12416 23902 12472
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 23386 10784 23442 10840
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 23294 6840 23350 6896
rect 23202 6296 23258 6352
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 23754 12144 23810 12200
rect 24122 17856 24178 17912
rect 24306 25336 24362 25392
rect 24582 23432 24638 23488
rect 24490 21664 24546 21720
rect 24490 20440 24546 20496
rect 24306 20304 24362 20360
rect 24490 18128 24546 18184
rect 24306 17040 24362 17096
rect 24122 16360 24178 16416
rect 24766 24404 24822 24440
rect 24766 24384 24768 24404
rect 24768 24384 24820 24404
rect 24820 24384 24822 24404
rect 25134 23840 25190 23896
rect 24766 22480 24822 22536
rect 24674 21120 24730 21176
rect 25042 22208 25098 22264
rect 25134 22092 25190 22128
rect 25134 22072 25136 22092
rect 25136 22072 25188 22092
rect 25188 22072 25190 22092
rect 25134 21412 25190 21448
rect 25134 21392 25136 21412
rect 25136 21392 25188 21412
rect 25188 21392 25190 21412
rect 24858 21120 24914 21176
rect 26054 24792 26110 24848
rect 25410 23024 25466 23080
rect 26054 23160 26110 23216
rect 26882 24928 26938 24984
rect 26238 24112 26294 24168
rect 26422 24112 26478 24168
rect 26146 23060 26148 23080
rect 26148 23060 26200 23080
rect 26200 23060 26202 23080
rect 26146 23024 26202 23060
rect 25318 22344 25374 22400
rect 24674 20748 24676 20768
rect 24676 20748 24728 20768
rect 24728 20748 24730 20768
rect 24674 20712 24730 20748
rect 24950 18400 25006 18456
rect 25318 18536 25374 18592
rect 24214 14728 24270 14784
rect 23846 11500 23848 11520
rect 23848 11500 23900 11520
rect 23900 11500 23902 11520
rect 23846 11464 23902 11500
rect 24030 10240 24086 10296
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 24582 15136 24638 15192
rect 24582 14864 24638 14920
rect 24490 14728 24546 14784
rect 24582 14592 24638 14648
rect 24950 16496 25006 16552
rect 24766 14320 24822 14376
rect 24674 12008 24730 12064
rect 24766 10920 24822 10976
rect 25134 13776 25190 13832
rect 25778 22888 25834 22944
rect 25778 22616 25834 22672
rect 25962 22516 25964 22536
rect 25964 22516 26016 22536
rect 26016 22516 26018 22536
rect 25962 22480 26018 22516
rect 25778 22344 25834 22400
rect 25778 21936 25834 21992
rect 25778 21664 25834 21720
rect 25686 20712 25742 20768
rect 25594 20576 25650 20632
rect 25594 18536 25650 18592
rect 25410 16768 25466 16824
rect 25502 15952 25558 16008
rect 26054 21936 26110 21992
rect 26330 23160 26386 23216
rect 26238 22072 26294 22128
rect 26422 22072 26478 22128
rect 26790 23976 26846 24032
rect 26606 23296 26662 23352
rect 26606 22616 26662 22672
rect 26606 22072 26662 22128
rect 26422 20848 26478 20904
rect 27158 24284 27160 24304
rect 27160 24284 27212 24304
rect 27212 24284 27214 24304
rect 27158 24248 27214 24284
rect 26974 22888 27030 22944
rect 26882 22616 26938 22672
rect 26514 19116 26516 19136
rect 26516 19116 26568 19136
rect 26568 19116 26570 19136
rect 26514 19080 26570 19116
rect 26054 18672 26110 18728
rect 26698 19624 26754 19680
rect 26422 17856 26478 17912
rect 25594 15272 25650 15328
rect 24858 7948 24914 7984
rect 24858 7928 24860 7948
rect 24860 7928 24912 7948
rect 24912 7928 24914 7948
rect 24398 7268 24454 7304
rect 24398 7248 24400 7268
rect 24400 7248 24452 7268
rect 24452 7248 24454 7268
rect 25502 14456 25558 14512
rect 25410 14048 25466 14104
rect 25686 14220 25688 14240
rect 25688 14220 25740 14240
rect 25740 14220 25742 14240
rect 25686 14184 25742 14220
rect 25410 13776 25466 13832
rect 25410 11056 25466 11112
rect 26238 16496 26294 16552
rect 26422 16360 26478 16416
rect 26790 18264 26846 18320
rect 27342 23432 27398 23488
rect 27802 23976 27858 24032
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 27802 23840 27858 23896
rect 27526 23296 27582 23352
rect 27802 23432 27858 23488
rect 27434 22888 27490 22944
rect 27250 22752 27306 22808
rect 26974 21528 27030 21584
rect 27066 21120 27122 21176
rect 26974 20984 27030 21040
rect 27618 22636 27674 22672
rect 27618 22616 27620 22636
rect 27620 22616 27672 22636
rect 27672 22616 27674 22636
rect 27710 22344 27766 22400
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27342 21528 27398 21584
rect 27066 18264 27122 18320
rect 26790 16496 26846 16552
rect 26422 15136 26478 15192
rect 26514 12416 26570 12472
rect 26146 10104 26202 10160
rect 25870 8744 25926 8800
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22098 1264 22154 1320
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 23386 2644 23442 2680
rect 23386 2624 23388 2644
rect 23388 2624 23440 2644
rect 23440 2624 23442 2644
rect 25962 8628 26018 8664
rect 25962 8608 25964 8628
rect 25964 8608 26016 8628
rect 26016 8608 26018 8628
rect 26238 9560 26294 9616
rect 26146 4528 26202 4584
rect 27710 21664 27766 21720
rect 28354 21800 28410 21856
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 28354 21684 28410 21720
rect 28354 21664 28356 21684
rect 28356 21664 28408 21684
rect 28408 21664 28410 21684
rect 27802 20984 27858 21040
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 28538 20032 28594 20088
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27342 15272 27398 15328
rect 27618 16360 27674 16416
rect 27526 15408 27582 15464
rect 27802 18572 27804 18592
rect 27804 18572 27856 18592
rect 27856 18572 27858 18592
rect 27802 18536 27858 18572
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27802 18400 27858 18456
rect 27802 18028 27804 18048
rect 27804 18028 27856 18048
rect 27856 18028 27858 18048
rect 27802 17992 27858 18028
rect 27894 17856 27950 17912
rect 28262 18128 28318 18184
rect 28998 24656 29054 24712
rect 28906 22208 28962 22264
rect 28906 22072 28962 22128
rect 28906 21664 28962 21720
rect 28630 19488 28686 19544
rect 27802 17448 27858 17504
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 28538 17448 28594 17504
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27802 16224 27858 16280
rect 27802 16088 27858 16144
rect 27986 16088 28042 16144
rect 27710 15952 27766 16008
rect 27986 15700 28042 15736
rect 27986 15680 27988 15700
rect 27988 15680 28040 15700
rect 28040 15680 28042 15700
rect 27710 15444 27712 15464
rect 27712 15444 27764 15464
rect 27764 15444 27766 15464
rect 27710 15408 27766 15444
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 29182 21528 29238 21584
rect 28998 19760 29054 19816
rect 28906 19488 28962 19544
rect 29090 19080 29146 19136
rect 29458 20712 29514 20768
rect 29182 18536 29238 18592
rect 29090 18400 29146 18456
rect 29458 18536 29514 18592
rect 28998 18128 29054 18184
rect 29550 17720 29606 17776
rect 28906 17312 28962 17368
rect 29274 17448 29330 17504
rect 30010 22072 30066 22128
rect 30562 22228 30618 22264
rect 30562 22208 30564 22228
rect 30564 22208 30616 22228
rect 30616 22208 30618 22228
rect 30378 22072 30434 22128
rect 30010 21120 30066 21176
rect 29918 20848 29974 20904
rect 29642 16788 29698 16824
rect 29642 16768 29644 16788
rect 29644 16768 29696 16788
rect 29696 16768 29698 16788
rect 29826 17856 29882 17912
rect 29918 16768 29974 16824
rect 28354 14864 28410 14920
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27894 13640 27950 13696
rect 27158 10512 27214 10568
rect 26606 992 26662 1048
rect 27342 11464 27398 11520
rect 27434 11228 27436 11248
rect 27436 11228 27488 11248
rect 27488 11228 27490 11248
rect 27434 11192 27490 11228
rect 27434 10784 27490 10840
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27802 11892 27858 11928
rect 27802 11872 27804 11892
rect 27804 11872 27856 11892
rect 27856 11872 27858 11892
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27710 9832 27766 9888
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 28722 15020 28778 15056
rect 28722 15000 28724 15020
rect 28724 15000 28776 15020
rect 28776 15000 28778 15020
rect 28722 14864 28778 14920
rect 28722 14592 28778 14648
rect 28906 13252 28962 13288
rect 28906 13232 28908 13252
rect 28908 13232 28960 13252
rect 28960 13232 28962 13252
rect 28906 12724 28908 12744
rect 28908 12724 28960 12744
rect 28960 12724 28962 12744
rect 28906 12688 28962 12724
rect 28354 9016 28410 9072
rect 27618 7792 27674 7848
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27618 3440 27674 3496
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 27250 856 27306 912
rect 28446 1808 28502 1864
rect 29182 16088 29238 16144
rect 30194 19660 30196 19680
rect 30196 19660 30248 19680
rect 30248 19660 30250 19680
rect 30194 19624 30250 19660
rect 30194 18572 30196 18592
rect 30196 18572 30248 18592
rect 30248 18572 30250 18592
rect 30194 18536 30250 18572
rect 30378 19760 30434 19816
rect 30746 20712 30802 20768
rect 30470 18264 30526 18320
rect 30102 17584 30158 17640
rect 30194 17040 30250 17096
rect 30654 17176 30710 17232
rect 29826 12552 29882 12608
rect 29182 8880 29238 8936
rect 30010 12280 30066 12336
rect 29642 7384 29698 7440
rect 30654 15544 30710 15600
rect 30562 11736 30618 11792
rect 31850 23432 31906 23488
rect 31482 22752 31538 22808
rect 31022 22616 31078 22672
rect 31114 21548 31170 21584
rect 31114 21528 31116 21548
rect 31116 21528 31168 21548
rect 31168 21528 31170 21548
rect 31114 20748 31116 20768
rect 31116 20748 31168 20768
rect 31168 20748 31170 20768
rect 31114 20712 31170 20748
rect 31022 18264 31078 18320
rect 31758 22380 31760 22400
rect 31760 22380 31812 22400
rect 31812 22380 31814 22400
rect 31758 22344 31814 22380
rect 31942 23296 31998 23352
rect 31574 21256 31630 21312
rect 31390 20576 31446 20632
rect 31482 18944 31538 19000
rect 31666 20884 31668 20904
rect 31668 20884 31720 20904
rect 31720 20884 31722 20904
rect 31666 20848 31722 20884
rect 31942 20712 31998 20768
rect 31758 19116 31760 19136
rect 31760 19116 31812 19136
rect 31812 19116 31814 19136
rect 31758 19080 31814 19116
rect 31666 18028 31668 18048
rect 31668 18028 31720 18048
rect 31720 18028 31722 18048
rect 31666 17992 31722 18028
rect 30838 13096 30894 13152
rect 31206 15000 31262 15056
rect 32586 24384 32642 24440
rect 32402 23160 32458 23216
rect 32494 18536 32550 18592
rect 31758 17584 31814 17640
rect 31666 16768 31722 16824
rect 31574 15952 31630 16008
rect 31758 15544 31814 15600
rect 31390 10240 31446 10296
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 33138 22480 33194 22536
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 33414 20576 33470 20632
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 32678 19896 32734 19952
rect 32770 19352 32826 19408
rect 31942 13504 31998 13560
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 33414 18944 33470 19000
rect 32862 18672 32918 18728
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 33690 8472 33746 8528
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32770 2896 32826 2952
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 34150 22616 34206 22672
rect 34058 19488 34114 19544
rect 34334 22772 34390 22808
rect 34334 22752 34336 22772
rect 34336 22752 34388 22772
rect 34388 22752 34390 22772
rect 34334 21664 34390 21720
rect 34518 21392 34574 21448
rect 34334 20340 34336 20360
rect 34336 20340 34388 20360
rect 34388 20340 34390 20360
rect 34334 20304 34390 20340
rect 34610 18944 34666 19000
rect 34426 17040 34482 17096
rect 34242 10648 34298 10704
rect 34058 6704 34114 6760
rect 34886 16088 34942 16144
rect 34794 14864 34850 14920
rect 33782 1944 33838 2000
rect 29090 584 29146 640
rect 35070 15136 35126 15192
rect 35254 13096 35310 13152
rect 36082 20984 36138 21040
rect 35806 18808 35862 18864
rect 35898 17856 35954 17912
rect 35530 17312 35586 17368
rect 36726 19624 36782 19680
rect 37094 23024 37150 23080
rect 36818 18264 36874 18320
rect 36910 17756 36912 17776
rect 36912 17756 36964 17776
rect 36964 17756 36966 17776
rect 36910 17720 36966 17756
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 37738 23568 37794 23624
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37370 17484 37372 17504
rect 37372 17484 37424 17504
rect 37424 17484 37426 17504
rect 37370 17448 37426 17484
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 38750 21936 38806 21992
rect 39026 20460 39082 20496
rect 39026 20440 39028 20460
rect 39028 20440 39080 20460
rect 39080 20440 39082 20460
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37462 12144 37518 12200
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 38658 15408 38714 15464
rect 41142 23160 41198 23216
rect 39946 12824 40002 12880
rect 40774 19216 40830 19272
rect 40958 11600 41014 11656
rect 41970 25744 42026 25800
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42706 23740 42708 23760
rect 42708 23740 42760 23760
rect 42760 23740 42762 23760
rect 42706 23704 42762 23740
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 41878 10512 41934 10568
rect 39578 8336 39634 8392
rect 38382 6840 38438 6896
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 43718 24792 43774 24848
rect 43350 20848 43406 20904
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 43350 5072 43406 5128
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 44086 21528 44142 21584
rect 44822 24112 44878 24168
rect 44730 19760 44786 19816
rect 43902 16496 43958 16552
rect 46202 24792 46258 24848
rect 46110 23196 46112 23216
rect 46112 23196 46164 23216
rect 46164 23196 46166 23216
rect 46110 23160 46166 23196
rect 46386 23704 46442 23760
rect 46754 22616 46810 22672
rect 46570 21936 46626 21992
rect 46386 14456 46442 14512
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 46570 14320 46626 14376
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 48962 9968 49018 10024
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 45190 9424 45246 9480
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 49238 22480 49294 22536
rect 49146 20984 49202 21040
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 43810 2352 43866 2408
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
<< metal3 >>
rect 15510 25740 15516 25804
rect 15580 25802 15586 25804
rect 41965 25802 42031 25805
rect 15580 25800 42031 25802
rect 15580 25744 41970 25800
rect 42026 25744 42031 25800
rect 15580 25742 42031 25744
rect 15580 25740 15586 25742
rect 41965 25739 42031 25742
rect 0 25666 800 25696
rect 4061 25666 4127 25669
rect 0 25664 4127 25666
rect 0 25608 4066 25664
rect 4122 25608 4127 25664
rect 0 25606 4127 25608
rect 0 25576 800 25606
rect 4061 25603 4127 25606
rect 6177 25530 6243 25533
rect 21398 25530 21404 25532
rect 6177 25528 21404 25530
rect 6177 25472 6182 25528
rect 6238 25472 21404 25528
rect 6177 25470 21404 25472
rect 6177 25467 6243 25470
rect 21398 25468 21404 25470
rect 21468 25468 21474 25532
rect 11973 25394 12039 25397
rect 24301 25394 24367 25397
rect 11973 25392 24367 25394
rect 11973 25336 11978 25392
rect 12034 25336 24306 25392
rect 24362 25336 24367 25392
rect 11973 25334 24367 25336
rect 11973 25331 12039 25334
rect 24301 25331 24367 25334
rect 0 25258 800 25288
rect 3325 25258 3391 25261
rect 0 25256 3391 25258
rect 0 25200 3330 25256
rect 3386 25200 3391 25256
rect 0 25198 3391 25200
rect 0 25168 800 25198
rect 3325 25195 3391 25198
rect 9857 25258 9923 25261
rect 27654 25258 27660 25260
rect 9857 25256 27660 25258
rect 9857 25200 9862 25256
rect 9918 25200 27660 25256
rect 9857 25198 27660 25200
rect 9857 25195 9923 25198
rect 27654 25196 27660 25198
rect 27724 25196 27730 25260
rect 4797 25122 4863 25125
rect 27470 25122 27476 25124
rect 4797 25120 27476 25122
rect 4797 25064 4802 25120
rect 4858 25064 27476 25120
rect 4797 25062 27476 25064
rect 4797 25059 4863 25062
rect 27470 25060 27476 25062
rect 27540 25060 27546 25124
rect 22461 24986 22527 24989
rect 26877 24986 26943 24989
rect 22461 24984 26943 24986
rect 22461 24928 22466 24984
rect 22522 24928 26882 24984
rect 26938 24928 26943 24984
rect 22461 24926 26943 24928
rect 22461 24923 22527 24926
rect 26877 24923 26943 24926
rect 0 24850 800 24880
rect 3969 24850 4035 24853
rect 0 24848 4035 24850
rect 0 24792 3974 24848
rect 4030 24792 4035 24848
rect 0 24790 4035 24792
rect 0 24760 800 24790
rect 3969 24787 4035 24790
rect 11053 24850 11119 24853
rect 16481 24850 16547 24853
rect 11053 24848 16547 24850
rect 11053 24792 11058 24848
rect 11114 24792 16486 24848
rect 16542 24792 16547 24848
rect 11053 24790 16547 24792
rect 11053 24787 11119 24790
rect 16481 24787 16547 24790
rect 22921 24850 22987 24853
rect 23606 24850 23612 24852
rect 22921 24848 23612 24850
rect 22921 24792 22926 24848
rect 22982 24792 23612 24848
rect 22921 24790 23612 24792
rect 22921 24787 22987 24790
rect 23606 24788 23612 24790
rect 23676 24788 23682 24852
rect 26049 24850 26115 24853
rect 43713 24850 43779 24853
rect 26049 24848 43779 24850
rect 26049 24792 26054 24848
rect 26110 24792 43718 24848
rect 43774 24792 43779 24848
rect 26049 24790 43779 24792
rect 26049 24787 26115 24790
rect 43713 24787 43779 24790
rect 46197 24850 46263 24853
rect 50200 24850 51000 24880
rect 46197 24848 51000 24850
rect 46197 24792 46202 24848
rect 46258 24792 51000 24848
rect 46197 24790 51000 24792
rect 46197 24787 46263 24790
rect 50200 24760 51000 24790
rect 12249 24714 12315 24717
rect 18597 24714 18663 24717
rect 28993 24714 29059 24717
rect 12249 24712 17050 24714
rect 12249 24656 12254 24712
rect 12310 24656 17050 24712
rect 12249 24654 17050 24656
rect 12249 24651 12315 24654
rect 16990 24578 17050 24654
rect 18597 24712 29059 24714
rect 18597 24656 18602 24712
rect 18658 24656 28998 24712
rect 29054 24656 29059 24712
rect 18597 24654 29059 24656
rect 18597 24651 18663 24654
rect 28993 24651 29059 24654
rect 20294 24578 20300 24580
rect 16990 24518 20300 24578
rect 20294 24516 20300 24518
rect 20364 24516 20370 24580
rect 23381 24578 23447 24581
rect 25446 24578 25452 24580
rect 23381 24576 25452 24578
rect 23381 24520 23386 24576
rect 23442 24520 25452 24576
rect 23381 24518 25452 24520
rect 23381 24515 23447 24518
rect 25446 24516 25452 24518
rect 25516 24516 25522 24580
rect 2946 24512 3262 24513
rect 0 24442 800 24472
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 2773 24442 2839 24445
rect 0 24440 2839 24442
rect 0 24384 2778 24440
rect 2834 24384 2839 24440
rect 0 24382 2839 24384
rect 0 24352 800 24382
rect 2773 24379 2839 24382
rect 15653 24442 15719 24445
rect 24761 24442 24827 24445
rect 32581 24442 32647 24445
rect 15653 24440 22110 24442
rect 15653 24384 15658 24440
rect 15714 24384 22110 24440
rect 15653 24382 22110 24384
rect 15653 24379 15719 24382
rect 2221 24306 2287 24309
rect 13537 24306 13603 24309
rect 2221 24304 13603 24306
rect 2221 24248 2226 24304
rect 2282 24248 13542 24304
rect 13598 24248 13603 24304
rect 2221 24246 13603 24248
rect 2221 24243 2287 24246
rect 13537 24243 13603 24246
rect 13905 24306 13971 24309
rect 14038 24306 14044 24308
rect 13905 24304 14044 24306
rect 13905 24248 13910 24304
rect 13966 24248 14044 24304
rect 13905 24246 14044 24248
rect 13905 24243 13971 24246
rect 14038 24244 14044 24246
rect 14108 24306 14114 24308
rect 18781 24306 18847 24309
rect 14108 24304 18847 24306
rect 14108 24248 18786 24304
rect 18842 24248 18847 24304
rect 14108 24246 18847 24248
rect 22050 24306 22110 24382
rect 24761 24440 32647 24442
rect 24761 24384 24766 24440
rect 24822 24384 32586 24440
rect 32642 24384 32647 24440
rect 24761 24382 32647 24384
rect 24761 24379 24827 24382
rect 32581 24379 32647 24382
rect 27153 24306 27219 24309
rect 22050 24304 27219 24306
rect 22050 24248 27158 24304
rect 27214 24248 27219 24304
rect 22050 24246 27219 24248
rect 14108 24244 14114 24246
rect 18781 24243 18847 24246
rect 27153 24243 27219 24246
rect 12525 24170 12591 24173
rect 12750 24170 12756 24172
rect 12525 24168 12756 24170
rect 12525 24112 12530 24168
rect 12586 24112 12756 24168
rect 12525 24110 12756 24112
rect 12525 24107 12591 24110
rect 12750 24108 12756 24110
rect 12820 24108 12826 24172
rect 14273 24170 14339 24173
rect 26233 24170 26299 24173
rect 14273 24168 26299 24170
rect 14273 24112 14278 24168
rect 14334 24112 26238 24168
rect 26294 24112 26299 24168
rect 14273 24110 26299 24112
rect 14273 24107 14339 24110
rect 26233 24107 26299 24110
rect 26417 24170 26483 24173
rect 44817 24170 44883 24173
rect 26417 24168 44883 24170
rect 26417 24112 26422 24168
rect 26478 24112 44822 24168
rect 44878 24112 44883 24168
rect 26417 24110 44883 24112
rect 26417 24107 26483 24110
rect 44817 24107 44883 24110
rect 0 24034 800 24064
rect 3693 24034 3759 24037
rect 0 24032 3759 24034
rect 0 23976 3698 24032
rect 3754 23976 3759 24032
rect 0 23974 3759 23976
rect 0 23944 800 23974
rect 3693 23971 3759 23974
rect 10869 24034 10935 24037
rect 15009 24034 15075 24037
rect 10869 24032 15075 24034
rect 10869 23976 10874 24032
rect 10930 23976 15014 24032
rect 15070 23976 15075 24032
rect 10869 23974 15075 23976
rect 10869 23971 10935 23974
rect 15009 23971 15075 23974
rect 18781 24034 18847 24037
rect 20478 24034 20484 24036
rect 18781 24032 20484 24034
rect 18781 23976 18786 24032
rect 18842 23976 20484 24032
rect 18781 23974 20484 23976
rect 18781 23971 18847 23974
rect 20478 23972 20484 23974
rect 20548 23972 20554 24036
rect 26785 24034 26851 24037
rect 27797 24034 27863 24037
rect 22050 24032 27863 24034
rect 22050 23976 26790 24032
rect 26846 23976 27802 24032
rect 27858 23976 27863 24032
rect 22050 23974 27863 23976
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 10593 23898 10659 23901
rect 16665 23898 16731 23901
rect 10593 23896 16731 23898
rect 10593 23840 10598 23896
rect 10654 23840 16670 23896
rect 16726 23840 16731 23896
rect 10593 23838 16731 23840
rect 10593 23835 10659 23838
rect 16665 23835 16731 23838
rect 16798 23836 16804 23900
rect 16868 23898 16874 23900
rect 17033 23898 17099 23901
rect 16868 23896 17099 23898
rect 16868 23840 17038 23896
rect 17094 23840 17099 23896
rect 16868 23838 17099 23840
rect 16868 23836 16874 23838
rect 17033 23835 17099 23838
rect 19701 23898 19767 23901
rect 22050 23898 22110 23974
rect 26785 23971 26851 23974
rect 27797 23971 27863 23974
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 47946 23903 48262 23904
rect 19701 23896 22110 23898
rect 19701 23840 19706 23896
rect 19762 23840 22110 23896
rect 19701 23838 22110 23840
rect 25129 23898 25195 23901
rect 27797 23898 27863 23901
rect 50200 23898 51000 23928
rect 25129 23896 27863 23898
rect 25129 23840 25134 23896
rect 25190 23840 27802 23896
rect 27858 23840 27863 23896
rect 25129 23838 27863 23840
rect 19701 23835 19767 23838
rect 25129 23835 25195 23838
rect 27797 23835 27863 23838
rect 48454 23838 51000 23898
rect 9673 23762 9739 23765
rect 15285 23762 15351 23765
rect 9673 23760 15351 23762
rect 9673 23704 9678 23760
rect 9734 23704 15290 23760
rect 15346 23704 15351 23760
rect 9673 23702 15351 23704
rect 9673 23699 9739 23702
rect 15285 23699 15351 23702
rect 17033 23762 17099 23765
rect 42701 23762 42767 23765
rect 17033 23760 42767 23762
rect 17033 23704 17038 23760
rect 17094 23704 42706 23760
rect 42762 23704 42767 23760
rect 17033 23702 42767 23704
rect 17033 23699 17099 23702
rect 42701 23699 42767 23702
rect 46381 23762 46447 23765
rect 48454 23762 48514 23838
rect 50200 23808 51000 23838
rect 46381 23760 48514 23762
rect 46381 23704 46386 23760
rect 46442 23704 48514 23760
rect 46381 23702 48514 23704
rect 46381 23699 46447 23702
rect 0 23626 800 23656
rect 4061 23626 4127 23629
rect 0 23624 4127 23626
rect 0 23568 4066 23624
rect 4122 23568 4127 23624
rect 0 23566 4127 23568
rect 0 23536 800 23566
rect 4061 23563 4127 23566
rect 10685 23626 10751 23629
rect 13670 23626 13676 23628
rect 10685 23624 13676 23626
rect 10685 23568 10690 23624
rect 10746 23568 13676 23624
rect 10685 23566 13676 23568
rect 10685 23563 10751 23566
rect 13670 23564 13676 23566
rect 13740 23564 13746 23628
rect 16389 23626 16455 23629
rect 37733 23626 37799 23629
rect 16389 23624 37799 23626
rect 16389 23568 16394 23624
rect 16450 23568 37738 23624
rect 37794 23568 37799 23624
rect 16389 23566 37799 23568
rect 16389 23563 16455 23566
rect 37733 23563 37799 23566
rect 4705 23490 4771 23493
rect 8477 23490 8543 23493
rect 4705 23488 8543 23490
rect 4705 23432 4710 23488
rect 4766 23432 8482 23488
rect 8538 23432 8543 23488
rect 4705 23430 8543 23432
rect 4705 23427 4771 23430
rect 8477 23427 8543 23430
rect 8886 23428 8892 23492
rect 8956 23490 8962 23492
rect 9765 23490 9831 23493
rect 8956 23488 9831 23490
rect 8956 23432 9770 23488
rect 9826 23432 9831 23488
rect 8956 23430 9831 23432
rect 8956 23428 8962 23430
rect 9765 23427 9831 23430
rect 11697 23490 11763 23493
rect 14917 23492 14983 23493
rect 15469 23492 15535 23493
rect 12382 23490 12388 23492
rect 11697 23488 12388 23490
rect 11697 23432 11702 23488
rect 11758 23432 12388 23488
rect 11697 23430 12388 23432
rect 11697 23427 11763 23430
rect 12382 23428 12388 23430
rect 12452 23428 12458 23492
rect 14917 23488 14964 23492
rect 15028 23490 15034 23492
rect 15469 23490 15516 23492
rect 14917 23432 14922 23488
rect 14917 23428 14964 23432
rect 15028 23430 15074 23490
rect 15424 23488 15516 23490
rect 15424 23432 15474 23488
rect 15424 23430 15516 23432
rect 15028 23428 15034 23430
rect 15469 23428 15516 23430
rect 15580 23428 15586 23492
rect 16481 23490 16547 23493
rect 22001 23490 22067 23493
rect 16481 23488 22067 23490
rect 16481 23432 16486 23488
rect 16542 23432 22006 23488
rect 22062 23432 22067 23488
rect 16481 23430 22067 23432
rect 14917 23427 14983 23428
rect 15469 23427 15535 23428
rect 16481 23427 16547 23430
rect 22001 23427 22067 23430
rect 24577 23490 24643 23493
rect 27337 23492 27403 23493
rect 24710 23490 24716 23492
rect 24577 23488 24716 23490
rect 24577 23432 24582 23488
rect 24638 23432 24716 23488
rect 24577 23430 24716 23432
rect 24577 23427 24643 23430
rect 24710 23428 24716 23430
rect 24780 23428 24786 23492
rect 27286 23490 27292 23492
rect 27246 23430 27292 23490
rect 27356 23488 27403 23492
rect 27398 23432 27403 23488
rect 27286 23428 27292 23430
rect 27356 23428 27403 23432
rect 27337 23427 27403 23428
rect 27797 23490 27863 23493
rect 31845 23490 31911 23493
rect 27797 23488 31911 23490
rect 27797 23432 27802 23488
rect 27858 23432 31850 23488
rect 31906 23432 31911 23488
rect 27797 23430 31911 23432
rect 27797 23427 27863 23430
rect 31845 23427 31911 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 13353 23354 13419 23357
rect 15510 23354 15516 23356
rect 13353 23352 15516 23354
rect 13353 23296 13358 23352
rect 13414 23296 15516 23352
rect 13353 23294 15516 23296
rect 13353 23291 13419 23294
rect 15510 23292 15516 23294
rect 15580 23292 15586 23356
rect 15837 23354 15903 23357
rect 18822 23354 18828 23356
rect 15837 23352 18828 23354
rect 15837 23296 15842 23352
rect 15898 23296 18828 23352
rect 15837 23294 18828 23296
rect 15837 23291 15903 23294
rect 18822 23292 18828 23294
rect 18892 23292 18898 23356
rect 19057 23354 19123 23357
rect 22461 23354 22527 23357
rect 19057 23352 22527 23354
rect 19057 23296 19062 23352
rect 19118 23296 22466 23352
rect 22522 23296 22527 23352
rect 19057 23294 22527 23296
rect 19057 23291 19123 23294
rect 22461 23291 22527 23294
rect 23749 23354 23815 23357
rect 26601 23354 26667 23357
rect 23749 23352 26667 23354
rect 23749 23296 23754 23352
rect 23810 23296 26606 23352
rect 26662 23296 26667 23352
rect 23749 23294 26667 23296
rect 23749 23291 23815 23294
rect 26601 23291 26667 23294
rect 27521 23354 27587 23357
rect 31937 23354 32003 23357
rect 27521 23352 32003 23354
rect 27521 23296 27526 23352
rect 27582 23296 31942 23352
rect 31998 23296 32003 23352
rect 27521 23294 32003 23296
rect 27521 23291 27587 23294
rect 31937 23291 32003 23294
rect 0 23218 800 23248
rect 3601 23218 3667 23221
rect 14365 23218 14431 23221
rect 14641 23218 14707 23221
rect 26049 23218 26115 23221
rect 0 23158 2790 23218
rect 0 23128 800 23158
rect 2730 23082 2790 23158
rect 3601 23216 14431 23218
rect 3601 23160 3606 23216
rect 3662 23160 14370 23216
rect 14426 23160 14431 23216
rect 3601 23158 14431 23160
rect 3601 23155 3667 23158
rect 14365 23155 14431 23158
rect 14598 23216 26115 23218
rect 14598 23160 14646 23216
rect 14702 23160 26054 23216
rect 26110 23160 26115 23216
rect 14598 23158 26115 23160
rect 14598 23155 14707 23158
rect 26049 23155 26115 23158
rect 26325 23218 26391 23221
rect 32397 23218 32463 23221
rect 26325 23216 32463 23218
rect 26325 23160 26330 23216
rect 26386 23160 32402 23216
rect 32458 23160 32463 23216
rect 26325 23158 32463 23160
rect 26325 23155 26391 23158
rect 32397 23155 32463 23158
rect 41137 23218 41203 23221
rect 46105 23218 46171 23221
rect 41137 23216 46171 23218
rect 41137 23160 41142 23216
rect 41198 23160 46110 23216
rect 46166 23160 46171 23216
rect 41137 23158 46171 23160
rect 41137 23155 41203 23158
rect 46105 23155 46171 23158
rect 3877 23082 3943 23085
rect 2730 23080 3943 23082
rect 2730 23024 3882 23080
rect 3938 23024 3943 23080
rect 2730 23022 3943 23024
rect 3877 23019 3943 23022
rect 11789 23082 11855 23085
rect 14598 23082 14658 23155
rect 11789 23080 14658 23082
rect 11789 23024 11794 23080
rect 11850 23024 14658 23080
rect 11789 23022 14658 23024
rect 17953 23082 18019 23085
rect 25405 23082 25471 23085
rect 17953 23080 25471 23082
rect 17953 23024 17958 23080
rect 18014 23024 25410 23080
rect 25466 23024 25471 23080
rect 17953 23022 25471 23024
rect 11789 23019 11855 23022
rect 17953 23019 18019 23022
rect 25405 23019 25471 23022
rect 26141 23082 26207 23085
rect 37089 23082 37155 23085
rect 26141 23080 37155 23082
rect 26141 23024 26146 23080
rect 26202 23024 37094 23080
rect 37150 23024 37155 23080
rect 26141 23022 37155 23024
rect 26141 23019 26207 23022
rect 37089 23019 37155 23022
rect 11973 22946 12039 22949
rect 14089 22946 14155 22949
rect 11973 22944 14155 22946
rect 11973 22888 11978 22944
rect 12034 22888 14094 22944
rect 14150 22888 14155 22944
rect 11973 22886 14155 22888
rect 11973 22883 12039 22886
rect 14089 22883 14155 22886
rect 14365 22946 14431 22949
rect 15561 22946 15627 22949
rect 14365 22944 15627 22946
rect 14365 22888 14370 22944
rect 14426 22888 15566 22944
rect 15622 22888 15627 22944
rect 14365 22886 15627 22888
rect 14365 22883 14431 22886
rect 15561 22883 15627 22886
rect 20989 22946 21055 22949
rect 25773 22946 25839 22949
rect 20989 22944 25839 22946
rect 20989 22888 20994 22944
rect 21050 22888 25778 22944
rect 25834 22888 25839 22944
rect 20989 22886 25839 22888
rect 20989 22883 21055 22886
rect 25773 22883 25839 22886
rect 26969 22946 27035 22949
rect 27429 22946 27495 22949
rect 50200 22946 51000 22976
rect 26969 22944 27495 22946
rect 26969 22888 26974 22944
rect 27030 22888 27434 22944
rect 27490 22888 27495 22944
rect 26969 22886 27495 22888
rect 26969 22883 27035 22886
rect 27429 22883 27495 22886
rect 48454 22886 51000 22946
rect 7946 22880 8262 22881
rect 0 22810 800 22840
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 3785 22810 3851 22813
rect 12525 22810 12591 22813
rect 0 22808 3851 22810
rect 0 22752 3790 22808
rect 3846 22752 3851 22808
rect 0 22750 3851 22752
rect 0 22720 800 22750
rect 3785 22747 3851 22750
rect 8342 22808 12591 22810
rect 8342 22752 12530 22808
rect 12586 22752 12591 22808
rect 8342 22750 12591 22752
rect 5533 22674 5599 22677
rect 8342 22674 8402 22750
rect 12525 22747 12591 22750
rect 12893 22810 12959 22813
rect 12893 22808 17832 22810
rect 12893 22752 12898 22808
rect 12954 22752 17832 22808
rect 12893 22750 17832 22752
rect 12893 22747 12959 22750
rect 5533 22672 8402 22674
rect 5533 22616 5538 22672
rect 5594 22616 8402 22672
rect 5533 22614 8402 22616
rect 11421 22674 11487 22677
rect 17534 22674 17540 22676
rect 11421 22672 17540 22674
rect 11421 22616 11426 22672
rect 11482 22616 17540 22672
rect 11421 22614 17540 22616
rect 5533 22611 5599 22614
rect 11421 22611 11487 22614
rect 17534 22612 17540 22614
rect 17604 22612 17610 22676
rect 17772 22674 17832 22750
rect 19374 22748 19380 22812
rect 19444 22810 19450 22812
rect 19609 22810 19675 22813
rect 19444 22808 19675 22810
rect 19444 22752 19614 22808
rect 19670 22752 19675 22808
rect 19444 22750 19675 22752
rect 19444 22748 19450 22750
rect 19609 22747 19675 22750
rect 20069 22810 20135 22813
rect 21265 22810 21331 22813
rect 20069 22808 21331 22810
rect 20069 22752 20074 22808
rect 20130 22752 21270 22808
rect 21326 22752 21331 22808
rect 20069 22750 21331 22752
rect 20069 22747 20135 22750
rect 21265 22747 21331 22750
rect 22461 22810 22527 22813
rect 24117 22810 24183 22813
rect 27245 22810 27311 22813
rect 22461 22808 27311 22810
rect 22461 22752 22466 22808
rect 22522 22752 24122 22808
rect 24178 22752 27250 22808
rect 27306 22752 27311 22808
rect 22461 22750 27311 22752
rect 22461 22747 22527 22750
rect 24117 22747 24183 22750
rect 27245 22747 27311 22750
rect 31477 22810 31543 22813
rect 34329 22810 34395 22813
rect 31477 22808 34395 22810
rect 31477 22752 31482 22808
rect 31538 22752 34334 22808
rect 34390 22752 34395 22808
rect 31477 22750 34395 22752
rect 31477 22747 31543 22750
rect 34329 22747 34395 22750
rect 25773 22674 25839 22677
rect 26601 22674 26667 22677
rect 17772 22614 25514 22674
rect 3325 22538 3391 22541
rect 12893 22538 12959 22541
rect 2270 22536 3391 22538
rect 2270 22480 3330 22536
rect 3386 22480 3391 22536
rect 2270 22478 3391 22480
rect 0 22402 800 22432
rect 2270 22402 2330 22478
rect 3325 22475 3391 22478
rect 12758 22536 12959 22538
rect 12758 22480 12898 22536
rect 12954 22480 12959 22536
rect 12758 22478 12959 22480
rect 0 22342 2330 22402
rect 12433 22402 12499 22405
rect 12758 22402 12818 22478
rect 12893 22475 12959 22478
rect 14273 22538 14339 22541
rect 20253 22538 20319 22541
rect 14273 22536 20319 22538
rect 14273 22480 14278 22536
rect 14334 22480 20258 22536
rect 20314 22480 20319 22536
rect 14273 22478 20319 22480
rect 14273 22475 14339 22478
rect 20253 22475 20319 22478
rect 22001 22538 22067 22541
rect 24761 22538 24827 22541
rect 22001 22536 24827 22538
rect 22001 22480 22006 22536
rect 22062 22480 24766 22536
rect 24822 22480 24827 22536
rect 22001 22478 24827 22480
rect 22001 22475 22067 22478
rect 24761 22475 24827 22478
rect 12433 22400 12818 22402
rect 12433 22344 12438 22400
rect 12494 22344 12818 22400
rect 12433 22342 12818 22344
rect 14825 22402 14891 22405
rect 20069 22402 20135 22405
rect 14825 22400 20135 22402
rect 14825 22344 14830 22400
rect 14886 22344 20074 22400
rect 20130 22344 20135 22400
rect 14825 22342 20135 22344
rect 0 22312 800 22342
rect 12433 22339 12499 22342
rect 14825 22339 14891 22342
rect 20069 22339 20135 22342
rect 20294 22340 20300 22404
rect 20364 22402 20370 22404
rect 21582 22402 21588 22404
rect 20364 22342 21588 22402
rect 20364 22340 20370 22342
rect 21582 22340 21588 22342
rect 21652 22340 21658 22404
rect 21725 22402 21791 22405
rect 22686 22402 22692 22404
rect 21725 22400 22692 22402
rect 21725 22344 21730 22400
rect 21786 22344 22692 22400
rect 21725 22342 22692 22344
rect 21725 22339 21791 22342
rect 22686 22340 22692 22342
rect 22756 22340 22762 22404
rect 23657 22402 23723 22405
rect 25313 22402 25379 22405
rect 23657 22400 25379 22402
rect 23657 22344 23662 22400
rect 23718 22344 25318 22400
rect 25374 22344 25379 22400
rect 23657 22342 25379 22344
rect 23657 22339 23723 22342
rect 25313 22339 25379 22342
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 9029 22266 9095 22269
rect 12709 22266 12775 22269
rect 9029 22264 12775 22266
rect 9029 22208 9034 22264
rect 9090 22208 12714 22264
rect 12770 22208 12775 22264
rect 9029 22206 12775 22208
rect 9029 22203 9095 22206
rect 12709 22203 12775 22206
rect 16665 22266 16731 22269
rect 21725 22266 21791 22269
rect 16665 22264 21791 22266
rect 16665 22208 16670 22264
rect 16726 22208 21730 22264
rect 21786 22208 21791 22264
rect 16665 22206 21791 22208
rect 16665 22203 16731 22206
rect 21725 22203 21791 22206
rect 22277 22266 22343 22269
rect 25037 22266 25103 22269
rect 25454 22266 25514 22614
rect 25773 22672 26667 22674
rect 25773 22616 25778 22672
rect 25834 22616 26606 22672
rect 26662 22616 26667 22672
rect 25773 22614 26667 22616
rect 25773 22611 25839 22614
rect 26601 22611 26667 22614
rect 26877 22674 26943 22677
rect 27613 22674 27679 22677
rect 31017 22674 31083 22677
rect 26877 22672 31083 22674
rect 26877 22616 26882 22672
rect 26938 22616 27618 22672
rect 27674 22616 31022 22672
rect 31078 22616 31083 22672
rect 26877 22614 31083 22616
rect 26877 22611 26943 22614
rect 27613 22611 27679 22614
rect 31017 22611 31083 22614
rect 34145 22674 34211 22677
rect 46749 22674 46815 22677
rect 48454 22674 48514 22886
rect 50200 22856 51000 22886
rect 34145 22672 45570 22674
rect 34145 22616 34150 22672
rect 34206 22616 45570 22672
rect 34145 22614 45570 22616
rect 34145 22611 34211 22614
rect 25957 22538 26023 22541
rect 33133 22538 33199 22541
rect 25957 22536 33199 22538
rect 25957 22480 25962 22536
rect 26018 22480 33138 22536
rect 33194 22480 33199 22536
rect 25957 22478 33199 22480
rect 45510 22538 45570 22614
rect 46749 22672 48514 22674
rect 46749 22616 46754 22672
rect 46810 22616 48514 22672
rect 46749 22614 48514 22616
rect 46749 22611 46815 22614
rect 49233 22538 49299 22541
rect 45510 22536 49299 22538
rect 45510 22480 49238 22536
rect 49294 22480 49299 22536
rect 45510 22478 49299 22480
rect 25957 22475 26023 22478
rect 33133 22475 33199 22478
rect 49233 22475 49299 22478
rect 25773 22402 25839 22405
rect 25998 22402 26004 22404
rect 25773 22400 26004 22402
rect 25773 22344 25778 22400
rect 25834 22344 26004 22400
rect 25773 22342 26004 22344
rect 25773 22339 25839 22342
rect 25998 22340 26004 22342
rect 26068 22340 26074 22404
rect 27705 22402 27771 22405
rect 31753 22402 31819 22405
rect 27705 22400 31819 22402
rect 27705 22344 27710 22400
rect 27766 22344 31758 22400
rect 31814 22344 31819 22400
rect 27705 22342 31819 22344
rect 27705 22339 27771 22342
rect 31753 22339 31819 22342
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 28758 22266 28764 22268
rect 22277 22264 22754 22266
rect 22277 22208 22282 22264
rect 22338 22208 22754 22264
rect 22277 22206 22754 22208
rect 22277 22203 22343 22206
rect 3601 22130 3667 22133
rect 9765 22130 9831 22133
rect 3601 22128 9831 22130
rect 3601 22072 3606 22128
rect 3662 22072 9770 22128
rect 9826 22072 9831 22128
rect 3601 22070 9831 22072
rect 3601 22067 3667 22070
rect 9765 22067 9831 22070
rect 10501 22130 10567 22133
rect 13721 22130 13787 22133
rect 10501 22128 13787 22130
rect 10501 22072 10506 22128
rect 10562 22072 13726 22128
rect 13782 22072 13787 22128
rect 10501 22070 13787 22072
rect 10501 22067 10567 22070
rect 13721 22067 13787 22070
rect 14917 22130 14983 22133
rect 16614 22130 16620 22132
rect 14917 22128 16620 22130
rect 14917 22072 14922 22128
rect 14978 22072 16620 22128
rect 14917 22070 16620 22072
rect 14917 22067 14983 22070
rect 16614 22068 16620 22070
rect 16684 22068 16690 22132
rect 16757 22130 16823 22133
rect 18689 22130 18755 22133
rect 16757 22128 18755 22130
rect 16757 22072 16762 22128
rect 16818 22072 18694 22128
rect 18750 22072 18755 22128
rect 16757 22070 18755 22072
rect 16757 22067 16823 22070
rect 18689 22067 18755 22070
rect 19425 22130 19491 22133
rect 19742 22130 19748 22132
rect 19425 22128 19748 22130
rect 19425 22072 19430 22128
rect 19486 22072 19748 22128
rect 19425 22070 19748 22072
rect 19425 22067 19491 22070
rect 19742 22068 19748 22070
rect 19812 22068 19818 22132
rect 19885 22130 19951 22133
rect 21357 22130 21423 22133
rect 19885 22128 21423 22130
rect 19885 22072 19890 22128
rect 19946 22072 21362 22128
rect 21418 22072 21423 22128
rect 19885 22070 21423 22072
rect 19885 22067 19951 22070
rect 21357 22067 21423 22070
rect 21633 22130 21699 22133
rect 22461 22130 22527 22133
rect 21633 22128 22527 22130
rect 21633 22072 21638 22128
rect 21694 22072 22466 22128
rect 22522 22072 22527 22128
rect 21633 22070 22527 22072
rect 22694 22130 22754 22206
rect 25037 22264 25330 22266
rect 25037 22208 25042 22264
rect 25098 22208 25330 22264
rect 25037 22206 25330 22208
rect 25454 22206 28764 22266
rect 25037 22203 25103 22206
rect 25129 22130 25195 22133
rect 22694 22128 25195 22130
rect 22694 22072 25134 22128
rect 25190 22072 25195 22128
rect 22694 22070 25195 22072
rect 25270 22130 25330 22206
rect 28758 22204 28764 22206
rect 28828 22204 28834 22268
rect 28901 22266 28967 22269
rect 30557 22266 30623 22269
rect 28901 22264 30623 22266
rect 28901 22208 28906 22264
rect 28962 22208 30562 22264
rect 30618 22208 30623 22264
rect 28901 22206 30623 22208
rect 28901 22203 28967 22206
rect 30557 22203 30623 22206
rect 26233 22130 26299 22133
rect 26417 22130 26483 22133
rect 25270 22070 26112 22130
rect 21633 22067 21699 22070
rect 22461 22067 22527 22070
rect 25129 22067 25195 22070
rect 0 21994 800 22024
rect 26052 21997 26112 22070
rect 26233 22128 26483 22130
rect 26233 22072 26238 22128
rect 26294 22072 26422 22128
rect 26478 22072 26483 22128
rect 26233 22070 26483 22072
rect 26233 22067 26299 22070
rect 26417 22067 26483 22070
rect 26601 22130 26667 22133
rect 28901 22130 28967 22133
rect 26601 22128 28967 22130
rect 26601 22072 26606 22128
rect 26662 22072 28906 22128
rect 28962 22072 28967 22128
rect 26601 22070 28967 22072
rect 26601 22067 26667 22070
rect 28901 22067 28967 22070
rect 30005 22130 30071 22133
rect 30373 22130 30439 22133
rect 30005 22128 30439 22130
rect 30005 22072 30010 22128
rect 30066 22072 30378 22128
rect 30434 22072 30439 22128
rect 30005 22070 30439 22072
rect 30005 22067 30071 22070
rect 30373 22067 30439 22070
rect 3325 21994 3391 21997
rect 0 21992 3391 21994
rect 0 21936 3330 21992
rect 3386 21936 3391 21992
rect 0 21934 3391 21936
rect 0 21904 800 21934
rect 3325 21931 3391 21934
rect 9029 21994 9095 21997
rect 14917 21994 14983 21997
rect 9029 21992 14983 21994
rect 9029 21936 9034 21992
rect 9090 21936 14922 21992
rect 14978 21936 14983 21992
rect 9029 21934 14983 21936
rect 9029 21931 9095 21934
rect 14917 21931 14983 21934
rect 15193 21994 15259 21997
rect 16573 21994 16639 21997
rect 20345 21994 20411 21997
rect 15193 21992 16498 21994
rect 15193 21936 15198 21992
rect 15254 21936 16498 21992
rect 15193 21934 16498 21936
rect 15193 21931 15259 21934
rect 8753 21858 8819 21861
rect 15377 21858 15443 21861
rect 8753 21856 15443 21858
rect 8753 21800 8758 21856
rect 8814 21800 15382 21856
rect 15438 21800 15443 21856
rect 8753 21798 15443 21800
rect 16438 21858 16498 21934
rect 16573 21992 20411 21994
rect 16573 21936 16578 21992
rect 16634 21936 20350 21992
rect 20406 21936 20411 21992
rect 16573 21934 20411 21936
rect 16573 21931 16639 21934
rect 20345 21931 20411 21934
rect 20478 21932 20484 21996
rect 20548 21994 20554 21996
rect 25773 21994 25839 21997
rect 20548 21992 25839 21994
rect 20548 21936 25778 21992
rect 25834 21936 25839 21992
rect 20548 21934 25839 21936
rect 20548 21932 20554 21934
rect 25773 21931 25839 21934
rect 26049 21992 26115 21997
rect 38745 21994 38811 21997
rect 26049 21936 26054 21992
rect 26110 21936 26115 21992
rect 26049 21931 26115 21936
rect 26926 21992 38811 21994
rect 26926 21936 38750 21992
rect 38806 21936 38811 21992
rect 26926 21934 38811 21936
rect 17401 21858 17467 21861
rect 16438 21856 17467 21858
rect 16438 21800 17406 21856
rect 17462 21800 17467 21856
rect 16438 21798 17467 21800
rect 8753 21795 8819 21798
rect 15377 21795 15443 21798
rect 17401 21795 17467 21798
rect 19333 21860 19399 21861
rect 19333 21856 19380 21860
rect 19444 21858 19450 21860
rect 21449 21858 21515 21861
rect 26926 21858 26986 21934
rect 38745 21931 38811 21934
rect 46565 21994 46631 21997
rect 50200 21994 51000 22024
rect 46565 21992 51000 21994
rect 46565 21936 46570 21992
rect 46626 21936 51000 21992
rect 46565 21934 51000 21936
rect 46565 21931 46631 21934
rect 50200 21904 51000 21934
rect 19333 21800 19338 21856
rect 19333 21796 19380 21800
rect 19444 21798 19490 21858
rect 21449 21856 26986 21858
rect 21449 21800 21454 21856
rect 21510 21800 26986 21856
rect 21449 21798 26986 21800
rect 28349 21858 28415 21861
rect 29494 21858 29500 21860
rect 28349 21856 29500 21858
rect 28349 21800 28354 21856
rect 28410 21800 29500 21856
rect 28349 21798 29500 21800
rect 19444 21796 19450 21798
rect 19333 21795 19399 21796
rect 21449 21795 21515 21798
rect 28349 21795 28415 21798
rect 29494 21796 29500 21798
rect 29564 21858 29570 21860
rect 29564 21798 31770 21858
rect 29564 21796 29570 21798
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 8702 21660 8708 21724
rect 8772 21722 8778 21724
rect 9305 21722 9371 21725
rect 8772 21720 9371 21722
rect 8772 21664 9310 21720
rect 9366 21664 9371 21720
rect 8772 21662 9371 21664
rect 8772 21660 8778 21662
rect 9305 21659 9371 21662
rect 11329 21722 11395 21725
rect 15929 21722 15995 21725
rect 11329 21720 15995 21722
rect 11329 21664 11334 21720
rect 11390 21664 15934 21720
rect 15990 21664 15995 21720
rect 11329 21662 15995 21664
rect 11329 21659 11395 21662
rect 15929 21659 15995 21662
rect 16297 21722 16363 21725
rect 17534 21722 17540 21724
rect 16297 21720 17540 21722
rect 16297 21664 16302 21720
rect 16358 21664 17540 21720
rect 16297 21662 17540 21664
rect 16297 21659 16363 21662
rect 17534 21660 17540 21662
rect 17604 21660 17610 21724
rect 18689 21722 18755 21725
rect 24485 21722 24551 21725
rect 18689 21720 24551 21722
rect 18689 21664 18694 21720
rect 18750 21664 24490 21720
rect 24546 21664 24551 21720
rect 18689 21662 24551 21664
rect 18689 21659 18755 21662
rect 24485 21659 24551 21662
rect 25773 21722 25839 21725
rect 27705 21722 27771 21725
rect 25773 21720 27771 21722
rect 25773 21664 25778 21720
rect 25834 21664 27710 21720
rect 27766 21664 27771 21720
rect 25773 21662 27771 21664
rect 25773 21659 25839 21662
rect 27705 21659 27771 21662
rect 28349 21722 28415 21725
rect 28901 21722 28967 21725
rect 28349 21720 28967 21722
rect 28349 21664 28354 21720
rect 28410 21664 28906 21720
rect 28962 21664 28967 21720
rect 28349 21662 28967 21664
rect 31710 21722 31770 21798
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 34329 21722 34395 21725
rect 31710 21720 34395 21722
rect 31710 21664 34334 21720
rect 34390 21664 34395 21720
rect 31710 21662 34395 21664
rect 28349 21659 28415 21662
rect 28901 21659 28967 21662
rect 34329 21659 34395 21662
rect 0 21586 800 21616
rect 2681 21586 2747 21589
rect 0 21584 2747 21586
rect 0 21528 2686 21584
rect 2742 21528 2747 21584
rect 0 21526 2747 21528
rect 0 21496 800 21526
rect 2681 21523 2747 21526
rect 3550 21524 3556 21588
rect 3620 21586 3626 21588
rect 3969 21586 4035 21589
rect 3620 21584 4035 21586
rect 3620 21528 3974 21584
rect 4030 21528 4035 21584
rect 3620 21526 4035 21528
rect 3620 21524 3626 21526
rect 3969 21523 4035 21526
rect 5809 21586 5875 21589
rect 14958 21586 14964 21588
rect 5809 21584 14964 21586
rect 5809 21528 5814 21584
rect 5870 21528 14964 21584
rect 5809 21526 14964 21528
rect 5809 21523 5875 21526
rect 14958 21524 14964 21526
rect 15028 21524 15034 21588
rect 15101 21586 15167 21589
rect 18873 21586 18939 21589
rect 15101 21584 18939 21586
rect 15101 21528 15106 21584
rect 15162 21528 18878 21584
rect 18934 21528 18939 21584
rect 15101 21526 18939 21528
rect 15101 21523 15167 21526
rect 18873 21523 18939 21526
rect 21081 21586 21147 21589
rect 26969 21586 27035 21589
rect 21081 21584 27035 21586
rect 21081 21528 21086 21584
rect 21142 21528 26974 21584
rect 27030 21528 27035 21584
rect 21081 21526 27035 21528
rect 21081 21523 21147 21526
rect 26969 21523 27035 21526
rect 27337 21586 27403 21589
rect 29177 21586 29243 21589
rect 27337 21584 29243 21586
rect 27337 21528 27342 21584
rect 27398 21528 29182 21584
rect 29238 21528 29243 21584
rect 27337 21526 29243 21528
rect 27337 21523 27403 21526
rect 29177 21523 29243 21526
rect 31109 21586 31175 21589
rect 44081 21586 44147 21589
rect 31109 21584 44147 21586
rect 31109 21528 31114 21584
rect 31170 21528 44086 21584
rect 44142 21528 44147 21584
rect 31109 21526 44147 21528
rect 31109 21523 31175 21526
rect 44081 21523 44147 21526
rect 9581 21450 9647 21453
rect 12249 21452 12315 21453
rect 12198 21450 12204 21452
rect 9581 21448 12204 21450
rect 12268 21448 12315 21452
rect 17125 21452 17191 21453
rect 17125 21450 17172 21452
rect 9581 21392 9586 21448
rect 9642 21392 12204 21448
rect 12310 21392 12315 21448
rect 9581 21390 12204 21392
rect 9581 21387 9647 21390
rect 12198 21388 12204 21390
rect 12268 21388 12315 21392
rect 17080 21448 17172 21450
rect 17080 21392 17130 21448
rect 17080 21390 17172 21392
rect 12249 21387 12315 21388
rect 17125 21388 17172 21390
rect 17236 21388 17242 21452
rect 17953 21450 18019 21453
rect 19149 21450 19215 21453
rect 25129 21450 25195 21453
rect 34513 21450 34579 21453
rect 17953 21448 24962 21450
rect 17953 21392 17958 21448
rect 18014 21392 19154 21448
rect 19210 21392 24962 21448
rect 17953 21390 24962 21392
rect 17125 21387 17191 21388
rect 17953 21387 18019 21390
rect 19149 21387 19215 21390
rect 3325 21314 3391 21317
rect 12525 21314 12591 21317
rect 3325 21312 12591 21314
rect 3325 21256 3330 21312
rect 3386 21256 12530 21312
rect 12586 21256 12591 21312
rect 3325 21254 12591 21256
rect 3325 21251 3391 21254
rect 12525 21251 12591 21254
rect 16297 21314 16363 21317
rect 21449 21314 21515 21317
rect 22737 21314 22803 21317
rect 16297 21312 21515 21314
rect 16297 21256 16302 21312
rect 16358 21256 21454 21312
rect 21510 21256 21515 21312
rect 16297 21254 21515 21256
rect 16297 21251 16363 21254
rect 21449 21251 21515 21254
rect 21820 21312 22803 21314
rect 21820 21256 22742 21312
rect 22798 21256 22803 21312
rect 21820 21254 22803 21256
rect 24902 21314 24962 21390
rect 25129 21448 34579 21450
rect 25129 21392 25134 21448
rect 25190 21392 34518 21448
rect 34574 21392 34579 21448
rect 25129 21390 34579 21392
rect 25129 21387 25195 21390
rect 34513 21387 34579 21390
rect 31569 21314 31635 21317
rect 24902 21312 31635 21314
rect 24902 21256 31574 21312
rect 31630 21256 31635 21312
rect 24902 21254 31635 21256
rect 2946 21248 3262 21249
rect 0 21178 800 21208
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 2221 21178 2287 21181
rect 6913 21178 6979 21181
rect 0 21176 2287 21178
rect 0 21120 2226 21176
rect 2282 21120 2287 21176
rect 0 21118 2287 21120
rect 0 21088 800 21118
rect 2221 21115 2287 21118
rect 3926 21176 6979 21178
rect 3926 21120 6918 21176
rect 6974 21120 6979 21176
rect 3926 21118 6979 21120
rect 974 20980 980 21044
rect 1044 21042 1050 21044
rect 3926 21042 3986 21118
rect 6913 21115 6979 21118
rect 14958 21116 14964 21180
rect 15028 21178 15034 21180
rect 17125 21178 17191 21181
rect 19149 21180 19215 21181
rect 15028 21176 17191 21178
rect 15028 21120 17130 21176
rect 17186 21120 17191 21176
rect 15028 21118 17191 21120
rect 15028 21116 15034 21118
rect 17125 21115 17191 21118
rect 17718 21116 17724 21180
rect 17788 21178 17794 21180
rect 19006 21178 19012 21180
rect 17788 21118 19012 21178
rect 17788 21116 17794 21118
rect 19006 21116 19012 21118
rect 19076 21116 19082 21180
rect 19149 21176 19196 21180
rect 19260 21178 19266 21180
rect 21081 21178 21147 21181
rect 21820 21178 21880 21254
rect 22737 21251 22803 21254
rect 31569 21251 31635 21254
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 42946 21183 43262 21184
rect 19149 21120 19154 21176
rect 19149 21116 19196 21120
rect 19260 21118 19306 21178
rect 21081 21176 21880 21178
rect 21081 21120 21086 21176
rect 21142 21120 21880 21176
rect 21081 21118 21880 21120
rect 23473 21178 23539 21181
rect 24669 21178 24735 21181
rect 23473 21176 24735 21178
rect 23473 21120 23478 21176
rect 23534 21120 24674 21176
rect 24730 21120 24735 21176
rect 23473 21118 24735 21120
rect 19260 21116 19266 21118
rect 19149 21115 19215 21116
rect 21081 21115 21147 21118
rect 23473 21115 23539 21118
rect 24669 21115 24735 21118
rect 24853 21178 24919 21181
rect 27061 21178 27127 21181
rect 30005 21178 30071 21181
rect 24853 21176 27127 21178
rect 24853 21120 24858 21176
rect 24914 21120 27066 21176
rect 27122 21120 27127 21176
rect 24853 21118 27127 21120
rect 24853 21115 24919 21118
rect 27061 21115 27127 21118
rect 27294 21176 30071 21178
rect 27294 21120 30010 21176
rect 30066 21120 30071 21176
rect 27294 21118 30071 21120
rect 1044 20982 3986 21042
rect 4061 21042 4127 21045
rect 13854 21042 13860 21044
rect 4061 21040 13860 21042
rect 4061 20984 4066 21040
rect 4122 20984 13860 21040
rect 4061 20982 13860 20984
rect 1044 20980 1050 20982
rect 4061 20979 4127 20982
rect 13854 20980 13860 20982
rect 13924 20980 13930 21044
rect 15101 21042 15167 21045
rect 26182 21042 26188 21044
rect 15101 21040 26188 21042
rect 15101 20984 15106 21040
rect 15162 20984 26188 21040
rect 15101 20982 26188 20984
rect 15101 20979 15167 20982
rect 26182 20980 26188 20982
rect 26252 20980 26258 21044
rect 26969 21042 27035 21045
rect 27294 21042 27354 21118
rect 30005 21115 30071 21118
rect 26969 21040 27354 21042
rect 26969 20984 26974 21040
rect 27030 20984 27354 21040
rect 26969 20982 27354 20984
rect 27797 21042 27863 21045
rect 36077 21042 36143 21045
rect 27797 21040 36143 21042
rect 27797 20984 27802 21040
rect 27858 20984 36082 21040
rect 36138 20984 36143 21040
rect 27797 20982 36143 20984
rect 26969 20979 27035 20982
rect 27797 20979 27863 20982
rect 36077 20979 36143 20982
rect 49141 21042 49207 21045
rect 50200 21042 51000 21072
rect 49141 21040 51000 21042
rect 49141 20984 49146 21040
rect 49202 20984 51000 21040
rect 49141 20982 51000 20984
rect 49141 20979 49207 20982
rect 50200 20952 51000 20982
rect 1669 20908 1735 20909
rect 1669 20904 1716 20908
rect 1780 20906 1786 20908
rect 1669 20848 1674 20904
rect 1669 20844 1716 20848
rect 1780 20846 1826 20906
rect 1780 20844 1786 20846
rect 5390 20844 5396 20908
rect 5460 20906 5466 20908
rect 8017 20906 8083 20909
rect 5460 20904 8083 20906
rect 5460 20848 8022 20904
rect 8078 20848 8083 20904
rect 5460 20846 8083 20848
rect 5460 20844 5466 20846
rect 1669 20843 1735 20844
rect 8017 20843 8083 20846
rect 11830 20844 11836 20908
rect 11900 20906 11906 20908
rect 16757 20906 16823 20909
rect 11900 20904 16823 20906
rect 11900 20848 16762 20904
rect 16818 20848 16823 20904
rect 11900 20846 16823 20848
rect 11900 20844 11906 20846
rect 16757 20843 16823 20846
rect 17217 20906 17283 20909
rect 19374 20906 19380 20908
rect 17217 20904 19380 20906
rect 17217 20848 17222 20904
rect 17278 20848 19380 20904
rect 17217 20846 19380 20848
rect 17217 20843 17283 20846
rect 19374 20844 19380 20846
rect 19444 20844 19450 20908
rect 19517 20906 19583 20909
rect 21817 20906 21883 20909
rect 23749 20906 23815 20909
rect 19517 20904 21883 20906
rect 19517 20848 19522 20904
rect 19578 20848 21822 20904
rect 21878 20848 21883 20904
rect 19517 20846 21883 20848
rect 19517 20843 19583 20846
rect 21817 20843 21883 20846
rect 21958 20904 23815 20906
rect 21958 20848 23754 20904
rect 23810 20848 23815 20904
rect 21958 20846 23815 20848
rect 0 20770 800 20800
rect 3785 20770 3851 20773
rect 0 20768 3851 20770
rect 0 20712 3790 20768
rect 3846 20712 3851 20768
rect 0 20710 3851 20712
rect 0 20680 800 20710
rect 3785 20707 3851 20710
rect 5625 20770 5691 20773
rect 6126 20770 6132 20772
rect 5625 20768 6132 20770
rect 5625 20712 5630 20768
rect 5686 20712 6132 20768
rect 5625 20710 6132 20712
rect 5625 20707 5691 20710
rect 6126 20708 6132 20710
rect 6196 20708 6202 20772
rect 6545 20770 6611 20773
rect 6862 20770 6868 20772
rect 6545 20768 6868 20770
rect 6545 20712 6550 20768
rect 6606 20712 6868 20768
rect 6545 20710 6868 20712
rect 6545 20707 6611 20710
rect 6862 20708 6868 20710
rect 6932 20708 6938 20772
rect 9673 20770 9739 20773
rect 10910 20770 10916 20772
rect 9673 20768 10916 20770
rect 9673 20712 9678 20768
rect 9734 20712 10916 20768
rect 9673 20710 10916 20712
rect 9673 20707 9739 20710
rect 10910 20708 10916 20710
rect 10980 20708 10986 20772
rect 11329 20770 11395 20773
rect 17401 20770 17467 20773
rect 18413 20772 18479 20773
rect 18413 20770 18460 20772
rect 11329 20768 17467 20770
rect 11329 20712 11334 20768
rect 11390 20712 17406 20768
rect 17462 20712 17467 20768
rect 11329 20710 17467 20712
rect 18368 20768 18460 20770
rect 18368 20712 18418 20768
rect 18368 20710 18460 20712
rect 11329 20707 11395 20710
rect 17401 20707 17467 20710
rect 18413 20708 18460 20710
rect 18524 20708 18530 20772
rect 19609 20770 19675 20773
rect 21958 20770 22018 20846
rect 23749 20843 23815 20846
rect 26417 20906 26483 20909
rect 29913 20906 29979 20909
rect 26417 20904 29979 20906
rect 26417 20848 26422 20904
rect 26478 20848 29918 20904
rect 29974 20848 29979 20904
rect 26417 20846 29979 20848
rect 26417 20843 26483 20846
rect 29913 20843 29979 20846
rect 31661 20906 31727 20909
rect 43345 20906 43411 20909
rect 31661 20904 43411 20906
rect 31661 20848 31666 20904
rect 31722 20848 43350 20904
rect 43406 20848 43411 20904
rect 31661 20846 43411 20848
rect 31661 20843 31727 20846
rect 43345 20843 43411 20846
rect 19609 20768 22018 20770
rect 19609 20712 19614 20768
rect 19670 20712 22018 20768
rect 19609 20710 22018 20712
rect 22185 20770 22251 20773
rect 22185 20768 22386 20770
rect 22185 20712 22190 20768
rect 22246 20712 22386 20768
rect 22185 20710 22386 20712
rect 18413 20707 18479 20708
rect 19609 20707 19675 20710
rect 22185 20707 22251 20710
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 2262 20572 2268 20636
rect 2332 20634 2338 20636
rect 6453 20634 6519 20637
rect 2332 20632 6519 20634
rect 2332 20576 6458 20632
rect 6514 20576 6519 20632
rect 2332 20574 6519 20576
rect 2332 20572 2338 20574
rect 6453 20571 6519 20574
rect 9029 20634 9095 20637
rect 14825 20634 14891 20637
rect 16573 20634 16639 20637
rect 9029 20632 16639 20634
rect 9029 20576 9034 20632
rect 9090 20576 14830 20632
rect 14886 20576 16578 20632
rect 16634 20576 16639 20632
rect 9029 20574 16639 20576
rect 9029 20571 9095 20574
rect 14825 20571 14891 20574
rect 16573 20571 16639 20574
rect 17534 20572 17540 20636
rect 17604 20634 17610 20636
rect 17677 20634 17743 20637
rect 19558 20634 19564 20636
rect 17604 20632 17743 20634
rect 17604 20576 17682 20632
rect 17738 20576 17743 20632
rect 17604 20574 17743 20576
rect 17604 20572 17610 20574
rect 17677 20571 17743 20574
rect 18462 20574 19564 20634
rect 5533 20498 5599 20501
rect 11789 20498 11855 20501
rect 5533 20496 11855 20498
rect 5533 20440 5538 20496
rect 5594 20440 11794 20496
rect 11850 20440 11855 20496
rect 5533 20438 11855 20440
rect 5533 20435 5599 20438
rect 11789 20435 11855 20438
rect 14365 20498 14431 20501
rect 16113 20498 16179 20501
rect 14365 20496 16179 20498
rect 14365 20440 14370 20496
rect 14426 20440 16118 20496
rect 16174 20440 16179 20496
rect 14365 20438 16179 20440
rect 14365 20435 14431 20438
rect 16113 20435 16179 20438
rect 16614 20436 16620 20500
rect 16684 20498 16690 20500
rect 18462 20498 18522 20574
rect 19558 20572 19564 20574
rect 19628 20572 19634 20636
rect 19742 20572 19748 20636
rect 19812 20634 19818 20636
rect 21541 20634 21607 20637
rect 19812 20632 21607 20634
rect 19812 20576 21546 20632
rect 21602 20576 21607 20632
rect 19812 20574 21607 20576
rect 19812 20572 19818 20574
rect 21541 20571 21607 20574
rect 21817 20634 21883 20637
rect 22326 20634 22386 20710
rect 24526 20708 24532 20772
rect 24596 20770 24602 20772
rect 24669 20770 24735 20773
rect 24596 20768 24735 20770
rect 24596 20712 24674 20768
rect 24730 20712 24735 20768
rect 24596 20710 24735 20712
rect 24596 20708 24602 20710
rect 24669 20707 24735 20710
rect 25681 20770 25747 20773
rect 25814 20770 25820 20772
rect 25681 20768 25820 20770
rect 25681 20712 25686 20768
rect 25742 20712 25820 20768
rect 25681 20710 25820 20712
rect 25681 20707 25747 20710
rect 25814 20708 25820 20710
rect 25884 20708 25890 20772
rect 29453 20770 29519 20773
rect 30741 20770 30807 20773
rect 29453 20768 30807 20770
rect 29453 20712 29458 20768
rect 29514 20712 30746 20768
rect 30802 20712 30807 20768
rect 29453 20710 30807 20712
rect 29453 20707 29519 20710
rect 30741 20707 30807 20710
rect 31109 20770 31175 20773
rect 31937 20770 32003 20773
rect 31109 20768 32003 20770
rect 31109 20712 31114 20768
rect 31170 20712 31942 20768
rect 31998 20712 32003 20768
rect 31109 20710 32003 20712
rect 31109 20707 31175 20710
rect 31937 20707 32003 20710
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 23565 20634 23631 20637
rect 25589 20634 25655 20637
rect 21817 20632 22248 20634
rect 21817 20576 21822 20632
rect 21878 20576 22248 20632
rect 21817 20574 22248 20576
rect 22326 20632 23631 20634
rect 22326 20576 23570 20632
rect 23626 20576 23631 20632
rect 22326 20574 23631 20576
rect 21817 20571 21883 20574
rect 16684 20438 18522 20498
rect 18965 20498 19031 20501
rect 21950 20498 21956 20500
rect 18965 20496 21956 20498
rect 18965 20440 18970 20496
rect 19026 20440 21956 20496
rect 18965 20438 21956 20440
rect 16684 20436 16690 20438
rect 18965 20435 19031 20438
rect 21950 20436 21956 20438
rect 22020 20436 22026 20500
rect 0 20362 800 20392
rect 1485 20362 1551 20365
rect 0 20360 1551 20362
rect 0 20304 1490 20360
rect 1546 20304 1551 20360
rect 0 20302 1551 20304
rect 0 20272 800 20302
rect 1485 20299 1551 20302
rect 5901 20362 5967 20365
rect 12985 20362 13051 20365
rect 5901 20360 13051 20362
rect 5901 20304 5906 20360
rect 5962 20304 12990 20360
rect 13046 20304 13051 20360
rect 5901 20302 13051 20304
rect 5901 20299 5967 20302
rect 12985 20299 13051 20302
rect 13813 20362 13879 20365
rect 15561 20362 15627 20365
rect 21081 20362 21147 20365
rect 13813 20360 15440 20362
rect 13813 20304 13818 20360
rect 13874 20304 15440 20360
rect 13813 20302 15440 20304
rect 13813 20299 13879 20302
rect 3969 20226 4035 20229
rect 12709 20226 12775 20229
rect 3969 20224 12775 20226
rect 3969 20168 3974 20224
rect 4030 20168 12714 20224
rect 12770 20168 12775 20224
rect 3969 20166 12775 20168
rect 3969 20163 4035 20166
rect 12709 20163 12775 20166
rect 13997 20226 14063 20229
rect 14825 20226 14891 20229
rect 13997 20224 14891 20226
rect 13997 20168 14002 20224
rect 14058 20168 14830 20224
rect 14886 20168 14891 20224
rect 13997 20166 14891 20168
rect 15380 20226 15440 20302
rect 15561 20360 21147 20362
rect 15561 20304 15566 20360
rect 15622 20304 21086 20360
rect 21142 20304 21147 20360
rect 15561 20302 21147 20304
rect 22188 20362 22248 20574
rect 23565 20571 23631 20574
rect 23752 20632 25655 20634
rect 23752 20576 25594 20632
rect 25650 20576 25655 20632
rect 23752 20574 25655 20576
rect 22318 20436 22324 20500
rect 22388 20498 22394 20500
rect 23752 20498 23812 20574
rect 25589 20571 25655 20574
rect 31385 20634 31451 20637
rect 33409 20634 33475 20637
rect 31385 20632 33475 20634
rect 31385 20576 31390 20632
rect 31446 20576 33414 20632
rect 33470 20576 33475 20632
rect 31385 20574 33475 20576
rect 31385 20571 31451 20574
rect 33409 20571 33475 20574
rect 22388 20438 23812 20498
rect 24485 20498 24551 20501
rect 39021 20498 39087 20501
rect 24485 20496 39087 20498
rect 24485 20440 24490 20496
rect 24546 20440 39026 20496
rect 39082 20440 39087 20496
rect 24485 20438 39087 20440
rect 22388 20436 22394 20438
rect 24485 20435 24551 20438
rect 39021 20435 39087 20438
rect 24158 20362 24164 20364
rect 22188 20302 24164 20362
rect 15561 20299 15627 20302
rect 21081 20299 21147 20302
rect 24158 20300 24164 20302
rect 24228 20300 24234 20364
rect 24301 20362 24367 20365
rect 30414 20362 30420 20364
rect 24301 20360 30420 20362
rect 24301 20304 24306 20360
rect 24362 20304 30420 20360
rect 24301 20302 30420 20304
rect 24301 20299 24367 20302
rect 30414 20300 30420 20302
rect 30484 20300 30490 20364
rect 34329 20362 34395 20365
rect 31710 20360 34395 20362
rect 31710 20304 34334 20360
rect 34390 20304 34395 20360
rect 31710 20302 34395 20304
rect 16113 20226 16179 20229
rect 16849 20226 16915 20229
rect 15380 20224 16915 20226
rect 15380 20168 16118 20224
rect 16174 20168 16854 20224
rect 16910 20168 16915 20224
rect 15380 20166 16915 20168
rect 13997 20163 14063 20166
rect 14825 20163 14891 20166
rect 16113 20163 16179 20166
rect 16849 20163 16915 20166
rect 17125 20226 17191 20229
rect 22737 20226 22803 20229
rect 17125 20224 22803 20226
rect 17125 20168 17130 20224
rect 17186 20168 22742 20224
rect 22798 20168 22803 20224
rect 17125 20166 22803 20168
rect 17125 20163 17191 20166
rect 22737 20163 22803 20166
rect 27470 20164 27476 20228
rect 27540 20226 27546 20228
rect 31710 20226 31770 20302
rect 34329 20299 34395 20302
rect 27540 20166 31770 20226
rect 27540 20164 27546 20166
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 14641 20090 14707 20093
rect 16481 20090 16547 20093
rect 14641 20088 16547 20090
rect 14641 20032 14646 20088
rect 14702 20032 16486 20088
rect 16542 20032 16547 20088
rect 14641 20030 16547 20032
rect 14641 20027 14707 20030
rect 16481 20027 16547 20030
rect 17217 20090 17283 20093
rect 17350 20090 17356 20092
rect 17217 20088 17356 20090
rect 17217 20032 17222 20088
rect 17278 20032 17356 20088
rect 17217 20030 17356 20032
rect 17217 20027 17283 20030
rect 17350 20028 17356 20030
rect 17420 20028 17426 20092
rect 17677 20090 17743 20093
rect 21449 20090 21515 20093
rect 17677 20088 21515 20090
rect 17677 20032 17682 20088
rect 17738 20032 21454 20088
rect 21510 20032 21515 20088
rect 17677 20030 21515 20032
rect 17677 20027 17743 20030
rect 21449 20027 21515 20030
rect 23749 20090 23815 20093
rect 28533 20090 28599 20093
rect 23749 20088 28599 20090
rect 23749 20032 23754 20088
rect 23810 20032 28538 20088
rect 28594 20032 28599 20088
rect 23749 20030 28599 20032
rect 23749 20027 23815 20030
rect 28533 20027 28599 20030
rect 0 19954 800 19984
rect 2773 19954 2839 19957
rect 0 19952 2839 19954
rect 0 19896 2778 19952
rect 2834 19896 2839 19952
rect 0 19894 2839 19896
rect 0 19864 800 19894
rect 2773 19891 2839 19894
rect 8385 19954 8451 19957
rect 13721 19954 13787 19957
rect 8385 19952 13787 19954
rect 8385 19896 8390 19952
rect 8446 19896 13726 19952
rect 13782 19896 13787 19952
rect 8385 19894 13787 19896
rect 8385 19891 8451 19894
rect 13721 19891 13787 19894
rect 15193 19954 15259 19957
rect 32673 19954 32739 19957
rect 15193 19952 32739 19954
rect 15193 19896 15198 19952
rect 15254 19896 32678 19952
rect 32734 19896 32739 19952
rect 15193 19894 32739 19896
rect 15193 19891 15259 19894
rect 32673 19891 32739 19894
rect 2589 19818 2655 19821
rect 10317 19818 10383 19821
rect 2589 19816 10383 19818
rect 2589 19760 2594 19816
rect 2650 19760 10322 19816
rect 10378 19760 10383 19816
rect 2589 19758 10383 19760
rect 2589 19755 2655 19758
rect 10317 19755 10383 19758
rect 12709 19818 12775 19821
rect 13813 19818 13879 19821
rect 12709 19816 13879 19818
rect 12709 19760 12714 19816
rect 12770 19760 13818 19816
rect 13874 19760 13879 19816
rect 12709 19758 13879 19760
rect 12709 19755 12775 19758
rect 13813 19755 13879 19758
rect 14273 19818 14339 19821
rect 28993 19818 29059 19821
rect 14273 19816 17464 19818
rect 14273 19760 14278 19816
rect 14334 19784 17464 19816
rect 17910 19816 29059 19818
rect 17910 19784 28998 19816
rect 14334 19760 28998 19784
rect 29054 19760 29059 19816
rect 14273 19758 29059 19760
rect 14273 19755 14339 19758
rect 6821 19682 6887 19685
rect 7557 19682 7623 19685
rect 6821 19680 7623 19682
rect 6821 19624 6826 19680
rect 6882 19624 7562 19680
rect 7618 19624 7623 19680
rect 6821 19622 7623 19624
rect 6821 19619 6887 19622
rect 7557 19619 7623 19622
rect 7946 19616 8262 19617
rect 0 19546 800 19576
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 2037 19546 2103 19549
rect 0 19544 2103 19546
rect 0 19488 2042 19544
rect 2098 19488 2103 19544
rect 0 19486 2103 19488
rect 0 19456 800 19486
rect 2037 19483 2103 19486
rect 11605 19546 11671 19549
rect 13816 19546 13876 19755
rect 17404 19724 17970 19758
rect 28993 19755 29059 19758
rect 30373 19818 30439 19821
rect 44725 19818 44791 19821
rect 30373 19816 44791 19818
rect 30373 19760 30378 19816
rect 30434 19760 44730 19816
rect 44786 19760 44791 19816
rect 30373 19758 44791 19760
rect 30373 19755 30439 19758
rect 44725 19755 44791 19758
rect 14641 19682 14707 19685
rect 14774 19682 14780 19684
rect 14641 19680 14780 19682
rect 14641 19624 14646 19680
rect 14702 19624 14780 19680
rect 14641 19622 14780 19624
rect 14641 19619 14707 19622
rect 14774 19620 14780 19622
rect 14844 19620 14850 19684
rect 15285 19682 15351 19685
rect 16849 19682 16915 19685
rect 15285 19680 16915 19682
rect 15285 19624 15290 19680
rect 15346 19624 16854 19680
rect 16910 19624 16915 19680
rect 15285 19622 16915 19624
rect 15285 19619 15351 19622
rect 16849 19619 16915 19622
rect 18505 19682 18571 19685
rect 19742 19682 19748 19684
rect 18505 19680 19748 19682
rect 18505 19624 18510 19680
rect 18566 19624 19748 19680
rect 18505 19622 19748 19624
rect 18505 19619 18571 19622
rect 19742 19620 19748 19622
rect 19812 19620 19818 19684
rect 20621 19682 20687 19685
rect 26693 19682 26759 19685
rect 20621 19680 26759 19682
rect 20621 19624 20626 19680
rect 20682 19624 26698 19680
rect 26754 19624 26759 19680
rect 20621 19622 26759 19624
rect 20621 19619 20687 19622
rect 26693 19619 26759 19622
rect 30189 19682 30255 19685
rect 36721 19682 36787 19685
rect 30189 19680 36787 19682
rect 30189 19624 30194 19680
rect 30250 19624 36726 19680
rect 36782 19624 36787 19680
rect 30189 19622 36787 19624
rect 30189 19619 30255 19622
rect 36721 19619 36787 19622
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 16297 19546 16363 19549
rect 11605 19544 13738 19546
rect 11605 19488 11610 19544
rect 11666 19488 13738 19544
rect 11605 19486 13738 19488
rect 13816 19544 16363 19546
rect 13816 19488 16302 19544
rect 16358 19488 16363 19544
rect 13816 19486 16363 19488
rect 11605 19483 11671 19486
rect 9489 19410 9555 19413
rect 9806 19410 9812 19412
rect 9489 19408 9812 19410
rect 9489 19352 9494 19408
rect 9550 19352 9812 19408
rect 9489 19350 9812 19352
rect 9489 19347 9555 19350
rect 9806 19348 9812 19350
rect 9876 19348 9882 19412
rect 13678 19410 13738 19486
rect 16297 19483 16363 19486
rect 16941 19548 17007 19549
rect 16941 19544 16988 19548
rect 17052 19546 17058 19548
rect 17493 19546 17559 19549
rect 17769 19546 17835 19549
rect 16941 19488 16946 19544
rect 16941 19484 16988 19488
rect 17052 19486 17098 19546
rect 17493 19544 17835 19546
rect 17493 19488 17498 19544
rect 17554 19488 17774 19544
rect 17830 19488 17835 19544
rect 17493 19486 17835 19488
rect 17052 19484 17058 19486
rect 16941 19483 17007 19484
rect 17493 19483 17559 19486
rect 17769 19483 17835 19486
rect 18597 19546 18663 19549
rect 21766 19546 21772 19548
rect 18597 19544 21772 19546
rect 18597 19488 18602 19544
rect 18658 19488 21772 19544
rect 18597 19486 21772 19488
rect 18597 19483 18663 19486
rect 21766 19484 21772 19486
rect 21836 19484 21842 19548
rect 22369 19546 22435 19549
rect 22502 19546 22508 19548
rect 22369 19544 22508 19546
rect 22369 19488 22374 19544
rect 22430 19488 22508 19544
rect 22369 19486 22508 19488
rect 22369 19483 22435 19486
rect 22502 19484 22508 19486
rect 22572 19484 22578 19548
rect 22737 19546 22803 19549
rect 28625 19548 28691 19549
rect 25630 19546 25636 19548
rect 22737 19544 25636 19546
rect 22737 19488 22742 19544
rect 22798 19488 25636 19544
rect 22737 19486 25636 19488
rect 22737 19483 22803 19486
rect 25630 19484 25636 19486
rect 25700 19484 25706 19548
rect 28574 19546 28580 19548
rect 28534 19486 28580 19546
rect 28644 19544 28691 19548
rect 28686 19488 28691 19544
rect 28574 19484 28580 19486
rect 28644 19484 28691 19488
rect 28625 19483 28691 19484
rect 28901 19546 28967 19549
rect 34053 19546 34119 19549
rect 28901 19544 34119 19546
rect 28901 19488 28906 19544
rect 28962 19488 34058 19544
rect 34114 19488 34119 19544
rect 28901 19486 34119 19488
rect 28901 19483 28967 19486
rect 34053 19483 34119 19486
rect 16481 19410 16547 19413
rect 13678 19408 16547 19410
rect 13678 19352 16486 19408
rect 16542 19352 16547 19408
rect 13678 19350 16547 19352
rect 17769 19410 17835 19413
rect 19057 19410 19123 19413
rect 17769 19408 19123 19410
rect 17769 19352 17774 19408
rect 17830 19352 19062 19408
rect 19118 19352 19123 19408
rect 17769 19350 19123 19352
rect 16481 19347 16547 19350
rect 16990 19308 17602 19350
rect 17769 19347 17835 19350
rect 19057 19347 19123 19350
rect 22645 19410 22711 19413
rect 22921 19410 22987 19413
rect 22645 19408 22987 19410
rect 22645 19352 22650 19408
rect 22706 19352 22926 19408
rect 22982 19352 22987 19408
rect 22645 19350 22987 19352
rect 22645 19347 22711 19350
rect 22921 19347 22987 19350
rect 23105 19410 23171 19413
rect 23565 19410 23631 19413
rect 32765 19410 32831 19413
rect 23105 19408 32831 19410
rect 23105 19352 23110 19408
rect 23166 19352 23570 19408
rect 23626 19352 32770 19408
rect 32826 19352 32831 19408
rect 23105 19350 32831 19352
rect 23105 19347 23171 19350
rect 23565 19347 23631 19350
rect 32765 19347 32831 19350
rect 16944 19290 17602 19308
rect 6310 19212 6316 19276
rect 6380 19274 6386 19276
rect 9673 19274 9739 19277
rect 6380 19272 9739 19274
rect 6380 19216 9678 19272
rect 9734 19216 9739 19272
rect 6380 19214 9739 19216
rect 6380 19212 6386 19214
rect 9673 19211 9739 19214
rect 10777 19274 10843 19277
rect 12617 19274 12683 19277
rect 13169 19274 13235 19277
rect 16944 19274 17050 19290
rect 10777 19272 12683 19274
rect 10777 19216 10782 19272
rect 10838 19216 12622 19272
rect 12678 19216 12683 19272
rect 10777 19214 12683 19216
rect 10777 19211 10843 19214
rect 12617 19211 12683 19214
rect 12758 19272 17050 19274
rect 12758 19216 13174 19272
rect 13230 19248 17050 19272
rect 17542 19274 17602 19290
rect 40769 19274 40835 19277
rect 17542 19272 40835 19274
rect 13230 19216 17004 19248
rect 12758 19214 17004 19216
rect 17542 19216 40774 19272
rect 40830 19216 40835 19272
rect 17542 19214 40835 19216
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 4889 19138 4955 19141
rect 8937 19138 9003 19141
rect 12758 19138 12818 19214
rect 13169 19211 13235 19214
rect 40769 19211 40835 19214
rect 4889 19136 12818 19138
rect 4889 19080 4894 19136
rect 4950 19080 8942 19136
rect 8998 19080 12818 19136
rect 4889 19078 12818 19080
rect 15653 19138 15719 19141
rect 17033 19138 17099 19141
rect 15653 19136 17099 19138
rect 15653 19080 15658 19136
rect 15714 19080 17038 19136
rect 17094 19080 17099 19136
rect 15653 19078 17099 19080
rect 4889 19075 4955 19078
rect 8937 19075 9003 19078
rect 15653 19075 15719 19078
rect 17033 19075 17099 19078
rect 17350 19076 17356 19140
rect 17420 19138 17426 19140
rect 18597 19138 18663 19141
rect 17420 19136 18663 19138
rect 17420 19080 18602 19136
rect 18658 19080 18663 19136
rect 17420 19078 18663 19080
rect 17420 19076 17426 19078
rect 18597 19075 18663 19078
rect 18822 19076 18828 19140
rect 18892 19138 18898 19140
rect 20989 19138 21055 19141
rect 18892 19136 21055 19138
rect 18892 19080 20994 19136
rect 21050 19080 21055 19136
rect 18892 19078 21055 19080
rect 18892 19076 18898 19078
rect 20989 19075 21055 19078
rect 23657 19136 23723 19141
rect 26509 19140 26575 19141
rect 26509 19138 26556 19140
rect 23657 19080 23662 19136
rect 23718 19080 23723 19136
rect 23657 19075 23723 19080
rect 26464 19136 26556 19138
rect 26464 19080 26514 19136
rect 26464 19078 26556 19080
rect 26509 19076 26556 19078
rect 26620 19076 26626 19140
rect 29085 19138 29151 19141
rect 31753 19138 31819 19141
rect 29085 19136 31819 19138
rect 29085 19080 29090 19136
rect 29146 19080 31758 19136
rect 31814 19080 31819 19136
rect 29085 19078 31819 19080
rect 26509 19075 26575 19076
rect 29085 19075 29151 19078
rect 31753 19075 31819 19078
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 4286 18940 4292 19004
rect 4356 19002 4362 19004
rect 10777 19002 10843 19005
rect 4356 19000 10843 19002
rect 4356 18944 10782 19000
rect 10838 18944 10843 19000
rect 4356 18942 10843 18944
rect 4356 18940 4362 18942
rect 10777 18939 10843 18942
rect 16113 19002 16179 19005
rect 21633 19002 21699 19005
rect 16113 19000 21699 19002
rect 16113 18944 16118 19000
rect 16174 18944 21638 19000
rect 21694 18944 21699 19000
rect 16113 18942 21699 18944
rect 23660 19002 23720 19075
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 31477 19004 31543 19005
rect 29126 19002 29132 19004
rect 23660 18942 29132 19002
rect 16113 18939 16179 18942
rect 21633 18939 21699 18942
rect 29126 18940 29132 18942
rect 29196 18940 29202 19004
rect 31477 19002 31524 19004
rect 31432 19000 31524 19002
rect 31432 18944 31482 19000
rect 31432 18942 31524 18944
rect 31477 18940 31524 18942
rect 31588 18940 31594 19004
rect 33409 19002 33475 19005
rect 34605 19002 34671 19005
rect 33409 19000 34671 19002
rect 33409 18944 33414 19000
rect 33470 18944 34610 19000
rect 34666 18944 34671 19000
rect 33409 18942 34671 18944
rect 31477 18939 31543 18940
rect 33409 18939 33475 18942
rect 34605 18939 34671 18942
rect 6126 18804 6132 18868
rect 6196 18866 6202 18868
rect 12709 18866 12775 18869
rect 14222 18866 14228 18868
rect 6196 18806 10242 18866
rect 6196 18804 6202 18806
rect 0 18730 800 18760
rect 1485 18730 1551 18733
rect 0 18728 1551 18730
rect 0 18672 1490 18728
rect 1546 18672 1551 18728
rect 0 18670 1551 18672
rect 0 18640 800 18670
rect 1485 18667 1551 18670
rect 8017 18730 8083 18733
rect 9990 18730 9996 18732
rect 8017 18728 9996 18730
rect 8017 18672 8022 18728
rect 8078 18672 9996 18728
rect 8017 18670 9996 18672
rect 8017 18667 8083 18670
rect 9990 18668 9996 18670
rect 10060 18668 10066 18732
rect 1158 18532 1164 18596
rect 1228 18594 1234 18596
rect 6085 18594 6151 18597
rect 1228 18592 6151 18594
rect 1228 18536 6090 18592
rect 6146 18536 6151 18592
rect 1228 18534 6151 18536
rect 1228 18532 1234 18534
rect 6085 18531 6151 18534
rect 9070 18532 9076 18596
rect 9140 18594 9146 18596
rect 9489 18594 9555 18597
rect 9140 18592 9555 18594
rect 9140 18536 9494 18592
rect 9550 18536 9555 18592
rect 9140 18534 9555 18536
rect 10182 18594 10242 18806
rect 12709 18864 14228 18866
rect 12709 18808 12714 18864
rect 12770 18808 14228 18864
rect 12709 18806 14228 18808
rect 12709 18803 12775 18806
rect 14222 18804 14228 18806
rect 14292 18804 14298 18868
rect 14457 18866 14523 18869
rect 16757 18866 16823 18869
rect 14457 18864 16823 18866
rect 14457 18808 14462 18864
rect 14518 18808 16762 18864
rect 16818 18808 16823 18864
rect 14457 18806 16823 18808
rect 14457 18803 14523 18806
rect 16757 18803 16823 18806
rect 17125 18866 17191 18869
rect 18045 18866 18111 18869
rect 17125 18864 18111 18866
rect 17125 18808 17130 18864
rect 17186 18808 18050 18864
rect 18106 18808 18111 18864
rect 17125 18806 18111 18808
rect 17125 18803 17191 18806
rect 18045 18803 18111 18806
rect 18229 18866 18295 18869
rect 18781 18866 18847 18869
rect 35801 18866 35867 18869
rect 18229 18864 35867 18866
rect 18229 18808 18234 18864
rect 18290 18808 18786 18864
rect 18842 18808 35806 18864
rect 35862 18808 35867 18864
rect 18229 18806 35867 18808
rect 18229 18803 18295 18806
rect 18781 18803 18847 18806
rect 35801 18803 35867 18806
rect 10593 18730 10659 18733
rect 13905 18730 13971 18733
rect 10593 18728 13971 18730
rect 10593 18672 10598 18728
rect 10654 18672 13910 18728
rect 13966 18672 13971 18728
rect 10593 18670 13971 18672
rect 10593 18667 10659 18670
rect 13905 18667 13971 18670
rect 14641 18730 14707 18733
rect 19149 18730 19215 18733
rect 20253 18730 20319 18733
rect 14641 18728 20319 18730
rect 14641 18672 14646 18728
rect 14702 18672 19154 18728
rect 19210 18672 20258 18728
rect 20314 18672 20319 18728
rect 14641 18670 20319 18672
rect 14641 18667 14707 18670
rect 19149 18667 19215 18670
rect 20253 18667 20319 18670
rect 21081 18730 21147 18733
rect 26049 18730 26115 18733
rect 21081 18728 26115 18730
rect 21081 18672 21086 18728
rect 21142 18672 26054 18728
rect 26110 18672 26115 18728
rect 21081 18670 26115 18672
rect 21081 18667 21147 18670
rect 26049 18667 26115 18670
rect 28942 18668 28948 18732
rect 29012 18730 29018 18732
rect 32857 18730 32923 18733
rect 29012 18728 32923 18730
rect 29012 18672 32862 18728
rect 32918 18672 32923 18728
rect 29012 18670 32923 18672
rect 29012 18668 29018 18670
rect 32857 18667 32923 18670
rect 16113 18594 16179 18597
rect 10182 18592 16179 18594
rect 10182 18536 16118 18592
rect 16174 18536 16179 18592
rect 10182 18534 16179 18536
rect 9140 18532 9146 18534
rect 9489 18531 9555 18534
rect 16113 18531 16179 18534
rect 16389 18594 16455 18597
rect 17585 18594 17651 18597
rect 16389 18592 17651 18594
rect 16389 18536 16394 18592
rect 16450 18536 17590 18592
rect 17646 18536 17651 18592
rect 16389 18534 17651 18536
rect 16389 18531 16455 18534
rect 17585 18531 17651 18534
rect 18454 18532 18460 18596
rect 18524 18594 18530 18596
rect 20294 18594 20300 18596
rect 18524 18534 20300 18594
rect 18524 18532 18530 18534
rect 20294 18532 20300 18534
rect 20364 18532 20370 18596
rect 20437 18594 20503 18597
rect 21030 18594 21036 18596
rect 20437 18592 21036 18594
rect 20437 18536 20442 18592
rect 20498 18536 21036 18592
rect 20437 18534 21036 18536
rect 20437 18531 20503 18534
rect 21030 18532 21036 18534
rect 21100 18532 21106 18596
rect 22553 18594 22619 18597
rect 25313 18594 25379 18597
rect 22553 18592 25379 18594
rect 22553 18536 22558 18592
rect 22614 18536 25318 18592
rect 25374 18536 25379 18592
rect 22553 18534 25379 18536
rect 22553 18531 22619 18534
rect 25313 18531 25379 18534
rect 25589 18594 25655 18597
rect 27797 18594 27863 18597
rect 25589 18592 27863 18594
rect 25589 18536 25594 18592
rect 25650 18536 27802 18592
rect 27858 18536 27863 18592
rect 25589 18534 27863 18536
rect 25589 18531 25655 18534
rect 27797 18531 27863 18534
rect 29177 18594 29243 18597
rect 29310 18594 29316 18596
rect 29177 18592 29316 18594
rect 29177 18536 29182 18592
rect 29238 18536 29316 18592
rect 29177 18534 29316 18536
rect 29177 18531 29243 18534
rect 29310 18532 29316 18534
rect 29380 18532 29386 18596
rect 29453 18594 29519 18597
rect 29678 18594 29684 18596
rect 29453 18592 29684 18594
rect 29453 18536 29458 18592
rect 29514 18536 29684 18592
rect 29453 18534 29684 18536
rect 29453 18531 29519 18534
rect 29678 18532 29684 18534
rect 29748 18532 29754 18596
rect 30189 18594 30255 18597
rect 32489 18594 32555 18597
rect 30189 18592 32555 18594
rect 30189 18536 30194 18592
rect 30250 18536 32494 18592
rect 32550 18536 32555 18592
rect 30189 18534 32555 18536
rect 30189 18531 30255 18534
rect 32489 18531 32555 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 47946 18463 48262 18464
rect 9857 18458 9923 18461
rect 13353 18458 13419 18461
rect 16849 18460 16915 18461
rect 9857 18456 13419 18458
rect 9857 18400 9862 18456
rect 9918 18400 13358 18456
rect 13414 18400 13419 18456
rect 9857 18398 13419 18400
rect 9857 18395 9923 18398
rect 13353 18395 13419 18398
rect 13854 18396 13860 18460
rect 13924 18458 13930 18460
rect 13924 18398 16268 18458
rect 13924 18396 13930 18398
rect 0 18322 800 18352
rect 2037 18322 2103 18325
rect 0 18320 2103 18322
rect 0 18264 2042 18320
rect 2098 18264 2103 18320
rect 0 18262 2103 18264
rect 0 18232 800 18262
rect 2037 18259 2103 18262
rect 3601 18322 3667 18325
rect 10685 18322 10751 18325
rect 11329 18322 11395 18325
rect 3601 18320 11395 18322
rect 3601 18264 3606 18320
rect 3662 18264 10690 18320
rect 10746 18264 11334 18320
rect 11390 18264 11395 18320
rect 3601 18262 11395 18264
rect 3601 18259 3667 18262
rect 10685 18259 10751 18262
rect 11329 18259 11395 18262
rect 11605 18322 11671 18325
rect 16021 18322 16087 18325
rect 11605 18320 16087 18322
rect 11605 18264 11610 18320
rect 11666 18264 16026 18320
rect 16082 18264 16087 18320
rect 11605 18262 16087 18264
rect 11605 18259 11671 18262
rect 16021 18259 16087 18262
rect 4061 18186 4127 18189
rect 8109 18186 8175 18189
rect 4061 18184 8175 18186
rect 4061 18128 4066 18184
rect 4122 18128 8114 18184
rect 8170 18128 8175 18184
rect 4061 18126 8175 18128
rect 4061 18123 4127 18126
rect 8109 18123 8175 18126
rect 8569 18186 8635 18189
rect 14181 18186 14247 18189
rect 15377 18188 15443 18189
rect 8569 18184 14247 18186
rect 8569 18128 8574 18184
rect 8630 18128 14186 18184
rect 14242 18128 14247 18184
rect 8569 18126 14247 18128
rect 8569 18123 8635 18126
rect 14181 18123 14247 18126
rect 15326 18124 15332 18188
rect 15396 18186 15443 18188
rect 16208 18186 16268 18398
rect 16798 18396 16804 18460
rect 16868 18458 16915 18460
rect 16868 18456 16960 18458
rect 16910 18400 16960 18456
rect 16868 18398 16960 18400
rect 16868 18396 16915 18398
rect 17534 18396 17540 18460
rect 17604 18458 17610 18460
rect 17677 18458 17743 18461
rect 17604 18456 17743 18458
rect 17604 18400 17682 18456
rect 17738 18400 17743 18456
rect 17604 18398 17743 18400
rect 17604 18396 17610 18398
rect 16849 18395 16915 18396
rect 17677 18395 17743 18398
rect 18505 18458 18571 18461
rect 18822 18458 18828 18460
rect 18505 18456 18828 18458
rect 18505 18400 18510 18456
rect 18566 18400 18828 18456
rect 18505 18398 18828 18400
rect 18505 18395 18571 18398
rect 18822 18396 18828 18398
rect 18892 18396 18898 18460
rect 18965 18458 19031 18461
rect 22553 18458 22619 18461
rect 18965 18456 22619 18458
rect 18965 18400 18970 18456
rect 19026 18400 22558 18456
rect 22614 18400 22619 18456
rect 18965 18398 22619 18400
rect 18965 18395 19031 18398
rect 22553 18395 22619 18398
rect 23841 18458 23907 18461
rect 24945 18458 25011 18461
rect 27797 18458 27863 18461
rect 23841 18456 24410 18458
rect 23841 18400 23846 18456
rect 23902 18400 24410 18456
rect 23841 18398 24410 18400
rect 23841 18395 23907 18398
rect 16573 18322 16639 18325
rect 17493 18322 17559 18325
rect 16573 18320 17559 18322
rect 16573 18264 16578 18320
rect 16634 18264 17498 18320
rect 17554 18264 17559 18320
rect 16573 18262 17559 18264
rect 16573 18259 16639 18262
rect 17493 18259 17559 18262
rect 17953 18322 18019 18325
rect 18822 18322 18828 18324
rect 17953 18320 18828 18322
rect 17953 18264 17958 18320
rect 18014 18264 18828 18320
rect 17953 18262 18828 18264
rect 17953 18259 18019 18262
rect 18822 18260 18828 18262
rect 18892 18260 18898 18324
rect 19517 18322 19583 18325
rect 20437 18322 20503 18325
rect 19517 18320 20503 18322
rect 19517 18264 19522 18320
rect 19578 18264 20442 18320
rect 20498 18264 20503 18320
rect 19517 18262 20503 18264
rect 19517 18259 19583 18262
rect 20437 18259 20503 18262
rect 20989 18322 21055 18325
rect 24117 18322 24183 18325
rect 20989 18320 24183 18322
rect 20989 18264 20994 18320
rect 21050 18264 24122 18320
rect 24178 18264 24183 18320
rect 20989 18262 24183 18264
rect 24350 18322 24410 18398
rect 24945 18456 27863 18458
rect 24945 18400 24950 18456
rect 25006 18400 27802 18456
rect 27858 18400 27863 18456
rect 24945 18398 27863 18400
rect 24945 18395 25011 18398
rect 27797 18395 27863 18398
rect 29085 18458 29151 18461
rect 29085 18456 30666 18458
rect 29085 18400 29090 18456
rect 29146 18400 30666 18456
rect 29085 18398 30666 18400
rect 29085 18395 29151 18398
rect 26785 18322 26851 18325
rect 24350 18320 26851 18322
rect 24350 18264 26790 18320
rect 26846 18264 26851 18320
rect 24350 18262 26851 18264
rect 20989 18259 21055 18262
rect 24117 18259 24183 18262
rect 26785 18259 26851 18262
rect 27061 18322 27127 18325
rect 30465 18322 30531 18325
rect 27061 18320 30531 18322
rect 27061 18264 27066 18320
rect 27122 18264 30470 18320
rect 30526 18264 30531 18320
rect 27061 18262 30531 18264
rect 30606 18322 30666 18398
rect 31017 18322 31083 18325
rect 36813 18322 36879 18325
rect 30606 18320 36879 18322
rect 30606 18264 31022 18320
rect 31078 18264 36818 18320
rect 36874 18264 36879 18320
rect 30606 18262 36879 18264
rect 27061 18259 27127 18262
rect 30465 18259 30531 18262
rect 31017 18259 31083 18262
rect 36813 18259 36879 18262
rect 24485 18186 24551 18189
rect 15396 18184 15488 18186
rect 15438 18128 15488 18184
rect 15396 18126 15488 18128
rect 16208 18184 24551 18186
rect 16208 18128 24490 18184
rect 24546 18128 24551 18184
rect 16208 18126 24551 18128
rect 15396 18124 15443 18126
rect 15377 18123 15443 18124
rect 24485 18123 24551 18126
rect 26182 18124 26188 18188
rect 26252 18186 26258 18188
rect 28257 18186 28323 18189
rect 28993 18186 29059 18189
rect 26252 18126 27538 18186
rect 26252 18124 26258 18126
rect 6821 18050 6887 18053
rect 9213 18050 9279 18053
rect 6821 18048 9279 18050
rect 6821 17992 6826 18048
rect 6882 17992 9218 18048
rect 9274 17992 9279 18048
rect 6821 17990 9279 17992
rect 6821 17987 6887 17990
rect 9213 17987 9279 17990
rect 9765 18050 9831 18053
rect 12014 18050 12020 18052
rect 9765 18048 12020 18050
rect 9765 17992 9770 18048
rect 9826 17992 12020 18048
rect 9765 17990 12020 17992
rect 9765 17987 9831 17990
rect 12014 17988 12020 17990
rect 12084 17988 12090 18052
rect 13353 18050 13419 18053
rect 15745 18050 15811 18053
rect 16205 18050 16271 18053
rect 13353 18048 16271 18050
rect 13353 17992 13358 18048
rect 13414 17992 15750 18048
rect 15806 17992 16210 18048
rect 16266 17992 16271 18048
rect 13353 17990 16271 17992
rect 13353 17987 13419 17990
rect 15745 17987 15811 17990
rect 16205 17987 16271 17990
rect 17033 18050 17099 18053
rect 18781 18050 18847 18053
rect 19241 18050 19307 18053
rect 17033 18048 19307 18050
rect 17033 17992 17038 18048
rect 17094 17992 18786 18048
rect 18842 17992 19246 18048
rect 19302 17992 19307 18048
rect 17033 17990 19307 17992
rect 17033 17987 17099 17990
rect 18781 17987 18847 17990
rect 19241 17987 19307 17990
rect 19609 18050 19675 18053
rect 19977 18050 20043 18053
rect 19609 18048 20043 18050
rect 19609 17992 19614 18048
rect 19670 17992 19982 18048
rect 20038 17992 20043 18048
rect 19609 17990 20043 17992
rect 19609 17987 19675 17990
rect 19977 17987 20043 17990
rect 20529 18050 20595 18053
rect 21817 18050 21883 18053
rect 20529 18048 21883 18050
rect 20529 17992 20534 18048
rect 20590 17992 21822 18048
rect 21878 17992 21883 18048
rect 20529 17990 21883 17992
rect 20529 17987 20595 17990
rect 21817 17987 21883 17990
rect 24025 18050 24091 18053
rect 26182 18050 26188 18052
rect 24025 18048 26188 18050
rect 24025 17992 24030 18048
rect 24086 17992 26188 18048
rect 24025 17990 26188 17992
rect 24025 17987 24091 17990
rect 26182 17988 26188 17990
rect 26252 17988 26258 18052
rect 2946 17984 3262 17985
rect 0 17914 800 17944
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 1393 17914 1459 17917
rect 0 17912 1459 17914
rect 0 17856 1398 17912
rect 1454 17856 1459 17912
rect 0 17854 1459 17856
rect 0 17824 800 17854
rect 1393 17851 1459 17854
rect 7833 17914 7899 17917
rect 8293 17914 8359 17917
rect 12525 17914 12591 17917
rect 7833 17912 8359 17914
rect 7833 17856 7838 17912
rect 7894 17856 8298 17912
rect 8354 17856 8359 17912
rect 7833 17854 8359 17856
rect 7833 17851 7899 17854
rect 8293 17851 8359 17854
rect 9630 17912 12591 17914
rect 9630 17856 12530 17912
rect 12586 17856 12591 17912
rect 9630 17854 12591 17856
rect 3601 17778 3667 17781
rect 7465 17778 7531 17781
rect 3601 17776 7531 17778
rect 3601 17720 3606 17776
rect 3662 17720 7470 17776
rect 7526 17720 7531 17776
rect 3601 17718 7531 17720
rect 3601 17715 3667 17718
rect 7465 17715 7531 17718
rect 8201 17778 8267 17781
rect 9397 17778 9463 17781
rect 8201 17776 9463 17778
rect 8201 17720 8206 17776
rect 8262 17720 9402 17776
rect 9458 17720 9463 17776
rect 8201 17718 9463 17720
rect 8201 17715 8267 17718
rect 9397 17715 9463 17718
rect 4337 17642 4403 17645
rect 5022 17642 5028 17644
rect 4337 17640 5028 17642
rect 4337 17584 4342 17640
rect 4398 17584 5028 17640
rect 4337 17582 5028 17584
rect 4337 17579 4403 17582
rect 5022 17580 5028 17582
rect 5092 17580 5098 17644
rect 7189 17642 7255 17645
rect 9630 17642 9690 17854
rect 12525 17851 12591 17854
rect 14365 17914 14431 17917
rect 20110 17914 20116 17916
rect 14365 17912 20116 17914
rect 14365 17856 14370 17912
rect 14426 17856 20116 17912
rect 14365 17854 20116 17856
rect 14365 17851 14431 17854
rect 20110 17852 20116 17854
rect 20180 17852 20186 17916
rect 24117 17914 24183 17917
rect 26417 17914 26483 17917
rect 24117 17912 26483 17914
rect 24117 17856 24122 17912
rect 24178 17856 26422 17912
rect 26478 17856 26483 17912
rect 24117 17854 26483 17856
rect 27478 17914 27538 18126
rect 28257 18184 28826 18186
rect 28257 18128 28262 18184
rect 28318 18128 28826 18184
rect 28257 18126 28826 18128
rect 28257 18123 28323 18126
rect 27654 17988 27660 18052
rect 27724 18050 27730 18052
rect 27797 18050 27863 18053
rect 28390 18050 28396 18052
rect 27724 18048 28396 18050
rect 27724 17992 27802 18048
rect 27858 17992 28396 18048
rect 27724 17990 28396 17992
rect 27724 17988 27730 17990
rect 27797 17987 27863 17990
rect 28390 17988 28396 17990
rect 28460 17988 28466 18052
rect 28766 18050 28826 18126
rect 28993 18184 33426 18186
rect 28993 18128 28998 18184
rect 29054 18128 33426 18184
rect 28993 18126 33426 18128
rect 28993 18123 29059 18126
rect 31661 18050 31727 18053
rect 28766 18048 31727 18050
rect 28766 17992 31666 18048
rect 31722 17992 31727 18048
rect 28766 17990 31727 17992
rect 31661 17987 31727 17990
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 27654 17914 27660 17916
rect 27478 17854 27660 17914
rect 24117 17851 24183 17854
rect 26417 17851 26483 17854
rect 27654 17852 27660 17854
rect 27724 17852 27730 17916
rect 27889 17914 27955 17917
rect 29821 17914 29887 17917
rect 27889 17912 29887 17914
rect 27889 17856 27894 17912
rect 27950 17856 29826 17912
rect 29882 17856 29887 17912
rect 27889 17854 29887 17856
rect 33366 17914 33426 18126
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 35893 17914 35959 17917
rect 33366 17912 35959 17914
rect 33366 17856 35898 17912
rect 35954 17856 35959 17912
rect 33366 17854 35959 17856
rect 27889 17851 27955 17854
rect 29821 17851 29887 17854
rect 35893 17851 35959 17854
rect 11329 17778 11395 17781
rect 14825 17778 14891 17781
rect 11329 17776 14891 17778
rect 11329 17720 11334 17776
rect 11390 17720 14830 17776
rect 14886 17720 14891 17776
rect 11329 17718 14891 17720
rect 11329 17715 11395 17718
rect 14825 17715 14891 17718
rect 15101 17778 15167 17781
rect 19609 17778 19675 17781
rect 19793 17780 19859 17781
rect 15101 17776 19675 17778
rect 15101 17720 15106 17776
rect 15162 17720 19614 17776
rect 19670 17720 19675 17776
rect 15101 17718 19675 17720
rect 15101 17715 15167 17718
rect 19609 17715 19675 17718
rect 19742 17716 19748 17780
rect 19812 17778 19859 17780
rect 19977 17778 20043 17781
rect 23197 17778 23263 17781
rect 29545 17778 29611 17781
rect 19812 17776 19904 17778
rect 19854 17720 19904 17776
rect 19812 17718 19904 17720
rect 19977 17776 23122 17778
rect 19977 17720 19982 17776
rect 20038 17720 23122 17776
rect 19977 17718 23122 17720
rect 19812 17716 19859 17718
rect 19793 17715 19859 17716
rect 19977 17715 20043 17718
rect 11513 17644 11579 17645
rect 7189 17640 9690 17642
rect 7189 17584 7194 17640
rect 7250 17584 9690 17640
rect 7189 17582 9690 17584
rect 7189 17579 7255 17582
rect 11462 17580 11468 17644
rect 11532 17642 11579 17644
rect 20713 17642 20779 17645
rect 11532 17640 11624 17642
rect 11574 17584 11624 17640
rect 11532 17582 11624 17584
rect 12390 17640 20779 17642
rect 12390 17584 20718 17640
rect 20774 17584 20779 17640
rect 12390 17582 20779 17584
rect 23062 17642 23122 17718
rect 23197 17776 29611 17778
rect 23197 17720 23202 17776
rect 23258 17720 29550 17776
rect 29606 17720 29611 17776
rect 23197 17718 29611 17720
rect 23197 17715 23263 17718
rect 29545 17715 29611 17718
rect 30414 17716 30420 17780
rect 30484 17778 30490 17780
rect 36905 17778 36971 17781
rect 30484 17776 36971 17778
rect 30484 17720 36910 17776
rect 36966 17720 36971 17776
rect 30484 17718 36971 17720
rect 30484 17716 30490 17718
rect 36905 17715 36971 17718
rect 23749 17642 23815 17645
rect 30097 17642 30163 17645
rect 31753 17642 31819 17645
rect 23062 17640 31819 17642
rect 23062 17584 23754 17640
rect 23810 17584 30102 17640
rect 30158 17584 31758 17640
rect 31814 17584 31819 17640
rect 23062 17582 31819 17584
rect 11532 17580 11579 17582
rect 11513 17579 11579 17580
rect 0 17506 800 17536
rect 2037 17506 2103 17509
rect 0 17504 2103 17506
rect 0 17448 2042 17504
rect 2098 17448 2103 17504
rect 0 17446 2103 17448
rect 0 17416 800 17446
rect 2037 17443 2103 17446
rect 10501 17506 10567 17509
rect 12390 17506 12450 17582
rect 20713 17579 20779 17582
rect 23749 17579 23815 17582
rect 30097 17579 30163 17582
rect 31753 17579 31819 17582
rect 10501 17504 12450 17506
rect 10501 17448 10506 17504
rect 10562 17448 12450 17504
rect 10501 17446 12450 17448
rect 14273 17506 14339 17509
rect 14641 17506 14707 17509
rect 14273 17504 14707 17506
rect 14273 17448 14278 17504
rect 14334 17448 14646 17504
rect 14702 17448 14707 17504
rect 14273 17446 14707 17448
rect 10501 17443 10567 17446
rect 14273 17443 14339 17446
rect 14641 17443 14707 17446
rect 14825 17506 14891 17509
rect 18597 17506 18663 17509
rect 22042 17506 22048 17508
rect 14825 17504 17602 17506
rect 14825 17448 14830 17504
rect 14886 17448 17602 17504
rect 14825 17446 17602 17448
rect 14825 17443 14891 17446
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 11789 17370 11855 17373
rect 15193 17370 15259 17373
rect 11789 17368 15259 17370
rect 11789 17312 11794 17368
rect 11850 17312 15198 17368
rect 15254 17312 15259 17368
rect 11789 17310 15259 17312
rect 11789 17307 11855 17310
rect 15193 17307 15259 17310
rect 8845 17236 8911 17237
rect 4102 17172 4108 17236
rect 4172 17234 4178 17236
rect 8845 17234 8892 17236
rect 4172 17174 8402 17234
rect 8800 17232 8892 17234
rect 8800 17176 8850 17232
rect 8800 17174 8892 17176
rect 4172 17172 4178 17174
rect 0 17098 800 17128
rect 1209 17098 1275 17101
rect 0 17096 1275 17098
rect 0 17040 1214 17096
rect 1270 17040 1275 17096
rect 0 17038 1275 17040
rect 0 17008 800 17038
rect 1209 17035 1275 17038
rect 6453 17098 6519 17101
rect 6678 17098 6684 17100
rect 6453 17096 6684 17098
rect 6453 17040 6458 17096
rect 6514 17040 6684 17096
rect 6453 17038 6684 17040
rect 6453 17035 6519 17038
rect 6678 17036 6684 17038
rect 6748 17098 6754 17100
rect 8201 17098 8267 17101
rect 6748 17096 8267 17098
rect 6748 17040 8206 17096
rect 8262 17040 8267 17096
rect 6748 17038 8267 17040
rect 8342 17098 8402 17174
rect 8845 17172 8892 17174
rect 8956 17172 8962 17236
rect 9305 17234 9371 17237
rect 9438 17234 9444 17236
rect 9305 17232 9444 17234
rect 9305 17176 9310 17232
rect 9366 17176 9444 17232
rect 9305 17174 9444 17176
rect 8845 17171 8911 17172
rect 9305 17171 9371 17174
rect 9438 17172 9444 17174
rect 9508 17172 9514 17236
rect 12750 17172 12756 17236
rect 12820 17234 12826 17236
rect 14590 17234 14596 17236
rect 12820 17174 14596 17234
rect 12820 17172 12826 17174
rect 14590 17172 14596 17174
rect 14660 17172 14666 17236
rect 14733 17234 14799 17237
rect 16614 17234 16620 17236
rect 14733 17232 16620 17234
rect 14733 17176 14738 17232
rect 14794 17176 16620 17232
rect 14733 17174 16620 17176
rect 14733 17171 14799 17174
rect 16614 17172 16620 17174
rect 16684 17172 16690 17236
rect 17542 17234 17602 17446
rect 18597 17504 22048 17506
rect 18597 17448 18602 17504
rect 18658 17448 22048 17504
rect 18597 17446 22048 17448
rect 18597 17443 18663 17446
rect 22042 17444 22048 17446
rect 22112 17444 22118 17508
rect 22185 17506 22251 17509
rect 23841 17506 23907 17509
rect 27797 17506 27863 17509
rect 28533 17508 28599 17509
rect 28533 17506 28580 17508
rect 22185 17504 27863 17506
rect 22185 17448 22190 17504
rect 22246 17448 23846 17504
rect 23902 17448 27802 17504
rect 27858 17448 27863 17504
rect 22185 17446 27863 17448
rect 28488 17504 28580 17506
rect 28488 17448 28538 17504
rect 28488 17446 28580 17448
rect 22185 17443 22251 17446
rect 23841 17443 23907 17446
rect 27797 17443 27863 17446
rect 28533 17444 28580 17446
rect 28644 17444 28650 17508
rect 29269 17506 29335 17509
rect 29678 17506 29684 17508
rect 29269 17504 29684 17506
rect 29269 17448 29274 17504
rect 29330 17448 29684 17504
rect 29269 17446 29684 17448
rect 28533 17443 28599 17444
rect 29269 17443 29335 17446
rect 29678 17444 29684 17446
rect 29748 17444 29754 17508
rect 32806 17444 32812 17508
rect 32876 17506 32882 17508
rect 37365 17506 37431 17509
rect 32876 17504 37431 17506
rect 32876 17448 37370 17504
rect 37426 17448 37431 17504
rect 32876 17446 37431 17448
rect 32876 17444 32882 17446
rect 37365 17443 37431 17446
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 20846 17370 20852 17372
rect 18416 17310 20852 17370
rect 18416 17234 18476 17310
rect 20846 17308 20852 17310
rect 20916 17308 20922 17372
rect 21398 17308 21404 17372
rect 21468 17370 21474 17372
rect 23422 17370 23428 17372
rect 21468 17310 23428 17370
rect 21468 17308 21474 17310
rect 23422 17308 23428 17310
rect 23492 17308 23498 17372
rect 28901 17370 28967 17373
rect 35525 17370 35591 17373
rect 28901 17368 35591 17370
rect 28901 17312 28906 17368
rect 28962 17312 35530 17368
rect 35586 17312 35591 17368
rect 28901 17310 35591 17312
rect 28901 17307 28967 17310
rect 35525 17307 35591 17310
rect 17542 17174 18476 17234
rect 19149 17234 19215 17237
rect 30649 17234 30715 17237
rect 19149 17232 30715 17234
rect 19149 17176 19154 17232
rect 19210 17176 30654 17232
rect 30710 17176 30715 17232
rect 19149 17174 30715 17176
rect 19149 17171 19215 17174
rect 30649 17171 30715 17174
rect 22093 17098 22159 17101
rect 8342 17096 22159 17098
rect 8342 17040 22098 17096
rect 22154 17040 22159 17096
rect 8342 17038 22159 17040
rect 6748 17036 6754 17038
rect 8201 17035 8267 17038
rect 22093 17035 22159 17038
rect 22737 17098 22803 17101
rect 24301 17098 24367 17101
rect 30189 17098 30255 17101
rect 34421 17098 34487 17101
rect 22737 17096 23490 17098
rect 22737 17040 22742 17096
rect 22798 17040 23490 17096
rect 22737 17038 23490 17040
rect 22737 17035 22803 17038
rect 3877 16962 3943 16965
rect 10317 16962 10383 16965
rect 3877 16960 10383 16962
rect 3877 16904 3882 16960
rect 3938 16904 10322 16960
rect 10378 16904 10383 16960
rect 3877 16902 10383 16904
rect 3877 16899 3943 16902
rect 10317 16899 10383 16902
rect 13997 16962 14063 16965
rect 15142 16962 15148 16964
rect 13997 16960 15148 16962
rect 13997 16904 14002 16960
rect 14058 16904 15148 16960
rect 13997 16902 15148 16904
rect 13997 16899 14063 16902
rect 15142 16900 15148 16902
rect 15212 16900 15218 16964
rect 17718 16900 17724 16964
rect 17788 16962 17794 16964
rect 18505 16962 18571 16965
rect 17788 16960 18571 16962
rect 17788 16904 18510 16960
rect 18566 16904 18571 16960
rect 17788 16902 18571 16904
rect 17788 16900 17794 16902
rect 18505 16899 18571 16902
rect 19006 16900 19012 16964
rect 19076 16962 19082 16964
rect 20529 16962 20595 16965
rect 19076 16960 20595 16962
rect 19076 16904 20534 16960
rect 20590 16904 20595 16960
rect 19076 16902 20595 16904
rect 23430 16962 23490 17038
rect 24301 17096 30255 17098
rect 24301 17040 24306 17096
rect 24362 17040 30194 17096
rect 30250 17040 30255 17096
rect 24301 17038 30255 17040
rect 24301 17035 24367 17038
rect 30189 17035 30255 17038
rect 31710 17096 34487 17098
rect 31710 17040 34426 17096
rect 34482 17040 34487 17096
rect 31710 17038 34487 17040
rect 31710 16962 31770 17038
rect 34421 17035 34487 17038
rect 23430 16902 31770 16962
rect 19076 16900 19082 16902
rect 20529 16899 20595 16902
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 5942 16764 5948 16828
rect 6012 16826 6018 16828
rect 6913 16826 6979 16829
rect 6012 16824 6979 16826
rect 6012 16768 6918 16824
rect 6974 16768 6979 16824
rect 6012 16766 6979 16768
rect 6012 16764 6018 16766
rect 6913 16763 6979 16766
rect 7046 16764 7052 16828
rect 7116 16826 7122 16828
rect 8017 16826 8083 16829
rect 7116 16824 8083 16826
rect 7116 16768 8022 16824
rect 8078 16768 8083 16824
rect 7116 16766 8083 16768
rect 7116 16764 7122 16766
rect 8017 16763 8083 16766
rect 8569 16826 8635 16829
rect 15377 16826 15443 16829
rect 18413 16826 18479 16829
rect 8569 16824 12450 16826
rect 8569 16768 8574 16824
rect 8630 16768 12450 16824
rect 8569 16766 12450 16768
rect 8569 16763 8635 16766
rect 0 16690 800 16720
rect 1301 16690 1367 16693
rect 0 16688 1367 16690
rect 0 16632 1306 16688
rect 1362 16632 1367 16688
rect 0 16630 1367 16632
rect 0 16600 800 16630
rect 1301 16627 1367 16630
rect 3417 16690 3483 16693
rect 7649 16690 7715 16693
rect 7833 16692 7899 16693
rect 3417 16688 7715 16690
rect 3417 16632 3422 16688
rect 3478 16632 7654 16688
rect 7710 16632 7715 16688
rect 3417 16630 7715 16632
rect 3417 16627 3483 16630
rect 7649 16627 7715 16630
rect 7782 16628 7788 16692
rect 7852 16690 7899 16692
rect 9213 16690 9279 16693
rect 9581 16690 9647 16693
rect 7852 16688 7944 16690
rect 7894 16632 7944 16688
rect 7852 16630 7944 16632
rect 9213 16688 9647 16690
rect 9213 16632 9218 16688
rect 9274 16632 9586 16688
rect 9642 16632 9647 16688
rect 9213 16630 9647 16632
rect 7852 16628 7899 16630
rect 7833 16627 7899 16628
rect 9213 16627 9279 16630
rect 9581 16627 9647 16630
rect 9949 16690 10015 16693
rect 11053 16690 11119 16693
rect 9949 16688 11119 16690
rect 9949 16632 9954 16688
rect 10010 16632 11058 16688
rect 11114 16632 11119 16688
rect 9949 16630 11119 16632
rect 12390 16690 12450 16766
rect 15377 16824 18479 16826
rect 15377 16768 15382 16824
rect 15438 16768 18418 16824
rect 18474 16768 18479 16824
rect 15377 16766 18479 16768
rect 15377 16763 15443 16766
rect 18413 16763 18479 16766
rect 18965 16826 19031 16829
rect 23565 16826 23631 16829
rect 25262 16826 25268 16828
rect 18965 16824 22754 16826
rect 18965 16768 18970 16824
rect 19026 16768 22754 16824
rect 18965 16766 22754 16768
rect 18965 16763 19031 16766
rect 14733 16690 14799 16693
rect 12390 16688 14799 16690
rect 12390 16632 14738 16688
rect 14794 16632 14799 16688
rect 12390 16630 14799 16632
rect 9949 16627 10015 16630
rect 11053 16627 11119 16630
rect 14733 16627 14799 16630
rect 16113 16690 16179 16693
rect 16430 16690 16436 16692
rect 16113 16688 16436 16690
rect 16113 16632 16118 16688
rect 16174 16632 16436 16688
rect 16113 16630 16436 16632
rect 16113 16627 16179 16630
rect 16430 16628 16436 16630
rect 16500 16628 16506 16692
rect 17769 16690 17835 16693
rect 22694 16690 22754 16766
rect 23565 16824 25268 16826
rect 23565 16768 23570 16824
rect 23626 16768 25268 16824
rect 23565 16766 25268 16768
rect 23565 16763 23631 16766
rect 25262 16764 25268 16766
rect 25332 16764 25338 16828
rect 25405 16826 25471 16829
rect 28942 16826 28948 16828
rect 25405 16824 28948 16826
rect 25405 16768 25410 16824
rect 25466 16768 28948 16824
rect 25405 16766 28948 16768
rect 25405 16763 25471 16766
rect 28942 16764 28948 16766
rect 29012 16764 29018 16828
rect 29310 16764 29316 16828
rect 29380 16826 29386 16828
rect 29637 16826 29703 16829
rect 29380 16824 29703 16826
rect 29380 16768 29642 16824
rect 29698 16768 29703 16824
rect 29380 16766 29703 16768
rect 29380 16764 29386 16766
rect 29637 16763 29703 16766
rect 29913 16826 29979 16829
rect 31661 16826 31727 16829
rect 29913 16824 31727 16826
rect 29913 16768 29918 16824
rect 29974 16768 31666 16824
rect 31722 16768 31727 16824
rect 29913 16766 31727 16768
rect 29913 16763 29979 16766
rect 31661 16763 31727 16766
rect 17769 16688 22570 16690
rect 17769 16632 17774 16688
rect 17830 16632 22570 16688
rect 17769 16630 22570 16632
rect 22694 16630 27676 16690
rect 17769 16627 17835 16630
rect 5022 16492 5028 16556
rect 5092 16554 5098 16556
rect 8109 16554 8175 16557
rect 5092 16552 8175 16554
rect 5092 16496 8114 16552
rect 8170 16496 8175 16552
rect 5092 16494 8175 16496
rect 5092 16492 5098 16494
rect 8109 16491 8175 16494
rect 8293 16554 8359 16557
rect 10174 16554 10180 16556
rect 8293 16552 10180 16554
rect 8293 16496 8298 16552
rect 8354 16496 10180 16552
rect 8293 16494 10180 16496
rect 8293 16491 8359 16494
rect 10174 16492 10180 16494
rect 10244 16492 10250 16556
rect 11646 16492 11652 16556
rect 11716 16554 11722 16556
rect 13353 16554 13419 16557
rect 11716 16552 13419 16554
rect 11716 16496 13358 16552
rect 13414 16496 13419 16552
rect 11716 16494 13419 16496
rect 11716 16492 11722 16494
rect 13353 16491 13419 16494
rect 16205 16554 16271 16557
rect 18689 16554 18755 16557
rect 21950 16554 21956 16556
rect 16205 16552 18755 16554
rect 16205 16496 16210 16552
rect 16266 16496 18694 16552
rect 18750 16496 18755 16552
rect 16205 16494 18755 16496
rect 16205 16491 16271 16494
rect 18689 16491 18755 16494
rect 18830 16494 21956 16554
rect 8569 16418 8635 16421
rect 12525 16418 12591 16421
rect 17401 16418 17467 16421
rect 8569 16416 9690 16418
rect 8569 16360 8574 16416
rect 8630 16360 9690 16416
rect 8569 16358 9690 16360
rect 8569 16355 8635 16358
rect 7946 16352 8262 16353
rect 0 16282 800 16312
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 1301 16282 1367 16285
rect 0 16280 1367 16282
rect 0 16224 1306 16280
rect 1362 16224 1367 16280
rect 0 16222 1367 16224
rect 0 16192 800 16222
rect 1301 16219 1367 16222
rect 1894 16220 1900 16284
rect 1964 16282 1970 16284
rect 8661 16282 8727 16285
rect 9397 16282 9463 16285
rect 1964 16222 7850 16282
rect 1964 16220 1970 16222
rect 5206 16084 5212 16148
rect 5276 16146 5282 16148
rect 5993 16146 6059 16149
rect 5276 16144 6059 16146
rect 5276 16088 5998 16144
rect 6054 16088 6059 16144
rect 5276 16086 6059 16088
rect 5276 16084 5282 16086
rect 5993 16083 6059 16086
rect 6637 16146 6703 16149
rect 7598 16146 7604 16148
rect 6637 16144 7604 16146
rect 6637 16088 6642 16144
rect 6698 16088 7604 16144
rect 6637 16086 7604 16088
rect 6637 16083 6703 16086
rect 7598 16084 7604 16086
rect 7668 16084 7674 16148
rect 7790 16146 7850 16222
rect 8661 16280 9463 16282
rect 8661 16224 8666 16280
rect 8722 16224 9402 16280
rect 9458 16224 9463 16280
rect 8661 16222 9463 16224
rect 9630 16282 9690 16358
rect 12525 16416 17467 16418
rect 12525 16360 12530 16416
rect 12586 16360 17406 16416
rect 17462 16360 17467 16416
rect 12525 16358 17467 16360
rect 12525 16355 12591 16358
rect 17401 16355 17467 16358
rect 18597 16418 18663 16421
rect 18830 16418 18890 16494
rect 21950 16492 21956 16494
rect 22020 16492 22026 16556
rect 22510 16554 22570 16630
rect 24945 16554 25011 16557
rect 22510 16552 25011 16554
rect 22510 16496 24950 16552
rect 25006 16496 25011 16552
rect 22510 16494 25011 16496
rect 24945 16491 25011 16494
rect 26233 16554 26299 16557
rect 26785 16554 26851 16557
rect 26233 16552 26851 16554
rect 26233 16496 26238 16552
rect 26294 16496 26790 16552
rect 26846 16496 26851 16552
rect 26233 16494 26851 16496
rect 27616 16554 27676 16630
rect 43897 16554 43963 16557
rect 27616 16552 43963 16554
rect 27616 16496 43902 16552
rect 43958 16496 43963 16552
rect 27616 16494 43963 16496
rect 26233 16491 26299 16494
rect 26785 16491 26851 16494
rect 43897 16491 43963 16494
rect 18597 16416 18890 16418
rect 18597 16360 18602 16416
rect 18658 16360 18890 16416
rect 18597 16358 18890 16360
rect 18965 16418 19031 16421
rect 19425 16420 19491 16421
rect 19190 16418 19196 16420
rect 18965 16416 19196 16418
rect 18965 16360 18970 16416
rect 19026 16360 19196 16416
rect 18965 16358 19196 16360
rect 18597 16355 18663 16358
rect 18965 16355 19031 16358
rect 19190 16356 19196 16358
rect 19260 16356 19266 16420
rect 19374 16356 19380 16420
rect 19444 16418 19491 16420
rect 19444 16416 19536 16418
rect 19486 16360 19536 16416
rect 19444 16358 19536 16360
rect 19444 16356 19491 16358
rect 22686 16356 22692 16420
rect 22756 16418 22762 16420
rect 23197 16418 23263 16421
rect 24117 16418 24183 16421
rect 22756 16416 24183 16418
rect 22756 16360 23202 16416
rect 23258 16360 24122 16416
rect 24178 16360 24183 16416
rect 22756 16358 24183 16360
rect 22756 16356 22762 16358
rect 19425 16355 19491 16356
rect 23197 16355 23263 16358
rect 24117 16355 24183 16358
rect 26417 16418 26483 16421
rect 27613 16418 27679 16421
rect 26417 16416 27679 16418
rect 26417 16360 26422 16416
rect 26478 16360 27618 16416
rect 27674 16360 27679 16416
rect 26417 16358 27679 16360
rect 26417 16355 26483 16358
rect 27613 16355 27679 16358
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 10685 16282 10751 16285
rect 11421 16282 11487 16285
rect 11830 16282 11836 16284
rect 9630 16280 11836 16282
rect 9630 16224 10690 16280
rect 10746 16224 11426 16280
rect 11482 16224 11836 16280
rect 9630 16222 11836 16224
rect 8661 16219 8727 16222
rect 9397 16219 9463 16222
rect 10685 16219 10751 16222
rect 11421 16219 11487 16222
rect 11830 16220 11836 16222
rect 11900 16220 11906 16284
rect 13721 16282 13787 16285
rect 16246 16282 16252 16284
rect 13721 16280 16252 16282
rect 13721 16224 13726 16280
rect 13782 16224 16252 16280
rect 13721 16222 16252 16224
rect 13721 16219 13787 16222
rect 16246 16220 16252 16222
rect 16316 16220 16322 16284
rect 17125 16282 17191 16285
rect 17585 16282 17651 16285
rect 22645 16282 22711 16285
rect 23565 16284 23631 16285
rect 23565 16282 23612 16284
rect 17125 16280 17651 16282
rect 17125 16224 17130 16280
rect 17186 16224 17590 16280
rect 17646 16224 17651 16280
rect 17125 16222 17651 16224
rect 17125 16219 17191 16222
rect 17585 16219 17651 16222
rect 18462 16280 22711 16282
rect 18462 16224 22650 16280
rect 22706 16224 22711 16280
rect 18462 16222 22711 16224
rect 23520 16280 23612 16282
rect 23676 16282 23682 16284
rect 25078 16282 25084 16284
rect 23520 16224 23570 16280
rect 23520 16222 23612 16224
rect 11053 16146 11119 16149
rect 7790 16144 11119 16146
rect 7790 16088 11058 16144
rect 11114 16088 11119 16144
rect 7790 16086 11119 16088
rect 11053 16083 11119 16086
rect 11513 16146 11579 16149
rect 12893 16146 12959 16149
rect 11513 16144 12959 16146
rect 11513 16088 11518 16144
rect 11574 16088 12898 16144
rect 12954 16088 12959 16144
rect 11513 16086 12959 16088
rect 11513 16083 11579 16086
rect 12893 16083 12959 16086
rect 13353 16146 13419 16149
rect 18462 16146 18522 16222
rect 22645 16219 22711 16222
rect 23565 16220 23612 16222
rect 23676 16222 25084 16282
rect 23676 16220 23682 16222
rect 25078 16220 25084 16222
rect 25148 16220 25154 16284
rect 25630 16220 25636 16284
rect 25700 16282 25706 16284
rect 27797 16282 27863 16285
rect 25700 16280 27863 16282
rect 25700 16224 27802 16280
rect 27858 16224 27863 16280
rect 25700 16222 27863 16224
rect 25700 16220 25706 16222
rect 23565 16219 23631 16220
rect 27797 16219 27863 16222
rect 13353 16144 18522 16146
rect 13353 16088 13358 16144
rect 13414 16088 18522 16144
rect 13353 16086 18522 16088
rect 18597 16146 18663 16149
rect 27797 16146 27863 16149
rect 18597 16144 27863 16146
rect 18597 16088 18602 16144
rect 18658 16088 27802 16144
rect 27858 16088 27863 16144
rect 18597 16086 27863 16088
rect 13353 16083 13419 16086
rect 18597 16083 18663 16086
rect 27797 16083 27863 16086
rect 27981 16146 28047 16149
rect 29177 16146 29243 16149
rect 34881 16146 34947 16149
rect 27981 16144 29243 16146
rect 27981 16088 27986 16144
rect 28042 16088 29182 16144
rect 29238 16088 29243 16144
rect 27981 16086 29243 16088
rect 27981 16083 28047 16086
rect 29177 16083 29243 16086
rect 31710 16144 34947 16146
rect 31710 16088 34886 16144
rect 34942 16088 34947 16144
rect 31710 16086 34947 16088
rect 974 15948 980 16012
rect 1044 16010 1050 16012
rect 8753 16010 8819 16013
rect 1044 16008 8819 16010
rect 1044 15952 8758 16008
rect 8814 15952 8819 16008
rect 1044 15950 8819 15952
rect 1044 15948 1050 15950
rect 8753 15947 8819 15950
rect 10317 16010 10383 16013
rect 14457 16010 14523 16013
rect 25497 16010 25563 16013
rect 10317 16008 13416 16010
rect 10317 15952 10322 16008
rect 10378 15952 13416 16008
rect 10317 15950 13416 15952
rect 10317 15947 10383 15950
rect 0 15874 800 15904
rect 1301 15874 1367 15877
rect 0 15872 1367 15874
rect 0 15816 1306 15872
rect 1362 15816 1367 15872
rect 0 15814 1367 15816
rect 0 15784 800 15814
rect 1301 15811 1367 15814
rect 7230 15812 7236 15876
rect 7300 15874 7306 15876
rect 13356 15874 13416 15950
rect 14457 16008 25563 16010
rect 14457 15952 14462 16008
rect 14518 15952 25502 16008
rect 25558 15952 25563 16008
rect 14457 15950 25563 15952
rect 14457 15947 14523 15950
rect 25497 15947 25563 15950
rect 27705 16010 27771 16013
rect 31569 16010 31635 16013
rect 27705 16008 31635 16010
rect 27705 15952 27710 16008
rect 27766 15952 31574 16008
rect 31630 15952 31635 16008
rect 27705 15950 31635 15952
rect 27705 15947 27771 15950
rect 31569 15947 31635 15950
rect 15561 15874 15627 15877
rect 7300 15814 12450 15874
rect 13356 15872 15627 15874
rect 13356 15816 15566 15872
rect 15622 15816 15627 15872
rect 13356 15814 15627 15816
rect 7300 15812 7306 15814
rect 2946 15808 3262 15809
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 7649 15738 7715 15741
rect 9029 15738 9095 15741
rect 10225 15738 10291 15741
rect 7649 15736 8770 15738
rect 7649 15680 7654 15736
rect 7710 15680 8770 15736
rect 7649 15678 8770 15680
rect 7649 15675 7715 15678
rect 3601 15602 3667 15605
rect 7649 15602 7715 15605
rect 3601 15600 7715 15602
rect 3601 15544 3606 15600
rect 3662 15544 7654 15600
rect 7710 15544 7715 15600
rect 3601 15542 7715 15544
rect 3601 15539 3667 15542
rect 7649 15539 7715 15542
rect 7925 15602 7991 15605
rect 8518 15602 8524 15604
rect 7925 15600 8524 15602
rect 7925 15544 7930 15600
rect 7986 15544 8524 15600
rect 7925 15542 8524 15544
rect 7925 15539 7991 15542
rect 8518 15540 8524 15542
rect 8588 15540 8594 15604
rect 8710 15602 8770 15678
rect 9029 15736 10291 15738
rect 9029 15680 9034 15736
rect 9090 15680 10230 15736
rect 10286 15680 10291 15736
rect 9029 15678 10291 15680
rect 12390 15738 12450 15814
rect 15561 15811 15627 15814
rect 17166 15812 17172 15876
rect 17236 15874 17242 15876
rect 19742 15874 19748 15876
rect 17236 15814 19748 15874
rect 17236 15812 17242 15814
rect 19742 15812 19748 15814
rect 19812 15812 19818 15876
rect 24158 15812 24164 15876
rect 24228 15874 24234 15876
rect 31710 15874 31770 16086
rect 34881 16083 34947 16086
rect 24228 15814 31770 15874
rect 24228 15812 24234 15814
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 42946 15743 43262 15744
rect 13997 15738 14063 15741
rect 14457 15738 14523 15741
rect 18781 15738 18847 15741
rect 12390 15678 12818 15738
rect 9029 15675 9095 15678
rect 10225 15675 10291 15678
rect 12525 15602 12591 15605
rect 8710 15600 12591 15602
rect 8710 15544 12530 15600
rect 12586 15544 12591 15600
rect 8710 15542 12591 15544
rect 12758 15602 12818 15678
rect 13997 15736 14290 15738
rect 13997 15680 14002 15736
rect 14058 15680 14290 15736
rect 13997 15678 14290 15680
rect 13997 15675 14063 15678
rect 14089 15602 14155 15605
rect 12758 15600 14155 15602
rect 12758 15544 14094 15600
rect 14150 15544 14155 15600
rect 12758 15542 14155 15544
rect 14230 15602 14290 15678
rect 14457 15736 18847 15738
rect 14457 15680 14462 15736
rect 14518 15680 18786 15736
rect 18842 15680 18847 15736
rect 14457 15678 18847 15680
rect 14457 15675 14523 15678
rect 18781 15675 18847 15678
rect 19558 15676 19564 15740
rect 19628 15738 19634 15740
rect 22318 15738 22324 15740
rect 19628 15678 22324 15738
rect 19628 15676 19634 15678
rect 22318 15676 22324 15678
rect 22388 15676 22394 15740
rect 27654 15676 27660 15740
rect 27724 15738 27730 15740
rect 27981 15738 28047 15741
rect 27724 15736 28047 15738
rect 27724 15680 27986 15736
rect 28042 15680 28047 15736
rect 27724 15678 28047 15680
rect 27724 15676 27730 15678
rect 27981 15675 28047 15678
rect 16665 15602 16731 15605
rect 14230 15600 16731 15602
rect 14230 15544 16670 15600
rect 16726 15544 16731 15600
rect 14230 15542 16731 15544
rect 12525 15539 12591 15542
rect 14089 15539 14155 15542
rect 16665 15539 16731 15542
rect 16849 15602 16915 15605
rect 17350 15602 17356 15604
rect 16849 15600 17356 15602
rect 16849 15544 16854 15600
rect 16910 15544 17356 15600
rect 16849 15542 17356 15544
rect 16849 15539 16915 15542
rect 17350 15540 17356 15542
rect 17420 15540 17426 15604
rect 17585 15602 17651 15605
rect 19006 15602 19012 15604
rect 17585 15600 19012 15602
rect 17585 15544 17590 15600
rect 17646 15544 19012 15600
rect 17585 15542 19012 15544
rect 17585 15539 17651 15542
rect 19006 15540 19012 15542
rect 19076 15540 19082 15604
rect 19885 15602 19951 15605
rect 20161 15602 20227 15605
rect 19885 15600 20227 15602
rect 19885 15544 19890 15600
rect 19946 15544 20166 15600
rect 20222 15544 20227 15600
rect 19885 15542 20227 15544
rect 19885 15539 19951 15542
rect 20161 15539 20227 15542
rect 20529 15602 20595 15605
rect 20662 15602 20668 15604
rect 20529 15600 20668 15602
rect 20529 15544 20534 15600
rect 20590 15544 20668 15600
rect 20529 15542 20668 15544
rect 20529 15539 20595 15542
rect 20662 15540 20668 15542
rect 20732 15540 20738 15604
rect 22134 15540 22140 15604
rect 22204 15602 22210 15604
rect 30649 15602 30715 15605
rect 22204 15600 30715 15602
rect 22204 15544 30654 15600
rect 30710 15544 30715 15600
rect 22204 15542 30715 15544
rect 22204 15540 22210 15542
rect 30649 15539 30715 15542
rect 31518 15540 31524 15604
rect 31588 15602 31594 15604
rect 31753 15602 31819 15605
rect 31588 15600 31819 15602
rect 31588 15544 31758 15600
rect 31814 15544 31819 15600
rect 31588 15542 31819 15544
rect 31588 15540 31594 15542
rect 31753 15539 31819 15542
rect 0 15466 800 15496
rect 1301 15466 1367 15469
rect 0 15464 1367 15466
rect 0 15408 1306 15464
rect 1362 15408 1367 15464
rect 0 15406 1367 15408
rect 0 15376 800 15406
rect 1301 15403 1367 15406
rect 3417 15466 3483 15469
rect 7925 15466 7991 15469
rect 3417 15464 7991 15466
rect 3417 15408 3422 15464
rect 3478 15408 7930 15464
rect 7986 15408 7991 15464
rect 3417 15406 7991 15408
rect 3417 15403 3483 15406
rect 7925 15403 7991 15406
rect 11145 15466 11211 15469
rect 14273 15466 14339 15469
rect 11145 15464 14339 15466
rect 11145 15408 11150 15464
rect 11206 15408 14278 15464
rect 14334 15408 14339 15464
rect 11145 15406 14339 15408
rect 11145 15403 11211 15406
rect 14273 15403 14339 15406
rect 15653 15466 15719 15469
rect 17125 15466 17191 15469
rect 27521 15466 27587 15469
rect 15653 15464 17050 15466
rect 15653 15408 15658 15464
rect 15714 15408 17050 15464
rect 15653 15406 17050 15408
rect 15653 15403 15719 15406
rect 9254 15268 9260 15332
rect 9324 15330 9330 15332
rect 11421 15330 11487 15333
rect 9324 15328 11487 15330
rect 9324 15272 11426 15328
rect 11482 15272 11487 15328
rect 9324 15270 11487 15272
rect 9324 15268 9330 15270
rect 11421 15267 11487 15270
rect 11973 15330 12039 15333
rect 16849 15330 16915 15333
rect 11973 15328 16915 15330
rect 11973 15272 11978 15328
rect 12034 15272 16854 15328
rect 16910 15272 16915 15328
rect 11973 15270 16915 15272
rect 16990 15330 17050 15406
rect 17125 15464 27587 15466
rect 17125 15408 17130 15464
rect 17186 15408 27526 15464
rect 27582 15408 27587 15464
rect 17125 15406 27587 15408
rect 17125 15403 17191 15406
rect 27521 15403 27587 15406
rect 27705 15466 27771 15469
rect 38653 15466 38719 15469
rect 27705 15464 38719 15466
rect 27705 15408 27710 15464
rect 27766 15408 38658 15464
rect 38714 15408 38719 15464
rect 27705 15406 38719 15408
rect 27705 15403 27771 15406
rect 38653 15403 38719 15406
rect 17677 15330 17743 15333
rect 18505 15332 18571 15333
rect 16990 15328 17743 15330
rect 16990 15272 17682 15328
rect 17738 15272 17743 15328
rect 16990 15270 17743 15272
rect 11973 15267 12039 15270
rect 16849 15267 16915 15270
rect 17677 15267 17743 15270
rect 18454 15268 18460 15332
rect 18524 15330 18571 15332
rect 18689 15330 18755 15333
rect 19374 15330 19380 15332
rect 18524 15328 18616 15330
rect 18566 15272 18616 15328
rect 18524 15270 18616 15272
rect 18689 15328 19380 15330
rect 18689 15272 18694 15328
rect 18750 15272 19380 15328
rect 18689 15270 19380 15272
rect 18524 15268 18571 15270
rect 18505 15267 18571 15268
rect 18689 15267 18755 15270
rect 19374 15268 19380 15270
rect 19444 15268 19450 15332
rect 19517 15330 19583 15333
rect 25589 15330 25655 15333
rect 27337 15330 27403 15333
rect 19517 15328 24824 15330
rect 19517 15272 19522 15328
rect 19578 15272 24824 15328
rect 19517 15270 24824 15272
rect 19517 15267 19583 15270
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 3366 15132 3372 15196
rect 3436 15194 3442 15196
rect 3693 15194 3759 15197
rect 3436 15192 3759 15194
rect 3436 15136 3698 15192
rect 3754 15136 3759 15192
rect 3436 15134 3759 15136
rect 3436 15132 3442 15134
rect 3693 15131 3759 15134
rect 5533 15194 5599 15197
rect 7649 15194 7715 15197
rect 5533 15192 7715 15194
rect 5533 15136 5538 15192
rect 5594 15136 7654 15192
rect 7710 15136 7715 15192
rect 5533 15134 7715 15136
rect 5533 15131 5599 15134
rect 7649 15131 7715 15134
rect 8569 15194 8635 15197
rect 9397 15194 9463 15197
rect 9857 15194 9923 15197
rect 8569 15192 9923 15194
rect 8569 15136 8574 15192
rect 8630 15136 9402 15192
rect 9458 15136 9862 15192
rect 9918 15136 9923 15192
rect 8569 15134 9923 15136
rect 8569 15131 8635 15134
rect 9397 15131 9463 15134
rect 9857 15131 9923 15134
rect 10501 15194 10567 15197
rect 12341 15194 12407 15197
rect 12525 15194 12591 15197
rect 10501 15192 12591 15194
rect 10501 15136 10506 15192
rect 10562 15136 12346 15192
rect 12402 15136 12530 15192
rect 12586 15136 12591 15192
rect 10501 15134 12591 15136
rect 10501 15131 10567 15134
rect 12341 15131 12407 15134
rect 12525 15131 12591 15134
rect 12750 15132 12756 15196
rect 12820 15194 12826 15196
rect 17166 15194 17172 15196
rect 12820 15134 17172 15194
rect 12820 15132 12826 15134
rect 17166 15132 17172 15134
rect 17236 15132 17242 15196
rect 18413 15194 18479 15197
rect 24577 15194 24643 15197
rect 18413 15192 24643 15194
rect 18413 15136 18418 15192
rect 18474 15136 24582 15192
rect 24638 15136 24643 15192
rect 18413 15134 24643 15136
rect 24764 15194 24824 15270
rect 25589 15328 27403 15330
rect 25589 15272 25594 15328
rect 25650 15272 27342 15328
rect 27398 15272 27403 15328
rect 25589 15270 27403 15272
rect 25589 15267 25655 15270
rect 27337 15267 27403 15270
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 26417 15194 26483 15197
rect 24764 15192 26483 15194
rect 24764 15136 26422 15192
rect 26478 15136 26483 15192
rect 24764 15134 26483 15136
rect 18413 15131 18479 15134
rect 24577 15131 24643 15134
rect 26417 15131 26483 15134
rect 28390 15132 28396 15196
rect 28460 15194 28466 15196
rect 35065 15194 35131 15197
rect 28460 15192 35131 15194
rect 28460 15136 35070 15192
rect 35126 15136 35131 15192
rect 28460 15134 35131 15136
rect 28460 15132 28466 15134
rect 35065 15131 35131 15134
rect 0 15058 800 15088
rect 1301 15058 1367 15061
rect 0 15056 1367 15058
rect 0 15000 1306 15056
rect 1362 15000 1367 15056
rect 0 14998 1367 15000
rect 0 14968 800 14998
rect 1301 14995 1367 14998
rect 3734 14996 3740 15060
rect 3804 15058 3810 15060
rect 3969 15058 4035 15061
rect 4102 15058 4108 15060
rect 3804 15056 4108 15058
rect 3804 15000 3974 15056
rect 4030 15000 4108 15056
rect 3804 14998 4108 15000
rect 3804 14996 3810 14998
rect 3969 14995 4035 14998
rect 4102 14996 4108 14998
rect 4172 14996 4178 15060
rect 6494 14996 6500 15060
rect 6564 15058 6570 15060
rect 7005 15058 7071 15061
rect 6564 15056 7071 15058
rect 6564 15000 7010 15056
rect 7066 15000 7071 15056
rect 6564 14998 7071 15000
rect 6564 14996 6570 14998
rect 7005 14995 7071 14998
rect 7373 15058 7439 15061
rect 13629 15058 13695 15061
rect 15745 15060 15811 15061
rect 7373 15056 13695 15058
rect 7373 15000 7378 15056
rect 7434 15000 13634 15056
rect 13690 15000 13695 15056
rect 7373 14998 13695 15000
rect 7373 14995 7439 14998
rect 13629 14995 13695 14998
rect 15694 14996 15700 15060
rect 15764 15058 15811 15060
rect 16297 15058 16363 15061
rect 28717 15058 28783 15061
rect 15764 15056 15856 15058
rect 15806 15000 15856 15056
rect 15764 14998 15856 15000
rect 16297 15056 28783 15058
rect 16297 15000 16302 15056
rect 16358 15000 28722 15056
rect 28778 15000 28783 15056
rect 16297 14998 28783 15000
rect 15764 14996 15811 14998
rect 15745 14995 15811 14996
rect 16297 14995 16363 14998
rect 28717 14995 28783 14998
rect 29126 14996 29132 15060
rect 29196 15058 29202 15060
rect 31201 15058 31267 15061
rect 29196 15056 31267 15058
rect 29196 15000 31206 15056
rect 31262 15000 31267 15056
rect 29196 14998 31267 15000
rect 29196 14996 29202 14998
rect 31201 14995 31267 14998
rect 3877 14922 3943 14925
rect 8017 14922 8083 14925
rect 3877 14920 8083 14922
rect 3877 14864 3882 14920
rect 3938 14864 8022 14920
rect 8078 14864 8083 14920
rect 3877 14862 8083 14864
rect 3877 14859 3943 14862
rect 8017 14859 8083 14862
rect 11237 14922 11303 14925
rect 16481 14922 16547 14925
rect 11237 14920 16547 14922
rect 11237 14864 11242 14920
rect 11298 14864 16486 14920
rect 16542 14864 16547 14920
rect 11237 14862 16547 14864
rect 11237 14859 11303 14862
rect 16481 14859 16547 14862
rect 16665 14922 16731 14925
rect 17125 14922 17191 14925
rect 16665 14920 17191 14922
rect 16665 14864 16670 14920
rect 16726 14864 17130 14920
rect 17186 14864 17191 14920
rect 16665 14862 17191 14864
rect 16665 14859 16731 14862
rect 17125 14859 17191 14862
rect 17401 14922 17467 14925
rect 23197 14922 23263 14925
rect 17401 14920 23263 14922
rect 17401 14864 17406 14920
rect 17462 14864 23202 14920
rect 23258 14864 23263 14920
rect 17401 14862 23263 14864
rect 17401 14859 17467 14862
rect 23197 14859 23263 14862
rect 24577 14922 24643 14925
rect 28349 14922 28415 14925
rect 24577 14920 28415 14922
rect 24577 14864 24582 14920
rect 24638 14864 28354 14920
rect 28410 14864 28415 14920
rect 24577 14862 28415 14864
rect 24577 14859 24643 14862
rect 28349 14859 28415 14862
rect 28717 14922 28783 14925
rect 34789 14922 34855 14925
rect 28717 14920 34855 14922
rect 28717 14864 28722 14920
rect 28778 14864 34794 14920
rect 34850 14864 34855 14920
rect 28717 14862 34855 14864
rect 28717 14859 28783 14862
rect 34789 14859 34855 14862
rect 4245 14786 4311 14789
rect 7097 14786 7163 14789
rect 4245 14784 7163 14786
rect 4245 14728 4250 14784
rect 4306 14728 7102 14784
rect 7158 14728 7163 14784
rect 4245 14726 7163 14728
rect 4245 14723 4311 14726
rect 7097 14723 7163 14726
rect 10961 14786 11027 14789
rect 11789 14788 11855 14789
rect 11789 14786 11836 14788
rect 10961 14784 11836 14786
rect 10961 14728 10966 14784
rect 11022 14728 11794 14784
rect 10961 14726 11836 14728
rect 10961 14723 11027 14726
rect 11789 14724 11836 14726
rect 11900 14724 11906 14788
rect 13813 14786 13879 14789
rect 20253 14786 20319 14789
rect 13813 14784 20319 14786
rect 13813 14728 13818 14784
rect 13874 14728 20258 14784
rect 20314 14728 20319 14784
rect 13813 14726 20319 14728
rect 11789 14723 11855 14724
rect 13813 14723 13879 14726
rect 20253 14723 20319 14726
rect 21582 14724 21588 14788
rect 21652 14786 21658 14788
rect 21725 14786 21791 14789
rect 22686 14786 22692 14788
rect 21652 14784 22692 14786
rect 21652 14728 21730 14784
rect 21786 14728 22692 14784
rect 21652 14726 22692 14728
rect 21652 14724 21658 14726
rect 21725 14723 21791 14726
rect 22686 14724 22692 14726
rect 22756 14724 22762 14788
rect 24209 14786 24275 14789
rect 24485 14786 24551 14789
rect 24209 14784 24551 14786
rect 24209 14728 24214 14784
rect 24270 14728 24490 14784
rect 24546 14728 24551 14784
rect 24209 14726 24551 14728
rect 24209 14723 24275 14726
rect 24485 14723 24551 14726
rect 25998 14724 26004 14788
rect 26068 14786 26074 14788
rect 32806 14786 32812 14788
rect 26068 14726 32812 14786
rect 26068 14724 26074 14726
rect 32806 14724 32812 14726
rect 32876 14724 32882 14788
rect 2946 14720 3262 14721
rect 0 14650 800 14680
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 1301 14650 1367 14653
rect 0 14648 1367 14650
rect 0 14592 1306 14648
rect 1362 14592 1367 14648
rect 0 14590 1367 14592
rect 0 14560 800 14590
rect 1301 14587 1367 14590
rect 9438 14588 9444 14652
rect 9508 14650 9514 14652
rect 10685 14650 10751 14653
rect 9508 14648 10751 14650
rect 9508 14592 10690 14648
rect 10746 14592 10751 14648
rect 9508 14590 10751 14592
rect 9508 14588 9514 14590
rect 10685 14587 10751 14590
rect 11697 14650 11763 14653
rect 12801 14650 12867 14653
rect 11697 14648 12867 14650
rect 11697 14592 11702 14648
rect 11758 14592 12806 14648
rect 12862 14592 12867 14648
rect 11697 14590 12867 14592
rect 11697 14587 11763 14590
rect 12801 14587 12867 14590
rect 15469 14650 15535 14653
rect 21582 14650 21588 14652
rect 15469 14648 21588 14650
rect 15469 14592 15474 14648
rect 15530 14592 21588 14648
rect 15469 14590 21588 14592
rect 15469 14587 15535 14590
rect 21582 14588 21588 14590
rect 21652 14588 21658 14652
rect 23422 14588 23428 14652
rect 23492 14650 23498 14652
rect 24342 14650 24348 14652
rect 23492 14590 24348 14650
rect 23492 14588 23498 14590
rect 24342 14588 24348 14590
rect 24412 14650 24418 14652
rect 24577 14650 24643 14653
rect 24412 14648 24643 14650
rect 24412 14592 24582 14648
rect 24638 14592 24643 14648
rect 24412 14590 24643 14592
rect 24412 14588 24418 14590
rect 24577 14587 24643 14590
rect 25446 14588 25452 14652
rect 25516 14650 25522 14652
rect 28717 14650 28783 14653
rect 25516 14648 28783 14650
rect 25516 14592 28722 14648
rect 28778 14592 28783 14648
rect 25516 14590 28783 14592
rect 25516 14588 25522 14590
rect 28717 14587 28783 14590
rect 7782 14452 7788 14516
rect 7852 14514 7858 14516
rect 13486 14514 13492 14516
rect 7852 14454 13492 14514
rect 7852 14452 7858 14454
rect 13486 14452 13492 14454
rect 13556 14452 13562 14516
rect 13721 14514 13787 14517
rect 13678 14512 13787 14514
rect 13678 14456 13726 14512
rect 13782 14456 13787 14512
rect 13678 14451 13787 14456
rect 15142 14452 15148 14516
rect 15212 14514 15218 14516
rect 16297 14514 16363 14517
rect 15212 14512 16363 14514
rect 15212 14456 16302 14512
rect 16358 14456 16363 14512
rect 15212 14454 16363 14456
rect 15212 14452 15218 14454
rect 16297 14451 16363 14454
rect 16614 14452 16620 14516
rect 16684 14514 16690 14516
rect 18597 14514 18663 14517
rect 16684 14512 18663 14514
rect 16684 14456 18602 14512
rect 18658 14456 18663 14512
rect 16684 14454 18663 14456
rect 16684 14452 16690 14454
rect 18597 14451 18663 14454
rect 20529 14514 20595 14517
rect 25497 14514 25563 14517
rect 46381 14514 46447 14517
rect 20529 14512 46447 14514
rect 20529 14456 20534 14512
rect 20590 14456 25502 14512
rect 25558 14456 46386 14512
rect 46442 14456 46447 14512
rect 20529 14454 46447 14456
rect 20529 14451 20595 14454
rect 25497 14451 25563 14454
rect 46381 14451 46447 14454
rect 6637 14378 6703 14381
rect 7281 14378 7347 14381
rect 7925 14378 7991 14381
rect 6637 14376 7347 14378
rect 6637 14320 6642 14376
rect 6698 14320 7286 14376
rect 7342 14320 7347 14376
rect 6637 14318 7347 14320
rect 6637 14315 6703 14318
rect 7281 14315 7347 14318
rect 7560 14376 7991 14378
rect 7560 14320 7930 14376
rect 7986 14320 7991 14376
rect 7560 14318 7991 14320
rect 0 14242 800 14272
rect 1301 14242 1367 14245
rect 0 14240 1367 14242
rect 0 14184 1306 14240
rect 1362 14184 1367 14240
rect 0 14182 1367 14184
rect 0 14152 800 14182
rect 1301 14179 1367 14182
rect 3601 14242 3667 14245
rect 7281 14242 7347 14245
rect 3601 14240 7347 14242
rect 3601 14184 3606 14240
rect 3662 14184 7286 14240
rect 7342 14184 7347 14240
rect 3601 14182 7347 14184
rect 3601 14179 3667 14182
rect 7281 14179 7347 14182
rect 7560 14109 7620 14318
rect 7925 14315 7991 14318
rect 8334 14316 8340 14380
rect 8404 14378 8410 14380
rect 8477 14378 8543 14381
rect 8404 14376 8543 14378
rect 8404 14320 8482 14376
rect 8538 14320 8543 14376
rect 8404 14318 8543 14320
rect 8404 14316 8410 14318
rect 8477 14315 8543 14318
rect 9029 14378 9095 14381
rect 9949 14378 10015 14381
rect 10869 14378 10935 14381
rect 9029 14376 10935 14378
rect 9029 14320 9034 14376
rect 9090 14320 9954 14376
rect 10010 14320 10874 14376
rect 10930 14320 10935 14376
rect 9029 14318 10935 14320
rect 9029 14315 9095 14318
rect 9949 14315 10015 14318
rect 10869 14315 10935 14318
rect 11881 14378 11947 14381
rect 13678 14378 13738 14451
rect 11881 14376 13738 14378
rect 11881 14320 11886 14376
rect 11942 14320 13738 14376
rect 11881 14318 13738 14320
rect 15285 14378 15351 14381
rect 20069 14378 20135 14381
rect 15285 14376 22110 14378
rect 15285 14320 15290 14376
rect 15346 14320 20074 14376
rect 20130 14320 22110 14376
rect 15285 14318 22110 14320
rect 11881 14315 11947 14318
rect 15285 14315 15351 14318
rect 20069 14315 20135 14318
rect 9806 14180 9812 14244
rect 9876 14242 9882 14244
rect 11278 14242 11284 14244
rect 9876 14182 11284 14242
rect 9876 14180 9882 14182
rect 11278 14180 11284 14182
rect 11348 14180 11354 14244
rect 11462 14180 11468 14244
rect 11532 14242 11538 14244
rect 16481 14242 16547 14245
rect 11532 14240 16547 14242
rect 11532 14184 16486 14240
rect 16542 14184 16547 14240
rect 11532 14182 16547 14184
rect 11532 14180 11538 14182
rect 16481 14179 16547 14182
rect 18505 14242 18571 14245
rect 19926 14242 19932 14244
rect 18505 14240 19932 14242
rect 18505 14184 18510 14240
rect 18566 14184 19932 14240
rect 18505 14182 19932 14184
rect 18505 14179 18571 14182
rect 19926 14180 19932 14182
rect 19996 14180 20002 14244
rect 22050 14242 22110 14318
rect 22318 14316 22324 14380
rect 22388 14378 22394 14380
rect 23841 14378 23907 14381
rect 22388 14376 23907 14378
rect 22388 14320 23846 14376
rect 23902 14320 23907 14376
rect 22388 14318 23907 14320
rect 22388 14316 22394 14318
rect 23841 14315 23907 14318
rect 24761 14378 24827 14381
rect 46565 14378 46631 14381
rect 24761 14376 46631 14378
rect 24761 14320 24766 14376
rect 24822 14320 46570 14376
rect 46626 14320 46631 14376
rect 24761 14318 46631 14320
rect 24761 14315 24827 14318
rect 46565 14315 46631 14318
rect 25681 14242 25747 14245
rect 22050 14240 25747 14242
rect 22050 14184 25686 14240
rect 25742 14184 25747 14240
rect 22050 14182 25747 14184
rect 25681 14179 25747 14182
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 4705 14106 4771 14109
rect 4981 14106 5047 14109
rect 6545 14108 6611 14109
rect 4705 14104 5047 14106
rect 4705 14048 4710 14104
rect 4766 14048 4986 14104
rect 5042 14048 5047 14104
rect 4705 14046 5047 14048
rect 4705 14043 4771 14046
rect 4981 14043 5047 14046
rect 6494 14044 6500 14108
rect 6564 14106 6611 14108
rect 6564 14104 6656 14106
rect 6606 14048 6656 14104
rect 6564 14046 6656 14048
rect 7557 14104 7623 14109
rect 7557 14048 7562 14104
rect 7618 14048 7623 14104
rect 6564 14044 6611 14046
rect 6545 14043 6611 14044
rect 7557 14043 7623 14048
rect 8477 14106 8543 14109
rect 9070 14106 9076 14108
rect 8477 14104 9076 14106
rect 8477 14048 8482 14104
rect 8538 14048 9076 14104
rect 8477 14046 9076 14048
rect 8477 14043 8543 14046
rect 9070 14044 9076 14046
rect 9140 14044 9146 14108
rect 11053 14106 11119 14109
rect 16665 14106 16731 14109
rect 11053 14104 16731 14106
rect 11053 14048 11058 14104
rect 11114 14048 16670 14104
rect 16726 14048 16731 14104
rect 11053 14046 16731 14048
rect 11053 14043 11119 14046
rect 16665 14043 16731 14046
rect 18822 14044 18828 14108
rect 18892 14106 18898 14108
rect 19793 14106 19859 14109
rect 18892 14104 19859 14106
rect 18892 14048 19798 14104
rect 19854 14048 19859 14104
rect 18892 14046 19859 14048
rect 18892 14044 18898 14046
rect 19793 14043 19859 14046
rect 21950 14044 21956 14108
rect 22020 14106 22026 14108
rect 25405 14106 25471 14109
rect 22020 14104 25471 14106
rect 22020 14048 25410 14104
rect 25466 14048 25471 14104
rect 22020 14046 25471 14048
rect 22020 14044 22026 14046
rect 25405 14043 25471 14046
rect 1577 13972 1643 13973
rect 1526 13908 1532 13972
rect 1596 13970 1643 13972
rect 1596 13968 1688 13970
rect 1638 13912 1688 13968
rect 1596 13910 1688 13912
rect 1596 13908 1643 13910
rect 7414 13908 7420 13972
rect 7484 13970 7490 13972
rect 7649 13970 7715 13973
rect 7484 13968 7715 13970
rect 7484 13912 7654 13968
rect 7710 13912 7715 13968
rect 7484 13910 7715 13912
rect 7484 13908 7490 13910
rect 1577 13907 1643 13908
rect 7649 13907 7715 13910
rect 7782 13908 7788 13972
rect 7852 13970 7858 13972
rect 8937 13970 9003 13973
rect 7852 13968 9003 13970
rect 7852 13912 8942 13968
rect 8998 13912 9003 13968
rect 7852 13910 9003 13912
rect 7852 13908 7858 13910
rect 8937 13907 9003 13910
rect 9673 13970 9739 13973
rect 12525 13970 12591 13973
rect 20897 13972 20963 13973
rect 9673 13968 12591 13970
rect 9673 13912 9678 13968
rect 9734 13912 12530 13968
rect 12586 13912 12591 13968
rect 9673 13910 12591 13912
rect 9673 13907 9739 13910
rect 12525 13907 12591 13910
rect 14774 13908 14780 13972
rect 14844 13970 14850 13972
rect 20846 13970 20852 13972
rect 14844 13910 18890 13970
rect 20806 13910 20852 13970
rect 20916 13968 20963 13972
rect 20958 13912 20963 13968
rect 14844 13908 14850 13910
rect 0 13834 800 13864
rect 2037 13834 2103 13837
rect 0 13832 2103 13834
rect 0 13776 2042 13832
rect 2098 13776 2103 13832
rect 0 13774 2103 13776
rect 0 13744 800 13774
rect 2037 13771 2103 13774
rect 3509 13834 3575 13837
rect 7465 13834 7531 13837
rect 18689 13834 18755 13837
rect 3509 13832 18755 13834
rect 3509 13776 3514 13832
rect 3570 13776 7470 13832
rect 7526 13776 18694 13832
rect 18750 13776 18755 13832
rect 3509 13774 18755 13776
rect 3509 13771 3575 13774
rect 7465 13771 7531 13774
rect 18689 13771 18755 13774
rect 3785 13698 3851 13701
rect 7598 13698 7604 13700
rect 3785 13696 7604 13698
rect 3785 13640 3790 13696
rect 3846 13640 7604 13696
rect 3785 13638 7604 13640
rect 3785 13635 3851 13638
rect 7598 13636 7604 13638
rect 7668 13636 7674 13700
rect 7833 13698 7899 13701
rect 11278 13698 11284 13700
rect 7833 13696 11284 13698
rect 7833 13640 7838 13696
rect 7894 13640 11284 13696
rect 7833 13638 11284 13640
rect 7833 13635 7899 13638
rect 11278 13636 11284 13638
rect 11348 13636 11354 13700
rect 11421 13698 11487 13701
rect 12566 13698 12572 13700
rect 11421 13696 12572 13698
rect 11421 13640 11426 13696
rect 11482 13640 12572 13696
rect 11421 13638 12572 13640
rect 11421 13635 11487 13638
rect 12566 13636 12572 13638
rect 12636 13636 12642 13700
rect 15878 13636 15884 13700
rect 15948 13698 15954 13700
rect 16665 13698 16731 13701
rect 18638 13698 18644 13700
rect 15948 13638 16498 13698
rect 15948 13636 15954 13638
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 4245 13562 4311 13565
rect 7046 13562 7052 13564
rect 4245 13560 7052 13562
rect 4245 13504 4250 13560
rect 4306 13504 7052 13560
rect 4245 13502 7052 13504
rect 4245 13499 4311 13502
rect 7046 13500 7052 13502
rect 7116 13500 7122 13564
rect 7373 13562 7439 13565
rect 11145 13562 11211 13565
rect 7373 13560 11211 13562
rect 7373 13504 7378 13560
rect 7434 13504 11150 13560
rect 11206 13504 11211 13560
rect 7373 13502 11211 13504
rect 7373 13499 7439 13502
rect 11145 13499 11211 13502
rect 15510 13500 15516 13564
rect 15580 13562 15586 13564
rect 16297 13562 16363 13565
rect 15580 13560 16363 13562
rect 15580 13504 16302 13560
rect 16358 13504 16363 13560
rect 15580 13502 16363 13504
rect 16438 13562 16498 13638
rect 16665 13696 18644 13698
rect 16665 13640 16670 13696
rect 16726 13640 18644 13696
rect 16665 13638 18644 13640
rect 16665 13635 16731 13638
rect 18638 13636 18644 13638
rect 18708 13636 18714 13700
rect 18830 13698 18890 13910
rect 20846 13908 20852 13910
rect 20916 13908 20963 13912
rect 20897 13907 20963 13908
rect 21449 13970 21515 13973
rect 22461 13970 22527 13973
rect 21449 13968 22527 13970
rect 21449 13912 21454 13968
rect 21510 13912 22466 13968
rect 22522 13912 22527 13968
rect 21449 13910 22527 13912
rect 21449 13907 21515 13910
rect 22461 13907 22527 13910
rect 22645 13970 22711 13973
rect 23790 13970 23796 13972
rect 22645 13968 23796 13970
rect 22645 13912 22650 13968
rect 22706 13912 23796 13968
rect 22645 13910 23796 13912
rect 22645 13907 22711 13910
rect 23790 13908 23796 13910
rect 23860 13908 23866 13972
rect 21081 13834 21147 13837
rect 22553 13834 22619 13837
rect 25129 13834 25195 13837
rect 25405 13834 25471 13837
rect 21081 13832 22619 13834
rect 21081 13776 21086 13832
rect 21142 13776 22558 13832
rect 22614 13776 22619 13832
rect 21081 13774 22619 13776
rect 21081 13771 21147 13774
rect 22553 13771 22619 13774
rect 22694 13774 23490 13834
rect 19793 13698 19859 13701
rect 18830 13696 19859 13698
rect 18830 13640 19798 13696
rect 19854 13640 19859 13696
rect 18830 13638 19859 13640
rect 19793 13635 19859 13638
rect 20713 13698 20779 13701
rect 22134 13698 22140 13700
rect 20713 13696 22140 13698
rect 20713 13640 20718 13696
rect 20774 13640 22140 13696
rect 20713 13638 22140 13640
rect 20713 13635 20779 13638
rect 22134 13636 22140 13638
rect 22204 13636 22210 13700
rect 16573 13562 16639 13565
rect 16438 13560 16639 13562
rect 16438 13504 16578 13560
rect 16634 13504 16639 13560
rect 16438 13502 16639 13504
rect 15580 13500 15586 13502
rect 16297 13499 16363 13502
rect 16573 13499 16639 13502
rect 16849 13562 16915 13565
rect 22694 13562 22754 13774
rect 23430 13698 23490 13774
rect 25129 13832 25471 13834
rect 25129 13776 25134 13832
rect 25190 13776 25410 13832
rect 25466 13776 25471 13832
rect 25129 13774 25471 13776
rect 25129 13771 25195 13774
rect 25405 13771 25471 13774
rect 27889 13698 27955 13701
rect 23430 13696 27955 13698
rect 23430 13640 27894 13696
rect 27950 13640 27955 13696
rect 23430 13638 27955 13640
rect 27889 13635 27955 13638
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 31937 13562 32003 13565
rect 16849 13560 22754 13562
rect 16849 13504 16854 13560
rect 16910 13504 22754 13560
rect 16849 13502 22754 13504
rect 31710 13560 32003 13562
rect 31710 13504 31942 13560
rect 31998 13504 32003 13560
rect 31710 13502 32003 13504
rect 16849 13499 16915 13502
rect 0 13426 800 13456
rect 1117 13426 1183 13429
rect 0 13424 1183 13426
rect 0 13368 1122 13424
rect 1178 13368 1183 13424
rect 0 13366 1183 13368
rect 0 13336 800 13366
rect 1117 13363 1183 13366
rect 3785 13426 3851 13429
rect 4248 13426 4308 13499
rect 8201 13426 8267 13429
rect 3785 13424 4308 13426
rect 3785 13368 3790 13424
rect 3846 13368 4308 13424
rect 3785 13366 4308 13368
rect 6686 13424 8267 13426
rect 6686 13368 8206 13424
rect 8262 13368 8267 13424
rect 6686 13366 8267 13368
rect 3785 13363 3851 13366
rect 1342 13228 1348 13292
rect 1412 13290 1418 13292
rect 1577 13290 1643 13293
rect 1412 13288 1643 13290
rect 1412 13232 1582 13288
rect 1638 13232 1643 13288
rect 1412 13230 1643 13232
rect 1412 13228 1418 13230
rect 1577 13227 1643 13230
rect 3509 13290 3575 13293
rect 6686 13290 6746 13366
rect 8201 13363 8267 13366
rect 8937 13426 9003 13429
rect 9489 13426 9555 13429
rect 8937 13424 9555 13426
rect 8937 13368 8942 13424
rect 8998 13368 9494 13424
rect 9550 13368 9555 13424
rect 8937 13366 9555 13368
rect 8937 13363 9003 13366
rect 9489 13363 9555 13366
rect 9765 13426 9831 13429
rect 11094 13426 11100 13428
rect 9765 13424 11100 13426
rect 9765 13368 9770 13424
rect 9826 13368 11100 13424
rect 9765 13366 11100 13368
rect 9765 13363 9831 13366
rect 11094 13364 11100 13366
rect 11164 13364 11170 13428
rect 11881 13426 11947 13429
rect 15837 13426 15903 13429
rect 31710 13426 31770 13502
rect 31937 13499 32003 13502
rect 11881 13424 15762 13426
rect 11881 13368 11886 13424
rect 11942 13368 15762 13424
rect 11881 13366 15762 13368
rect 11881 13363 11947 13366
rect 3509 13288 6746 13290
rect 3509 13232 3514 13288
rect 3570 13232 6746 13288
rect 3509 13230 6746 13232
rect 7189 13290 7255 13293
rect 15702 13290 15762 13366
rect 15837 13424 31770 13426
rect 15837 13368 15842 13424
rect 15898 13368 31770 13424
rect 15837 13366 31770 13368
rect 15837 13363 15903 13366
rect 18689 13290 18755 13293
rect 18873 13290 18939 13293
rect 7189 13288 15394 13290
rect 7189 13232 7194 13288
rect 7250 13232 15394 13288
rect 7189 13230 15394 13232
rect 15702 13230 18522 13290
rect 3509 13227 3575 13230
rect 7189 13227 7255 13230
rect 2865 13154 2931 13157
rect 7373 13154 7439 13157
rect 2865 13152 7439 13154
rect 2865 13096 2870 13152
rect 2926 13096 7378 13152
rect 7434 13096 7439 13152
rect 2865 13094 7439 13096
rect 2865 13091 2931 13094
rect 7373 13091 7439 13094
rect 9070 13092 9076 13156
rect 9140 13154 9146 13156
rect 9765 13154 9831 13157
rect 9140 13152 9831 13154
rect 9140 13096 9770 13152
rect 9826 13096 9831 13152
rect 9140 13094 9831 13096
rect 9140 13092 9146 13094
rect 9765 13091 9831 13094
rect 10777 13154 10843 13157
rect 12750 13154 12756 13156
rect 10777 13152 12756 13154
rect 10777 13096 10782 13152
rect 10838 13096 12756 13152
rect 10777 13094 12756 13096
rect 10777 13091 10843 13094
rect 12750 13092 12756 13094
rect 12820 13092 12826 13156
rect 15334 13154 15394 13230
rect 16205 13154 16271 13157
rect 15334 13152 16271 13154
rect 15334 13096 16210 13152
rect 16266 13096 16271 13152
rect 15334 13094 16271 13096
rect 16205 13091 16271 13094
rect 16481 13154 16547 13157
rect 17769 13154 17835 13157
rect 16481 13152 17835 13154
rect 16481 13096 16486 13152
rect 16542 13096 17774 13152
rect 17830 13096 17835 13152
rect 16481 13094 17835 13096
rect 18462 13154 18522 13230
rect 18689 13288 18939 13290
rect 18689 13232 18694 13288
rect 18750 13232 18878 13288
rect 18934 13232 18939 13288
rect 18689 13230 18939 13232
rect 18689 13227 18755 13230
rect 18873 13227 18939 13230
rect 19241 13290 19307 13293
rect 28901 13290 28967 13293
rect 19241 13288 28967 13290
rect 19241 13232 19246 13288
rect 19302 13232 28906 13288
rect 28962 13232 28967 13288
rect 19241 13230 28967 13232
rect 19241 13227 19307 13230
rect 28901 13227 28967 13230
rect 19333 13154 19399 13157
rect 18462 13152 19399 13154
rect 18462 13096 19338 13152
rect 19394 13096 19399 13152
rect 18462 13094 19399 13096
rect 16481 13091 16547 13094
rect 17769 13091 17835 13094
rect 19333 13091 19399 13094
rect 20662 13092 20668 13156
rect 20732 13154 20738 13156
rect 20732 13094 26986 13154
rect 20732 13092 20738 13094
rect 7946 13088 8262 13089
rect 0 13018 800 13048
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 2865 13018 2931 13021
rect 0 13016 2931 13018
rect 0 12960 2870 13016
rect 2926 12960 2931 13016
rect 0 12958 2931 12960
rect 0 12928 800 12958
rect 2865 12955 2931 12958
rect 3233 13018 3299 13021
rect 6729 13018 6795 13021
rect 3233 13016 6795 13018
rect 3233 12960 3238 13016
rect 3294 12960 6734 13016
rect 6790 12960 6795 13016
rect 3233 12958 6795 12960
rect 3233 12955 3299 12958
rect 6729 12955 6795 12958
rect 7046 12956 7052 13020
rect 7116 13018 7122 13020
rect 7281 13018 7347 13021
rect 7116 13016 7347 13018
rect 7116 12960 7286 13016
rect 7342 12960 7347 13016
rect 7116 12958 7347 12960
rect 7116 12956 7122 12958
rect 7281 12955 7347 12958
rect 9581 13018 9647 13021
rect 17718 13018 17724 13020
rect 9581 13016 17724 13018
rect 9581 12960 9586 13016
rect 9642 12960 17724 13016
rect 9581 12958 17724 12960
rect 9581 12955 9647 12958
rect 17718 12956 17724 12958
rect 17788 12956 17794 13020
rect 18454 12956 18460 13020
rect 18524 13018 18530 13020
rect 18689 13018 18755 13021
rect 18524 13016 18755 13018
rect 18524 12960 18694 13016
rect 18750 12960 18755 13016
rect 18524 12958 18755 12960
rect 18524 12956 18530 12958
rect 18689 12955 18755 12958
rect 19793 13018 19859 13021
rect 19793 13016 22110 13018
rect 19793 12960 19798 13016
rect 19854 12960 22110 13016
rect 19793 12958 22110 12960
rect 19793 12955 19859 12958
rect 5073 12882 5139 12885
rect 5574 12882 5580 12884
rect 5073 12880 5580 12882
rect 5073 12824 5078 12880
rect 5134 12824 5580 12880
rect 5073 12822 5580 12824
rect 5073 12819 5139 12822
rect 5574 12820 5580 12822
rect 5644 12820 5650 12884
rect 6545 12882 6611 12885
rect 11697 12882 11763 12885
rect 13905 12882 13971 12885
rect 6545 12880 11763 12882
rect 6545 12824 6550 12880
rect 6606 12824 11702 12880
rect 11758 12824 11763 12880
rect 6545 12822 11763 12824
rect 6545 12819 6611 12822
rect 11697 12819 11763 12822
rect 12390 12880 13971 12882
rect 12390 12824 13910 12880
rect 13966 12824 13971 12880
rect 12390 12822 13971 12824
rect 10542 12746 10548 12748
rect 2730 12686 10548 12746
rect 0 12610 800 12640
rect 2730 12610 2790 12686
rect 10542 12684 10548 12686
rect 10612 12684 10618 12748
rect 12390 12746 12450 12822
rect 13905 12819 13971 12822
rect 16430 12820 16436 12884
rect 16500 12882 16506 12884
rect 21398 12882 21404 12884
rect 16500 12822 21404 12882
rect 16500 12820 16506 12822
rect 21398 12820 21404 12822
rect 21468 12820 21474 12884
rect 22050 12882 22110 12958
rect 22686 12956 22692 13020
rect 22756 13018 22762 13020
rect 24894 13018 24900 13020
rect 22756 12958 24900 13018
rect 22756 12956 22762 12958
rect 24894 12956 24900 12958
rect 24964 12956 24970 13020
rect 26926 12882 26986 13094
rect 28942 13092 28948 13156
rect 29012 13154 29018 13156
rect 30833 13154 30899 13157
rect 35249 13154 35315 13157
rect 29012 13152 35315 13154
rect 29012 13096 30838 13152
rect 30894 13096 35254 13152
rect 35310 13096 35315 13152
rect 29012 13094 35315 13096
rect 29012 13092 29018 13094
rect 30833 13091 30899 13094
rect 35249 13091 35315 13094
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 47946 13023 48262 13024
rect 39941 12882 40007 12885
rect 22050 12822 25514 12882
rect 26926 12880 40007 12882
rect 26926 12824 39946 12880
rect 40002 12824 40007 12880
rect 26926 12822 40007 12824
rect 10734 12686 12450 12746
rect 13169 12746 13235 12749
rect 25454 12746 25514 12822
rect 39941 12819 40007 12822
rect 28901 12746 28967 12749
rect 13169 12744 25330 12746
rect 13169 12688 13174 12744
rect 13230 12688 25330 12744
rect 13169 12686 25330 12688
rect 25454 12744 28967 12746
rect 25454 12688 28906 12744
rect 28962 12688 28967 12744
rect 25454 12686 28967 12688
rect 0 12550 2790 12610
rect 5073 12608 5139 12613
rect 5073 12552 5078 12608
rect 5134 12552 5139 12608
rect 0 12520 800 12550
rect 5073 12547 5139 12552
rect 6637 12610 6703 12613
rect 7230 12610 7236 12612
rect 6637 12608 7236 12610
rect 6637 12552 6642 12608
rect 6698 12552 7236 12608
rect 6637 12550 7236 12552
rect 6637 12547 6703 12550
rect 7230 12548 7236 12550
rect 7300 12548 7306 12612
rect 8201 12610 8267 12613
rect 10734 12610 10794 12686
rect 13169 12683 13235 12686
rect 8201 12608 10794 12610
rect 8201 12552 8206 12608
rect 8262 12552 10794 12608
rect 8201 12550 10794 12552
rect 11789 12610 11855 12613
rect 11789 12608 12634 12610
rect 11789 12552 11794 12608
rect 11850 12552 12634 12608
rect 11789 12550 12634 12552
rect 8201 12547 8267 12550
rect 11789 12547 11855 12550
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 3366 12412 3372 12476
rect 3436 12474 3442 12476
rect 3877 12474 3943 12477
rect 3436 12472 3943 12474
rect 3436 12416 3882 12472
rect 3938 12416 3943 12472
rect 3436 12414 3943 12416
rect 3436 12412 3442 12414
rect 3877 12411 3943 12414
rect 5076 12341 5136 12547
rect 5993 12474 6059 12477
rect 6361 12474 6427 12477
rect 5993 12472 6427 12474
rect 5993 12416 5998 12472
rect 6054 12416 6366 12472
rect 6422 12416 6427 12472
rect 5993 12414 6427 12416
rect 5993 12411 6059 12414
rect 6361 12411 6427 12414
rect 9254 12412 9260 12476
rect 9324 12474 9330 12476
rect 12198 12474 12204 12476
rect 9324 12414 12204 12474
rect 9324 12412 9330 12414
rect 12198 12412 12204 12414
rect 12268 12412 12274 12476
rect 3325 12340 3391 12341
rect 3325 12338 3372 12340
rect 3280 12336 3372 12338
rect 3280 12280 3330 12336
rect 3280 12278 3372 12280
rect 3325 12276 3372 12278
rect 3436 12276 3442 12340
rect 5073 12336 5139 12341
rect 5073 12280 5078 12336
rect 5134 12280 5139 12336
rect 3325 12275 3391 12276
rect 5073 12275 5139 12280
rect 6269 12338 6335 12341
rect 9581 12338 9647 12341
rect 6269 12336 9647 12338
rect 6269 12280 6274 12336
rect 6330 12280 9586 12336
rect 9642 12280 9647 12336
rect 6269 12278 9647 12280
rect 6269 12275 6335 12278
rect 9581 12275 9647 12278
rect 10726 12276 10732 12340
rect 10796 12338 10802 12340
rect 11237 12338 11303 12341
rect 10796 12336 11303 12338
rect 10796 12280 11242 12336
rect 11298 12280 11303 12336
rect 10796 12278 11303 12280
rect 12574 12338 12634 12550
rect 13670 12548 13676 12612
rect 13740 12610 13746 12612
rect 14406 12610 14412 12612
rect 13740 12550 14412 12610
rect 13740 12548 13746 12550
rect 14406 12548 14412 12550
rect 14476 12548 14482 12612
rect 14733 12608 14799 12613
rect 14733 12552 14738 12608
rect 14794 12552 14799 12608
rect 14733 12547 14799 12552
rect 16297 12610 16363 12613
rect 19558 12610 19564 12612
rect 16297 12608 19564 12610
rect 16297 12552 16302 12608
rect 16358 12552 19564 12608
rect 16297 12550 19564 12552
rect 16297 12547 16363 12550
rect 19558 12548 19564 12550
rect 19628 12548 19634 12612
rect 20897 12610 20963 12613
rect 21909 12610 21975 12613
rect 20897 12608 21975 12610
rect 20897 12552 20902 12608
rect 20958 12552 21914 12608
rect 21970 12552 21975 12608
rect 20897 12550 21975 12552
rect 20897 12547 20963 12550
rect 21909 12547 21975 12550
rect 22277 12612 22343 12613
rect 22277 12608 22324 12612
rect 22388 12610 22394 12612
rect 25270 12610 25330 12686
rect 28901 12683 28967 12686
rect 29821 12610 29887 12613
rect 22277 12552 22282 12608
rect 22277 12548 22324 12552
rect 22388 12550 22434 12610
rect 25270 12608 29887 12610
rect 25270 12552 29826 12608
rect 29882 12552 29887 12608
rect 25270 12550 29887 12552
rect 22388 12548 22394 12550
rect 22277 12547 22343 12548
rect 29821 12547 29887 12550
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 14736 12474 14796 12547
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 17953 12474 18019 12477
rect 14736 12472 18019 12474
rect 14736 12416 17958 12472
rect 18014 12416 18019 12472
rect 14736 12414 18019 12416
rect 17953 12411 18019 12414
rect 18137 12474 18203 12477
rect 18454 12474 18460 12476
rect 18137 12472 18460 12474
rect 18137 12416 18142 12472
rect 18198 12416 18460 12472
rect 18137 12414 18460 12416
rect 18137 12411 18203 12414
rect 18454 12412 18460 12414
rect 18524 12412 18530 12476
rect 18873 12474 18939 12477
rect 19190 12474 19196 12476
rect 18873 12472 19196 12474
rect 18873 12416 18878 12472
rect 18934 12416 19196 12472
rect 18873 12414 19196 12416
rect 18873 12411 18939 12414
rect 19190 12412 19196 12414
rect 19260 12412 19266 12476
rect 23841 12474 23907 12477
rect 26509 12474 26575 12477
rect 23841 12472 26575 12474
rect 23841 12416 23846 12472
rect 23902 12416 26514 12472
rect 26570 12416 26575 12472
rect 23841 12414 26575 12416
rect 23841 12411 23907 12414
rect 26509 12411 26575 12414
rect 15142 12338 15148 12340
rect 12574 12278 15148 12338
rect 10796 12276 10802 12278
rect 11237 12275 11303 12278
rect 15142 12276 15148 12278
rect 15212 12276 15218 12340
rect 16481 12338 16547 12341
rect 16798 12338 16804 12340
rect 16481 12336 16804 12338
rect 16481 12280 16486 12336
rect 16542 12280 16804 12336
rect 16481 12278 16804 12280
rect 16481 12275 16547 12278
rect 16798 12276 16804 12278
rect 16868 12276 16874 12340
rect 17718 12276 17724 12340
rect 17788 12338 17794 12340
rect 23289 12338 23355 12341
rect 17788 12336 23355 12338
rect 17788 12280 23294 12336
rect 23350 12280 23355 12336
rect 17788 12278 23355 12280
rect 17788 12276 17794 12278
rect 23289 12275 23355 12278
rect 23790 12276 23796 12340
rect 23860 12338 23866 12340
rect 30005 12338 30071 12341
rect 23860 12336 30071 12338
rect 23860 12280 30010 12336
rect 30066 12280 30071 12336
rect 23860 12278 30071 12280
rect 23860 12276 23866 12278
rect 30005 12275 30071 12278
rect 0 12202 800 12232
rect 1393 12202 1459 12205
rect 0 12200 1459 12202
rect 0 12144 1398 12200
rect 1454 12144 1459 12200
rect 0 12142 1459 12144
rect 0 12112 800 12142
rect 1393 12139 1459 12142
rect 4981 12202 5047 12205
rect 7465 12202 7531 12205
rect 4981 12200 7531 12202
rect 4981 12144 4986 12200
rect 5042 12144 7470 12200
rect 7526 12144 7531 12200
rect 4981 12142 7531 12144
rect 4981 12139 5047 12142
rect 7465 12139 7531 12142
rect 7598 12140 7604 12204
rect 7668 12202 7674 12204
rect 7668 12142 8402 12202
rect 7668 12140 7674 12142
rect 3693 12066 3759 12069
rect 6729 12066 6795 12069
rect 3693 12064 6795 12066
rect 3693 12008 3698 12064
rect 3754 12008 6734 12064
rect 6790 12008 6795 12064
rect 3693 12006 6795 12008
rect 3693 12003 3759 12006
rect 6729 12003 6795 12006
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 5165 11930 5231 11933
rect 5993 11930 6059 11933
rect 6269 11930 6335 11933
rect 5165 11928 5274 11930
rect 5165 11872 5170 11928
rect 5226 11872 5274 11928
rect 5165 11867 5274 11872
rect 5993 11928 6335 11930
rect 5993 11872 5998 11928
rect 6054 11872 6274 11928
rect 6330 11872 6335 11928
rect 5993 11870 6335 11872
rect 8342 11930 8402 12142
rect 8518 12140 8524 12204
rect 8588 12202 8594 12204
rect 23749 12202 23815 12205
rect 8588 12200 23815 12202
rect 8588 12144 23754 12200
rect 23810 12144 23815 12200
rect 8588 12142 23815 12144
rect 8588 12140 8594 12142
rect 23749 12139 23815 12142
rect 27286 12140 27292 12204
rect 27356 12202 27362 12204
rect 37457 12202 37523 12205
rect 27356 12200 37523 12202
rect 27356 12144 37462 12200
rect 37518 12144 37523 12200
rect 27356 12142 37523 12144
rect 27356 12140 27362 12142
rect 37457 12139 37523 12142
rect 9857 12068 9923 12069
rect 9806 12066 9812 12068
rect 9766 12006 9812 12066
rect 9876 12064 9923 12068
rect 9918 12008 9923 12064
rect 9806 12004 9812 12006
rect 9876 12004 9923 12008
rect 9857 12003 9923 12004
rect 11421 12066 11487 12069
rect 12382 12066 12388 12068
rect 11421 12064 12388 12066
rect 11421 12008 11426 12064
rect 11482 12008 12388 12064
rect 11421 12006 12388 12008
rect 11421 12003 11487 12006
rect 12382 12004 12388 12006
rect 12452 12004 12458 12068
rect 12566 12004 12572 12068
rect 12636 12004 12642 12068
rect 13537 12066 13603 12069
rect 13854 12066 13860 12068
rect 13537 12064 13860 12066
rect 13537 12008 13542 12064
rect 13598 12008 13860 12064
rect 13537 12006 13860 12008
rect 12433 11930 12499 11933
rect 8342 11928 12499 11930
rect 8342 11872 12438 11928
rect 12494 11872 12499 11928
rect 8342 11870 12499 11872
rect 12574 11930 12634 12004
rect 13537 12003 13603 12006
rect 13854 12004 13860 12006
rect 13924 12004 13930 12068
rect 15469 12066 15535 12069
rect 17769 12066 17835 12069
rect 15469 12064 17835 12066
rect 15469 12008 15474 12064
rect 15530 12008 17774 12064
rect 17830 12008 17835 12064
rect 15469 12006 17835 12008
rect 15469 12003 15535 12006
rect 17769 12003 17835 12006
rect 18597 12066 18663 12069
rect 19926 12066 19932 12068
rect 18597 12064 19932 12066
rect 18597 12008 18602 12064
rect 18658 12008 19932 12064
rect 18597 12006 19932 12008
rect 18597 12003 18663 12006
rect 19926 12004 19932 12006
rect 19996 12004 20002 12068
rect 20621 12066 20687 12069
rect 24669 12066 24735 12069
rect 20621 12064 24735 12066
rect 20621 12008 20626 12064
rect 20682 12008 24674 12064
rect 24730 12008 24735 12064
rect 20621 12006 24735 12008
rect 20621 12003 20687 12006
rect 24669 12003 24735 12006
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 13486 11930 13492 11932
rect 12574 11870 13492 11930
rect 5993 11867 6059 11870
rect 6269 11867 6335 11870
rect 12433 11867 12499 11870
rect 13486 11868 13492 11870
rect 13556 11868 13562 11932
rect 13905 11930 13971 11933
rect 13905 11928 14106 11930
rect 13905 11872 13910 11928
rect 13966 11872 14106 11928
rect 13905 11870 14106 11872
rect 13905 11867 13971 11870
rect 0 11794 800 11824
rect 3233 11794 3299 11797
rect 0 11792 3299 11794
rect 0 11736 3238 11792
rect 3294 11736 3299 11792
rect 0 11734 3299 11736
rect 5214 11794 5274 11867
rect 11237 11794 11303 11797
rect 5214 11792 11303 11794
rect 5214 11736 11242 11792
rect 11298 11736 11303 11792
rect 5214 11734 11303 11736
rect 0 11704 800 11734
rect 3233 11731 3299 11734
rect 11237 11731 11303 11734
rect 11421 11794 11487 11797
rect 11646 11794 11652 11796
rect 11421 11792 11652 11794
rect 11421 11736 11426 11792
rect 11482 11736 11652 11792
rect 11421 11734 11652 11736
rect 11421 11731 11487 11734
rect 11646 11732 11652 11734
rect 11716 11732 11722 11796
rect 12198 11732 12204 11796
rect 12268 11794 12274 11796
rect 13813 11794 13879 11797
rect 12268 11792 13879 11794
rect 12268 11736 13818 11792
rect 13874 11736 13879 11792
rect 12268 11734 13879 11736
rect 12268 11732 12274 11734
rect 13813 11731 13879 11734
rect 14046 11658 14106 11870
rect 14774 11868 14780 11932
rect 14844 11930 14850 11932
rect 15285 11930 15351 11933
rect 14844 11928 15351 11930
rect 14844 11872 15290 11928
rect 15346 11872 15351 11928
rect 14844 11870 15351 11872
rect 14844 11868 14850 11870
rect 15285 11867 15351 11870
rect 15837 11928 15903 11933
rect 15837 11872 15842 11928
rect 15898 11872 15903 11928
rect 15837 11867 15903 11872
rect 19241 11930 19307 11933
rect 20161 11930 20227 11933
rect 19241 11928 20227 11930
rect 19241 11872 19246 11928
rect 19302 11872 20166 11928
rect 20222 11872 20227 11928
rect 19241 11870 20227 11872
rect 19241 11867 19307 11870
rect 20161 11867 20227 11870
rect 21909 11930 21975 11933
rect 27797 11930 27863 11933
rect 21909 11928 27863 11930
rect 21909 11872 21914 11928
rect 21970 11872 27802 11928
rect 27858 11872 27863 11928
rect 21909 11870 27863 11872
rect 21909 11867 21975 11870
rect 27797 11867 27863 11870
rect 14365 11796 14431 11797
rect 14365 11794 14412 11796
rect 14320 11792 14412 11794
rect 14320 11736 14370 11792
rect 14320 11734 14412 11736
rect 14365 11732 14412 11734
rect 14476 11732 14482 11796
rect 14549 11794 14615 11797
rect 15840 11794 15900 11867
rect 14549 11792 15900 11794
rect 14549 11736 14554 11792
rect 14610 11736 15900 11792
rect 14549 11734 15900 11736
rect 16113 11794 16179 11797
rect 22829 11794 22895 11797
rect 16113 11792 22895 11794
rect 16113 11736 16118 11792
rect 16174 11736 22834 11792
rect 22890 11736 22895 11792
rect 16113 11734 22895 11736
rect 14365 11731 14431 11732
rect 14549 11731 14615 11734
rect 16113 11731 16179 11734
rect 22829 11731 22895 11734
rect 23289 11794 23355 11797
rect 30557 11794 30623 11797
rect 23289 11792 30623 11794
rect 23289 11736 23294 11792
rect 23350 11736 30562 11792
rect 30618 11736 30623 11792
rect 23289 11734 30623 11736
rect 23289 11731 23355 11734
rect 30557 11731 30623 11734
rect 22093 11658 22159 11661
rect 23197 11658 23263 11661
rect 2730 11598 13600 11658
rect 14046 11656 22159 11658
rect 14046 11600 22098 11656
rect 22154 11600 22159 11656
rect 14046 11598 22159 11600
rect 0 11386 800 11416
rect 2730 11386 2790 11598
rect 8886 11460 8892 11524
rect 8956 11522 8962 11524
rect 11513 11522 11579 11525
rect 8956 11520 11579 11522
rect 8956 11464 11518 11520
rect 11574 11464 11579 11520
rect 8956 11462 11579 11464
rect 8956 11460 8962 11462
rect 11513 11459 11579 11462
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 8569 11388 8635 11389
rect 0 11326 2790 11386
rect 0 11296 800 11326
rect 8518 11324 8524 11388
rect 8588 11386 8635 11388
rect 10961 11386 11027 11389
rect 11237 11386 11303 11389
rect 8588 11384 8680 11386
rect 8630 11328 8680 11384
rect 8588 11326 8680 11328
rect 8848 11384 11303 11386
rect 8848 11328 10966 11384
rect 11022 11328 11242 11384
rect 11298 11328 11303 11384
rect 8848 11326 11303 11328
rect 13540 11386 13600 11598
rect 22093 11595 22159 11598
rect 22740 11656 23263 11658
rect 22740 11600 23202 11656
rect 23258 11600 23263 11656
rect 22740 11598 23263 11600
rect 14181 11522 14247 11525
rect 19926 11522 19932 11524
rect 14181 11520 19932 11522
rect 14181 11464 14186 11520
rect 14242 11464 19932 11520
rect 14181 11462 19932 11464
rect 14181 11459 14247 11462
rect 19926 11460 19932 11462
rect 19996 11460 20002 11524
rect 20897 11522 20963 11525
rect 22740 11522 22800 11598
rect 23197 11595 23263 11598
rect 25078 11596 25084 11660
rect 25148 11658 25154 11660
rect 40953 11658 41019 11661
rect 25148 11656 41019 11658
rect 25148 11600 40958 11656
rect 41014 11600 41019 11656
rect 25148 11598 41019 11600
rect 25148 11596 25154 11598
rect 40953 11595 41019 11598
rect 20897 11520 22800 11522
rect 20897 11464 20902 11520
rect 20958 11464 22800 11520
rect 20897 11462 22800 11464
rect 23841 11522 23907 11525
rect 27337 11522 27403 11525
rect 23841 11520 27403 11522
rect 23841 11464 23846 11520
rect 23902 11464 27342 11520
rect 27398 11464 27403 11520
rect 23841 11462 27403 11464
rect 20897 11459 20963 11462
rect 23841 11459 23907 11462
rect 27337 11459 27403 11462
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 16389 11386 16455 11389
rect 13540 11384 16455 11386
rect 13540 11328 16394 11384
rect 16450 11328 16455 11384
rect 13540 11326 16455 11328
rect 8588 11324 8635 11326
rect 8569 11323 8635 11324
rect 3366 11188 3372 11252
rect 3436 11250 3442 11252
rect 3785 11250 3851 11253
rect 8848 11250 8908 11326
rect 10961 11323 11027 11326
rect 11237 11323 11303 11326
rect 16389 11323 16455 11326
rect 17166 11324 17172 11388
rect 17236 11386 17242 11388
rect 18873 11386 18939 11389
rect 17236 11384 18939 11386
rect 17236 11328 18878 11384
rect 18934 11328 18939 11384
rect 17236 11326 18939 11328
rect 17236 11324 17242 11326
rect 18873 11323 18939 11326
rect 3436 11248 8908 11250
rect 3436 11192 3790 11248
rect 3846 11192 8908 11248
rect 3436 11190 8908 11192
rect 3436 11188 3442 11190
rect 3785 11187 3851 11190
rect 9622 11188 9628 11252
rect 9692 11250 9698 11252
rect 10593 11250 10659 11253
rect 9692 11248 10659 11250
rect 9692 11192 10598 11248
rect 10654 11192 10659 11248
rect 9692 11190 10659 11192
rect 9692 11188 9698 11190
rect 10593 11187 10659 11190
rect 11513 11250 11579 11253
rect 13537 11250 13603 11253
rect 11513 11248 13603 11250
rect 11513 11192 11518 11248
rect 11574 11192 13542 11248
rect 13598 11192 13603 11248
rect 11513 11190 13603 11192
rect 11513 11187 11579 11190
rect 13537 11187 13603 11190
rect 13813 11250 13879 11253
rect 14774 11250 14780 11252
rect 13813 11248 14780 11250
rect 13813 11192 13818 11248
rect 13874 11192 14780 11248
rect 13813 11190 14780 11192
rect 13813 11187 13879 11190
rect 14774 11188 14780 11190
rect 14844 11188 14850 11252
rect 14917 11250 14983 11253
rect 27429 11250 27495 11253
rect 14917 11248 27495 11250
rect 14917 11192 14922 11248
rect 14978 11192 27434 11248
rect 27490 11192 27495 11248
rect 14917 11190 27495 11192
rect 14917 11187 14983 11190
rect 27429 11187 27495 11190
rect 1761 11116 1827 11117
rect 1710 11052 1716 11116
rect 1780 11114 1827 11116
rect 4797 11114 4863 11117
rect 6494 11114 6500 11116
rect 1780 11112 1872 11114
rect 1822 11056 1872 11112
rect 1780 11054 1872 11056
rect 4797 11112 6500 11114
rect 4797 11056 4802 11112
rect 4858 11056 6500 11112
rect 4797 11054 6500 11056
rect 1780 11052 1827 11054
rect 1761 11051 1827 11052
rect 4797 11051 4863 11054
rect 6494 11052 6500 11054
rect 6564 11052 6570 11116
rect 7925 11114 7991 11117
rect 12198 11114 12204 11116
rect 7925 11112 12204 11114
rect 7925 11056 7930 11112
rect 7986 11056 12204 11112
rect 7925 11054 12204 11056
rect 7925 11051 7991 11054
rect 12198 11052 12204 11054
rect 12268 11052 12274 11116
rect 12382 11052 12388 11116
rect 12452 11114 12458 11116
rect 13261 11114 13327 11117
rect 12452 11112 13327 11114
rect 12452 11056 13266 11112
rect 13322 11056 13327 11112
rect 12452 11054 13327 11056
rect 12452 11052 12458 11054
rect 13261 11051 13327 11054
rect 13670 11052 13676 11116
rect 13740 11114 13746 11116
rect 14774 11114 14780 11116
rect 13740 11054 14780 11114
rect 13740 11052 13746 11054
rect 14774 11052 14780 11054
rect 14844 11052 14850 11116
rect 16941 11114 17007 11117
rect 25405 11114 25471 11117
rect 16941 11112 25471 11114
rect 16941 11056 16946 11112
rect 17002 11056 25410 11112
rect 25466 11056 25471 11112
rect 16941 11054 25471 11056
rect 16941 11051 17007 11054
rect 25405 11051 25471 11054
rect 0 10978 800 11008
rect 7097 10980 7163 10981
rect 9857 10980 9923 10981
rect 0 10918 1042 10978
rect 0 10888 800 10918
rect 982 10842 1042 10918
rect 7046 10916 7052 10980
rect 7116 10978 7163 10980
rect 7116 10976 7208 10978
rect 7158 10920 7208 10976
rect 7116 10918 7208 10920
rect 7116 10916 7163 10918
rect 9806 10916 9812 10980
rect 9876 10978 9923 10980
rect 10041 10978 10107 10981
rect 11094 10978 11100 10980
rect 9876 10976 9968 10978
rect 9918 10920 9968 10976
rect 9876 10918 9968 10920
rect 10041 10976 11100 10978
rect 10041 10920 10046 10976
rect 10102 10920 11100 10976
rect 10041 10918 11100 10920
rect 9876 10916 9923 10918
rect 7097 10915 7163 10916
rect 9857 10915 9923 10916
rect 10041 10915 10107 10918
rect 11094 10916 11100 10918
rect 11164 10916 11170 10980
rect 13813 10978 13879 10981
rect 11838 10976 13879 10978
rect 11838 10920 13818 10976
rect 13874 10920 13879 10976
rect 11838 10918 13879 10920
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 1761 10842 1827 10845
rect 982 10840 1827 10842
rect 982 10784 1766 10840
rect 1822 10784 1827 10840
rect 982 10782 1827 10784
rect 1761 10779 1827 10782
rect 1945 10842 2011 10845
rect 2957 10842 3023 10845
rect 5574 10842 5580 10844
rect 1945 10840 2790 10842
rect 1945 10784 1950 10840
rect 2006 10784 2790 10840
rect 1945 10782 2790 10784
rect 1945 10779 2011 10782
rect 2730 10706 2790 10782
rect 2957 10840 5580 10842
rect 2957 10784 2962 10840
rect 3018 10784 5580 10840
rect 2957 10782 5580 10784
rect 2957 10779 3023 10782
rect 5574 10780 5580 10782
rect 5644 10842 5650 10844
rect 6545 10842 6611 10845
rect 5644 10840 6611 10842
rect 5644 10784 6550 10840
rect 6606 10784 6611 10840
rect 5644 10782 6611 10784
rect 5644 10780 5650 10782
rect 6545 10779 6611 10782
rect 8569 10842 8635 10845
rect 11838 10842 11898 10918
rect 13813 10915 13879 10918
rect 14038 10916 14044 10980
rect 14108 10978 14114 10980
rect 14549 10978 14615 10981
rect 14108 10976 14615 10978
rect 14108 10920 14554 10976
rect 14610 10920 14615 10976
rect 14108 10918 14615 10920
rect 14108 10916 14114 10918
rect 14549 10915 14615 10918
rect 18454 10916 18460 10980
rect 18524 10978 18530 10980
rect 18873 10978 18939 10981
rect 18524 10976 18939 10978
rect 18524 10920 18878 10976
rect 18934 10920 18939 10976
rect 18524 10918 18939 10920
rect 18524 10916 18530 10918
rect 18873 10915 18939 10918
rect 21582 10916 21588 10980
rect 21652 10978 21658 10980
rect 21950 10978 21956 10980
rect 21652 10918 21956 10978
rect 21652 10916 21658 10918
rect 21950 10916 21956 10918
rect 22020 10916 22026 10980
rect 22134 10916 22140 10980
rect 22204 10978 22210 10980
rect 24761 10978 24827 10981
rect 22204 10976 24827 10978
rect 22204 10920 24766 10976
rect 24822 10920 24827 10976
rect 22204 10918 24827 10920
rect 22204 10916 22210 10918
rect 24761 10915 24827 10918
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 8569 10840 11898 10842
rect 8569 10784 8574 10840
rect 8630 10784 11898 10840
rect 8569 10782 11898 10784
rect 8569 10779 8635 10782
rect 12198 10780 12204 10844
rect 12268 10842 12274 10844
rect 13813 10842 13879 10845
rect 14958 10842 14964 10844
rect 12268 10840 13879 10842
rect 12268 10784 13818 10840
rect 13874 10784 13879 10840
rect 12268 10782 13879 10784
rect 12268 10780 12274 10782
rect 13813 10779 13879 10782
rect 14046 10782 14964 10842
rect 8293 10706 8359 10709
rect 2730 10704 8359 10706
rect 2730 10648 8298 10704
rect 8354 10648 8359 10704
rect 2730 10646 8359 10648
rect 8293 10643 8359 10646
rect 10542 10644 10548 10708
rect 10612 10706 10618 10708
rect 14046 10706 14106 10782
rect 14958 10780 14964 10782
rect 15028 10780 15034 10844
rect 23381 10842 23447 10845
rect 27429 10844 27495 10845
rect 27429 10842 27476 10844
rect 19290 10840 23447 10842
rect 19290 10784 23386 10840
rect 23442 10784 23447 10840
rect 19290 10782 23447 10784
rect 27384 10840 27476 10842
rect 27384 10784 27434 10840
rect 27384 10782 27476 10784
rect 10612 10646 14106 10706
rect 14365 10706 14431 10709
rect 19290 10706 19350 10782
rect 23381 10779 23447 10782
rect 27429 10780 27476 10782
rect 27540 10780 27546 10844
rect 27429 10779 27495 10780
rect 14365 10704 19350 10706
rect 14365 10648 14370 10704
rect 14426 10648 19350 10704
rect 14365 10646 19350 10648
rect 10612 10644 10618 10646
rect 14365 10643 14431 10646
rect 21398 10644 21404 10708
rect 21468 10706 21474 10708
rect 34237 10706 34303 10709
rect 21468 10704 34303 10706
rect 21468 10648 34242 10704
rect 34298 10648 34303 10704
rect 21468 10646 34303 10648
rect 21468 10644 21474 10646
rect 34237 10643 34303 10646
rect 0 10570 800 10600
rect 1945 10570 2011 10573
rect 0 10568 2011 10570
rect 0 10512 1950 10568
rect 2006 10512 2011 10568
rect 0 10510 2011 10512
rect 0 10480 800 10510
rect 1945 10507 2011 10510
rect 3049 10570 3115 10573
rect 10409 10570 10475 10573
rect 3049 10568 10475 10570
rect 3049 10512 3054 10568
rect 3110 10512 10414 10568
rect 10470 10512 10475 10568
rect 3049 10510 10475 10512
rect 3049 10507 3115 10510
rect 10409 10507 10475 10510
rect 11145 10570 11211 10573
rect 11697 10570 11763 10573
rect 27153 10570 27219 10573
rect 41873 10570 41939 10573
rect 11145 10568 27219 10570
rect 11145 10512 11150 10568
rect 11206 10512 11702 10568
rect 11758 10512 27158 10568
rect 27214 10512 27219 10568
rect 11145 10510 27219 10512
rect 11145 10507 11211 10510
rect 11697 10507 11763 10510
rect 27153 10507 27219 10510
rect 31710 10568 41939 10570
rect 31710 10512 41878 10568
rect 41934 10512 41939 10568
rect 31710 10510 41939 10512
rect 4061 10434 4127 10437
rect 8385 10434 8451 10437
rect 4061 10432 8451 10434
rect 4061 10376 4066 10432
rect 4122 10376 8390 10432
rect 8446 10376 8451 10432
rect 4061 10374 8451 10376
rect 4061 10371 4127 10374
rect 8385 10371 8451 10374
rect 8845 10434 8911 10437
rect 12801 10434 12867 10437
rect 8845 10432 12867 10434
rect 8845 10376 8850 10432
rect 8906 10376 12806 10432
rect 12862 10376 12867 10432
rect 8845 10374 12867 10376
rect 8845 10371 8911 10374
rect 12801 10371 12867 10374
rect 13486 10372 13492 10436
rect 13556 10434 13562 10436
rect 13556 10374 14658 10434
rect 13556 10372 13562 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 6729 10298 6795 10301
rect 9949 10298 10015 10301
rect 6729 10296 10015 10298
rect 6729 10240 6734 10296
rect 6790 10240 9954 10296
rect 10010 10240 10015 10296
rect 6729 10238 10015 10240
rect 6729 10235 6795 10238
rect 9949 10235 10015 10238
rect 11237 10298 11303 10301
rect 11462 10298 11468 10300
rect 11237 10296 11468 10298
rect 11237 10240 11242 10296
rect 11298 10240 11468 10296
rect 11237 10238 11468 10240
rect 11237 10235 11303 10238
rect 11462 10236 11468 10238
rect 11532 10236 11538 10300
rect 12157 10298 12223 10301
rect 12382 10298 12388 10300
rect 12157 10296 12388 10298
rect 12157 10240 12162 10296
rect 12218 10240 12388 10296
rect 12157 10238 12388 10240
rect 12157 10235 12223 10238
rect 12382 10236 12388 10238
rect 12452 10236 12458 10300
rect 14038 10298 14044 10300
rect 13448 10238 14044 10298
rect 0 10162 800 10192
rect 2313 10162 2379 10165
rect 0 10160 2379 10162
rect 0 10104 2318 10160
rect 2374 10104 2379 10160
rect 0 10102 2379 10104
rect 0 10072 800 10102
rect 2313 10099 2379 10102
rect 3141 10162 3207 10165
rect 11094 10162 11100 10164
rect 3141 10160 11100 10162
rect 3141 10104 3146 10160
rect 3202 10104 11100 10160
rect 3141 10102 11100 10104
rect 3141 10099 3207 10102
rect 11094 10100 11100 10102
rect 11164 10100 11170 10164
rect 11973 10162 12039 10165
rect 13448 10162 13508 10238
rect 14038 10236 14044 10238
rect 14108 10236 14114 10300
rect 14598 10298 14658 10374
rect 14774 10372 14780 10436
rect 14844 10434 14850 10436
rect 14844 10374 20224 10434
rect 14844 10372 14850 10374
rect 18229 10298 18295 10301
rect 19977 10298 20043 10301
rect 14598 10296 20043 10298
rect 14598 10240 18234 10296
rect 18290 10240 19982 10296
rect 20038 10240 20043 10296
rect 14598 10238 20043 10240
rect 20164 10298 20224 10374
rect 20294 10372 20300 10436
rect 20364 10434 20370 10436
rect 20364 10374 22754 10434
rect 20364 10372 20370 10374
rect 20345 10298 20411 10301
rect 20164 10296 20411 10298
rect 20164 10240 20350 10296
rect 20406 10240 20411 10296
rect 20164 10238 20411 10240
rect 18229 10235 18295 10238
rect 19977 10235 20043 10238
rect 20345 10235 20411 10238
rect 11973 10160 13508 10162
rect 11973 10104 11978 10160
rect 12034 10104 13508 10160
rect 11973 10102 13508 10104
rect 13813 10162 13879 10165
rect 22277 10162 22343 10165
rect 13813 10160 22343 10162
rect 13813 10104 13818 10160
rect 13874 10104 22282 10160
rect 22338 10104 22343 10160
rect 13813 10102 22343 10104
rect 22694 10162 22754 10374
rect 24894 10372 24900 10436
rect 24964 10434 24970 10436
rect 31710 10434 31770 10510
rect 41873 10507 41939 10510
rect 24964 10374 31770 10434
rect 24964 10372 24970 10374
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 42946 10303 43262 10304
rect 24025 10298 24091 10301
rect 31385 10298 31451 10301
rect 24025 10296 31451 10298
rect 24025 10240 24030 10296
rect 24086 10240 31390 10296
rect 31446 10240 31451 10296
rect 24025 10238 31451 10240
rect 24025 10235 24091 10238
rect 31385 10235 31451 10238
rect 26141 10162 26207 10165
rect 22694 10160 26207 10162
rect 22694 10104 26146 10160
rect 26202 10104 26207 10160
rect 22694 10102 26207 10104
rect 11973 10099 12039 10102
rect 13813 10099 13879 10102
rect 22277 10099 22343 10102
rect 26141 10099 26207 10102
rect 4337 10026 4403 10029
rect 5942 10026 5948 10028
rect 4337 10024 5948 10026
rect 4337 9968 4342 10024
rect 4398 9968 5948 10024
rect 4337 9966 5948 9968
rect 4337 9963 4403 9966
rect 5942 9964 5948 9966
rect 6012 9964 6018 10028
rect 8334 10026 8340 10028
rect 7790 9966 8340 10026
rect 1945 9890 2011 9893
rect 5758 9890 5764 9892
rect 1945 9888 5764 9890
rect 1945 9832 1950 9888
rect 2006 9832 5764 9888
rect 1945 9830 5764 9832
rect 1945 9827 2011 9830
rect 5758 9828 5764 9830
rect 5828 9828 5834 9892
rect 7230 9828 7236 9892
rect 7300 9890 7306 9892
rect 7373 9890 7439 9893
rect 7790 9890 7850 9966
rect 8334 9964 8340 9966
rect 8404 9964 8410 10028
rect 9029 10026 9095 10029
rect 9397 10026 9463 10029
rect 9029 10024 9463 10026
rect 9029 9968 9034 10024
rect 9090 9968 9402 10024
rect 9458 9968 9463 10024
rect 9029 9966 9463 9968
rect 9029 9963 9095 9966
rect 9397 9963 9463 9966
rect 9765 10026 9831 10029
rect 10593 10026 10659 10029
rect 9765 10024 10659 10026
rect 9765 9968 9770 10024
rect 9826 9968 10598 10024
rect 10654 9968 10659 10024
rect 9765 9966 10659 9968
rect 9765 9963 9831 9966
rect 10593 9963 10659 9966
rect 12065 10026 12131 10029
rect 13813 10026 13879 10029
rect 14549 10028 14615 10029
rect 14549 10026 14596 10028
rect 12065 10024 13879 10026
rect 12065 9968 12070 10024
rect 12126 9968 13818 10024
rect 13874 9968 13879 10024
rect 12065 9966 13879 9968
rect 14508 10024 14596 10026
rect 14660 10026 14666 10028
rect 15510 10026 15516 10028
rect 14508 9968 14554 10024
rect 14508 9966 14596 9968
rect 12065 9963 12131 9966
rect 13813 9963 13879 9966
rect 14549 9964 14596 9966
rect 14660 9966 15516 10026
rect 14660 9964 14666 9966
rect 15510 9964 15516 9966
rect 15580 9964 15586 10028
rect 17350 9964 17356 10028
rect 17420 10026 17426 10028
rect 18781 10026 18847 10029
rect 17420 10024 18847 10026
rect 17420 9968 18786 10024
rect 18842 9968 18847 10024
rect 17420 9966 18847 9968
rect 17420 9964 17426 9966
rect 14549 9963 14615 9964
rect 18781 9963 18847 9966
rect 19977 10026 20043 10029
rect 48957 10026 49023 10029
rect 19977 10024 49023 10026
rect 19977 9968 19982 10024
rect 20038 9968 48962 10024
rect 49018 9968 49023 10024
rect 19977 9966 49023 9968
rect 19977 9963 20043 9966
rect 48957 9963 49023 9966
rect 7300 9888 7850 9890
rect 7300 9832 7378 9888
rect 7434 9832 7850 9888
rect 7300 9830 7850 9832
rect 8342 9830 11346 9890
rect 7300 9828 7306 9830
rect 7373 9827 7439 9830
rect 7946 9824 8262 9825
rect 0 9754 800 9784
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 0 9694 7850 9754
rect 0 9664 800 9694
rect 1526 9556 1532 9620
rect 1596 9618 1602 9620
rect 1669 9618 1735 9621
rect 3785 9620 3851 9621
rect 3734 9618 3740 9620
rect 1596 9616 1735 9618
rect 1596 9560 1674 9616
rect 1730 9560 1735 9616
rect 1596 9558 1735 9560
rect 3694 9558 3740 9618
rect 3804 9616 3851 9620
rect 3846 9560 3851 9616
rect 1596 9556 1602 9558
rect 1669 9555 1735 9558
rect 3734 9556 3740 9558
rect 3804 9556 3851 9560
rect 3785 9555 3851 9556
rect 4245 9620 4311 9621
rect 4245 9616 4292 9620
rect 4356 9618 4362 9620
rect 5625 9618 5691 9621
rect 6637 9618 6703 9621
rect 4245 9560 4250 9616
rect 4245 9556 4292 9560
rect 4356 9558 4402 9618
rect 5625 9616 6703 9618
rect 5625 9560 5630 9616
rect 5686 9560 6642 9616
rect 6698 9560 6703 9616
rect 5625 9558 6703 9560
rect 4356 9556 4362 9558
rect 4245 9555 4311 9556
rect 5625 9555 5691 9558
rect 6637 9555 6703 9558
rect 7097 9618 7163 9621
rect 7598 9618 7604 9620
rect 7097 9616 7604 9618
rect 7097 9560 7102 9616
rect 7158 9560 7604 9616
rect 7097 9558 7604 9560
rect 7097 9555 7163 9558
rect 7598 9556 7604 9558
rect 7668 9556 7674 9620
rect 7790 9618 7850 9694
rect 8342 9618 8402 9830
rect 10409 9754 10475 9757
rect 11145 9754 11211 9757
rect 10409 9752 11211 9754
rect 10409 9696 10414 9752
rect 10470 9696 11150 9752
rect 11206 9696 11211 9752
rect 10409 9694 11211 9696
rect 11286 9754 11346 9830
rect 12014 9828 12020 9892
rect 12084 9890 12090 9892
rect 13486 9890 13492 9892
rect 12084 9830 13492 9890
rect 12084 9828 12090 9830
rect 13486 9828 13492 9830
rect 13556 9828 13562 9892
rect 14089 9890 14155 9893
rect 15694 9890 15700 9892
rect 14089 9888 15700 9890
rect 14089 9832 14094 9888
rect 14150 9832 15700 9888
rect 14089 9830 15700 9832
rect 14089 9827 14155 9830
rect 15694 9828 15700 9830
rect 15764 9828 15770 9892
rect 17401 9890 17467 9893
rect 17769 9890 17835 9893
rect 17401 9888 17835 9890
rect 17401 9832 17406 9888
rect 17462 9832 17774 9888
rect 17830 9832 17835 9888
rect 17401 9830 17835 9832
rect 17401 9827 17467 9830
rect 17769 9827 17835 9830
rect 18638 9828 18644 9892
rect 18708 9890 18714 9892
rect 18708 9830 21650 9890
rect 18708 9828 18714 9830
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 12341 9754 12407 9757
rect 13670 9754 13676 9756
rect 11286 9694 12266 9754
rect 10409 9691 10475 9694
rect 11145 9691 11211 9694
rect 7790 9558 8402 9618
rect 8845 9618 8911 9621
rect 10409 9618 10475 9621
rect 11881 9618 11947 9621
rect 8845 9616 11947 9618
rect 8845 9560 8850 9616
rect 8906 9560 10414 9616
rect 10470 9560 11886 9616
rect 11942 9560 11947 9616
rect 8845 9558 11947 9560
rect 12206 9618 12266 9694
rect 12341 9752 13676 9754
rect 12341 9696 12346 9752
rect 12402 9696 13676 9752
rect 12341 9694 13676 9696
rect 12341 9691 12407 9694
rect 13670 9692 13676 9694
rect 13740 9692 13746 9756
rect 19057 9754 19123 9757
rect 21398 9754 21404 9756
rect 19057 9752 21404 9754
rect 19057 9696 19062 9752
rect 19118 9696 21404 9752
rect 19057 9694 21404 9696
rect 19057 9691 19123 9694
rect 21398 9692 21404 9694
rect 21468 9692 21474 9756
rect 21590 9754 21650 9830
rect 21950 9828 21956 9892
rect 22020 9890 22026 9892
rect 27705 9890 27771 9893
rect 22020 9888 27771 9890
rect 22020 9832 27710 9888
rect 27766 9832 27771 9888
rect 22020 9830 27771 9832
rect 22020 9828 22026 9830
rect 27705 9827 27771 9830
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 22277 9754 22343 9757
rect 21590 9752 22343 9754
rect 21590 9696 22282 9752
rect 22338 9696 22343 9752
rect 21590 9694 22343 9696
rect 22277 9691 22343 9694
rect 12382 9618 12388 9620
rect 12206 9558 12388 9618
rect 8845 9555 8911 9558
rect 10409 9555 10475 9558
rect 11881 9555 11947 9558
rect 12382 9556 12388 9558
rect 12452 9556 12458 9620
rect 12525 9618 12591 9621
rect 14733 9618 14799 9621
rect 26233 9618 26299 9621
rect 12525 9616 12634 9618
rect 12525 9560 12530 9616
rect 12586 9560 12634 9616
rect 12525 9555 12634 9560
rect 14733 9616 26299 9618
rect 14733 9560 14738 9616
rect 14794 9560 26238 9616
rect 26294 9560 26299 9616
rect 14733 9558 26299 9560
rect 14733 9555 14799 9558
rect 26233 9555 26299 9558
rect 933 9482 999 9485
rect 2078 9482 2084 9484
rect 933 9480 2084 9482
rect 933 9424 938 9480
rect 994 9424 2084 9480
rect 933 9422 2084 9424
rect 933 9419 999 9422
rect 2078 9420 2084 9422
rect 2148 9420 2154 9484
rect 2957 9482 3023 9485
rect 4102 9482 4108 9484
rect 2957 9480 4108 9482
rect 2957 9424 2962 9480
rect 3018 9424 4108 9480
rect 2957 9422 4108 9424
rect 2957 9419 3023 9422
rect 4102 9420 4108 9422
rect 4172 9420 4178 9484
rect 5073 9482 5139 9485
rect 6821 9482 6887 9485
rect 5073 9480 6887 9482
rect 5073 9424 5078 9480
rect 5134 9424 6826 9480
rect 6882 9424 6887 9480
rect 5073 9422 6887 9424
rect 5073 9419 5139 9422
rect 6821 9419 6887 9422
rect 7557 9482 7623 9485
rect 12433 9482 12499 9485
rect 12574 9482 12634 9555
rect 7557 9480 11760 9482
rect 7557 9424 7562 9480
rect 7618 9424 11760 9480
rect 7557 9422 11760 9424
rect 7557 9419 7623 9422
rect 0 9346 800 9376
rect 11700 9349 11760 9422
rect 12433 9480 12634 9482
rect 12433 9424 12438 9480
rect 12494 9424 12634 9480
rect 12433 9422 12634 9424
rect 17401 9482 17467 9485
rect 19374 9482 19380 9484
rect 17401 9480 19380 9482
rect 17401 9424 17406 9480
rect 17462 9424 19380 9480
rect 17401 9422 19380 9424
rect 12433 9419 12499 9422
rect 17401 9419 17467 9422
rect 19374 9420 19380 9422
rect 19444 9420 19450 9484
rect 21030 9420 21036 9484
rect 21100 9482 21106 9484
rect 45185 9482 45251 9485
rect 21100 9480 45251 9482
rect 21100 9424 45190 9480
rect 45246 9424 45251 9480
rect 21100 9422 45251 9424
rect 21100 9420 21106 9422
rect 45185 9419 45251 9422
rect 1393 9346 1459 9349
rect 0 9344 1459 9346
rect 0 9288 1398 9344
rect 1454 9288 1459 9344
rect 0 9286 1459 9288
rect 0 9256 800 9286
rect 1393 9283 1459 9286
rect 6545 9346 6611 9349
rect 11462 9346 11468 9348
rect 6545 9344 11468 9346
rect 6545 9288 6550 9344
rect 6606 9288 11468 9344
rect 6545 9286 11468 9288
rect 6545 9283 6611 9286
rect 11462 9284 11468 9286
rect 11532 9284 11538 9348
rect 11697 9344 11763 9349
rect 14181 9348 14247 9349
rect 14181 9346 14228 9348
rect 11697 9288 11702 9344
rect 11758 9288 11763 9344
rect 11697 9283 11763 9288
rect 14136 9344 14228 9346
rect 14136 9288 14186 9344
rect 14136 9286 14228 9288
rect 14181 9284 14228 9286
rect 14292 9284 14298 9348
rect 16798 9284 16804 9348
rect 16868 9346 16874 9348
rect 17493 9346 17559 9349
rect 16868 9344 17559 9346
rect 16868 9288 17498 9344
rect 17554 9288 17559 9344
rect 16868 9286 17559 9288
rect 16868 9284 16874 9286
rect 14181 9283 14247 9284
rect 17493 9283 17559 9286
rect 17861 9346 17927 9349
rect 19609 9346 19675 9349
rect 17861 9344 19675 9346
rect 17861 9288 17866 9344
rect 17922 9288 19614 9344
rect 19670 9288 19675 9344
rect 17861 9286 19675 9288
rect 17861 9283 17927 9286
rect 19609 9283 19675 9286
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 6637 9210 6703 9213
rect 8385 9210 8451 9213
rect 6637 9208 8451 9210
rect 6637 9152 6642 9208
rect 6698 9152 8390 9208
rect 8446 9152 8451 9208
rect 6637 9150 8451 9152
rect 6637 9147 6703 9150
rect 8385 9147 8451 9150
rect 10225 9210 10291 9213
rect 11329 9210 11395 9213
rect 10225 9208 11395 9210
rect 10225 9152 10230 9208
rect 10286 9152 11334 9208
rect 11390 9152 11395 9208
rect 10225 9150 11395 9152
rect 10225 9147 10291 9150
rect 11329 9147 11395 9150
rect 11513 9210 11579 9213
rect 11646 9210 11652 9212
rect 11513 9208 11652 9210
rect 11513 9152 11518 9208
rect 11574 9152 11652 9208
rect 11513 9150 11652 9152
rect 11513 9147 11579 9150
rect 11646 9148 11652 9150
rect 11716 9148 11722 9212
rect 14917 9210 14983 9213
rect 16481 9210 16547 9213
rect 14917 9208 16547 9210
rect 14917 9152 14922 9208
rect 14978 9152 16486 9208
rect 16542 9152 16547 9208
rect 14917 9150 16547 9152
rect 14917 9147 14983 9150
rect 16481 9147 16547 9150
rect 17585 9210 17651 9213
rect 21081 9210 21147 9213
rect 17585 9208 21147 9210
rect 17585 9152 17590 9208
rect 17646 9152 21086 9208
rect 21142 9152 21147 9208
rect 17585 9150 21147 9152
rect 17585 9147 17651 9150
rect 21081 9147 21147 9150
rect 7782 9012 7788 9076
rect 7852 9074 7858 9076
rect 11973 9074 12039 9077
rect 15878 9074 15884 9076
rect 7852 9014 11852 9074
rect 7852 9012 7858 9014
rect 0 8938 800 8968
rect 3734 8938 3740 8940
rect 0 8878 3740 8938
rect 0 8848 800 8878
rect 3734 8876 3740 8878
rect 3804 8876 3810 8940
rect 10777 8938 10843 8941
rect 11513 8938 11579 8941
rect 7790 8936 11579 8938
rect 7790 8880 10782 8936
rect 10838 8880 11518 8936
rect 11574 8880 11579 8936
rect 7790 8878 11579 8880
rect 1577 8802 1643 8805
rect 7790 8802 7850 8878
rect 10777 8875 10843 8878
rect 11513 8875 11579 8878
rect 1577 8800 7850 8802
rect 1577 8744 1582 8800
rect 1638 8744 7850 8800
rect 1577 8742 7850 8744
rect 8845 8802 8911 8805
rect 9121 8802 9187 8805
rect 11145 8802 11211 8805
rect 8845 8800 11211 8802
rect 8845 8744 8850 8800
rect 8906 8744 9126 8800
rect 9182 8744 11150 8800
rect 11206 8744 11211 8800
rect 8845 8742 11211 8744
rect 11792 8802 11852 9014
rect 11973 9072 15884 9074
rect 11973 9016 11978 9072
rect 12034 9016 15884 9072
rect 11973 9014 15884 9016
rect 11973 9011 12039 9014
rect 15878 9012 15884 9014
rect 15948 9012 15954 9076
rect 22001 9074 22067 9077
rect 28349 9074 28415 9077
rect 22001 9072 28415 9074
rect 22001 9016 22006 9072
rect 22062 9016 28354 9072
rect 28410 9016 28415 9072
rect 22001 9014 28415 9016
rect 22001 9011 22067 9014
rect 28349 9011 28415 9014
rect 12198 8876 12204 8940
rect 12268 8938 12274 8940
rect 13261 8938 13327 8941
rect 12268 8936 13327 8938
rect 12268 8880 13266 8936
rect 13322 8880 13327 8936
rect 12268 8878 13327 8880
rect 12268 8876 12274 8878
rect 13261 8875 13327 8878
rect 13537 8938 13603 8941
rect 17585 8938 17651 8941
rect 13537 8936 17651 8938
rect 13537 8880 13542 8936
rect 13598 8880 17590 8936
rect 17646 8880 17651 8936
rect 13537 8878 17651 8880
rect 13537 8875 13603 8878
rect 17585 8875 17651 8878
rect 17861 8938 17927 8941
rect 29177 8938 29243 8941
rect 17861 8936 29243 8938
rect 17861 8880 17866 8936
rect 17922 8880 29182 8936
rect 29238 8880 29243 8936
rect 17861 8878 29243 8880
rect 17861 8875 17927 8878
rect 29177 8875 29243 8878
rect 11792 8742 14474 8802
rect 1577 8739 1643 8742
rect 8845 8739 8911 8742
rect 9121 8739 9187 8742
rect 11145 8739 11211 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 9673 8666 9739 8669
rect 9857 8666 9923 8669
rect 10041 8668 10107 8669
rect 9673 8664 9923 8666
rect 9673 8608 9678 8664
rect 9734 8608 9862 8664
rect 9918 8608 9923 8664
rect 9673 8606 9923 8608
rect 9673 8603 9739 8606
rect 9857 8603 9923 8606
rect 9990 8604 9996 8668
rect 10060 8666 10107 8668
rect 10060 8664 10152 8666
rect 10102 8608 10152 8664
rect 10060 8606 10152 8608
rect 10060 8604 10107 8606
rect 11094 8604 11100 8668
rect 11164 8666 11170 8668
rect 11164 8606 13922 8666
rect 11164 8604 11170 8606
rect 10041 8603 10107 8604
rect 0 8530 800 8560
rect 2630 8530 2636 8532
rect 0 8470 2636 8530
rect 0 8440 800 8470
rect 2630 8468 2636 8470
rect 2700 8468 2706 8532
rect 4245 8530 4311 8533
rect 9029 8530 9095 8533
rect 4245 8528 9095 8530
rect 4245 8472 4250 8528
rect 4306 8472 9034 8528
rect 9090 8472 9095 8528
rect 4245 8470 9095 8472
rect 4245 8467 4311 8470
rect 9029 8467 9095 8470
rect 9857 8530 9923 8533
rect 10961 8530 11027 8533
rect 9857 8528 11027 8530
rect 9857 8472 9862 8528
rect 9918 8472 10966 8528
rect 11022 8472 11027 8528
rect 9857 8470 11027 8472
rect 9857 8467 9923 8470
rect 10961 8467 11027 8470
rect 11237 8530 11303 8533
rect 13537 8530 13603 8533
rect 11237 8528 13603 8530
rect 11237 8472 11242 8528
rect 11298 8472 13542 8528
rect 13598 8472 13603 8528
rect 11237 8470 13603 8472
rect 13862 8530 13922 8606
rect 14089 8530 14155 8533
rect 13862 8528 14155 8530
rect 13862 8472 14094 8528
rect 14150 8472 14155 8528
rect 13862 8470 14155 8472
rect 11237 8467 11303 8470
rect 13537 8467 13603 8470
rect 14089 8467 14155 8470
rect 2957 8394 3023 8397
rect 5809 8394 5875 8397
rect 6637 8394 6703 8397
rect 2957 8392 5274 8394
rect 2957 8336 2962 8392
rect 3018 8336 5274 8392
rect 2957 8334 5274 8336
rect 2957 8331 3023 8334
rect 1342 8196 1348 8260
rect 1412 8258 1418 8260
rect 1485 8258 1551 8261
rect 1412 8256 1551 8258
rect 1412 8200 1490 8256
rect 1546 8200 1551 8256
rect 1412 8198 1551 8200
rect 1412 8196 1418 8198
rect 1485 8195 1551 8198
rect 4981 8260 5047 8261
rect 4981 8256 5028 8260
rect 5092 8258 5098 8260
rect 5214 8258 5274 8334
rect 5809 8392 6703 8394
rect 5809 8336 5814 8392
rect 5870 8336 6642 8392
rect 6698 8336 6703 8392
rect 5809 8334 6703 8336
rect 5809 8331 5875 8334
rect 6637 8331 6703 8334
rect 10041 8394 10107 8397
rect 10174 8394 10180 8396
rect 10041 8392 10180 8394
rect 10041 8336 10046 8392
rect 10102 8336 10180 8392
rect 10041 8334 10180 8336
rect 10041 8331 10107 8334
rect 10174 8332 10180 8334
rect 10244 8332 10250 8396
rect 10777 8394 10843 8397
rect 14181 8394 14247 8397
rect 10777 8392 14247 8394
rect 10777 8336 10782 8392
rect 10838 8336 14186 8392
rect 14242 8336 14247 8392
rect 10777 8334 14247 8336
rect 14414 8394 14474 8742
rect 20110 8740 20116 8804
rect 20180 8802 20186 8804
rect 25865 8802 25931 8805
rect 20180 8800 25931 8802
rect 20180 8744 25870 8800
rect 25926 8744 25931 8800
rect 20180 8742 25931 8744
rect 20180 8740 20186 8742
rect 25865 8739 25931 8742
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 16389 8668 16455 8669
rect 16389 8664 16436 8668
rect 16500 8666 16506 8668
rect 16389 8608 16394 8664
rect 16389 8604 16436 8608
rect 16500 8606 16546 8666
rect 16500 8604 16506 8606
rect 25262 8604 25268 8668
rect 25332 8666 25338 8668
rect 25957 8666 26023 8669
rect 25332 8664 26023 8666
rect 25332 8608 25962 8664
rect 26018 8608 26023 8664
rect 25332 8606 26023 8608
rect 25332 8604 25338 8606
rect 16389 8603 16455 8604
rect 25957 8603 26023 8606
rect 14641 8530 14707 8533
rect 33685 8530 33751 8533
rect 14641 8528 33751 8530
rect 14641 8472 14646 8528
rect 14702 8472 33690 8528
rect 33746 8472 33751 8528
rect 14641 8470 33751 8472
rect 14641 8467 14707 8470
rect 33685 8467 33751 8470
rect 18045 8394 18111 8397
rect 14414 8392 18111 8394
rect 14414 8336 18050 8392
rect 18106 8336 18111 8392
rect 14414 8334 18111 8336
rect 10777 8331 10843 8334
rect 14181 8331 14247 8334
rect 18045 8331 18111 8334
rect 19558 8332 19564 8396
rect 19628 8394 19634 8396
rect 39573 8394 39639 8397
rect 19628 8392 39639 8394
rect 19628 8336 39578 8392
rect 39634 8336 39639 8392
rect 19628 8334 39639 8336
rect 19628 8332 19634 8334
rect 39573 8331 39639 8334
rect 9121 8258 9187 8261
rect 4981 8200 4986 8256
rect 4981 8196 5028 8200
rect 5092 8198 5138 8258
rect 5214 8256 9187 8258
rect 5214 8200 9126 8256
rect 9182 8200 9187 8256
rect 5214 8198 9187 8200
rect 5092 8196 5098 8198
rect 4981 8195 5047 8196
rect 9121 8195 9187 8198
rect 10593 8258 10659 8261
rect 10910 8258 10916 8260
rect 10593 8256 10916 8258
rect 10593 8200 10598 8256
rect 10654 8200 10916 8256
rect 10593 8198 10916 8200
rect 10593 8195 10659 8198
rect 10910 8196 10916 8198
rect 10980 8196 10986 8260
rect 15510 8196 15516 8260
rect 15580 8258 15586 8260
rect 16113 8258 16179 8261
rect 15580 8256 16179 8258
rect 15580 8200 16118 8256
rect 16174 8200 16179 8256
rect 15580 8198 16179 8200
rect 15580 8196 15586 8198
rect 16113 8195 16179 8198
rect 2946 8192 3262 8193
rect 0 8122 800 8152
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 2313 8124 2379 8125
rect 0 8062 1410 8122
rect 0 8032 800 8062
rect 1350 7986 1410 8062
rect 2262 8060 2268 8124
rect 2332 8122 2379 8124
rect 4521 8122 4587 8125
rect 12157 8122 12223 8125
rect 2332 8120 2424 8122
rect 2374 8064 2424 8120
rect 2332 8062 2424 8064
rect 4521 8120 12223 8122
rect 4521 8064 4526 8120
rect 4582 8064 12162 8120
rect 12218 8064 12223 8120
rect 4521 8062 12223 8064
rect 2332 8060 2379 8062
rect 2313 8059 2379 8060
rect 4521 8059 4587 8062
rect 12157 8059 12223 8062
rect 13905 8122 13971 8125
rect 18822 8122 18828 8124
rect 13905 8120 18828 8122
rect 13905 8064 13910 8120
rect 13966 8064 18828 8120
rect 13905 8062 18828 8064
rect 13905 8059 13971 8062
rect 18822 8060 18828 8062
rect 18892 8060 18898 8124
rect 2405 7986 2471 7989
rect 1350 7984 2471 7986
rect 1350 7928 2410 7984
rect 2466 7928 2471 7984
rect 1350 7926 2471 7928
rect 2405 7923 2471 7926
rect 3734 7924 3740 7988
rect 3804 7986 3810 7988
rect 4797 7986 4863 7989
rect 3804 7984 4863 7986
rect 3804 7928 4802 7984
rect 4858 7928 4863 7984
rect 3804 7926 4863 7928
rect 3804 7924 3810 7926
rect 4797 7923 4863 7926
rect 5073 7986 5139 7989
rect 13486 7986 13492 7988
rect 5073 7984 13492 7986
rect 5073 7928 5078 7984
rect 5134 7928 13492 7984
rect 5073 7926 13492 7928
rect 5073 7923 5139 7926
rect 13486 7924 13492 7926
rect 13556 7986 13562 7988
rect 24853 7986 24919 7989
rect 13556 7984 24919 7986
rect 13556 7928 24858 7984
rect 24914 7928 24919 7984
rect 13556 7926 24919 7928
rect 13556 7924 13562 7926
rect 24853 7923 24919 7926
rect 7373 7850 7439 7853
rect 11329 7850 11395 7853
rect 27613 7850 27679 7853
rect 7373 7848 11395 7850
rect 7373 7792 7378 7848
rect 7434 7792 11334 7848
rect 11390 7792 11395 7848
rect 7373 7790 11395 7792
rect 7373 7787 7439 7790
rect 11329 7787 11395 7790
rect 11838 7848 27679 7850
rect 11838 7792 27618 7848
rect 27674 7792 27679 7848
rect 11838 7790 27679 7792
rect 0 7714 800 7744
rect 3509 7714 3575 7717
rect 0 7712 3575 7714
rect 0 7656 3514 7712
rect 3570 7656 3575 7712
rect 0 7654 3575 7656
rect 0 7624 800 7654
rect 3509 7651 3575 7654
rect 6821 7714 6887 7717
rect 7281 7714 7347 7717
rect 6821 7712 7347 7714
rect 6821 7656 6826 7712
rect 6882 7656 7286 7712
rect 7342 7656 7347 7712
rect 6821 7654 7347 7656
rect 6821 7651 6887 7654
rect 7281 7651 7347 7654
rect 11145 7714 11211 7717
rect 11278 7714 11284 7716
rect 11145 7712 11284 7714
rect 11145 7656 11150 7712
rect 11206 7656 11284 7712
rect 11145 7654 11284 7656
rect 11145 7651 11211 7654
rect 11278 7652 11284 7654
rect 11348 7652 11354 7716
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 1209 7578 1275 7581
rect 11237 7578 11303 7581
rect 11838 7578 11898 7790
rect 27613 7787 27679 7790
rect 12157 7714 12223 7717
rect 17585 7714 17651 7717
rect 12157 7712 17651 7714
rect 12157 7656 12162 7712
rect 12218 7656 17590 7712
rect 17646 7656 17651 7712
rect 12157 7654 17651 7656
rect 12157 7651 12223 7654
rect 17585 7651 17651 7654
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 47946 7583 48262 7584
rect 1209 7576 2790 7578
rect 1209 7520 1214 7576
rect 1270 7520 2790 7576
rect 1209 7518 2790 7520
rect 1209 7515 1275 7518
rect 2730 7442 2790 7518
rect 11237 7576 11898 7578
rect 11237 7520 11242 7576
rect 11298 7520 11898 7576
rect 11237 7518 11898 7520
rect 11237 7515 11303 7518
rect 12750 7516 12756 7580
rect 12820 7578 12826 7580
rect 12893 7578 12959 7581
rect 12820 7576 12959 7578
rect 12820 7520 12898 7576
rect 12954 7520 12959 7576
rect 12820 7518 12959 7520
rect 12820 7516 12826 7518
rect 12893 7515 12959 7518
rect 15142 7516 15148 7580
rect 15212 7578 15218 7580
rect 16757 7578 16823 7581
rect 21449 7580 21515 7581
rect 15212 7576 16823 7578
rect 15212 7520 16762 7576
rect 16818 7520 16823 7576
rect 15212 7518 16823 7520
rect 15212 7516 15218 7518
rect 16757 7515 16823 7518
rect 21398 7516 21404 7580
rect 21468 7578 21515 7580
rect 21468 7576 21560 7578
rect 21510 7520 21560 7576
rect 21468 7518 21560 7520
rect 21468 7516 21515 7518
rect 21449 7515 21515 7516
rect 5349 7442 5415 7445
rect 14273 7442 14339 7445
rect 29637 7442 29703 7445
rect 2730 7440 14339 7442
rect 2730 7384 5354 7440
rect 5410 7384 14278 7440
rect 14334 7384 14339 7440
rect 2730 7382 14339 7384
rect 5349 7379 5415 7382
rect 14273 7379 14339 7382
rect 14414 7440 29703 7442
rect 14414 7384 29642 7440
rect 29698 7384 29703 7440
rect 14414 7382 29703 7384
rect 0 7306 800 7336
rect 12157 7306 12223 7309
rect 13721 7306 13787 7309
rect 14414 7306 14474 7382
rect 29637 7379 29703 7382
rect 0 7304 12223 7306
rect 0 7248 12162 7304
rect 12218 7248 12223 7304
rect 0 7246 12223 7248
rect 0 7216 800 7246
rect 12157 7243 12223 7246
rect 12390 7246 13600 7306
rect 6729 7170 6795 7173
rect 7046 7170 7052 7172
rect 6729 7168 7052 7170
rect 6729 7112 6734 7168
rect 6790 7112 7052 7168
rect 6729 7110 7052 7112
rect 6729 7107 6795 7110
rect 7046 7108 7052 7110
rect 7116 7170 7122 7172
rect 10041 7170 10107 7173
rect 7116 7168 10107 7170
rect 7116 7112 10046 7168
rect 10102 7112 10107 7168
rect 7116 7110 10107 7112
rect 7116 7108 7122 7110
rect 10041 7107 10107 7110
rect 12157 7172 12223 7173
rect 12157 7168 12204 7172
rect 12268 7170 12274 7172
rect 12157 7112 12162 7168
rect 12157 7108 12204 7112
rect 12268 7110 12314 7170
rect 12268 7108 12274 7110
rect 12157 7107 12223 7108
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 4102 6972 4108 7036
rect 4172 7034 4178 7036
rect 4429 7034 4495 7037
rect 12390 7034 12450 7246
rect 13540 7170 13600 7246
rect 13721 7304 14474 7306
rect 13721 7248 13726 7304
rect 13782 7248 14474 7304
rect 13721 7246 14474 7248
rect 18321 7306 18387 7309
rect 24393 7306 24459 7309
rect 18321 7304 24459 7306
rect 18321 7248 18326 7304
rect 18382 7248 24398 7304
rect 24454 7248 24459 7304
rect 18321 7246 24459 7248
rect 13721 7243 13787 7246
rect 18321 7243 18387 7246
rect 24393 7243 24459 7246
rect 19701 7170 19767 7173
rect 13540 7168 19767 7170
rect 13540 7112 19706 7168
rect 19762 7112 19767 7168
rect 13540 7110 19767 7112
rect 19701 7107 19767 7110
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 4172 7032 12450 7034
rect 4172 6976 4434 7032
rect 4490 6976 12450 7032
rect 4172 6974 12450 6976
rect 4172 6972 4178 6974
rect 4429 6971 4495 6974
rect 0 6898 800 6928
rect 22185 6898 22251 6901
rect 0 6896 22251 6898
rect 0 6840 22190 6896
rect 22246 6840 22251 6896
rect 0 6838 22251 6840
rect 0 6808 800 6838
rect 22185 6835 22251 6838
rect 23289 6898 23355 6901
rect 38377 6898 38443 6901
rect 23289 6896 38443 6898
rect 23289 6840 23294 6896
rect 23350 6840 38382 6896
rect 38438 6840 38443 6896
rect 23289 6838 38443 6840
rect 23289 6835 23355 6838
rect 38377 6835 38443 6838
rect 1761 6764 1827 6765
rect 1710 6762 1716 6764
rect 1670 6702 1716 6762
rect 1780 6760 1827 6764
rect 1822 6704 1827 6760
rect 1710 6700 1716 6702
rect 1780 6700 1827 6704
rect 1761 6699 1827 6700
rect 2129 6762 2195 6765
rect 6729 6762 6795 6765
rect 9029 6764 9095 6765
rect 9029 6762 9076 6764
rect 2129 6760 6795 6762
rect 2129 6704 2134 6760
rect 2190 6704 6734 6760
rect 6790 6704 6795 6760
rect 2129 6702 6795 6704
rect 8984 6760 9076 6762
rect 8984 6704 9034 6760
rect 8984 6702 9076 6704
rect 2129 6699 2195 6702
rect 6729 6699 6795 6702
rect 9029 6700 9076 6702
rect 9140 6700 9146 6764
rect 10225 6762 10291 6765
rect 10869 6762 10935 6765
rect 10225 6760 10935 6762
rect 10225 6704 10230 6760
rect 10286 6704 10874 6760
rect 10930 6704 10935 6760
rect 10225 6702 10935 6704
rect 9029 6699 9095 6700
rect 10225 6699 10291 6702
rect 10869 6699 10935 6702
rect 11830 6700 11836 6764
rect 11900 6762 11906 6764
rect 12065 6762 12131 6765
rect 11900 6760 12131 6762
rect 11900 6704 12070 6760
rect 12126 6704 12131 6760
rect 11900 6702 12131 6704
rect 11900 6700 11906 6702
rect 12065 6699 12131 6702
rect 12433 6762 12499 6765
rect 13445 6762 13511 6765
rect 12433 6760 13511 6762
rect 12433 6704 12438 6760
rect 12494 6704 13450 6760
rect 13506 6704 13511 6760
rect 12433 6702 13511 6704
rect 12433 6699 12499 6702
rect 13445 6699 13511 6702
rect 15193 6762 15259 6765
rect 15326 6762 15332 6764
rect 15193 6760 15332 6762
rect 15193 6704 15198 6760
rect 15254 6704 15332 6760
rect 15193 6702 15332 6704
rect 15193 6699 15259 6702
rect 15326 6700 15332 6702
rect 15396 6700 15402 6764
rect 15469 6762 15535 6765
rect 19701 6764 19767 6765
rect 15469 6760 19626 6762
rect 15469 6704 15474 6760
rect 15530 6704 19626 6760
rect 15469 6702 19626 6704
rect 15469 6699 15535 6702
rect 1894 6564 1900 6628
rect 1964 6626 1970 6628
rect 3509 6626 3575 6629
rect 7414 6626 7420 6628
rect 1964 6624 3575 6626
rect 1964 6568 3514 6624
rect 3570 6568 3575 6624
rect 1964 6566 3575 6568
rect 1964 6564 1970 6566
rect 3509 6563 3575 6566
rect 5076 6566 7420 6626
rect 0 6490 800 6520
rect 3233 6490 3299 6493
rect 5076 6490 5136 6566
rect 7414 6564 7420 6566
rect 7484 6626 7490 6628
rect 7741 6626 7807 6629
rect 7484 6624 7807 6626
rect 7484 6568 7746 6624
rect 7802 6568 7807 6624
rect 7484 6566 7807 6568
rect 7484 6564 7490 6566
rect 7741 6563 7807 6566
rect 10225 6626 10291 6629
rect 13629 6626 13695 6629
rect 10225 6624 13695 6626
rect 10225 6568 10230 6624
rect 10286 6568 13634 6624
rect 13690 6568 13695 6624
rect 10225 6566 13695 6568
rect 10225 6563 10291 6566
rect 13629 6563 13695 6566
rect 14089 6626 14155 6629
rect 15745 6626 15811 6629
rect 14089 6624 15811 6626
rect 14089 6568 14094 6624
rect 14150 6568 15750 6624
rect 15806 6568 15811 6624
rect 14089 6566 15811 6568
rect 19566 6626 19626 6702
rect 19701 6760 19748 6764
rect 19812 6762 19818 6764
rect 34053 6762 34119 6765
rect 19701 6704 19706 6760
rect 19701 6700 19748 6704
rect 19812 6702 19858 6762
rect 22050 6760 34119 6762
rect 22050 6704 34058 6760
rect 34114 6704 34119 6760
rect 22050 6702 34119 6704
rect 19812 6700 19818 6702
rect 19701 6699 19767 6700
rect 22050 6626 22110 6702
rect 34053 6699 34119 6702
rect 19566 6566 22110 6626
rect 14089 6563 14155 6566
rect 15745 6563 15811 6566
rect 7946 6560 8262 6561
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 0 6430 2790 6490
rect 0 6400 800 6430
rect 2730 6354 2790 6430
rect 3233 6488 5136 6490
rect 3233 6432 3238 6488
rect 3294 6432 5136 6488
rect 3233 6430 5136 6432
rect 3233 6427 3299 6430
rect 5206 6428 5212 6492
rect 5276 6490 5282 6492
rect 7741 6490 7807 6493
rect 5276 6488 7807 6490
rect 5276 6432 7746 6488
rect 7802 6432 7807 6488
rect 5276 6430 7807 6432
rect 5276 6428 5282 6430
rect 7741 6427 7807 6430
rect 8385 6490 8451 6493
rect 9622 6490 9628 6492
rect 8385 6488 9628 6490
rect 8385 6432 8390 6488
rect 8446 6432 9628 6488
rect 8385 6430 9628 6432
rect 8385 6427 8451 6430
rect 9622 6428 9628 6430
rect 9692 6428 9698 6492
rect 10777 6490 10843 6493
rect 16665 6490 16731 6493
rect 10777 6488 16731 6490
rect 10777 6432 10782 6488
rect 10838 6432 16670 6488
rect 16726 6432 16731 6488
rect 10777 6430 16731 6432
rect 10777 6427 10843 6430
rect 16665 6427 16731 6430
rect 4153 6354 4219 6357
rect 2730 6352 4219 6354
rect 2730 6296 4158 6352
rect 4214 6296 4219 6352
rect 2730 6294 4219 6296
rect 4153 6291 4219 6294
rect 4613 6354 4679 6357
rect 5717 6354 5783 6357
rect 4613 6352 6194 6354
rect 4613 6296 4618 6352
rect 4674 6296 5722 6352
rect 5778 6296 6194 6352
rect 4613 6294 6194 6296
rect 4613 6291 4679 6294
rect 5717 6291 5783 6294
rect 1158 6156 1164 6220
rect 1228 6218 1234 6220
rect 5533 6218 5599 6221
rect 1228 6216 5599 6218
rect 1228 6160 5538 6216
rect 5594 6160 5599 6216
rect 1228 6158 5599 6160
rect 6134 6218 6194 6294
rect 6310 6292 6316 6356
rect 6380 6354 6386 6356
rect 7925 6354 7991 6357
rect 6380 6352 7991 6354
rect 6380 6296 7930 6352
rect 7986 6296 7991 6352
rect 6380 6294 7991 6296
rect 6380 6292 6386 6294
rect 7925 6291 7991 6294
rect 9673 6354 9739 6357
rect 18321 6354 18387 6357
rect 9673 6352 18387 6354
rect 9673 6296 9678 6352
rect 9734 6296 18326 6352
rect 18382 6296 18387 6352
rect 9673 6294 18387 6296
rect 9673 6291 9739 6294
rect 18321 6291 18387 6294
rect 23197 6354 23263 6357
rect 29494 6354 29500 6356
rect 23197 6352 29500 6354
rect 23197 6296 23202 6352
rect 23258 6296 29500 6352
rect 23197 6294 29500 6296
rect 23197 6291 23263 6294
rect 29494 6292 29500 6294
rect 29564 6292 29570 6356
rect 8845 6218 8911 6221
rect 6134 6216 8911 6218
rect 6134 6160 8850 6216
rect 8906 6160 8911 6216
rect 6134 6158 8911 6160
rect 1228 6156 1234 6158
rect 5533 6155 5599 6158
rect 8845 6155 8911 6158
rect 9029 6218 9095 6221
rect 10174 6218 10180 6220
rect 9029 6216 10180 6218
rect 9029 6160 9034 6216
rect 9090 6160 10180 6216
rect 9029 6158 10180 6160
rect 9029 6155 9095 6158
rect 10174 6156 10180 6158
rect 10244 6156 10250 6220
rect 11329 6218 11395 6221
rect 19333 6218 19399 6221
rect 11329 6216 19399 6218
rect 11329 6160 11334 6216
rect 11390 6160 19338 6216
rect 19394 6160 19399 6216
rect 11329 6158 19399 6160
rect 11329 6155 11395 6158
rect 19333 6155 19399 6158
rect 0 6082 800 6112
rect 1301 6082 1367 6085
rect 0 6080 1367 6082
rect 0 6024 1306 6080
rect 1362 6024 1367 6080
rect 0 6022 1367 6024
rect 0 5992 800 6022
rect 1301 6019 1367 6022
rect 3785 6082 3851 6085
rect 6085 6082 6151 6085
rect 3785 6080 6151 6082
rect 3785 6024 3790 6080
rect 3846 6024 6090 6080
rect 6146 6024 6151 6080
rect 3785 6022 6151 6024
rect 3785 6019 3851 6022
rect 6085 6019 6151 6022
rect 6361 6082 6427 6085
rect 6862 6082 6868 6084
rect 6361 6080 6868 6082
rect 6361 6024 6366 6080
rect 6422 6024 6868 6080
rect 6361 6022 6868 6024
rect 6361 6019 6427 6022
rect 6862 6020 6868 6022
rect 6932 6082 6938 6084
rect 12709 6082 12775 6085
rect 6932 6080 12775 6082
rect 6932 6024 12714 6080
rect 12770 6024 12775 6080
rect 6932 6022 12775 6024
rect 6932 6020 6938 6022
rect 12709 6019 12775 6022
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 5441 5946 5507 5949
rect 6126 5946 6132 5948
rect 5441 5944 6132 5946
rect 606 5850 612 5914
rect 676 5912 682 5914
rect 676 5852 1042 5912
rect 5441 5888 5446 5944
rect 5502 5888 6132 5944
rect 5441 5886 6132 5888
rect 5441 5883 5507 5886
rect 6126 5884 6132 5886
rect 6196 5884 6202 5948
rect 7598 5884 7604 5948
rect 7668 5946 7674 5948
rect 10225 5946 10291 5949
rect 11605 5948 11671 5949
rect 11605 5946 11652 5948
rect 7668 5944 10291 5946
rect 7668 5888 10230 5944
rect 10286 5888 10291 5944
rect 7668 5886 10291 5888
rect 11560 5944 11652 5946
rect 11560 5888 11610 5944
rect 11560 5886 11652 5888
rect 7668 5884 7674 5886
rect 10225 5883 10291 5886
rect 11605 5884 11652 5886
rect 11716 5884 11722 5948
rect 11605 5883 11671 5884
rect 676 5850 682 5852
rect 982 5810 1042 5852
rect 7833 5810 7899 5813
rect 982 5808 7899 5810
rect 982 5752 7838 5808
rect 7894 5752 7899 5808
rect 982 5750 7899 5752
rect 7833 5747 7899 5750
rect 12709 5810 12775 5813
rect 13854 5810 13860 5812
rect 12709 5808 13860 5810
rect 12709 5752 12714 5808
rect 12770 5752 13860 5808
rect 12709 5750 13860 5752
rect 12709 5747 12775 5750
rect 13854 5748 13860 5750
rect 13924 5748 13930 5812
rect 14958 5748 14964 5812
rect 15028 5810 15034 5812
rect 15929 5810 15995 5813
rect 15028 5808 15995 5810
rect 15028 5752 15934 5808
rect 15990 5752 15995 5808
rect 15028 5750 15995 5752
rect 15028 5748 15034 5750
rect 15929 5747 15995 5750
rect 16430 5748 16436 5812
rect 16500 5810 16506 5812
rect 19241 5810 19307 5813
rect 16500 5808 19307 5810
rect 16500 5752 19246 5808
rect 19302 5752 19307 5808
rect 16500 5750 19307 5752
rect 16500 5748 16506 5750
rect 19241 5747 19307 5750
rect 0 5674 800 5704
rect 1301 5674 1367 5677
rect 0 5672 1367 5674
rect 0 5616 1306 5672
rect 1362 5616 1367 5672
rect 0 5614 1367 5616
rect 0 5584 800 5614
rect 1301 5611 1367 5614
rect 6085 5674 6151 5677
rect 11329 5674 11395 5677
rect 6085 5672 11395 5674
rect 6085 5616 6090 5672
rect 6146 5616 11334 5672
rect 11390 5616 11395 5672
rect 6085 5614 11395 5616
rect 6085 5611 6151 5614
rect 11329 5611 11395 5614
rect 11697 5674 11763 5677
rect 22502 5674 22508 5676
rect 11697 5672 22508 5674
rect 11697 5616 11702 5672
rect 11758 5616 22508 5672
rect 11697 5614 22508 5616
rect 11697 5611 11763 5614
rect 22502 5612 22508 5614
rect 22572 5612 22578 5676
rect 2589 5538 2655 5541
rect 6545 5538 6611 5541
rect 2589 5536 6611 5538
rect 2589 5480 2594 5536
rect 2650 5480 6550 5536
rect 6606 5480 6611 5536
rect 2589 5478 6611 5480
rect 2589 5475 2655 5478
rect 6545 5475 6611 5478
rect 11053 5538 11119 5541
rect 16614 5538 16620 5540
rect 11053 5536 16620 5538
rect 11053 5480 11058 5536
rect 11114 5480 16620 5536
rect 11053 5478 16620 5480
rect 11053 5475 11119 5478
rect 16614 5476 16620 5478
rect 16684 5476 16690 5540
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 974 5340 980 5404
rect 1044 5402 1050 5404
rect 5165 5402 5231 5405
rect 1044 5400 5231 5402
rect 1044 5344 5170 5400
rect 5226 5344 5231 5400
rect 1044 5342 5231 5344
rect 1044 5340 1050 5342
rect 5165 5339 5231 5342
rect 5390 5340 5396 5404
rect 5460 5402 5466 5404
rect 7741 5402 7807 5405
rect 5460 5400 7807 5402
rect 5460 5344 7746 5400
rect 7802 5344 7807 5400
rect 5460 5342 7807 5344
rect 5460 5340 5466 5342
rect 7741 5339 7807 5342
rect 9990 5340 9996 5404
rect 10060 5402 10066 5404
rect 10060 5342 12450 5402
rect 10060 5340 10066 5342
rect 0 5266 800 5296
rect 1301 5266 1367 5269
rect 0 5264 1367 5266
rect 0 5208 1306 5264
rect 1362 5208 1367 5264
rect 0 5206 1367 5208
rect 0 5176 800 5206
rect 1301 5203 1367 5206
rect 2957 5266 3023 5269
rect 11697 5266 11763 5269
rect 2957 5264 11763 5266
rect 2957 5208 2962 5264
rect 3018 5208 11702 5264
rect 11758 5208 11763 5264
rect 2957 5206 11763 5208
rect 12390 5266 12450 5342
rect 19977 5266 20043 5269
rect 12390 5264 20043 5266
rect 12390 5208 19982 5264
rect 20038 5208 20043 5264
rect 12390 5206 20043 5208
rect 2957 5203 3023 5206
rect 11697 5203 11763 5206
rect 19977 5203 20043 5206
rect 6269 5130 6335 5133
rect 9949 5130 10015 5133
rect 2730 5070 3388 5130
rect 0 4858 800 4888
rect 1485 4858 1551 4861
rect 0 4856 1551 4858
rect 0 4800 1490 4856
rect 1546 4800 1551 4856
rect 0 4798 1551 4800
rect 0 4768 800 4798
rect 1485 4795 1551 4798
rect 2730 4725 2790 5070
rect 3328 4994 3388 5070
rect 6269 5128 10015 5130
rect 6269 5072 6274 5128
rect 6330 5072 9954 5128
rect 10010 5072 10015 5128
rect 6269 5070 10015 5072
rect 6269 5067 6335 5070
rect 9949 5067 10015 5070
rect 10961 5130 11027 5133
rect 12566 5130 12572 5132
rect 10961 5128 12572 5130
rect 10961 5072 10966 5128
rect 11022 5072 12572 5128
rect 10961 5070 12572 5072
rect 10961 5067 11027 5070
rect 12566 5068 12572 5070
rect 12636 5068 12642 5132
rect 18321 5130 18387 5133
rect 43345 5130 43411 5133
rect 12758 5070 18154 5130
rect 10726 4994 10732 4996
rect 3328 4934 10732 4994
rect 10726 4932 10732 4934
rect 10796 4932 10802 4996
rect 12382 4932 12388 4996
rect 12452 4994 12458 4996
rect 12758 4994 12818 5070
rect 12452 4934 12818 4994
rect 18094 4994 18154 5070
rect 18321 5128 43411 5130
rect 18321 5072 18326 5128
rect 18382 5072 43350 5128
rect 43406 5072 43411 5128
rect 18321 5070 43411 5072
rect 18321 5067 18387 5070
rect 43345 5067 43411 5070
rect 18873 4994 18939 4997
rect 18094 4992 18939 4994
rect 18094 4936 18878 4992
rect 18934 4936 18939 4992
rect 18094 4934 18939 4936
rect 12452 4932 12458 4934
rect 18873 4931 18939 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 42946 4863 43262 4864
rect 6453 4858 6519 4861
rect 9397 4858 9463 4861
rect 6453 4856 9463 4858
rect 6453 4800 6458 4856
rect 6514 4800 9402 4856
rect 9458 4800 9463 4856
rect 6453 4798 9463 4800
rect 6453 4795 6519 4798
rect 9397 4795 9463 4798
rect 2681 4720 2790 4725
rect 2681 4664 2686 4720
rect 2742 4664 2790 4720
rect 2681 4662 2790 4664
rect 3141 4722 3207 4725
rect 3550 4722 3556 4724
rect 3141 4720 3556 4722
rect 3141 4664 3146 4720
rect 3202 4664 3556 4720
rect 3141 4662 3556 4664
rect 2681 4659 2747 4662
rect 3141 4659 3207 4662
rect 3550 4660 3556 4662
rect 3620 4660 3626 4724
rect 5533 4722 5599 4725
rect 17309 4722 17375 4725
rect 19006 4722 19012 4724
rect 5533 4720 17234 4722
rect 5533 4664 5538 4720
rect 5594 4664 17234 4720
rect 5533 4662 17234 4664
rect 5533 4659 5599 4662
rect 2957 4586 3023 4589
rect 9029 4586 9095 4589
rect 2957 4584 9095 4586
rect 2957 4528 2962 4584
rect 3018 4528 9034 4584
rect 9090 4528 9095 4584
rect 2957 4526 9095 4528
rect 2957 4523 3023 4526
rect 9029 4523 9095 4526
rect 11462 4524 11468 4588
rect 11532 4586 11538 4588
rect 13813 4586 13879 4589
rect 11532 4584 13879 4586
rect 11532 4528 13818 4584
rect 13874 4528 13879 4584
rect 11532 4526 13879 4528
rect 17174 4586 17234 4662
rect 17309 4720 19012 4722
rect 17309 4664 17314 4720
rect 17370 4664 19012 4720
rect 17309 4662 19012 4664
rect 17309 4659 17375 4662
rect 19006 4660 19012 4662
rect 19076 4660 19082 4724
rect 21766 4660 21772 4724
rect 21836 4722 21842 4724
rect 21909 4722 21975 4725
rect 21836 4720 21975 4722
rect 21836 4664 21914 4720
rect 21970 4664 21975 4720
rect 21836 4662 21975 4664
rect 21836 4660 21842 4662
rect 21909 4659 21975 4662
rect 26141 4586 26207 4589
rect 17174 4584 26207 4586
rect 17174 4528 26146 4584
rect 26202 4528 26207 4584
rect 17174 4526 26207 4528
rect 11532 4524 11538 4526
rect 13813 4523 13879 4526
rect 26141 4523 26207 4526
rect 0 4450 800 4480
rect 3693 4450 3759 4453
rect 0 4448 3759 4450
rect 0 4392 3698 4448
rect 3754 4392 3759 4448
rect 0 4390 3759 4392
rect 0 4360 800 4390
rect 3693 4387 3759 4390
rect 9673 4450 9739 4453
rect 17309 4450 17375 4453
rect 9673 4448 17375 4450
rect 9673 4392 9678 4448
rect 9734 4392 17314 4448
rect 17370 4392 17375 4448
rect 9673 4390 17375 4392
rect 9673 4387 9739 4390
rect 17309 4387 17375 4390
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 12433 4314 12499 4317
rect 16982 4314 16988 4316
rect 12433 4312 16988 4314
rect 12433 4256 12438 4312
rect 12494 4256 16988 4312
rect 12433 4254 16988 4256
rect 12433 4251 12499 4254
rect 16982 4252 16988 4254
rect 17052 4252 17058 4316
rect 5349 4178 5415 4181
rect 24342 4178 24348 4180
rect 5349 4176 24348 4178
rect 5349 4120 5354 4176
rect 5410 4120 24348 4176
rect 5349 4118 24348 4120
rect 5349 4115 5415 4118
rect 24342 4116 24348 4118
rect 24412 4116 24418 4180
rect 0 4042 800 4072
rect 3785 4042 3851 4045
rect 0 4040 3851 4042
rect 0 3984 3790 4040
rect 3846 3984 3851 4040
rect 0 3982 3851 3984
rect 0 3952 800 3982
rect 3785 3979 3851 3982
rect 6545 4042 6611 4045
rect 9305 4044 9371 4045
rect 6678 4042 6684 4044
rect 6545 4040 6684 4042
rect 6545 3984 6550 4040
rect 6606 3984 6684 4040
rect 6545 3982 6684 3984
rect 6545 3979 6611 3982
rect 6678 3980 6684 3982
rect 6748 3980 6754 4044
rect 9254 3980 9260 4044
rect 9324 4042 9371 4044
rect 11145 4042 11211 4045
rect 9324 4040 9416 4042
rect 9366 3984 9416 4040
rect 9324 3982 9416 3984
rect 11145 4040 14106 4042
rect 11145 3984 11150 4040
rect 11206 3984 14106 4040
rect 11145 3982 14106 3984
rect 9324 3980 9371 3982
rect 9305 3979 9371 3980
rect 11145 3979 11211 3982
rect 5993 3906 6059 3909
rect 7230 3906 7236 3908
rect 5993 3904 7236 3906
rect 5993 3848 5998 3904
rect 6054 3848 7236 3904
rect 5993 3846 7236 3848
rect 5993 3843 6059 3846
rect 7230 3844 7236 3846
rect 7300 3844 7306 3908
rect 14046 3906 14106 3982
rect 14222 3980 14228 4044
rect 14292 4042 14298 4044
rect 15009 4042 15075 4045
rect 14292 4040 15075 4042
rect 14292 3984 15014 4040
rect 15070 3984 15075 4040
rect 14292 3982 15075 3984
rect 14292 3980 14298 3982
rect 15009 3979 15075 3982
rect 19333 4042 19399 4045
rect 24526 4042 24532 4044
rect 19333 4040 24532 4042
rect 19333 3984 19338 4040
rect 19394 3984 24532 4040
rect 19333 3982 24532 3984
rect 19333 3979 19399 3982
rect 24526 3980 24532 3982
rect 24596 3980 24602 4044
rect 18321 3906 18387 3909
rect 14046 3904 18387 3906
rect 14046 3848 18326 3904
rect 18382 3848 18387 3904
rect 14046 3846 18387 3848
rect 18321 3843 18387 3846
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 14549 3770 14615 3773
rect 22093 3770 22159 3773
rect 14549 3768 22159 3770
rect 14549 3712 14554 3768
rect 14610 3712 22098 3768
rect 22154 3712 22159 3768
rect 14549 3710 22159 3712
rect 14549 3707 14615 3710
rect 22093 3707 22159 3710
rect 0 3634 800 3664
rect 3601 3634 3667 3637
rect 0 3632 3667 3634
rect 0 3576 3606 3632
rect 3662 3576 3667 3632
rect 0 3574 3667 3576
rect 0 3544 800 3574
rect 3601 3571 3667 3574
rect 5809 3634 5875 3637
rect 15285 3634 15351 3637
rect 5809 3632 15351 3634
rect 5809 3576 5814 3632
rect 5870 3576 15290 3632
rect 15346 3576 15351 3632
rect 5809 3574 15351 3576
rect 5809 3571 5875 3574
rect 15285 3571 15351 3574
rect 20805 3634 20871 3637
rect 26182 3634 26188 3636
rect 20805 3632 26188 3634
rect 20805 3576 20810 3632
rect 20866 3576 26188 3632
rect 20805 3574 26188 3576
rect 20805 3571 20871 3574
rect 26182 3572 26188 3574
rect 26252 3572 26258 3636
rect 3049 3498 3115 3501
rect 8569 3498 8635 3501
rect 27613 3498 27679 3501
rect 3049 3496 8402 3498
rect 3049 3440 3054 3496
rect 3110 3440 8402 3496
rect 3049 3438 8402 3440
rect 3049 3435 3115 3438
rect 8342 3362 8402 3438
rect 8569 3496 27679 3498
rect 8569 3440 8574 3496
rect 8630 3440 27618 3496
rect 27674 3440 27679 3496
rect 8569 3438 27679 3440
rect 8569 3435 8635 3438
rect 27613 3435 27679 3438
rect 8342 3302 8770 3362
rect 7946 3296 8262 3297
rect 0 3226 800 3256
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 4061 3226 4127 3229
rect 8710 3228 8770 3302
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 0 3224 4127 3226
rect 0 3168 4066 3224
rect 4122 3168 4127 3224
rect 0 3166 4127 3168
rect 0 3136 800 3166
rect 4061 3163 4127 3166
rect 8702 3164 8708 3228
rect 8772 3226 8778 3228
rect 10869 3226 10935 3229
rect 8772 3224 10935 3226
rect 8772 3168 10874 3224
rect 10930 3168 10935 3224
rect 8772 3166 10935 3168
rect 8772 3164 8778 3166
rect 10869 3163 10935 3166
rect 13077 3226 13143 3229
rect 13353 3226 13419 3229
rect 13077 3224 15026 3226
rect 13077 3168 13082 3224
rect 13138 3168 13358 3224
rect 13414 3168 15026 3224
rect 13077 3166 15026 3168
rect 13077 3163 13143 3166
rect 13353 3163 13419 3166
rect 5257 3090 5323 3093
rect 14825 3090 14891 3093
rect 5257 3088 14891 3090
rect 5257 3032 5262 3088
rect 5318 3032 14830 3088
rect 14886 3032 14891 3088
rect 5257 3030 14891 3032
rect 14966 3090 15026 3166
rect 24710 3090 24716 3092
rect 14966 3030 24716 3090
rect 5257 3027 5323 3030
rect 14825 3027 14891 3030
rect 24710 3028 24716 3030
rect 24780 3028 24786 3092
rect 8753 2954 8819 2957
rect 32765 2954 32831 2957
rect 8753 2952 32831 2954
rect 8753 2896 8758 2952
rect 8814 2896 32770 2952
rect 32826 2896 32831 2952
rect 8753 2894 32831 2896
rect 8753 2891 8819 2894
rect 32765 2891 32831 2894
rect 0 2818 800 2848
rect 1577 2818 1643 2821
rect 0 2816 1643 2818
rect 0 2760 1582 2816
rect 1638 2760 1643 2816
rect 0 2758 1643 2760
rect 0 2728 800 2758
rect 1577 2755 1643 2758
rect 13353 2818 13419 2821
rect 13670 2818 13676 2820
rect 13353 2816 13676 2818
rect 13353 2760 13358 2816
rect 13414 2760 13676 2816
rect 13353 2758 13676 2760
rect 13353 2755 13419 2758
rect 13670 2756 13676 2758
rect 13740 2756 13746 2820
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 3325 2682 3391 2685
rect 8886 2682 8892 2684
rect 3325 2680 8892 2682
rect 3325 2624 3330 2680
rect 3386 2624 8892 2680
rect 3325 2622 8892 2624
rect 3325 2619 3391 2622
rect 8886 2620 8892 2622
rect 8956 2620 8962 2684
rect 9489 2682 9555 2685
rect 12433 2682 12499 2685
rect 9489 2680 12499 2682
rect 9489 2624 9494 2680
rect 9550 2624 12438 2680
rect 12494 2624 12499 2680
rect 9489 2622 12499 2624
rect 9489 2619 9555 2622
rect 12433 2619 12499 2622
rect 13445 2682 13511 2685
rect 13445 2680 17786 2682
rect 13445 2624 13450 2680
rect 13506 2624 17786 2680
rect 13445 2622 17786 2624
rect 13445 2619 13511 2622
rect 2773 2546 2839 2549
rect 17585 2546 17651 2549
rect 2773 2544 17651 2546
rect 2773 2488 2778 2544
rect 2834 2488 17590 2544
rect 17646 2488 17651 2544
rect 2773 2486 17651 2488
rect 17726 2546 17786 2622
rect 19926 2620 19932 2684
rect 19996 2682 20002 2684
rect 22001 2682 22067 2685
rect 19996 2680 22067 2682
rect 19996 2624 22006 2680
rect 22062 2624 22067 2680
rect 19996 2622 22067 2624
rect 19996 2620 20002 2622
rect 22001 2619 22067 2622
rect 23381 2682 23447 2685
rect 25814 2682 25820 2684
rect 23381 2680 25820 2682
rect 23381 2624 23386 2680
rect 23442 2624 25820 2680
rect 23381 2622 25820 2624
rect 23381 2619 23447 2622
rect 25814 2620 25820 2622
rect 25884 2620 25890 2684
rect 20161 2546 20227 2549
rect 17726 2544 20227 2546
rect 17726 2488 20166 2544
rect 20222 2488 20227 2544
rect 17726 2486 20227 2488
rect 2773 2483 2839 2486
rect 17585 2483 17651 2486
rect 20161 2483 20227 2486
rect 0 2410 800 2440
rect 1301 2410 1367 2413
rect 0 2408 1367 2410
rect 0 2352 1306 2408
rect 1362 2352 1367 2408
rect 0 2350 1367 2352
rect 0 2320 800 2350
rect 1301 2347 1367 2350
rect 5809 2410 5875 2413
rect 43805 2410 43871 2413
rect 5809 2408 43871 2410
rect 5809 2352 5814 2408
rect 5870 2352 43810 2408
rect 43866 2352 43871 2408
rect 5809 2350 43871 2352
rect 5809 2347 5875 2350
rect 43805 2347 43871 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 2002 800 2032
rect 3509 2002 3575 2005
rect 0 2000 3575 2002
rect 0 1944 3514 2000
rect 3570 1944 3575 2000
rect 0 1942 3575 1944
rect 0 1912 800 1942
rect 3509 1939 3575 1942
rect 14038 1940 14044 2004
rect 14108 2002 14114 2004
rect 33777 2002 33843 2005
rect 14108 2000 33843 2002
rect 14108 1944 33782 2000
rect 33838 1944 33843 2000
rect 14108 1942 33843 1944
rect 14108 1940 14114 1942
rect 33777 1939 33843 1942
rect 933 1866 999 1869
rect 10961 1866 11027 1869
rect 933 1864 11027 1866
rect 933 1808 938 1864
rect 994 1808 10966 1864
rect 11022 1808 11027 1864
rect 933 1806 11027 1808
rect 933 1803 999 1806
rect 10961 1803 11027 1806
rect 13721 1866 13787 1869
rect 28441 1866 28507 1869
rect 13721 1864 28507 1866
rect 13721 1808 13726 1864
rect 13782 1808 28446 1864
rect 28502 1808 28507 1864
rect 13721 1806 28507 1808
rect 13721 1803 13787 1806
rect 28441 1803 28507 1806
rect 0 1594 800 1624
rect 3417 1594 3483 1597
rect 0 1592 3483 1594
rect 0 1536 3422 1592
rect 3478 1536 3483 1592
rect 0 1534 3483 1536
rect 0 1504 800 1534
rect 3417 1531 3483 1534
rect 1853 1458 1919 1461
rect 14181 1458 14247 1461
rect 1853 1456 14247 1458
rect 1853 1400 1858 1456
rect 1914 1400 14186 1456
rect 14242 1400 14247 1456
rect 1853 1398 14247 1400
rect 1853 1395 1919 1398
rect 14181 1395 14247 1398
rect 6085 1322 6151 1325
rect 22093 1322 22159 1325
rect 6085 1320 22159 1322
rect 6085 1264 6090 1320
rect 6146 1264 22098 1320
rect 22154 1264 22159 1320
rect 6085 1262 22159 1264
rect 6085 1259 6151 1262
rect 22093 1259 22159 1262
rect 2630 1124 2636 1188
rect 2700 1186 2706 1188
rect 13905 1186 13971 1189
rect 2700 1184 13971 1186
rect 2700 1128 13910 1184
rect 13966 1128 13971 1184
rect 2700 1126 13971 1128
rect 2700 1124 2706 1126
rect 13905 1123 13971 1126
rect 15193 1186 15259 1189
rect 22318 1186 22324 1188
rect 15193 1184 22324 1186
rect 15193 1128 15198 1184
rect 15254 1128 22324 1184
rect 15193 1126 22324 1128
rect 15193 1123 15259 1126
rect 22318 1124 22324 1126
rect 22388 1124 22394 1188
rect 5758 988 5764 1052
rect 5828 1050 5834 1052
rect 26601 1050 26667 1053
rect 5828 1048 26667 1050
rect 5828 992 26606 1048
rect 26662 992 26667 1048
rect 5828 990 26667 992
rect 5828 988 5834 990
rect 26601 987 26667 990
rect 3877 914 3943 917
rect 9121 914 9187 917
rect 27245 914 27311 917
rect 3877 912 3986 914
rect 3877 856 3882 912
rect 3938 856 3986 912
rect 3877 851 3986 856
rect 9121 912 27311 914
rect 9121 856 9126 912
rect 9182 856 27250 912
rect 27306 856 27311 912
rect 9121 854 27311 856
rect 9121 851 9187 854
rect 27245 851 27311 854
rect 3926 642 3986 851
rect 5441 778 5507 781
rect 26550 778 26556 780
rect 5441 776 26556 778
rect 5441 720 5446 776
rect 5502 720 26556 776
rect 5441 718 26556 720
rect 5441 715 5507 718
rect 26550 716 26556 718
rect 26620 716 26626 780
rect 29085 642 29151 645
rect 3926 640 29151 642
rect 3926 584 29090 640
rect 29146 584 29151 640
rect 3926 582 29151 584
rect 29085 579 29151 582
<< via3 >>
rect 15516 25740 15580 25804
rect 21404 25468 21468 25532
rect 27660 25196 27724 25260
rect 27476 25060 27540 25124
rect 23612 24788 23676 24852
rect 20300 24516 20364 24580
rect 25452 24516 25516 24580
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 14044 24244 14108 24308
rect 12756 24108 12820 24172
rect 20484 23972 20548 24036
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 16804 23836 16868 23900
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 13676 23564 13740 23628
rect 8892 23428 8956 23492
rect 12388 23428 12452 23492
rect 14964 23488 15028 23492
rect 14964 23432 14978 23488
rect 14978 23432 15028 23488
rect 14964 23428 15028 23432
rect 15516 23488 15580 23492
rect 15516 23432 15530 23488
rect 15530 23432 15580 23488
rect 15516 23428 15580 23432
rect 24716 23428 24780 23492
rect 27292 23488 27356 23492
rect 27292 23432 27342 23488
rect 27342 23432 27356 23488
rect 27292 23428 27356 23432
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 15516 23292 15580 23356
rect 18828 23292 18892 23356
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 17540 22612 17604 22676
rect 19380 22748 19444 22812
rect 20300 22340 20364 22404
rect 21588 22340 21652 22404
rect 22692 22340 22756 22404
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 26004 22340 26068 22404
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 16620 22068 16684 22132
rect 19748 22068 19812 22132
rect 28764 22204 28828 22268
rect 20484 21932 20548 21996
rect 19380 21856 19444 21860
rect 19380 21800 19394 21856
rect 19394 21800 19444 21856
rect 19380 21796 19444 21800
rect 29500 21796 29564 21860
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 8708 21660 8772 21724
rect 17540 21660 17604 21724
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 3556 21524 3620 21588
rect 14964 21524 15028 21588
rect 12204 21448 12268 21452
rect 12204 21392 12254 21448
rect 12254 21392 12268 21448
rect 12204 21388 12268 21392
rect 17172 21448 17236 21452
rect 17172 21392 17186 21448
rect 17186 21392 17236 21448
rect 17172 21388 17236 21392
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 980 20980 1044 21044
rect 14964 21116 15028 21180
rect 17724 21116 17788 21180
rect 19012 21116 19076 21180
rect 19196 21176 19260 21180
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 19196 21120 19210 21176
rect 19210 21120 19260 21176
rect 19196 21116 19260 21120
rect 13860 20980 13924 21044
rect 26188 20980 26252 21044
rect 1716 20904 1780 20908
rect 1716 20848 1730 20904
rect 1730 20848 1780 20904
rect 1716 20844 1780 20848
rect 5396 20844 5460 20908
rect 11836 20844 11900 20908
rect 19380 20844 19444 20908
rect 6132 20708 6196 20772
rect 6868 20708 6932 20772
rect 10916 20708 10980 20772
rect 18460 20768 18524 20772
rect 18460 20712 18474 20768
rect 18474 20712 18524 20768
rect 18460 20708 18524 20712
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 2268 20572 2332 20636
rect 17540 20572 17604 20636
rect 16620 20436 16684 20500
rect 19564 20572 19628 20636
rect 19748 20572 19812 20636
rect 24532 20708 24596 20772
rect 25820 20708 25884 20772
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 21956 20436 22020 20500
rect 22324 20436 22388 20500
rect 24164 20300 24228 20364
rect 30420 20300 30484 20364
rect 27476 20164 27540 20228
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 17356 20028 17420 20092
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 14780 19620 14844 19684
rect 19748 19620 19812 19684
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 9812 19348 9876 19412
rect 16988 19544 17052 19548
rect 16988 19488 17002 19544
rect 17002 19488 17052 19544
rect 16988 19484 17052 19488
rect 21772 19484 21836 19548
rect 22508 19484 22572 19548
rect 25636 19484 25700 19548
rect 28580 19544 28644 19548
rect 28580 19488 28630 19544
rect 28630 19488 28644 19544
rect 28580 19484 28644 19488
rect 6316 19212 6380 19276
rect 17356 19076 17420 19140
rect 18828 19076 18892 19140
rect 26556 19136 26620 19140
rect 26556 19080 26570 19136
rect 26570 19080 26620 19136
rect 26556 19076 26620 19080
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 4292 18940 4356 19004
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 29132 18940 29196 19004
rect 31524 19000 31588 19004
rect 31524 18944 31538 19000
rect 31538 18944 31588 19000
rect 31524 18940 31588 18944
rect 6132 18804 6196 18868
rect 9996 18668 10060 18732
rect 1164 18532 1228 18596
rect 9076 18532 9140 18596
rect 14228 18804 14292 18868
rect 28948 18668 29012 18732
rect 18460 18532 18524 18596
rect 20300 18532 20364 18596
rect 21036 18532 21100 18596
rect 29316 18532 29380 18596
rect 29684 18532 29748 18596
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 13860 18396 13924 18460
rect 15332 18184 15396 18188
rect 16804 18456 16868 18460
rect 16804 18400 16854 18456
rect 16854 18400 16868 18456
rect 16804 18396 16868 18400
rect 17540 18396 17604 18460
rect 18828 18396 18892 18460
rect 18828 18260 18892 18324
rect 15332 18128 15382 18184
rect 15382 18128 15396 18184
rect 15332 18124 15396 18128
rect 26188 18124 26252 18188
rect 12020 17988 12084 18052
rect 26188 17988 26252 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 5028 17580 5092 17644
rect 20116 17852 20180 17916
rect 27660 17988 27724 18052
rect 28396 17988 28460 18052
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 27660 17852 27724 17916
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 19748 17776 19812 17780
rect 19748 17720 19798 17776
rect 19798 17720 19812 17776
rect 19748 17716 19812 17720
rect 11468 17640 11532 17644
rect 11468 17584 11518 17640
rect 11518 17584 11532 17640
rect 11468 17580 11532 17584
rect 30420 17716 30484 17780
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 4108 17172 4172 17236
rect 8892 17232 8956 17236
rect 8892 17176 8906 17232
rect 8906 17176 8956 17232
rect 6684 17036 6748 17100
rect 8892 17172 8956 17176
rect 9444 17172 9508 17236
rect 12756 17172 12820 17236
rect 14596 17172 14660 17236
rect 16620 17172 16684 17236
rect 22048 17444 22112 17508
rect 28580 17504 28644 17508
rect 28580 17448 28594 17504
rect 28594 17448 28644 17504
rect 28580 17444 28644 17448
rect 29684 17444 29748 17508
rect 32812 17444 32876 17508
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 20852 17308 20916 17372
rect 21404 17308 21468 17372
rect 23428 17308 23492 17372
rect 15148 16900 15212 16964
rect 17724 16900 17788 16964
rect 19012 16900 19076 16964
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 5948 16764 6012 16828
rect 7052 16764 7116 16828
rect 7788 16688 7852 16692
rect 7788 16632 7838 16688
rect 7838 16632 7852 16688
rect 7788 16628 7852 16632
rect 16436 16628 16500 16692
rect 25268 16764 25332 16828
rect 28948 16764 29012 16828
rect 29316 16764 29380 16828
rect 5028 16492 5092 16556
rect 10180 16492 10244 16556
rect 11652 16492 11716 16556
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 1900 16220 1964 16284
rect 5212 16084 5276 16148
rect 7604 16084 7668 16148
rect 21956 16492 22020 16556
rect 19196 16356 19260 16420
rect 19380 16416 19444 16420
rect 19380 16360 19430 16416
rect 19430 16360 19444 16416
rect 19380 16356 19444 16360
rect 22692 16356 22756 16420
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 11836 16220 11900 16284
rect 16252 16220 16316 16284
rect 23612 16280 23676 16284
rect 23612 16224 23626 16280
rect 23626 16224 23676 16280
rect 23612 16220 23676 16224
rect 25084 16220 25148 16284
rect 25636 16220 25700 16284
rect 980 15948 1044 16012
rect 7236 15812 7300 15876
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 8524 15540 8588 15604
rect 17172 15812 17236 15876
rect 19748 15812 19812 15876
rect 24164 15812 24228 15876
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 19564 15676 19628 15740
rect 22324 15676 22388 15740
rect 27660 15676 27724 15740
rect 17356 15540 17420 15604
rect 19012 15540 19076 15604
rect 20668 15540 20732 15604
rect 22140 15540 22204 15604
rect 31524 15540 31588 15604
rect 9260 15268 9324 15332
rect 18460 15328 18524 15332
rect 18460 15272 18510 15328
rect 18510 15272 18524 15328
rect 18460 15268 18524 15272
rect 19380 15268 19444 15332
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 3372 15132 3436 15196
rect 12756 15132 12820 15196
rect 17172 15132 17236 15196
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 28396 15132 28460 15196
rect 3740 14996 3804 15060
rect 4108 14996 4172 15060
rect 6500 14996 6564 15060
rect 15700 15056 15764 15060
rect 15700 15000 15750 15056
rect 15750 15000 15764 15056
rect 15700 14996 15764 15000
rect 29132 14996 29196 15060
rect 11836 14784 11900 14788
rect 11836 14728 11850 14784
rect 11850 14728 11900 14784
rect 11836 14724 11900 14728
rect 21588 14724 21652 14788
rect 22692 14724 22756 14788
rect 26004 14724 26068 14788
rect 32812 14724 32876 14788
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 9444 14588 9508 14652
rect 21588 14588 21652 14652
rect 23428 14588 23492 14652
rect 24348 14588 24412 14652
rect 25452 14588 25516 14652
rect 7788 14452 7852 14516
rect 13492 14452 13556 14516
rect 15148 14452 15212 14516
rect 16620 14452 16684 14516
rect 8340 14316 8404 14380
rect 9812 14180 9876 14244
rect 11284 14180 11348 14244
rect 11468 14180 11532 14244
rect 19932 14180 19996 14244
rect 22324 14316 22388 14380
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 6500 14104 6564 14108
rect 6500 14048 6550 14104
rect 6550 14048 6564 14104
rect 6500 14044 6564 14048
rect 9076 14044 9140 14108
rect 18828 14044 18892 14108
rect 21956 14044 22020 14108
rect 1532 13968 1596 13972
rect 1532 13912 1582 13968
rect 1582 13912 1596 13968
rect 1532 13908 1596 13912
rect 7420 13908 7484 13972
rect 7788 13908 7852 13972
rect 14780 13908 14844 13972
rect 20852 13968 20916 13972
rect 20852 13912 20902 13968
rect 20902 13912 20916 13968
rect 7604 13636 7668 13700
rect 11284 13636 11348 13700
rect 12572 13636 12636 13700
rect 15884 13636 15948 13700
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 7052 13500 7116 13564
rect 15516 13500 15580 13564
rect 18644 13636 18708 13700
rect 20852 13908 20916 13912
rect 23796 13908 23860 13972
rect 22140 13636 22204 13700
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 1348 13228 1412 13292
rect 11100 13364 11164 13428
rect 9076 13092 9140 13156
rect 12756 13092 12820 13156
rect 20668 13092 20732 13156
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 7052 12956 7116 13020
rect 17724 12956 17788 13020
rect 18460 12956 18524 13020
rect 5580 12820 5644 12884
rect 10548 12684 10612 12748
rect 16436 12820 16500 12884
rect 21404 12820 21468 12884
rect 22692 12956 22756 13020
rect 24900 12956 24964 13020
rect 28948 13092 29012 13156
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 7236 12548 7300 12612
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 3372 12412 3436 12476
rect 9260 12412 9324 12476
rect 12204 12412 12268 12476
rect 3372 12336 3436 12340
rect 3372 12280 3386 12336
rect 3386 12280 3436 12336
rect 3372 12276 3436 12280
rect 10732 12276 10796 12340
rect 13676 12548 13740 12612
rect 14412 12548 14476 12612
rect 19564 12548 19628 12612
rect 22324 12608 22388 12612
rect 22324 12552 22338 12608
rect 22338 12552 22388 12608
rect 22324 12548 22388 12552
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 18460 12412 18524 12476
rect 19196 12412 19260 12476
rect 15148 12276 15212 12340
rect 16804 12276 16868 12340
rect 17724 12276 17788 12340
rect 23796 12276 23860 12340
rect 7604 12140 7668 12204
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 8524 12140 8588 12204
rect 27292 12140 27356 12204
rect 9812 12064 9876 12068
rect 9812 12008 9862 12064
rect 9862 12008 9876 12064
rect 9812 12004 9876 12008
rect 12388 12004 12452 12068
rect 12572 12004 12636 12068
rect 13860 12004 13924 12068
rect 19932 12004 19996 12068
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 13492 11868 13556 11932
rect 11652 11732 11716 11796
rect 12204 11732 12268 11796
rect 14780 11868 14844 11932
rect 14412 11792 14476 11796
rect 14412 11736 14426 11792
rect 14426 11736 14476 11792
rect 14412 11732 14476 11736
rect 8892 11460 8956 11524
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 8524 11384 8588 11388
rect 8524 11328 8574 11384
rect 8574 11328 8588 11384
rect 8524 11324 8588 11328
rect 19932 11460 19996 11524
rect 25084 11596 25148 11660
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 3372 11188 3436 11252
rect 17172 11324 17236 11388
rect 9628 11188 9692 11252
rect 14780 11188 14844 11252
rect 1716 11112 1780 11116
rect 1716 11056 1766 11112
rect 1766 11056 1780 11112
rect 1716 11052 1780 11056
rect 6500 11052 6564 11116
rect 12204 11052 12268 11116
rect 12388 11052 12452 11116
rect 13676 11052 13740 11116
rect 14780 11052 14844 11116
rect 7052 10976 7116 10980
rect 7052 10920 7102 10976
rect 7102 10920 7116 10976
rect 7052 10916 7116 10920
rect 9812 10976 9876 10980
rect 9812 10920 9862 10976
rect 9862 10920 9876 10976
rect 9812 10916 9876 10920
rect 11100 10916 11164 10980
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 5580 10780 5644 10844
rect 14044 10916 14108 10980
rect 18460 10916 18524 10980
rect 21588 10916 21652 10980
rect 21956 10916 22020 10980
rect 22140 10916 22204 10980
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 12204 10780 12268 10844
rect 10548 10644 10612 10708
rect 14964 10780 15028 10844
rect 27476 10840 27540 10844
rect 27476 10784 27490 10840
rect 27490 10784 27540 10840
rect 27476 10780 27540 10784
rect 21404 10644 21468 10708
rect 13492 10372 13556 10436
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 11468 10236 11532 10300
rect 12388 10236 12452 10300
rect 11100 10100 11164 10164
rect 14044 10236 14108 10300
rect 14780 10372 14844 10436
rect 20300 10372 20364 10436
rect 24900 10372 24964 10436
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 5948 9964 6012 10028
rect 5764 9828 5828 9892
rect 7236 9828 7300 9892
rect 8340 9964 8404 10028
rect 14596 10024 14660 10028
rect 14596 9968 14610 10024
rect 14610 9968 14660 10024
rect 14596 9964 14660 9968
rect 15516 9964 15580 10028
rect 17356 9964 17420 10028
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 1532 9556 1596 9620
rect 3740 9616 3804 9620
rect 3740 9560 3790 9616
rect 3790 9560 3804 9616
rect 3740 9556 3804 9560
rect 4292 9616 4356 9620
rect 4292 9560 4306 9616
rect 4306 9560 4356 9616
rect 4292 9556 4356 9560
rect 7604 9556 7668 9620
rect 12020 9828 12084 9892
rect 13492 9828 13556 9892
rect 15700 9828 15764 9892
rect 18644 9828 18708 9892
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 13676 9692 13740 9756
rect 21404 9692 21468 9756
rect 21956 9828 22020 9892
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 12388 9556 12452 9620
rect 2084 9420 2148 9484
rect 4108 9420 4172 9484
rect 19380 9420 19444 9484
rect 21036 9420 21100 9484
rect 11468 9284 11532 9348
rect 14228 9344 14292 9348
rect 14228 9288 14242 9344
rect 14242 9288 14292 9344
rect 14228 9284 14292 9288
rect 16804 9284 16868 9348
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 11652 9148 11716 9212
rect 7788 9012 7852 9076
rect 3740 8876 3804 8940
rect 15884 9012 15948 9076
rect 12204 8876 12268 8940
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 9996 8664 10060 8668
rect 9996 8608 10046 8664
rect 10046 8608 10060 8664
rect 9996 8604 10060 8608
rect 11100 8604 11164 8668
rect 2636 8468 2700 8532
rect 1348 8196 1412 8260
rect 5028 8256 5092 8260
rect 10180 8332 10244 8396
rect 20116 8740 20180 8804
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 16436 8664 16500 8668
rect 16436 8608 16450 8664
rect 16450 8608 16500 8664
rect 16436 8604 16500 8608
rect 25268 8604 25332 8668
rect 19564 8332 19628 8396
rect 5028 8200 5042 8256
rect 5042 8200 5092 8256
rect 5028 8196 5092 8200
rect 10916 8196 10980 8260
rect 15516 8196 15580 8260
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 2268 8120 2332 8124
rect 2268 8064 2318 8120
rect 2318 8064 2332 8120
rect 2268 8060 2332 8064
rect 18828 8060 18892 8124
rect 3740 7924 3804 7988
rect 13492 7924 13556 7988
rect 11284 7652 11348 7716
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 12756 7516 12820 7580
rect 15148 7516 15212 7580
rect 21404 7576 21468 7580
rect 21404 7520 21454 7576
rect 21454 7520 21468 7576
rect 21404 7516 21468 7520
rect 7052 7108 7116 7172
rect 12204 7168 12268 7172
rect 12204 7112 12218 7168
rect 12218 7112 12268 7168
rect 12204 7108 12268 7112
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 4108 6972 4172 7036
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 1716 6760 1780 6764
rect 1716 6704 1766 6760
rect 1766 6704 1780 6760
rect 1716 6700 1780 6704
rect 9076 6760 9140 6764
rect 9076 6704 9090 6760
rect 9090 6704 9140 6760
rect 9076 6700 9140 6704
rect 11836 6700 11900 6764
rect 15332 6700 15396 6764
rect 1900 6564 1964 6628
rect 7420 6564 7484 6628
rect 19748 6760 19812 6764
rect 19748 6704 19762 6760
rect 19762 6704 19812 6760
rect 19748 6700 19812 6704
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 5212 6428 5276 6492
rect 9628 6428 9692 6492
rect 1164 6156 1228 6220
rect 6316 6292 6380 6356
rect 29500 6292 29564 6356
rect 10180 6156 10244 6220
rect 6868 6020 6932 6084
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 612 5850 676 5914
rect 6132 5884 6196 5948
rect 7604 5884 7668 5948
rect 11652 5944 11716 5948
rect 11652 5888 11666 5944
rect 11666 5888 11716 5944
rect 11652 5884 11716 5888
rect 13860 5748 13924 5812
rect 14964 5748 15028 5812
rect 16436 5748 16500 5812
rect 22508 5612 22572 5676
rect 16620 5476 16684 5540
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 980 5340 1044 5404
rect 5396 5340 5460 5404
rect 9996 5340 10060 5404
rect 12572 5068 12636 5132
rect 10732 4932 10796 4996
rect 12388 4932 12452 4996
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 3556 4660 3620 4724
rect 11468 4524 11532 4588
rect 19012 4660 19076 4724
rect 21772 4660 21836 4724
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 16988 4252 17052 4316
rect 24348 4116 24412 4180
rect 6684 3980 6748 4044
rect 9260 4040 9324 4044
rect 9260 3984 9310 4040
rect 9310 3984 9324 4040
rect 9260 3980 9324 3984
rect 7236 3844 7300 3908
rect 14228 3980 14292 4044
rect 24532 3980 24596 4044
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 26188 3572 26252 3636
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 8708 3164 8772 3228
rect 24716 3028 24780 3092
rect 13676 2756 13740 2820
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 8892 2620 8956 2684
rect 19932 2620 19996 2684
rect 25820 2620 25884 2684
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
rect 14044 1940 14108 2004
rect 2636 1124 2700 1188
rect 22324 1124 22388 1188
rect 5764 988 5828 1052
rect 26556 716 26620 780
<< metal4 >>
rect 15515 25804 15581 25805
rect 15515 25740 15516 25804
rect 15580 25740 15581 25804
rect 15515 25739 15581 25740
rect 2944 24512 3264 24528
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 7944 23968 8264 24528
rect 12944 24512 13264 24528
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12755 24172 12821 24173
rect 12755 24108 12756 24172
rect 12820 24108 12821 24172
rect 12755 24107 12821 24108
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 8891 23492 8957 23493
rect 8891 23428 8892 23492
rect 8956 23428 8957 23492
rect 8891 23427 8957 23428
rect 12387 23492 12453 23493
rect 12387 23428 12388 23492
rect 12452 23490 12453 23492
rect 12452 23430 12634 23490
rect 12452 23428 12453 23430
rect 12387 23427 12453 23428
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 3555 21588 3621 21589
rect 3555 21524 3556 21588
rect 3620 21524 3621 21588
rect 3555 21523 3621 21524
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 979 21044 1045 21045
rect 979 20980 980 21044
rect 1044 20980 1045 21044
rect 979 20979 1045 20980
rect 982 16590 1042 20979
rect 1715 20908 1781 20909
rect 1715 20844 1716 20908
rect 1780 20844 1781 20908
rect 1715 20843 1781 20844
rect 1163 18596 1229 18597
rect 1163 18532 1164 18596
rect 1228 18532 1229 18596
rect 1163 18531 1229 18532
rect 614 16530 1042 16590
rect 614 5915 674 16530
rect 979 16012 1045 16013
rect 979 15948 980 16012
rect 1044 15948 1045 16012
rect 979 15947 1045 15948
rect 611 5914 677 5915
rect 611 5850 612 5914
rect 676 5850 677 5914
rect 611 5849 677 5850
rect 982 5405 1042 15947
rect 1166 6221 1226 18531
rect 1531 13972 1597 13973
rect 1531 13908 1532 13972
rect 1596 13908 1597 13972
rect 1531 13907 1597 13908
rect 1347 13292 1413 13293
rect 1347 13228 1348 13292
rect 1412 13228 1413 13292
rect 1347 13227 1413 13228
rect 1350 8261 1410 13227
rect 1534 9621 1594 13907
rect 1718 11250 1778 20843
rect 2267 20636 2333 20637
rect 2267 20572 2268 20636
rect 2332 20572 2333 20636
rect 2267 20571 2333 20572
rect 1899 16284 1965 16285
rect 1899 16220 1900 16284
rect 1964 16220 1965 16284
rect 1899 16219 1965 16220
rect 1902 12450 1962 16219
rect 1902 12390 2146 12450
rect 1718 11190 1962 11250
rect 1715 11116 1781 11117
rect 1715 11052 1716 11116
rect 1780 11052 1781 11116
rect 1715 11051 1781 11052
rect 1531 9620 1597 9621
rect 1531 9556 1532 9620
rect 1596 9556 1597 9620
rect 1531 9555 1597 9556
rect 1347 8260 1413 8261
rect 1347 8196 1348 8260
rect 1412 8196 1413 8260
rect 1347 8195 1413 8196
rect 1718 6765 1778 11051
rect 1715 6764 1781 6765
rect 1715 6700 1716 6764
rect 1780 6700 1781 6764
rect 1715 6699 1781 6700
rect 1902 6629 1962 11190
rect 2086 9485 2146 12390
rect 2083 9484 2149 9485
rect 2083 9420 2084 9484
rect 2148 9420 2149 9484
rect 2083 9419 2149 9420
rect 2270 8125 2330 20571
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 3371 15196 3437 15197
rect 3371 15132 3372 15196
rect 3436 15132 3437 15196
rect 3371 15131 3437 15132
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 3374 12477 3434 15131
rect 3371 12476 3437 12477
rect 3371 12412 3372 12476
rect 3436 12412 3437 12476
rect 3371 12411 3437 12412
rect 3371 12340 3437 12341
rect 3371 12276 3372 12340
rect 3436 12276 3437 12340
rect 3371 12275 3437 12276
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 3374 11253 3434 12275
rect 3371 11252 3437 11253
rect 3371 11188 3372 11252
rect 3436 11188 3437 11252
rect 3371 11187 3437 11188
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2635 8532 2701 8533
rect 2635 8468 2636 8532
rect 2700 8468 2701 8532
rect 2635 8467 2701 8468
rect 2267 8124 2333 8125
rect 2267 8060 2268 8124
rect 2332 8060 2333 8124
rect 2267 8059 2333 8060
rect 1899 6628 1965 6629
rect 1899 6564 1900 6628
rect 1964 6564 1965 6628
rect 1899 6563 1965 6564
rect 1163 6220 1229 6221
rect 1163 6156 1164 6220
rect 1228 6156 1229 6220
rect 1163 6155 1229 6156
rect 979 5404 1045 5405
rect 979 5340 980 5404
rect 1044 5340 1045 5404
rect 979 5339 1045 5340
rect 2638 1189 2698 8467
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 3558 4725 3618 21523
rect 5395 20908 5461 20909
rect 5395 20844 5396 20908
rect 5460 20844 5461 20908
rect 5395 20843 5461 20844
rect 4291 19004 4357 19005
rect 4291 18940 4292 19004
rect 4356 18940 4357 19004
rect 4291 18939 4357 18940
rect 4107 17236 4173 17237
rect 4107 17172 4108 17236
rect 4172 17172 4173 17236
rect 4107 17171 4173 17172
rect 4110 15061 4170 17171
rect 3739 15060 3805 15061
rect 3739 14996 3740 15060
rect 3804 14996 3805 15060
rect 3739 14995 3805 14996
rect 4107 15060 4173 15061
rect 4107 14996 4108 15060
rect 4172 14996 4173 15060
rect 4107 14995 4173 14996
rect 3742 9621 3802 14995
rect 4294 9621 4354 18939
rect 5027 17644 5093 17645
rect 5027 17580 5028 17644
rect 5092 17580 5093 17644
rect 5027 17579 5093 17580
rect 5030 16557 5090 17579
rect 5027 16556 5093 16557
rect 5027 16492 5028 16556
rect 5092 16492 5093 16556
rect 5027 16491 5093 16492
rect 3739 9620 3805 9621
rect 3739 9556 3740 9620
rect 3804 9556 3805 9620
rect 3739 9555 3805 9556
rect 4291 9620 4357 9621
rect 4291 9556 4292 9620
rect 4356 9556 4357 9620
rect 4291 9555 4357 9556
rect 4107 9484 4173 9485
rect 4107 9420 4108 9484
rect 4172 9420 4173 9484
rect 4107 9419 4173 9420
rect 3739 8940 3805 8941
rect 3739 8876 3740 8940
rect 3804 8876 3805 8940
rect 3739 8875 3805 8876
rect 3742 7989 3802 8875
rect 3739 7988 3805 7989
rect 3739 7924 3740 7988
rect 3804 7924 3805 7988
rect 3739 7923 3805 7924
rect 4110 7037 4170 9419
rect 5030 8261 5090 16491
rect 5211 16148 5277 16149
rect 5211 16084 5212 16148
rect 5276 16084 5277 16148
rect 5211 16083 5277 16084
rect 5027 8260 5093 8261
rect 5027 8196 5028 8260
rect 5092 8196 5093 8260
rect 5027 8195 5093 8196
rect 4107 7036 4173 7037
rect 4107 6972 4108 7036
rect 4172 6972 4173 7036
rect 4107 6971 4173 6972
rect 5214 6493 5274 16083
rect 5211 6492 5277 6493
rect 5211 6428 5212 6492
rect 5276 6428 5277 6492
rect 5211 6427 5277 6428
rect 5398 5405 5458 20843
rect 6131 20772 6197 20773
rect 6131 20708 6132 20772
rect 6196 20708 6197 20772
rect 6131 20707 6197 20708
rect 6867 20772 6933 20773
rect 6867 20708 6868 20772
rect 6932 20708 6933 20772
rect 6867 20707 6933 20708
rect 6134 18869 6194 20707
rect 6315 19276 6381 19277
rect 6315 19212 6316 19276
rect 6380 19212 6381 19276
rect 6315 19211 6381 19212
rect 6131 18868 6197 18869
rect 6131 18804 6132 18868
rect 6196 18804 6197 18868
rect 6131 18803 6197 18804
rect 5947 16828 6013 16829
rect 5947 16764 5948 16828
rect 6012 16764 6013 16828
rect 5947 16763 6013 16764
rect 5579 12884 5645 12885
rect 5579 12820 5580 12884
rect 5644 12820 5645 12884
rect 5579 12819 5645 12820
rect 5582 10845 5642 12819
rect 5579 10844 5645 10845
rect 5579 10780 5580 10844
rect 5644 10780 5645 10844
rect 5579 10779 5645 10780
rect 5950 10029 6010 16763
rect 5947 10028 6013 10029
rect 5947 9964 5948 10028
rect 6012 9964 6013 10028
rect 5947 9963 6013 9964
rect 5763 9892 5829 9893
rect 5763 9828 5764 9892
rect 5828 9828 5829 9892
rect 5763 9827 5829 9828
rect 5395 5404 5461 5405
rect 5395 5340 5396 5404
rect 5460 5340 5461 5404
rect 5395 5339 5461 5340
rect 3555 4724 3621 4725
rect 3555 4660 3556 4724
rect 3620 4660 3621 4724
rect 3555 4659 3621 4660
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 2635 1188 2701 1189
rect 2635 1124 2636 1188
rect 2700 1124 2701 1188
rect 2635 1123 2701 1124
rect 5766 1053 5826 9827
rect 6134 5949 6194 18803
rect 6318 6357 6378 19211
rect 6683 17100 6749 17101
rect 6683 17036 6684 17100
rect 6748 17036 6749 17100
rect 6683 17035 6749 17036
rect 6499 15060 6565 15061
rect 6499 14996 6500 15060
rect 6564 14996 6565 15060
rect 6499 14995 6565 14996
rect 6502 14109 6562 14995
rect 6499 14108 6565 14109
rect 6499 14044 6500 14108
rect 6564 14044 6565 14108
rect 6499 14043 6565 14044
rect 6502 11117 6562 14043
rect 6499 11116 6565 11117
rect 6499 11052 6500 11116
rect 6564 11052 6565 11116
rect 6499 11051 6565 11052
rect 6315 6356 6381 6357
rect 6315 6292 6316 6356
rect 6380 6292 6381 6356
rect 6315 6291 6381 6292
rect 6131 5948 6197 5949
rect 6131 5884 6132 5948
rect 6196 5884 6197 5948
rect 6131 5883 6197 5884
rect 6686 4045 6746 17035
rect 6870 6085 6930 20707
rect 7944 20704 8264 21728
rect 8707 21724 8773 21725
rect 8707 21660 8708 21724
rect 8772 21660 8773 21724
rect 8707 21659 8773 21660
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7051 16828 7117 16829
rect 7051 16764 7052 16828
rect 7116 16764 7117 16828
rect 7051 16763 7117 16764
rect 7054 13565 7114 16763
rect 7787 16692 7853 16693
rect 7787 16628 7788 16692
rect 7852 16628 7853 16692
rect 7787 16627 7853 16628
rect 7603 16148 7669 16149
rect 7603 16084 7604 16148
rect 7668 16084 7669 16148
rect 7603 16083 7669 16084
rect 7235 15876 7301 15877
rect 7235 15812 7236 15876
rect 7300 15812 7301 15876
rect 7235 15811 7301 15812
rect 7051 13564 7117 13565
rect 7051 13500 7052 13564
rect 7116 13500 7117 13564
rect 7051 13499 7117 13500
rect 7051 13020 7117 13021
rect 7051 12956 7052 13020
rect 7116 12956 7117 13020
rect 7051 12955 7117 12956
rect 7054 10981 7114 12955
rect 7238 12613 7298 15811
rect 7419 13972 7485 13973
rect 7419 13908 7420 13972
rect 7484 13908 7485 13972
rect 7419 13907 7485 13908
rect 7235 12612 7301 12613
rect 7235 12548 7236 12612
rect 7300 12548 7301 12612
rect 7235 12547 7301 12548
rect 7051 10980 7117 10981
rect 7051 10916 7052 10980
rect 7116 10916 7117 10980
rect 7051 10915 7117 10916
rect 7054 7173 7114 10915
rect 7235 9892 7301 9893
rect 7235 9828 7236 9892
rect 7300 9828 7301 9892
rect 7235 9827 7301 9828
rect 7051 7172 7117 7173
rect 7051 7108 7052 7172
rect 7116 7108 7117 7172
rect 7051 7107 7117 7108
rect 6867 6084 6933 6085
rect 6867 6020 6868 6084
rect 6932 6020 6933 6084
rect 6867 6019 6933 6020
rect 6683 4044 6749 4045
rect 6683 3980 6684 4044
rect 6748 3980 6749 4044
rect 6683 3979 6749 3980
rect 7238 3909 7298 9827
rect 7422 6629 7482 13907
rect 7606 13701 7666 16083
rect 7790 14517 7850 16627
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 8523 15604 8589 15605
rect 8523 15540 8524 15604
rect 8588 15540 8589 15604
rect 8523 15539 8589 15540
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7787 14516 7853 14517
rect 7787 14452 7788 14516
rect 7852 14452 7853 14516
rect 7787 14451 7853 14452
rect 7944 14176 8264 15200
rect 8339 14380 8405 14381
rect 8339 14316 8340 14380
rect 8404 14316 8405 14380
rect 8339 14315 8405 14316
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7787 13972 7853 13973
rect 7787 13908 7788 13972
rect 7852 13908 7853 13972
rect 7787 13907 7853 13908
rect 7603 13700 7669 13701
rect 7603 13636 7604 13700
rect 7668 13636 7669 13700
rect 7603 13635 7669 13636
rect 7606 12205 7666 13635
rect 7603 12204 7669 12205
rect 7603 12140 7604 12204
rect 7668 12140 7669 12204
rect 7603 12139 7669 12140
rect 7603 9620 7669 9621
rect 7603 9556 7604 9620
rect 7668 9556 7669 9620
rect 7603 9555 7669 9556
rect 7419 6628 7485 6629
rect 7419 6564 7420 6628
rect 7484 6564 7485 6628
rect 7419 6563 7485 6564
rect 7606 5949 7666 9555
rect 7790 9077 7850 13907
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 8342 10029 8402 14315
rect 8526 12205 8586 15539
rect 8523 12204 8589 12205
rect 8523 12140 8524 12204
rect 8588 12140 8589 12204
rect 8523 12139 8589 12140
rect 8526 11389 8586 12139
rect 8523 11388 8589 11389
rect 8523 11324 8524 11388
rect 8588 11324 8589 11388
rect 8523 11323 8589 11324
rect 8339 10028 8405 10029
rect 8339 9964 8340 10028
rect 8404 9964 8405 10028
rect 8339 9963 8405 9964
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7787 9076 7853 9077
rect 7787 9012 7788 9076
rect 7852 9012 7853 9076
rect 7787 9011 7853 9012
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7603 5948 7669 5949
rect 7603 5884 7604 5948
rect 7668 5884 7669 5948
rect 7603 5883 7669 5884
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7235 3908 7301 3909
rect 7235 3844 7236 3908
rect 7300 3844 7301 3908
rect 7235 3843 7301 3844
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 8710 3229 8770 21659
rect 8894 17237 8954 23427
rect 12203 21452 12269 21453
rect 12203 21388 12204 21452
rect 12268 21388 12269 21452
rect 12203 21387 12269 21388
rect 11835 20908 11901 20909
rect 11835 20844 11836 20908
rect 11900 20844 11901 20908
rect 11835 20843 11901 20844
rect 10915 20772 10981 20773
rect 10915 20708 10916 20772
rect 10980 20708 10981 20772
rect 10915 20707 10981 20708
rect 9811 19412 9877 19413
rect 9811 19348 9812 19412
rect 9876 19348 9877 19412
rect 9811 19347 9877 19348
rect 9075 18596 9141 18597
rect 9075 18532 9076 18596
rect 9140 18532 9141 18596
rect 9075 18531 9141 18532
rect 8891 17236 8957 17237
rect 8891 17172 8892 17236
rect 8956 17172 8957 17236
rect 8891 17171 8957 17172
rect 9078 14109 9138 18531
rect 9443 17236 9509 17237
rect 9443 17172 9444 17236
rect 9508 17172 9509 17236
rect 9443 17171 9509 17172
rect 9259 15332 9325 15333
rect 9259 15268 9260 15332
rect 9324 15268 9325 15332
rect 9259 15267 9325 15268
rect 9075 14108 9141 14109
rect 9075 14044 9076 14108
rect 9140 14044 9141 14108
rect 9075 14043 9141 14044
rect 9078 13157 9138 14043
rect 9075 13156 9141 13157
rect 9075 13092 9076 13156
rect 9140 13092 9141 13156
rect 9075 13091 9141 13092
rect 9262 13018 9322 15267
rect 9446 14653 9506 17171
rect 9443 14652 9509 14653
rect 9443 14588 9444 14652
rect 9508 14588 9509 14652
rect 9443 14587 9509 14588
rect 9814 14245 9874 19347
rect 9995 18732 10061 18733
rect 9995 18668 9996 18732
rect 10060 18668 10061 18732
rect 9995 18667 10061 18668
rect 9998 18594 10058 18667
rect 9998 18534 10426 18594
rect 10179 16556 10245 16557
rect 10179 16492 10180 16556
rect 10244 16492 10245 16556
rect 10179 16491 10245 16492
rect 9811 14244 9877 14245
rect 9811 14180 9812 14244
rect 9876 14180 9877 14244
rect 9811 14179 9877 14180
rect 9078 12958 9322 13018
rect 8891 11524 8957 11525
rect 8891 11460 8892 11524
rect 8956 11460 8957 11524
rect 8891 11459 8957 11460
rect 8707 3228 8773 3229
rect 8707 3164 8708 3228
rect 8772 3164 8773 3228
rect 8707 3163 8773 3164
rect 8894 2685 8954 11459
rect 9078 6765 9138 12958
rect 9259 12476 9325 12477
rect 9259 12412 9260 12476
rect 9324 12412 9325 12476
rect 10182 12474 10242 16491
rect 9259 12411 9325 12412
rect 9998 12414 10242 12474
rect 9075 6764 9141 6765
rect 9075 6700 9076 6764
rect 9140 6700 9141 6764
rect 9075 6699 9141 6700
rect 9262 4045 9322 12411
rect 9811 12068 9877 12069
rect 9811 12004 9812 12068
rect 9876 12004 9877 12068
rect 9811 12003 9877 12004
rect 9627 11252 9693 11253
rect 9627 11188 9628 11252
rect 9692 11188 9693 11252
rect 9627 11187 9693 11188
rect 9630 6493 9690 11187
rect 9814 10981 9874 12003
rect 9811 10980 9877 10981
rect 9811 10916 9812 10980
rect 9876 10916 9877 10980
rect 9811 10915 9877 10916
rect 9998 8669 10058 12414
rect 10366 12338 10426 18534
rect 10547 12748 10613 12749
rect 10547 12684 10548 12748
rect 10612 12684 10613 12748
rect 10547 12683 10613 12684
rect 10182 12278 10426 12338
rect 9995 8668 10061 8669
rect 9995 8604 9996 8668
rect 10060 8604 10061 8668
rect 9995 8603 10061 8604
rect 9627 6492 9693 6493
rect 9627 6428 9628 6492
rect 9692 6428 9693 6492
rect 9627 6427 9693 6428
rect 9998 5405 10058 8603
rect 10182 8397 10242 12278
rect 10550 10709 10610 12683
rect 10731 12340 10797 12341
rect 10731 12276 10732 12340
rect 10796 12276 10797 12340
rect 10731 12275 10797 12276
rect 10547 10708 10613 10709
rect 10547 10644 10548 10708
rect 10612 10644 10613 10708
rect 10547 10643 10613 10644
rect 10179 8396 10245 8397
rect 10179 8332 10180 8396
rect 10244 8332 10245 8396
rect 10179 8331 10245 8332
rect 10182 6221 10242 8331
rect 10179 6220 10245 6221
rect 10179 6156 10180 6220
rect 10244 6156 10245 6220
rect 10179 6155 10245 6156
rect 9995 5404 10061 5405
rect 9995 5340 9996 5404
rect 10060 5340 10061 5404
rect 9995 5339 10061 5340
rect 10734 4997 10794 12275
rect 10918 8261 10978 20707
rect 11467 17644 11533 17645
rect 11467 17580 11468 17644
rect 11532 17580 11533 17644
rect 11467 17579 11533 17580
rect 11470 14245 11530 17579
rect 11651 16556 11717 16557
rect 11651 16492 11652 16556
rect 11716 16492 11717 16556
rect 11651 16491 11717 16492
rect 11283 14244 11349 14245
rect 11283 14180 11284 14244
rect 11348 14180 11349 14244
rect 11283 14179 11349 14180
rect 11467 14244 11533 14245
rect 11467 14180 11468 14244
rect 11532 14180 11533 14244
rect 11467 14179 11533 14180
rect 11286 13970 11346 14179
rect 11286 13910 11530 13970
rect 11283 13700 11349 13701
rect 11283 13636 11284 13700
rect 11348 13636 11349 13700
rect 11283 13635 11349 13636
rect 11099 13428 11165 13429
rect 11099 13364 11100 13428
rect 11164 13364 11165 13428
rect 11099 13363 11165 13364
rect 11102 10981 11162 13363
rect 11099 10980 11165 10981
rect 11099 10916 11100 10980
rect 11164 10916 11165 10980
rect 11099 10915 11165 10916
rect 11099 10164 11165 10165
rect 11099 10100 11100 10164
rect 11164 10100 11165 10164
rect 11099 10099 11165 10100
rect 11102 8669 11162 10099
rect 11099 8668 11165 8669
rect 11099 8604 11100 8668
rect 11164 8604 11165 8668
rect 11099 8603 11165 8604
rect 10915 8260 10981 8261
rect 10915 8196 10916 8260
rect 10980 8196 10981 8260
rect 10915 8195 10981 8196
rect 11286 7717 11346 13635
rect 11470 10301 11530 13910
rect 11654 11797 11714 16491
rect 11838 16285 11898 20843
rect 12019 18052 12085 18053
rect 12019 17988 12020 18052
rect 12084 17988 12085 18052
rect 12019 17987 12085 17988
rect 11835 16284 11901 16285
rect 11835 16220 11836 16284
rect 11900 16220 11901 16284
rect 11835 16219 11901 16220
rect 11835 14788 11901 14789
rect 11835 14724 11836 14788
rect 11900 14724 11901 14788
rect 11835 14723 11901 14724
rect 11651 11796 11717 11797
rect 11651 11732 11652 11796
rect 11716 11732 11717 11796
rect 11651 11731 11717 11732
rect 11467 10300 11533 10301
rect 11467 10236 11468 10300
rect 11532 10236 11533 10300
rect 11467 10235 11533 10236
rect 11467 9348 11533 9349
rect 11467 9284 11468 9348
rect 11532 9284 11533 9348
rect 11467 9283 11533 9284
rect 11283 7716 11349 7717
rect 11283 7652 11284 7716
rect 11348 7652 11349 7716
rect 11283 7651 11349 7652
rect 10731 4996 10797 4997
rect 10731 4932 10732 4996
rect 10796 4932 10797 4996
rect 10731 4931 10797 4932
rect 11470 4589 11530 9283
rect 11651 9212 11717 9213
rect 11651 9148 11652 9212
rect 11716 9148 11717 9212
rect 11651 9147 11717 9148
rect 11654 5949 11714 9147
rect 11838 6765 11898 14723
rect 12022 9893 12082 17987
rect 12206 12477 12266 21387
rect 12574 16418 12634 23430
rect 12758 17237 12818 24107
rect 12944 23424 13264 24448
rect 14043 24308 14109 24309
rect 14043 24244 14044 24308
rect 14108 24244 14109 24308
rect 14043 24243 14109 24244
rect 13675 23628 13741 23629
rect 13675 23564 13676 23628
rect 13740 23564 13741 23628
rect 13675 23563 13741 23564
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12755 17236 12821 17237
rect 12755 17172 12756 17236
rect 12820 17172 12821 17236
rect 12755 17171 12821 17172
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12574 16358 12818 16418
rect 12758 15197 12818 16358
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12755 15196 12821 15197
rect 12755 15132 12756 15196
rect 12820 15132 12821 15196
rect 12755 15131 12821 15132
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12571 13700 12637 13701
rect 12571 13636 12572 13700
rect 12636 13636 12637 13700
rect 12571 13635 12637 13636
rect 12203 12476 12269 12477
rect 12203 12412 12204 12476
rect 12268 12412 12269 12476
rect 12203 12411 12269 12412
rect 12206 11797 12266 12411
rect 12574 12069 12634 13635
rect 12944 13632 13264 14656
rect 13491 14516 13557 14517
rect 13491 14452 13492 14516
rect 13556 14452 13557 14516
rect 13491 14451 13557 14452
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12755 13156 12821 13157
rect 12755 13092 12756 13156
rect 12820 13092 12821 13156
rect 12755 13091 12821 13092
rect 12387 12068 12453 12069
rect 12387 12004 12388 12068
rect 12452 12004 12453 12068
rect 12387 12003 12453 12004
rect 12571 12068 12637 12069
rect 12571 12004 12572 12068
rect 12636 12004 12637 12068
rect 12571 12003 12637 12004
rect 12390 11930 12450 12003
rect 12390 11870 12634 11930
rect 12203 11796 12269 11797
rect 12203 11732 12204 11796
rect 12268 11732 12269 11796
rect 12203 11731 12269 11732
rect 12203 11116 12269 11117
rect 12203 11052 12204 11116
rect 12268 11052 12269 11116
rect 12203 11051 12269 11052
rect 12387 11116 12453 11117
rect 12387 11052 12388 11116
rect 12452 11052 12453 11116
rect 12387 11051 12453 11052
rect 12206 10845 12266 11051
rect 12203 10844 12269 10845
rect 12203 10780 12204 10844
rect 12268 10780 12269 10844
rect 12203 10779 12269 10780
rect 12390 10301 12450 11051
rect 12387 10300 12453 10301
rect 12387 10236 12388 10300
rect 12452 10236 12453 10300
rect 12387 10235 12453 10236
rect 12019 9892 12085 9893
rect 12019 9828 12020 9892
rect 12084 9828 12085 9892
rect 12019 9827 12085 9828
rect 12387 9620 12453 9621
rect 12387 9556 12388 9620
rect 12452 9556 12453 9620
rect 12387 9555 12453 9556
rect 12203 8940 12269 8941
rect 12203 8876 12204 8940
rect 12268 8876 12269 8940
rect 12203 8875 12269 8876
rect 12206 7173 12266 8875
rect 12203 7172 12269 7173
rect 12203 7108 12204 7172
rect 12268 7108 12269 7172
rect 12203 7107 12269 7108
rect 11835 6764 11901 6765
rect 11835 6700 11836 6764
rect 11900 6700 11901 6764
rect 11835 6699 11901 6700
rect 11651 5948 11717 5949
rect 11651 5884 11652 5948
rect 11716 5884 11717 5948
rect 11651 5883 11717 5884
rect 12390 4997 12450 9555
rect 12574 5133 12634 11870
rect 12758 7581 12818 13091
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 13494 12450 13554 14451
rect 13678 12613 13738 23563
rect 13859 21044 13925 21045
rect 13859 20980 13860 21044
rect 13924 20980 13925 21044
rect 13859 20979 13925 20980
rect 13862 18461 13922 20979
rect 13859 18460 13925 18461
rect 13859 18396 13860 18460
rect 13924 18396 13925 18460
rect 13859 18395 13925 18396
rect 13675 12612 13741 12613
rect 13675 12548 13676 12612
rect 13740 12548 13741 12612
rect 13675 12547 13741 12548
rect 13494 12390 13738 12450
rect 13491 11932 13557 11933
rect 13491 11868 13492 11932
rect 13556 11868 13557 11932
rect 13491 11867 13557 11868
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 13494 10437 13554 11867
rect 13678 11117 13738 12390
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13675 11116 13741 11117
rect 13675 11052 13676 11116
rect 13740 11052 13741 11116
rect 13675 11051 13741 11052
rect 13491 10436 13557 10437
rect 13491 10372 13492 10436
rect 13556 10372 13557 10436
rect 13491 10371 13557 10372
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 13491 9892 13557 9893
rect 13491 9828 13492 9892
rect 13556 9828 13557 9892
rect 13491 9827 13557 9828
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12755 7580 12821 7581
rect 12755 7516 12756 7580
rect 12820 7516 12821 7580
rect 12755 7515 12821 7516
rect 12944 7104 13264 8128
rect 13494 7989 13554 9827
rect 13675 9756 13741 9757
rect 13675 9692 13676 9756
rect 13740 9692 13741 9756
rect 13675 9691 13741 9692
rect 13491 7988 13557 7989
rect 13491 7924 13492 7988
rect 13556 7924 13557 7988
rect 13491 7923 13557 7924
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12571 5132 12637 5133
rect 12571 5068 12572 5132
rect 12636 5068 12637 5132
rect 12571 5067 12637 5068
rect 12387 4996 12453 4997
rect 12387 4932 12388 4996
rect 12452 4932 12453 4996
rect 12387 4931 12453 4932
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 11467 4588 11533 4589
rect 11467 4524 11468 4588
rect 11532 4524 11533 4588
rect 11467 4523 11533 4524
rect 9259 4044 9325 4045
rect 9259 3980 9260 4044
rect 9324 3980 9325 4044
rect 9259 3979 9325 3980
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 13678 2821 13738 9691
rect 13862 5813 13922 12003
rect 14046 10981 14106 24243
rect 15518 23493 15578 25739
rect 21403 25532 21469 25533
rect 21403 25468 21404 25532
rect 21468 25468 21469 25532
rect 21403 25467 21469 25468
rect 20299 24580 20365 24581
rect 17944 23968 18264 24528
rect 20299 24516 20300 24580
rect 20364 24516 20365 24580
rect 20299 24515 20365 24516
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 16803 23900 16869 23901
rect 16803 23836 16804 23900
rect 16868 23836 16869 23900
rect 16803 23835 16869 23836
rect 14963 23492 15029 23493
rect 14963 23428 14964 23492
rect 15028 23428 15029 23492
rect 14963 23427 15029 23428
rect 15515 23492 15581 23493
rect 15515 23428 15516 23492
rect 15580 23428 15581 23492
rect 15515 23427 15581 23428
rect 14966 21589 15026 23427
rect 15515 23356 15581 23357
rect 15515 23292 15516 23356
rect 15580 23292 15581 23356
rect 15515 23291 15581 23292
rect 14963 21588 15029 21589
rect 14963 21524 14964 21588
rect 15028 21524 15029 21588
rect 14963 21523 15029 21524
rect 14966 21181 15026 21523
rect 14963 21180 15029 21181
rect 14963 21116 14964 21180
rect 15028 21116 15029 21180
rect 14963 21115 15029 21116
rect 14779 19684 14845 19685
rect 14779 19620 14780 19684
rect 14844 19620 14845 19684
rect 14779 19619 14845 19620
rect 14227 18868 14293 18869
rect 14227 18804 14228 18868
rect 14292 18804 14293 18868
rect 14227 18803 14293 18804
rect 14043 10980 14109 10981
rect 14043 10916 14044 10980
rect 14108 10916 14109 10980
rect 14043 10915 14109 10916
rect 14043 10300 14109 10301
rect 14043 10236 14044 10300
rect 14108 10236 14109 10300
rect 14043 10235 14109 10236
rect 13859 5812 13925 5813
rect 13859 5748 13860 5812
rect 13924 5748 13925 5812
rect 13859 5747 13925 5748
rect 13675 2820 13741 2821
rect 13675 2756 13676 2820
rect 13740 2756 13741 2820
rect 13675 2755 13741 2756
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 8891 2684 8957 2685
rect 8891 2620 8892 2684
rect 8956 2620 8957 2684
rect 8891 2619 8957 2620
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 2128 13264 2688
rect 14046 2005 14106 10235
rect 14230 9349 14290 18803
rect 14595 17236 14661 17237
rect 14595 17172 14596 17236
rect 14660 17172 14661 17236
rect 14595 17171 14661 17172
rect 14411 12612 14477 12613
rect 14411 12548 14412 12612
rect 14476 12548 14477 12612
rect 14411 12547 14477 12548
rect 14414 11797 14474 12547
rect 14411 11796 14477 11797
rect 14411 11732 14412 11796
rect 14476 11732 14477 11796
rect 14411 11731 14477 11732
rect 14598 10029 14658 17171
rect 14782 13973 14842 19619
rect 15331 18188 15397 18189
rect 15331 18124 15332 18188
rect 15396 18124 15397 18188
rect 15331 18123 15397 18124
rect 15147 16964 15213 16965
rect 15147 16900 15148 16964
rect 15212 16900 15213 16964
rect 15147 16899 15213 16900
rect 15150 14517 15210 16899
rect 15147 14516 15213 14517
rect 15147 14452 15148 14516
rect 15212 14452 15213 14516
rect 15147 14451 15213 14452
rect 14779 13972 14845 13973
rect 14779 13908 14780 13972
rect 14844 13908 14845 13972
rect 14779 13907 14845 13908
rect 15147 12340 15213 12341
rect 15147 12276 15148 12340
rect 15212 12276 15213 12340
rect 15147 12275 15213 12276
rect 14779 11932 14845 11933
rect 14779 11868 14780 11932
rect 14844 11868 14845 11932
rect 14779 11867 14845 11868
rect 14782 11253 14842 11867
rect 14779 11252 14845 11253
rect 14779 11188 14780 11252
rect 14844 11188 14845 11252
rect 14779 11187 14845 11188
rect 14779 11116 14845 11117
rect 14779 11052 14780 11116
rect 14844 11052 14845 11116
rect 14779 11051 14845 11052
rect 14782 10437 14842 11051
rect 14963 10844 15029 10845
rect 14963 10780 14964 10844
rect 15028 10780 15029 10844
rect 14963 10779 15029 10780
rect 14779 10436 14845 10437
rect 14779 10372 14780 10436
rect 14844 10372 14845 10436
rect 14779 10371 14845 10372
rect 14595 10028 14661 10029
rect 14595 9964 14596 10028
rect 14660 9964 14661 10028
rect 14595 9963 14661 9964
rect 14227 9348 14293 9349
rect 14227 9284 14228 9348
rect 14292 9284 14293 9348
rect 14227 9283 14293 9284
rect 14230 4045 14290 9283
rect 14966 5813 15026 10779
rect 15150 7581 15210 12275
rect 15147 7580 15213 7581
rect 15147 7516 15148 7580
rect 15212 7516 15213 7580
rect 15147 7515 15213 7516
rect 15334 6765 15394 18123
rect 15518 13565 15578 23291
rect 16619 22132 16685 22133
rect 16619 22068 16620 22132
rect 16684 22068 16685 22132
rect 16619 22067 16685 22068
rect 16622 20501 16682 22067
rect 16619 20500 16685 20501
rect 16619 20436 16620 20500
rect 16684 20436 16685 20500
rect 16619 20435 16685 20436
rect 16806 18461 16866 23835
rect 17944 22880 18264 23904
rect 18827 23356 18893 23357
rect 18827 23292 18828 23356
rect 18892 23292 18893 23356
rect 18827 23291 18893 23292
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17539 22676 17605 22677
rect 17539 22612 17540 22676
rect 17604 22612 17605 22676
rect 17539 22611 17605 22612
rect 17542 22110 17602 22611
rect 17542 22050 17786 22110
rect 17539 21724 17605 21725
rect 17539 21660 17540 21724
rect 17604 21660 17605 21724
rect 17539 21659 17605 21660
rect 17171 21452 17237 21453
rect 17171 21388 17172 21452
rect 17236 21388 17237 21452
rect 17171 21387 17237 21388
rect 16987 19548 17053 19549
rect 16987 19484 16988 19548
rect 17052 19484 17053 19548
rect 16987 19483 17053 19484
rect 16803 18460 16869 18461
rect 16803 18396 16804 18460
rect 16868 18396 16869 18460
rect 16803 18395 16869 18396
rect 16619 17236 16685 17237
rect 16619 17172 16620 17236
rect 16684 17172 16685 17236
rect 16619 17171 16685 17172
rect 16435 16692 16501 16693
rect 16435 16628 16436 16692
rect 16500 16628 16501 16692
rect 16435 16627 16501 16628
rect 16251 16284 16317 16285
rect 16251 16220 16252 16284
rect 16316 16220 16317 16284
rect 16251 16219 16317 16220
rect 15699 15060 15765 15061
rect 15699 14996 15700 15060
rect 15764 14996 15765 15060
rect 15699 14995 15765 14996
rect 15515 13564 15581 13565
rect 15515 13500 15516 13564
rect 15580 13500 15581 13564
rect 15515 13499 15581 13500
rect 15515 10028 15581 10029
rect 15515 9964 15516 10028
rect 15580 9964 15581 10028
rect 15515 9963 15581 9964
rect 15518 8261 15578 9963
rect 15702 9893 15762 14995
rect 15883 13700 15949 13701
rect 15883 13636 15884 13700
rect 15948 13636 15949 13700
rect 15883 13635 15949 13636
rect 15699 9892 15765 9893
rect 15699 9828 15700 9892
rect 15764 9828 15765 9892
rect 15699 9827 15765 9828
rect 15886 9077 15946 13635
rect 16254 9690 16314 16219
rect 16438 12885 16498 16627
rect 16622 14517 16682 17171
rect 16619 14516 16685 14517
rect 16619 14452 16620 14516
rect 16684 14452 16685 14516
rect 16619 14451 16685 14452
rect 16435 12884 16501 12885
rect 16435 12820 16436 12884
rect 16500 12820 16501 12884
rect 16435 12819 16501 12820
rect 16803 12340 16869 12341
rect 16803 12276 16804 12340
rect 16868 12276 16869 12340
rect 16803 12275 16869 12276
rect 16254 9630 16682 9690
rect 15883 9076 15949 9077
rect 15883 9012 15884 9076
rect 15948 9012 15949 9076
rect 15883 9011 15949 9012
rect 16435 8668 16501 8669
rect 16435 8604 16436 8668
rect 16500 8604 16501 8668
rect 16435 8603 16501 8604
rect 15515 8260 15581 8261
rect 15515 8196 15516 8260
rect 15580 8196 15581 8260
rect 15515 8195 15581 8196
rect 15331 6764 15397 6765
rect 15331 6700 15332 6764
rect 15396 6700 15397 6764
rect 15331 6699 15397 6700
rect 16438 5813 16498 8603
rect 14963 5812 15029 5813
rect 14963 5748 14964 5812
rect 15028 5748 15029 5812
rect 14963 5747 15029 5748
rect 16435 5812 16501 5813
rect 16435 5748 16436 5812
rect 16500 5748 16501 5812
rect 16435 5747 16501 5748
rect 16622 5541 16682 9630
rect 16806 9349 16866 12275
rect 16803 9348 16869 9349
rect 16803 9284 16804 9348
rect 16868 9284 16869 9348
rect 16803 9283 16869 9284
rect 16619 5540 16685 5541
rect 16619 5476 16620 5540
rect 16684 5476 16685 5540
rect 16619 5475 16685 5476
rect 16990 4317 17050 19483
rect 17174 15877 17234 21387
rect 17542 20770 17602 21659
rect 17726 21181 17786 22050
rect 17944 21792 18264 22816
rect 18830 22110 18890 23291
rect 19379 22812 19445 22813
rect 19379 22748 19380 22812
rect 19444 22748 19445 22812
rect 19379 22747 19445 22748
rect 18830 22050 19258 22110
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17723 21180 17789 21181
rect 17723 21116 17724 21180
rect 17788 21116 17789 21180
rect 17723 21115 17789 21116
rect 17542 20710 17786 20770
rect 17539 20636 17605 20637
rect 17539 20572 17540 20636
rect 17604 20572 17605 20636
rect 17539 20571 17605 20572
rect 17355 20092 17421 20093
rect 17355 20028 17356 20092
rect 17420 20028 17421 20092
rect 17355 20027 17421 20028
rect 17358 19141 17418 20027
rect 17355 19140 17421 19141
rect 17355 19076 17356 19140
rect 17420 19076 17421 19140
rect 17355 19075 17421 19076
rect 17542 18461 17602 20571
rect 17539 18460 17605 18461
rect 17539 18396 17540 18460
rect 17604 18396 17605 18460
rect 17539 18395 17605 18396
rect 17726 16965 17786 20710
rect 17944 20704 18264 21728
rect 19198 21181 19258 22050
rect 19382 21861 19442 22747
rect 20302 22405 20362 24515
rect 20483 24036 20549 24037
rect 20483 23972 20484 24036
rect 20548 23972 20549 24036
rect 20483 23971 20549 23972
rect 20299 22404 20365 22405
rect 20299 22340 20300 22404
rect 20364 22340 20365 22404
rect 20299 22339 20365 22340
rect 19747 22132 19813 22133
rect 19747 22068 19748 22132
rect 19812 22068 19813 22132
rect 19747 22067 19813 22068
rect 19379 21860 19445 21861
rect 19379 21796 19380 21860
rect 19444 21796 19445 21860
rect 19379 21795 19445 21796
rect 19011 21180 19077 21181
rect 19011 21116 19012 21180
rect 19076 21116 19077 21180
rect 19011 21115 19077 21116
rect 19195 21180 19261 21181
rect 19195 21116 19196 21180
rect 19260 21116 19261 21180
rect 19195 21115 19261 21116
rect 18459 20772 18525 20773
rect 18459 20708 18460 20772
rect 18524 20708 18525 20772
rect 18459 20707 18525 20708
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 18462 18597 18522 20707
rect 18827 19140 18893 19141
rect 18827 19076 18828 19140
rect 18892 19076 18893 19140
rect 18827 19075 18893 19076
rect 18459 18596 18525 18597
rect 18459 18532 18460 18596
rect 18524 18532 18525 18596
rect 18459 18531 18525 18532
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 18830 18461 18890 19075
rect 18827 18460 18893 18461
rect 18827 18396 18828 18460
rect 18892 18396 18893 18460
rect 18827 18395 18893 18396
rect 18827 18324 18893 18325
rect 18827 18260 18828 18324
rect 18892 18260 18893 18324
rect 18827 18259 18893 18260
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17723 16964 17789 16965
rect 17723 16900 17724 16964
rect 17788 16900 17789 16964
rect 17723 16899 17789 16900
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17171 15876 17237 15877
rect 17171 15812 17172 15876
rect 17236 15812 17237 15876
rect 17171 15811 17237 15812
rect 17355 15604 17421 15605
rect 17355 15540 17356 15604
rect 17420 15540 17421 15604
rect 17355 15539 17421 15540
rect 17171 15196 17237 15197
rect 17171 15132 17172 15196
rect 17236 15132 17237 15196
rect 17171 15131 17237 15132
rect 17174 11389 17234 15131
rect 17171 11388 17237 11389
rect 17171 11324 17172 11388
rect 17236 11324 17237 11388
rect 17171 11323 17237 11324
rect 17358 10029 17418 15539
rect 17944 15264 18264 16288
rect 18459 15332 18525 15333
rect 18459 15268 18460 15332
rect 18524 15268 18525 15332
rect 18459 15267 18525 15268
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17723 13020 17789 13021
rect 17723 12956 17724 13020
rect 17788 12956 17789 13020
rect 17723 12955 17789 12956
rect 17726 12341 17786 12955
rect 17723 12340 17789 12341
rect 17723 12276 17724 12340
rect 17788 12276 17789 12340
rect 17723 12275 17789 12276
rect 17944 12000 18264 13024
rect 18462 13021 18522 15267
rect 18830 14109 18890 18259
rect 19014 16965 19074 21115
rect 19379 20908 19445 20909
rect 19379 20844 19380 20908
rect 19444 20844 19445 20908
rect 19379 20843 19445 20844
rect 19011 16964 19077 16965
rect 19011 16900 19012 16964
rect 19076 16900 19077 16964
rect 19011 16899 19077 16900
rect 19382 16421 19442 20843
rect 19750 20637 19810 22067
rect 20486 21997 20546 23971
rect 20483 21996 20549 21997
rect 20483 21932 20484 21996
rect 20548 21932 20549 21996
rect 20483 21931 20549 21932
rect 19563 20636 19629 20637
rect 19563 20572 19564 20636
rect 19628 20572 19629 20636
rect 19563 20571 19629 20572
rect 19747 20636 19813 20637
rect 19747 20572 19748 20636
rect 19812 20572 19813 20636
rect 19747 20571 19813 20572
rect 19195 16420 19261 16421
rect 19195 16356 19196 16420
rect 19260 16356 19261 16420
rect 19195 16355 19261 16356
rect 19379 16420 19445 16421
rect 19379 16356 19380 16420
rect 19444 16356 19445 16420
rect 19379 16355 19445 16356
rect 19011 15604 19077 15605
rect 19011 15540 19012 15604
rect 19076 15540 19077 15604
rect 19011 15539 19077 15540
rect 18827 14108 18893 14109
rect 18827 14044 18828 14108
rect 18892 14044 18893 14108
rect 18827 14043 18893 14044
rect 18643 13700 18709 13701
rect 18643 13636 18644 13700
rect 18708 13636 18709 13700
rect 18643 13635 18709 13636
rect 18459 13020 18525 13021
rect 18459 12956 18460 13020
rect 18524 12956 18525 13020
rect 18459 12955 18525 12956
rect 18459 12476 18525 12477
rect 18459 12412 18460 12476
rect 18524 12412 18525 12476
rect 18459 12411 18525 12412
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 18462 10981 18522 12411
rect 18459 10980 18525 10981
rect 18459 10916 18460 10980
rect 18524 10916 18525 10980
rect 18459 10915 18525 10916
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17355 10028 17421 10029
rect 17355 9964 17356 10028
rect 17420 9964 17421 10028
rect 17355 9963 17421 9964
rect 17944 9824 18264 10848
rect 18646 9893 18706 13635
rect 18643 9892 18709 9893
rect 18643 9828 18644 9892
rect 18708 9828 18709 9892
rect 18643 9827 18709 9828
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 18830 8125 18890 14043
rect 18827 8124 18893 8125
rect 18827 8060 18828 8124
rect 18892 8060 18893 8124
rect 18827 8059 18893 8060
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 19014 4725 19074 15539
rect 19198 12477 19258 16355
rect 19566 15741 19626 20571
rect 19747 19684 19813 19685
rect 19747 19620 19748 19684
rect 19812 19620 19813 19684
rect 19747 19619 19813 19620
rect 19750 17781 19810 19619
rect 20299 18596 20365 18597
rect 20299 18532 20300 18596
rect 20364 18532 20365 18596
rect 20299 18531 20365 18532
rect 21035 18596 21101 18597
rect 21035 18532 21036 18596
rect 21100 18532 21101 18596
rect 21035 18531 21101 18532
rect 20115 17916 20181 17917
rect 20115 17852 20116 17916
rect 20180 17852 20181 17916
rect 20115 17851 20181 17852
rect 19747 17780 19813 17781
rect 19747 17716 19748 17780
rect 19812 17716 19813 17780
rect 19747 17715 19813 17716
rect 19747 15876 19813 15877
rect 19747 15812 19748 15876
rect 19812 15812 19813 15876
rect 19747 15811 19813 15812
rect 19563 15740 19629 15741
rect 19563 15676 19564 15740
rect 19628 15676 19629 15740
rect 19563 15675 19629 15676
rect 19379 15332 19445 15333
rect 19379 15268 19380 15332
rect 19444 15268 19445 15332
rect 19379 15267 19445 15268
rect 19195 12476 19261 12477
rect 19195 12412 19196 12476
rect 19260 12412 19261 12476
rect 19195 12411 19261 12412
rect 19382 9485 19442 15267
rect 19563 12612 19629 12613
rect 19563 12548 19564 12612
rect 19628 12548 19629 12612
rect 19563 12547 19629 12548
rect 19379 9484 19445 9485
rect 19379 9420 19380 9484
rect 19444 9420 19445 9484
rect 19379 9419 19445 9420
rect 19566 8397 19626 12547
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19750 6765 19810 15811
rect 19931 14244 19997 14245
rect 19931 14180 19932 14244
rect 19996 14180 19997 14244
rect 19931 14179 19997 14180
rect 19934 12069 19994 14179
rect 19931 12068 19997 12069
rect 19931 12004 19932 12068
rect 19996 12004 19997 12068
rect 19931 12003 19997 12004
rect 19931 11524 19997 11525
rect 19931 11460 19932 11524
rect 19996 11460 19997 11524
rect 19931 11459 19997 11460
rect 19747 6764 19813 6765
rect 19747 6700 19748 6764
rect 19812 6700 19813 6764
rect 19747 6699 19813 6700
rect 19011 4724 19077 4725
rect 19011 4660 19012 4724
rect 19076 4660 19077 4724
rect 19011 4659 19077 4660
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 16987 4316 17053 4317
rect 16987 4252 16988 4316
rect 17052 4252 17053 4316
rect 16987 4251 17053 4252
rect 14227 4044 14293 4045
rect 14227 3980 14228 4044
rect 14292 3980 14293 4044
rect 14227 3979 14293 3980
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 19934 2685 19994 11459
rect 20118 8805 20178 17851
rect 20302 10437 20362 18531
rect 20851 17372 20917 17373
rect 20851 17308 20852 17372
rect 20916 17308 20917 17372
rect 20851 17307 20917 17308
rect 20667 15604 20733 15605
rect 20667 15540 20668 15604
rect 20732 15540 20733 15604
rect 20667 15539 20733 15540
rect 20670 13157 20730 15539
rect 20854 13973 20914 17307
rect 20851 13972 20917 13973
rect 20851 13908 20852 13972
rect 20916 13908 20917 13972
rect 20851 13907 20917 13908
rect 20667 13156 20733 13157
rect 20667 13092 20668 13156
rect 20732 13092 20733 13156
rect 20667 13091 20733 13092
rect 20299 10436 20365 10437
rect 20299 10372 20300 10436
rect 20364 10372 20365 10436
rect 20299 10371 20365 10372
rect 21038 9485 21098 18531
rect 21406 17373 21466 25467
rect 27659 25260 27725 25261
rect 27659 25196 27660 25260
rect 27724 25196 27725 25260
rect 27659 25195 27725 25196
rect 27475 25124 27541 25125
rect 27475 25060 27476 25124
rect 27540 25060 27541 25124
rect 27475 25059 27541 25060
rect 23611 24852 23677 24853
rect 23611 24788 23612 24852
rect 23676 24788 23677 24852
rect 23611 24787 23677 24788
rect 22944 24512 23264 24528
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 21587 22404 21653 22405
rect 21587 22340 21588 22404
rect 21652 22340 21653 22404
rect 21587 22339 21653 22340
rect 22691 22404 22757 22405
rect 22691 22340 22692 22404
rect 22756 22340 22757 22404
rect 22691 22339 22757 22340
rect 21403 17372 21469 17373
rect 21403 17308 21404 17372
rect 21468 17308 21469 17372
rect 21403 17307 21469 17308
rect 21590 14789 21650 22339
rect 21958 20574 22386 20634
rect 21958 20501 22018 20574
rect 22326 20501 22386 20574
rect 21955 20500 22021 20501
rect 21955 20436 21956 20500
rect 22020 20436 22021 20500
rect 21955 20435 22021 20436
rect 22323 20500 22389 20501
rect 22323 20436 22324 20500
rect 22388 20436 22389 20500
rect 22323 20435 22389 20436
rect 21771 19548 21837 19549
rect 21771 19484 21772 19548
rect 21836 19484 21837 19548
rect 21771 19483 21837 19484
rect 22507 19548 22573 19549
rect 22507 19484 22508 19548
rect 22572 19484 22573 19548
rect 22507 19483 22573 19484
rect 21587 14788 21653 14789
rect 21587 14724 21588 14788
rect 21652 14724 21653 14788
rect 21587 14723 21653 14724
rect 21587 14652 21653 14653
rect 21587 14588 21588 14652
rect 21652 14588 21653 14652
rect 21587 14587 21653 14588
rect 21403 12884 21469 12885
rect 21403 12820 21404 12884
rect 21468 12820 21469 12884
rect 21403 12819 21469 12820
rect 21406 10709 21466 12819
rect 21590 10981 21650 14587
rect 21587 10980 21653 10981
rect 21587 10916 21588 10980
rect 21652 10916 21653 10980
rect 21587 10915 21653 10916
rect 21403 10708 21469 10709
rect 21403 10644 21404 10708
rect 21468 10644 21469 10708
rect 21403 10643 21469 10644
rect 21403 9756 21469 9757
rect 21403 9692 21404 9756
rect 21468 9692 21469 9756
rect 21403 9691 21469 9692
rect 21035 9484 21101 9485
rect 21035 9420 21036 9484
rect 21100 9420 21101 9484
rect 21035 9419 21101 9420
rect 20115 8804 20181 8805
rect 20115 8740 20116 8804
rect 20180 8740 20181 8804
rect 20115 8739 20181 8740
rect 21406 7581 21466 9691
rect 21403 7580 21469 7581
rect 21403 7516 21404 7580
rect 21468 7516 21469 7580
rect 21403 7515 21469 7516
rect 21774 4725 21834 19483
rect 22047 17508 22113 17509
rect 22047 17444 22048 17508
rect 22112 17444 22113 17508
rect 22047 17443 22113 17444
rect 22050 17370 22110 17443
rect 22050 17310 22202 17370
rect 21955 16556 22021 16557
rect 21955 16492 21956 16556
rect 22020 16492 22021 16556
rect 21955 16491 22021 16492
rect 21958 14109 22018 16491
rect 22142 15605 22202 17310
rect 22323 15740 22389 15741
rect 22323 15676 22324 15740
rect 22388 15676 22389 15740
rect 22323 15675 22389 15676
rect 22139 15604 22205 15605
rect 22139 15540 22140 15604
rect 22204 15540 22205 15604
rect 22139 15539 22205 15540
rect 22326 14381 22386 15675
rect 22323 14380 22389 14381
rect 22323 14316 22324 14380
rect 22388 14316 22389 14380
rect 22323 14315 22389 14316
rect 21955 14108 22021 14109
rect 21955 14044 21956 14108
rect 22020 14044 22021 14108
rect 21955 14043 22021 14044
rect 22139 13700 22205 13701
rect 22139 13636 22140 13700
rect 22204 13636 22205 13700
rect 22139 13635 22205 13636
rect 22142 10981 22202 13635
rect 22323 12612 22389 12613
rect 22323 12548 22324 12612
rect 22388 12548 22389 12612
rect 22323 12547 22389 12548
rect 21955 10980 22021 10981
rect 21955 10916 21956 10980
rect 22020 10916 22021 10980
rect 21955 10915 22021 10916
rect 22139 10980 22205 10981
rect 22139 10916 22140 10980
rect 22204 10916 22205 10980
rect 22139 10915 22205 10916
rect 21958 9893 22018 10915
rect 21955 9892 22021 9893
rect 21955 9828 21956 9892
rect 22020 9828 22021 9892
rect 21955 9827 22021 9828
rect 21771 4724 21837 4725
rect 21771 4660 21772 4724
rect 21836 4660 21837 4724
rect 21771 4659 21837 4660
rect 19931 2684 19997 2685
rect 19931 2620 19932 2684
rect 19996 2620 19997 2684
rect 19931 2619 19997 2620
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 14043 2004 14109 2005
rect 14043 1940 14044 2004
rect 14108 1940 14109 2004
rect 14043 1939 14109 1940
rect 22326 1189 22386 12547
rect 22510 5677 22570 19483
rect 22694 16421 22754 22339
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 23427 17372 23493 17373
rect 23427 17308 23428 17372
rect 23492 17308 23493 17372
rect 23427 17307 23493 17308
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22691 16420 22757 16421
rect 22691 16356 22692 16420
rect 22756 16356 22757 16420
rect 22691 16355 22757 16356
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22691 14788 22757 14789
rect 22691 14724 22692 14788
rect 22756 14724 22757 14788
rect 22691 14723 22757 14724
rect 22694 13021 22754 14723
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 23430 14653 23490 17307
rect 23614 16285 23674 24787
rect 25451 24580 25517 24581
rect 25451 24516 25452 24580
rect 25516 24516 25517 24580
rect 25451 24515 25517 24516
rect 24715 23492 24781 23493
rect 24715 23428 24716 23492
rect 24780 23428 24781 23492
rect 24715 23427 24781 23428
rect 24531 20772 24597 20773
rect 24531 20708 24532 20772
rect 24596 20708 24597 20772
rect 24531 20707 24597 20708
rect 24163 20364 24229 20365
rect 24163 20300 24164 20364
rect 24228 20300 24229 20364
rect 24163 20299 24229 20300
rect 23611 16284 23677 16285
rect 23611 16220 23612 16284
rect 23676 16220 23677 16284
rect 23611 16219 23677 16220
rect 24166 15877 24226 20299
rect 24163 15876 24229 15877
rect 24163 15812 24164 15876
rect 24228 15812 24229 15876
rect 24163 15811 24229 15812
rect 23427 14652 23493 14653
rect 23427 14588 23428 14652
rect 23492 14588 23493 14652
rect 23427 14587 23493 14588
rect 24347 14652 24413 14653
rect 24347 14588 24348 14652
rect 24412 14588 24413 14652
rect 24347 14587 24413 14588
rect 23795 13972 23861 13973
rect 23795 13908 23796 13972
rect 23860 13908 23861 13972
rect 23795 13907 23861 13908
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22691 13020 22757 13021
rect 22691 12956 22692 13020
rect 22756 12956 22757 13020
rect 22691 12955 22757 12956
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 23798 12341 23858 13907
rect 23795 12340 23861 12341
rect 23795 12276 23796 12340
rect 23860 12276 23861 12340
rect 23795 12275 23861 12276
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22507 5676 22573 5677
rect 22507 5612 22508 5676
rect 22572 5612 22573 5676
rect 22507 5611 22573 5612
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 24350 4181 24410 14587
rect 24347 4180 24413 4181
rect 24347 4116 24348 4180
rect 24412 4116 24413 4180
rect 24347 4115 24413 4116
rect 24534 4045 24594 20707
rect 24531 4044 24597 4045
rect 24531 3980 24532 4044
rect 24596 3980 24597 4044
rect 24531 3979 24597 3980
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 24718 3093 24778 23427
rect 25267 16828 25333 16829
rect 25267 16764 25268 16828
rect 25332 16764 25333 16828
rect 25267 16763 25333 16764
rect 25083 16284 25149 16285
rect 25083 16220 25084 16284
rect 25148 16220 25149 16284
rect 25083 16219 25149 16220
rect 24899 13020 24965 13021
rect 24899 12956 24900 13020
rect 24964 12956 24965 13020
rect 24899 12955 24965 12956
rect 24902 10437 24962 12955
rect 25086 11661 25146 16219
rect 25083 11660 25149 11661
rect 25083 11596 25084 11660
rect 25148 11596 25149 11660
rect 25083 11595 25149 11596
rect 24899 10436 24965 10437
rect 24899 10372 24900 10436
rect 24964 10372 24965 10436
rect 24899 10371 24965 10372
rect 25270 8669 25330 16763
rect 25454 14653 25514 24515
rect 27291 23492 27357 23493
rect 27291 23428 27292 23492
rect 27356 23428 27357 23492
rect 27291 23427 27357 23428
rect 26003 22404 26069 22405
rect 26003 22340 26004 22404
rect 26068 22340 26069 22404
rect 26003 22339 26069 22340
rect 25819 20772 25885 20773
rect 25819 20708 25820 20772
rect 25884 20708 25885 20772
rect 25819 20707 25885 20708
rect 25635 19548 25701 19549
rect 25635 19484 25636 19548
rect 25700 19484 25701 19548
rect 25635 19483 25701 19484
rect 25638 16285 25698 19483
rect 25635 16284 25701 16285
rect 25635 16220 25636 16284
rect 25700 16220 25701 16284
rect 25635 16219 25701 16220
rect 25451 14652 25517 14653
rect 25451 14588 25452 14652
rect 25516 14588 25517 14652
rect 25451 14587 25517 14588
rect 25267 8668 25333 8669
rect 25267 8604 25268 8668
rect 25332 8604 25333 8668
rect 25267 8603 25333 8604
rect 24715 3092 24781 3093
rect 24715 3028 24716 3092
rect 24780 3028 24781 3092
rect 24715 3027 24781 3028
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22944 2128 23264 2688
rect 25822 2685 25882 20707
rect 26006 14789 26066 22339
rect 26187 21044 26253 21045
rect 26187 20980 26188 21044
rect 26252 20980 26253 21044
rect 26187 20979 26253 20980
rect 26190 18189 26250 20979
rect 26555 19140 26621 19141
rect 26555 19076 26556 19140
rect 26620 19076 26621 19140
rect 26555 19075 26621 19076
rect 26187 18188 26253 18189
rect 26187 18124 26188 18188
rect 26252 18124 26253 18188
rect 26187 18123 26253 18124
rect 26187 18052 26253 18053
rect 26187 17988 26188 18052
rect 26252 17988 26253 18052
rect 26187 17987 26253 17988
rect 26003 14788 26069 14789
rect 26003 14724 26004 14788
rect 26068 14724 26069 14788
rect 26003 14723 26069 14724
rect 26190 3637 26250 17987
rect 26187 3636 26253 3637
rect 26187 3572 26188 3636
rect 26252 3572 26253 3636
rect 26187 3571 26253 3572
rect 25819 2684 25885 2685
rect 25819 2620 25820 2684
rect 25884 2620 25885 2684
rect 25819 2619 25885 2620
rect 22323 1188 22389 1189
rect 22323 1124 22324 1188
rect 22388 1124 22389 1188
rect 22323 1123 22389 1124
rect 5763 1052 5829 1053
rect 5763 988 5764 1052
rect 5828 988 5829 1052
rect 5763 987 5829 988
rect 26558 781 26618 19075
rect 27294 12205 27354 23427
rect 27478 20229 27538 25059
rect 27475 20228 27541 20229
rect 27475 20164 27476 20228
rect 27540 20164 27541 20228
rect 27475 20163 27541 20164
rect 27291 12204 27357 12205
rect 27291 12140 27292 12204
rect 27356 12140 27357 12204
rect 27291 12139 27357 12140
rect 27478 10845 27538 20163
rect 27662 18053 27722 25195
rect 27944 23968 28264 24528
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 32944 24512 33264 24528
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 28763 22268 28829 22269
rect 28763 22204 28764 22268
rect 28828 22204 28829 22268
rect 28763 22203 28829 22204
rect 28766 22110 28826 22203
rect 28766 22050 29010 22110
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 28579 19548 28645 19549
rect 28579 19484 28580 19548
rect 28644 19484 28645 19548
rect 28579 19483 28645 19484
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27659 18052 27725 18053
rect 27659 17988 27660 18052
rect 27724 17988 27725 18052
rect 27659 17987 27725 17988
rect 27659 17916 27725 17917
rect 27659 17852 27660 17916
rect 27724 17852 27725 17916
rect 27659 17851 27725 17852
rect 27662 15741 27722 17851
rect 27944 17440 28264 18464
rect 28395 18052 28461 18053
rect 28395 17988 28396 18052
rect 28460 17988 28461 18052
rect 28395 17987 28461 17988
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27659 15740 27725 15741
rect 27659 15676 27660 15740
rect 27724 15676 27725 15740
rect 27659 15675 27725 15676
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 28398 15197 28458 17987
rect 28582 17509 28642 19483
rect 28950 18733 29010 22050
rect 29499 21860 29565 21861
rect 29499 21796 29500 21860
rect 29564 21796 29565 21860
rect 29499 21795 29565 21796
rect 29131 19004 29197 19005
rect 29131 18940 29132 19004
rect 29196 18940 29197 19004
rect 29131 18939 29197 18940
rect 28947 18732 29013 18733
rect 28947 18668 28948 18732
rect 29012 18668 29013 18732
rect 28947 18667 29013 18668
rect 28579 17508 28645 17509
rect 28579 17444 28580 17508
rect 28644 17444 28645 17508
rect 28579 17443 28645 17444
rect 28947 16828 29013 16829
rect 28947 16764 28948 16828
rect 29012 16764 29013 16828
rect 28947 16763 29013 16764
rect 28395 15196 28461 15197
rect 28395 15132 28396 15196
rect 28460 15132 28461 15196
rect 28395 15131 28461 15132
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 28950 13157 29010 16763
rect 29134 15061 29194 18939
rect 29315 18596 29381 18597
rect 29315 18532 29316 18596
rect 29380 18532 29381 18596
rect 29315 18531 29381 18532
rect 29318 16829 29378 18531
rect 29315 16828 29381 16829
rect 29315 16764 29316 16828
rect 29380 16764 29381 16828
rect 29315 16763 29381 16764
rect 29131 15060 29197 15061
rect 29131 14996 29132 15060
rect 29196 14996 29197 15060
rect 29131 14995 29197 14996
rect 28947 13156 29013 13157
rect 28947 13092 28948 13156
rect 29012 13092 29013 13156
rect 28947 13091 29013 13092
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27475 10844 27541 10845
rect 27475 10780 27476 10844
rect 27540 10780 27541 10844
rect 27475 10779 27541 10780
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 29502 6357 29562 21795
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 30419 20364 30485 20365
rect 30419 20300 30420 20364
rect 30484 20300 30485 20364
rect 30419 20299 30485 20300
rect 29683 18596 29749 18597
rect 29683 18532 29684 18596
rect 29748 18532 29749 18596
rect 29683 18531 29749 18532
rect 29686 17509 29746 18531
rect 30422 17781 30482 20299
rect 32944 20160 33264 21184
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 31523 19004 31589 19005
rect 31523 18940 31524 19004
rect 31588 18940 31589 19004
rect 31523 18939 31589 18940
rect 30419 17780 30485 17781
rect 30419 17716 30420 17780
rect 30484 17716 30485 17780
rect 30419 17715 30485 17716
rect 29683 17508 29749 17509
rect 29683 17444 29684 17508
rect 29748 17444 29749 17508
rect 29683 17443 29749 17444
rect 31526 15605 31586 18939
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32811 17508 32877 17509
rect 32811 17444 32812 17508
rect 32876 17444 32877 17508
rect 32811 17443 32877 17444
rect 31523 15604 31589 15605
rect 31523 15540 31524 15604
rect 31588 15540 31589 15604
rect 31523 15539 31589 15540
rect 32814 14789 32874 17443
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32811 14788 32877 14789
rect 32811 14724 32812 14788
rect 32876 14724 32877 14788
rect 32811 14723 32877 14724
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 29499 6356 29565 6357
rect 29499 6292 29500 6356
rect 29564 6292 29565 6356
rect 29499 6291 29565 6292
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 23968 38264 24528
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 24512 43264 24528
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 23968 48264 24528
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
rect 26555 780 26621 781
rect 26555 716 26556 780
rect 26620 716 26621 780
rect 26555 715 26621 716
use sky130_fd_sc_hd__clkbuf_2  _096_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23368 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _097_
timestamp 1679235063
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _098_
timestamp 1679235063
transform 1 0 4232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _099_
timestamp 1679235063
transform 1 0 7084 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _100_
timestamp 1679235063
transform 1 0 3956 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _101_
timestamp 1679235063
transform 1 0 6532 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _102_
timestamp 1679235063
transform 1 0 5888 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _103_
timestamp 1679235063
transform 1 0 6808 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _104_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 4140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _105_
timestamp 1679235063
transform 1 0 3128 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1679235063
transform 1 0 3956 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _107_
timestamp 1679235063
transform 1 0 16836 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _108_
timestamp 1679235063
transform 1 0 2392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _109_
timestamp 1679235063
transform 1 0 10764 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1679235063
transform 1 0 2024 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _111_
timestamp 1679235063
transform 1 0 3128 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1679235063
transform 1 0 5060 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1679235063
transform 1 0 26312 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1679235063
transform 1 0 18308 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1679235063
transform 1 0 24564 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1679235063
transform 1 0 2852 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _117_
timestamp 1679235063
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1679235063
transform 1 0 10856 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1679235063
transform 1 0 13432 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1679235063
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1679235063
transform 1 0 10672 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1679235063
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1679235063
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1679235063
transform 1 0 8280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1679235063
transform 1 0 14444 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1679235063
transform 1 0 24564 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1679235063
transform 1 0 14260 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1679235063
transform 1 0 24564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1679235063
transform 1 0 10856 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1679235063
transform 1 0 3496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1679235063
transform 1 0 5060 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _132_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24196 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1679235063
transform 1 0 27140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1679235063
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _135_
timestamp 1679235063
transform 1 0 22908 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1679235063
transform 1 0 5796 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _137_
timestamp 1679235063
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1679235063
transform 1 0 40756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _139_
timestamp 1679235063
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1679235063
transform 1 0 36616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1679235063
transform 1 0 34868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1679235063
transform 1 0 40020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1679235063
transform 1 0 34500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1679235063
transform 1 0 42596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1679235063
transform 1 0 37444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1679235063
transform 1 0 43332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1679235063
transform 1 0 25300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _148_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1679235063
transform 1 0 41124 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1679235063
transform 1 0 34040 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1679235063
transform 1 0 28244 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _152_
timestamp 1679235063
transform 1 0 20424 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _153_
timestamp 1679235063
transform 1 0 6532 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _154_
timestamp 1679235063
transform 1 0 3956 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _155_
timestamp 1679235063
transform 1 0 30820 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1679235063
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1679235063
transform 1 0 12420 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1679235063
transform 1 0 13984 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1679235063
transform 1 0 15732 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1679235063
transform 1 0 21620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1679235063
transform 1 0 16744 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1679235063
transform 1 0 23092 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1679235063
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1679235063
transform 1 0 14168 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1679235063
transform 1 0 26128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1679235063
transform 1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1679235063
transform 1 0 13340 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1679235063
transform 1 0 11500 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1679235063
transform 1 0 12512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1679235063
transform 1 0 5060 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1679235063
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1679235063
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1679235063
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1679235063
transform 1 0 11684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1679235063
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1679235063
transform 1 0 3220 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1679235063
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1679235063
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1679235063
transform 1 0 11500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1679235063
transform 1 0 5060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1679235063
transform 1 0 4232 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1679235063
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1679235063
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1679235063
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1679235063
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1679235063
transform 1 0 14168 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1679235063
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1679235063
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1679235063
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1679235063
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1679235063
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1679235063
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1679235063
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1679235063
transform 1 0 19228 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1679235063
transform 1 0 22448 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1679235063
transform 1 0 16560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__A
timestamp 1679235063
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1679235063
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1679235063
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1679235063
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1679235063
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1679235063
transform 1 0 18676 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1679235063
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1679235063
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1679235063
transform 1 0 2668 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1679235063
transform 1 0 5980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1679235063
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1679235063
transform 1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1679235063
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1679235063
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1679235063
transform 1 0 3312 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1679235063
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1679235063
transform 1 0 11684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1679235063
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1679235063
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1679235063
transform 1 0 15456 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1679235063
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1679235063
transform 1 0 25116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1679235063
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A
timestamp 1679235063
transform 1 0 24196 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1679235063
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1679235063
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1679235063
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A
timestamp 1679235063
transform 1 0 24748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A
timestamp 1679235063
transform 1 0 35420 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__A
timestamp 1679235063
transform 1 0 40756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A
timestamp 1679235063
transform 1 0 42504 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A
timestamp 1679235063
transform 1 0 36984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A
timestamp 1679235063
transform 1 0 43608 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1679235063
transform 1 0 42044 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A
timestamp 1679235063
transform 1 0 34316 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A
timestamp 1679235063
transform 1 0 28796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1679235063
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__156__A
timestamp 1679235063
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 9936 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 6440 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 8648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 11868 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 11776 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25944 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 1472 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 11500 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 9016 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__A0
timestamp 1679235063
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 34500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3864 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 1656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 15272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 4048 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 27140 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21988 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 34500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1679235063
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1679235063
transform 1 0 9660 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2__S
timestamp 1679235063
transform 1 0 3864 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A0
timestamp 1679235063
transform 1 0 3312 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__A1
timestamp 1679235063
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3__S
timestamp 1679235063
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A0
timestamp 1679235063
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__A1
timestamp 1679235063
transform 1 0 8648 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4__S
timestamp 1679235063
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 1564 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 5244 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1679235063
transform 1 0 1564 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2__S
timestamp 1679235063
transform 1 0 1472 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1679235063
transform 1 0 8832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__S
timestamp 1679235063
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0__S
timestamp 1679235063
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1__S
timestamp 1679235063
transform 1 0 16468 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 21528 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 21804 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 22356 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 23644 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23828 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR_A
timestamp 1679235063
transform 1 0 23736 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_A
timestamp 1679235063
transform 1 0 28152 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE_B_N
timestamp 1679235063
transform 1 0 27968 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE_TE_B
timestamp 1679235063
transform 1 0 16376 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 32016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_A
timestamp 1679235063
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_prog_clk_A
timestamp 1679235063
transform 1 0 13524 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_prog_clk_A
timestamp 1679235063
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_prog_clk_A
timestamp 1679235063
transform 1 0 16284 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_prog_clk_A
timestamp 1679235063
transform 1 0 14352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_prog_clk_A
timestamp 1679235063
transform 1 0 3312 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_prog_clk_A
timestamp 1679235063
transform 1 0 3312 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_prog_clk_A
timestamp 1679235063
transform 1 0 11868 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_prog_clk_A
timestamp 1679235063
transform 1 0 10304 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_prog_clk_A
timestamp 1679235063
transform 1 0 20976 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_prog_clk_A
timestamp 1679235063
transform 1 0 26312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_prog_clk_A
timestamp 1679235063
transform 1 0 22080 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_prog_clk_A
timestamp 1679235063
transform 1 0 18952 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_prog_clk_A
timestamp 1679235063
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_prog_clk_A
timestamp 1679235063
transform 1 0 23920 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_prog_clk_A
timestamp 1679235063
transform 1 0 25116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout143_A
timestamp 1679235063
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout144_A
timestamp 1679235063
transform 1 0 22540 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout145_A
timestamp 1679235063
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout146_A
timestamp 1679235063
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout148_A
timestamp 1679235063
transform 1 0 16744 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout149_A
timestamp 1679235063
transform 1 0 15180 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout150_A
timestamp 1679235063
transform 1 0 34316 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout151_A
timestamp 1679235063
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout152_A
timestamp 1679235063
transform 1 0 41308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold28_A
timestamp 1679235063
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold31_A
timestamp 1679235063
transform 1 0 36984 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold42_A
timestamp 1679235063
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold43_A
timestamp 1679235063
transform 1 0 34040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold82_A
timestamp 1679235063
transform 1 0 46092 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold88_A
timestamp 1679235063
transform 1 0 14168 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold95_A
timestamp 1679235063
transform 1 0 6164 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold113_A
timestamp 1679235063
transform 1 0 16284 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold137_A
timestamp 1679235063
transform 1 0 34224 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold139_A
timestamp 1679235063
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold147_A
timestamp 1679235063
transform 1 0 39468 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold151_A
timestamp 1679235063
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold157_A
timestamp 1679235063
transform 1 0 47012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold161_A
timestamp 1679235063
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold175_A
timestamp 1679235063
transform 1 0 31648 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold177_A
timestamp 1679235063
transform 1 0 11960 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold178_A
timestamp 1679235063
transform 1 0 47196 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold181_A
timestamp 1679235063
transform 1 0 39468 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold186_A
timestamp 1679235063
transform 1 0 29256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold190_A
timestamp 1679235063
transform 1 0 31004 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold211_A
timestamp 1679235063
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold217_A
timestamp 1679235063
transform 1 0 34408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold221_A
timestamp 1679235063
transform 1 0 32568 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold235_A
timestamp 1679235063
transform 1 0 9200 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold253_A
timestamp 1679235063
transform 1 0 36892 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold265_A
timestamp 1679235063
transform 1 0 3864 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold267_A
timestamp 1679235063
transform 1 0 37076 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold271_A
timestamp 1679235063
transform 1 0 41492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold285_A
timestamp 1679235063
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold286_A
timestamp 1679235063
transform 1 0 37076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold288_A
timestamp 1679235063
transform 1 0 45172 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold290_A
timestamp 1679235063
transform 1 0 30820 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold293_A
timestamp 1679235063
transform 1 0 32476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold305_A
timestamp 1679235063
transform 1 0 36708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold309_A
timestamp 1679235063
transform 1 0 44620 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold311_A
timestamp 1679235063
transform 1 0 11868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold312_A
timestamp 1679235063
transform 1 0 2668 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold314_A
timestamp 1679235063
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold315_A
timestamp 1679235063
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold316_A
timestamp 1679235063
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold317_A
timestamp 1679235063
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold322_A
timestamp 1679235063
transform 1 0 48300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1679235063
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1679235063
transform 1 0 10212 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1679235063
transform 1 0 10488 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1679235063
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1679235063
transform 1 0 22448 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1679235063
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1679235063
transform 1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1679235063
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1679235063
transform 1 0 18032 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1679235063
transform 1 0 20516 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1679235063
transform 1 0 21804 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1679235063
transform 1 0 18768 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1679235063
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1679235063
transform 1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1679235063
transform 1 0 26588 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1679235063
transform 1 0 14168 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1679235063
transform 1 0 19044 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1679235063
transform 1 0 29164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1679235063
transform 1 0 13064 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1679235063
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1679235063
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1679235063
transform 1 0 3404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1679235063
transform 1 0 8464 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1679235063
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1679235063
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1679235063
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1679235063
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1679235063
transform 1 0 18768 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1679235063
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1679235063
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1679235063
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1679235063
transform 1 0 43240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1679235063
transform 1 0 34500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1679235063
transform 1 0 35420 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1679235063
transform 1 0 34040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1679235063
transform 1 0 47196 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1679235063
transform 1 0 44436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1679235063
transform 1 0 45356 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1679235063
transform 1 0 32660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1679235063
transform 1 0 49220 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1679235063
transform 1 0 39836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1679235063
transform 1 0 29624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1679235063
transform 1 0 45724 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1679235063
transform 1 0 40020 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1679235063
transform 1 0 44620 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1679235063
transform 1 0 39376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1679235063
transform 1 0 40204 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1679235063
transform 1 0 40112 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1679235063
transform 1 0 41124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1679235063
transform 1 0 41952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1679235063
transform 1 0 42136 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1679235063
transform 1 0 43424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1679235063
transform 1 0 30728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1679235063
transform 1 0 36984 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1679235063
transform 1 0 32752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1679235063
transform 1 0 1656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1679235063
transform 1 0 32384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1679235063
transform 1 0 36892 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1679235063
transform 1 0 37812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1679235063
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1679235063
transform 1 0 25944 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1679235063
transform 1 0 28612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1679235063
transform 1 0 31280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1679235063
transform 1 0 33948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1679235063
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1679235063
transform 1 0 47012 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1679235063
transform 1 0 48300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1679235063
transform 1 0 46644 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1679235063
transform 1 0 46828 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1679235063
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1679235063
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1679235063
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1679235063
transform 1 0 46460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1679235063
transform 1 0 45540 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output77_A
timestamp 1679235063
transform 1 0 47748 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output79_A
timestamp 1679235063
transform 1 0 1472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1679235063
transform 1 0 14260 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output87_A
timestamp 1679235063
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1679235063
transform 1 0 27784 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1679235063
transform 1 0 9016 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1679235063
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output91_A
timestamp 1679235063
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1679235063
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1679235063
transform 1 0 34408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1679235063
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1679235063
transform 1 0 23368 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1679235063
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output114_A
timestamp 1679235063
transform 1 0 3496 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output115_A
timestamp 1679235063
transform 1 0 27600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output116_A
timestamp 1679235063
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output117_A
timestamp 1679235063
transform 1 0 13708 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1679235063
transform 1 0 14260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1679235063
transform 1 0 11500 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1679235063
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1679235063
transform 1 0 16284 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1679235063
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1679235063
transform 1 0 8648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1679235063
transform 1 0 5704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output126_A
timestamp 1679235063
transform 1 0 3496 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output131_A
timestamp 1679235063
transform 1 0 16744 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output133_A
timestamp 1679235063
transform 1 0 29072 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output134_A
timestamp 1679235063
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output135_A
timestamp 1679235063
transform 1 0 9568 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output136_A
timestamp 1679235063
transform 1 0 34316 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output137_A
timestamp 1679235063
transform 1 0 14076 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output138_A
timestamp 1679235063
transform 1 0 34316 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23092 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 14996 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 19136 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 14352 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 13616 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 11868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 14536 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 14168 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 34316 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 24012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 24104 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29072 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 29256 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 30452 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 31924 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 34500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31832 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 29072 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31648 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__CLK
timestamp 1679235063
transform 1 0 28980 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 31648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 31464 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 29072 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26496 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__CLK
timestamp 1679235063
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 43148 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 26956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 24472 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 23000 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1__RESET_B
timestamp 1679235063
transform 1 0 26496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2__RESET_B
timestamp 1679235063
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0__RESET_B
timestamp 1679235063
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 20516 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 3312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1__D
timestamp 1679235063
transform 1 0 9844 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0__D
timestamp 1679235063
transform 1 0 11592 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_1.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 12328 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 9108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26496 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 22264 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_5.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13616 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_7.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 23368 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11408 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 10856 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11500 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 27692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26956 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21804 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34316 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 31740 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 8924 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 8280 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 27968 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26588 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 20976 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_15.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_17.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 14168 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_19.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26312 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 11592 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29256 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 28888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_31.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 21344 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_33.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31648 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34316 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 22448 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 34316 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 31832 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 17296 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 31924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 31740 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 32292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_0.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 20148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 27416 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 27600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26680 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 3312 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23920 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 22264 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 23736 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 21896 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 23000 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23184 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16100 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_6.mux_l2_in_1__S
timestamp 1679235063
transform 1 0 16652 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 25760 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 26220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_8.mux_l2_in_1__A1
timestamp 1679235063
transform 1 0 16560 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 24288 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 24472 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 24840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_10.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 24656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 20608 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_12.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_14.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19228 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_16.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 21712 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 23000 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16836 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_20.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14168 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_22.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_24.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_26.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_28.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11592 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 11592 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 41860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 39928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 43056 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 10856 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 10856 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3312 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 22448 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 3864 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 12144 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 11684 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 1472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__A0
timestamp 1679235063
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 14168 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 15640 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 10488 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 35788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.mux_l2_in_0__S
timestamp 1679235063
transform 1 0 5796 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 19320 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A0
timestamp 1679235063
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 11408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 11592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 42320 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A0
timestamp 1679235063
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__A1
timestamp 1679235063
transform 1 0 20424 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_0__S
timestamp 1679235063
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__A1
timestamp 1679235063
transform 1 0 13984 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.mux_l1_in_1__S
timestamp 1679235063
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0__A
timestamp 1679235063
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9292 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 8464 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 3956 0 -1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4140 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4784 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 5428 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 5796 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 6808 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 7176 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7636 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 4968 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 4784 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.cbx_8__0_.mem_top_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1679235063
transform 1 0 4232 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10028 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_2_
timestamp 1679235063
transform 1 0 8740 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l1_in_4_
timestamp 1679235063
transform 1 0 12144 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7820 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3_
timestamp 1679235063
transform 1 0 10396 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l2_in_3__192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 9108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 9476 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9844 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.mux_l4_in_0_
timestamp 1679235063
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 3404 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 2944 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_2_
timestamp 1679235063
transform 1 0 10396 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_3_
timestamp 1679235063
transform 1 0 9200 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 4048 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_2_
timestamp 1679235063
transform 1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3_
timestamp 1679235063
transform 1 0 4416 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l2_in_3__193
timestamp 1679235063
transform 1 0 28244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_0_
timestamp 1679235063
transform 1 0 4600 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l3_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.mux_l4_in_0_
timestamp 1679235063
transform 1 0 6532 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_2_
timestamp 1679235063
transform 1 0 6624 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7544 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_2_
timestamp 1679235063
transform 1 0 9384 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3_
timestamp 1679235063
transform 1 0 14260 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l2_in_3__194
timestamp 1679235063
transform 1 0 6532 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 5612 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l3_in_1_
timestamp 1679235063
transform 1 0 10304 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 8832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_1_
timestamp 1679235063
transform 1 0 1564 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_2_
timestamp 1679235063
transform 1 0 7636 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_3_
timestamp 1679235063
transform 1 0 7544 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l1_in_4_
timestamp 1679235063
transform 1 0 10396 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_1_
timestamp 1679235063
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_2_
timestamp 1679235063
transform 1 0 8096 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3_
timestamp 1679235063
transform 1 0 12696 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l2_in_3__195
timestamp 1679235063
transform 1 0 16836 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_0_
timestamp 1679235063
transform 1 0 10488 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l3_in_1_
timestamp 1679235063
transform 1 0 9108 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.mux_l4_in_0_
timestamp 1679235063
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 20424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 29440 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 18492 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 8832 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 27140 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22908 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 20884 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 16836 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 25668 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22172 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 22816 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 15640 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1679235063
transform 1 0 24748 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1679235063
transform 1 0 22632 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1679235063
transform 1 0 27140 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1679235063
transform 1 0 14260 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 17204 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 10212 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1679235063
transform 1 0 9384 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1679235063
transform 1 0 14904 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1679235063
transform 1 0 14720 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1679235063
transform 1 0 9108 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1679235063
transform 1 0 8924 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1679235063
transform 1 0 13432 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1679235063
transform 1 0 12788 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1679235063
transform 1 0 19412 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1679235063
transform 1 0 25116 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1679235063
transform 1 0 22540 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1679235063
transform 1 0 19596 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1679235063
transform 1 0 21988 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1679235063
transform 1 0 24932 0 -1 19584
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1679235063
transform 1 0 25300 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout143
timestamp 1679235063
transform 1 0 10212 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout144
timestamp 1679235063
transform 1 0 22448 0 1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout145
timestamp 1679235063
transform 1 0 10212 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout146
timestamp 1679235063
transform 1 0 6072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout147 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout148
timestamp 1679235063
transform 1 0 21988 0 -1 21760
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  fanout149 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20976 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout150
timestamp 1679235063
transform 1 0 30820 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout151
timestamp 1679235063
transform 1 0 29808 0 1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  fanout152
timestamp 1679235063
transform 1 0 40020 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1679235063
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1679235063
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1679235063
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31
timestamp 1679235063
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1679235063
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 6532 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_78
timestamp 1679235063
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_89
timestamp 1679235063
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_107
timestamp 1679235063
transform 1 0 10948 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1679235063
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_115 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1679235063
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_136
timestamp 1679235063
transform 1 0 13616 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 1679235063
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1679235063
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_152
timestamp 1679235063
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1679235063
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 1679235063
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1679235063
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_182
timestamp 1679235063
transform 1 0 17848 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_189
timestamp 1679235063
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1679235063
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_202
timestamp 1679235063
transform 1 0 19688 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1679235063
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_216 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 20976 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1679235063
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_230
timestamp 1679235063
transform 1 0 22264 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_234 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 22632 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1679235063
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_268
timestamp 1679235063
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1679235063
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1679235063
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_293
timestamp 1679235063
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_297
timestamp 1679235063
transform 1 0 28428 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_301
timestamp 1679235063
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1679235063
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1679235063
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_321
timestamp 1679235063
transform 1 0 30636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_326
timestamp 1679235063
transform 1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_330
timestamp 1679235063
transform 1 0 31464 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1679235063
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_349
timestamp 1679235063
transform 1 0 33212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_355
timestamp 1679235063
transform 1 0 33764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_359
timestamp 1679235063
transform 1 0 34132 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1679235063
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1679235063
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_377
timestamp 1679235063
transform 1 0 35788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_390
timestamp 1679235063
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_395
timestamp 1679235063
transform 1 0 37444 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_407
timestamp 1679235063
transform 1 0 38548 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1679235063
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_421
timestamp 1679235063
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_433
timestamp 1679235063
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1679235063
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_449
timestamp 1679235063
transform 1 0 42412 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_461
timestamp 1679235063
transform 1 0 43516 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_473
timestamp 1679235063
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_477
timestamp 1679235063
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_489
timestamp 1679235063
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_501
timestamp 1679235063
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_505
timestamp 1679235063
transform 1 0 47564 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_517
timestamp 1679235063
transform 1 0 48668 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_525
timestamp 1679235063
transform 1 0 49404 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1679235063
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1679235063
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_22
timestamp 1679235063
transform 1 0 3128 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1679235063
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_46
timestamp 1679235063
transform 1 0 5336 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_50
timestamp 1679235063
transform 1 0 5704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1679235063
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1679235063
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_67
timestamp 1679235063
transform 1 0 7268 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_71
timestamp 1679235063
transform 1 0 7636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_80
timestamp 1679235063
transform 1 0 8464 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_104
timestamp 1679235063
transform 1 0 10672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_108
timestamp 1679235063
transform 1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_113
timestamp 1679235063
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1679235063
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_127
timestamp 1679235063
transform 1 0 12788 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1679235063
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1679235063
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_144
timestamp 1679235063
transform 1 0 14352 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_152
timestamp 1679235063
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157
timestamp 1679235063
transform 1 0 15548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_163
timestamp 1679235063
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1679235063
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_182
timestamp 1679235063
transform 1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_186
timestamp 1679235063
transform 1 0 18216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_210
timestamp 1679235063
transform 1 0 20424 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1679235063
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1679235063
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1679235063
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_230
timestamp 1679235063
transform 1 0 22264 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_234
timestamp 1679235063
transform 1 0 22632 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_246
timestamp 1679235063
transform 1 0 23736 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_258
timestamp 1679235063
transform 1 0 24840 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_270
timestamp 1679235063
transform 1 0 25944 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_278
timestamp 1679235063
transform 1 0 26680 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1679235063
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1679235063
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1679235063
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1679235063
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1679235063
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1679235063
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1679235063
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1679235063
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1679235063
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1679235063
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1679235063
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1679235063
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1679235063
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_405
timestamp 1679235063
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_417
timestamp 1679235063
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_429
timestamp 1679235063
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_441
timestamp 1679235063
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1679235063
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_449
timestamp 1679235063
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_461
timestamp 1679235063
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_473
timestamp 1679235063
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_485
timestamp 1679235063
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1679235063
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1679235063
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_505
timestamp 1679235063
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_517
timestamp 1679235063
transform 1 0 48668 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1679235063
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 1679235063
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_14
timestamp 1679235063
transform 1 0 2392 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1679235063
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1679235063
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_34
timestamp 1679235063
transform 1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_46
timestamp 1679235063
transform 1 0 5336 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_60
timestamp 1679235063
transform 1 0 6624 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_67
timestamp 1679235063
transform 1 0 7268 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_74
timestamp 1679235063
transform 1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1679235063
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_89
timestamp 1679235063
transform 1 0 9292 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_99
timestamp 1679235063
transform 1 0 10212 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_111
timestamp 1679235063
transform 1 0 11316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_118
timestamp 1679235063
transform 1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1679235063
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1679235063
transform 1 0 13432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1679235063
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1679235063
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_147
timestamp 1679235063
transform 1 0 14628 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_155
timestamp 1679235063
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_163
timestamp 1679235063
transform 1 0 16100 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_175
timestamp 1679235063
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_2_189
timestamp 1679235063
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1679235063
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_202
timestamp 1679235063
transform 1 0 19688 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_209
timestamp 1679235063
transform 1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_216
timestamp 1679235063
transform 1 0 20976 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_228
timestamp 1679235063
transform 1 0 22080 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_240
timestamp 1679235063
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1679235063
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1679235063
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1679235063
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1679235063
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1679235063
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1679235063
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1679235063
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1679235063
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1679235063
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1679235063
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1679235063
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1679235063
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1679235063
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1679235063
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1679235063
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_401
timestamp 1679235063
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_413
timestamp 1679235063
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1679235063
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_421
timestamp 1679235063
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_433
timestamp 1679235063
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1679235063
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_457
timestamp 1679235063
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_469
timestamp 1679235063
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1679235063
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_477
timestamp 1679235063
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_489
timestamp 1679235063
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_501
timestamp 1679235063
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_513
timestamp 1679235063
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1679235063
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_3
timestamp 1679235063
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1679235063
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_27
timestamp 1679235063
transform 1 0 3588 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_39
timestamp 1679235063
transform 1 0 4692 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_47
timestamp 1679235063
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1679235063
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1679235063
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_67
timestamp 1679235063
transform 1 0 7268 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_74
timestamp 1679235063
transform 1 0 7912 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_82
timestamp 1679235063
transform 1 0 8648 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 1679235063
transform 1 0 9384 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_100
timestamp 1679235063
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_104
timestamp 1679235063
transform 1 0 10672 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1679235063
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_113
timestamp 1679235063
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_123
timestamp 1679235063
transform 1 0 12420 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_127
timestamp 1679235063
transform 1 0 12788 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1679235063
transform 1 0 13156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_143
timestamp 1679235063
transform 1 0 14260 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_155
timestamp 1679235063
transform 1 0 15364 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1679235063
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1679235063
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_169
timestamp 1679235063
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_192
timestamp 1679235063
transform 1 0 18768 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1679235063
transform 1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_206
timestamp 1679235063
transform 1 0 20056 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1679235063
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_220
timestamp 1679235063
transform 1 0 21344 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_227
timestamp 1679235063
transform 1 0 21988 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_239
timestamp 1679235063
transform 1 0 23092 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_251
timestamp 1679235063
transform 1 0 24196 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_263
timestamp 1679235063
transform 1 0 25300 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_275
timestamp 1679235063
transform 1 0 26404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1679235063
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1679235063
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1679235063
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1679235063
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1679235063
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1679235063
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1679235063
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1679235063
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1679235063
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1679235063
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1679235063
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1679235063
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1679235063
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1679235063
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_405
timestamp 1679235063
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_417
timestamp 1679235063
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1679235063
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1679235063
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1679235063
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1679235063
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_461
timestamp 1679235063
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_473
timestamp 1679235063
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_485
timestamp 1679235063
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_497
timestamp 1679235063
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1679235063
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1679235063
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_517
timestamp 1679235063
transform 1 0 48668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_525
timestamp 1679235063
transform 1 0 49404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_3
timestamp 1679235063
transform 1 0 1380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1679235063
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 1679235063
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1679235063
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1679235063
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_39
timestamp 1679235063
transform 1 0 4692 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_47
timestamp 1679235063
transform 1 0 5428 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_55
timestamp 1679235063
transform 1 0 6164 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1679235063
transform 1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_70
timestamp 1679235063
transform 1 0 7544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1679235063
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1679235063
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_97
timestamp 1679235063
transform 1 0 10028 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_101
timestamp 1679235063
transform 1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 1679235063
transform 1 0 11592 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_120
timestamp 1679235063
transform 1 0 12144 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_131
timestamp 1679235063
transform 1 0 13156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1679235063
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1679235063
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_4_151
timestamp 1679235063
transform 1 0 14996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_157
timestamp 1679235063
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_179
timestamp 1679235063
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_191
timestamp 1679235063
transform 1 0 18676 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1679235063
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1679235063
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1679235063
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_222
timestamp 1679235063
transform 1 0 21528 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_229
timestamp 1679235063
transform 1 0 22172 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_233
timestamp 1679235063
transform 1 0 22540 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_240
timestamp 1679235063
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 1679235063
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_258
timestamp 1679235063
transform 1 0 24840 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_266
timestamp 1679235063
transform 1 0 25576 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_288
timestamp 1679235063
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1679235063
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1679235063
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1679235063
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1679235063
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1679235063
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1679235063
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1679235063
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1679235063
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1679235063
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1679235063
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1679235063
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1679235063
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1679235063
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1679235063
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1679235063
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1679235063
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1679235063
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1679235063
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1679235063
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1679235063
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1679235063
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_501
timestamp 1679235063
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_513
timestamp 1679235063
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1679235063
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1679235063
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_14
timestamp 1679235063
transform 1 0 2392 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1679235063
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1679235063
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1679235063
transform 1 0 5336 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1679235063
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1679235063
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_62
timestamp 1679235063
transform 1 0 6808 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_74
timestamp 1679235063
transform 1 0 7912 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_86
timestamp 1679235063
transform 1 0 9016 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_98
timestamp 1679235063
transform 1 0 10120 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1679235063
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_117
timestamp 1679235063
transform 1 0 11868 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_128
timestamp 1679235063
transform 1 0 12880 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_132
timestamp 1679235063
transform 1 0 13248 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_141
timestamp 1679235063
transform 1 0 14076 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_145
timestamp 1679235063
transform 1 0 14444 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1679235063
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1679235063
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1679235063
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_179
timestamp 1679235063
transform 1 0 17572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_183
timestamp 1679235063
transform 1 0 17940 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_186
timestamp 1679235063
transform 1 0 18216 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_198
timestamp 1679235063
transform 1 0 19320 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_212
timestamp 1679235063
transform 1 0 20608 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_220
timestamp 1679235063
transform 1 0 21344 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_227
timestamp 1679235063
transform 1 0 21988 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_232
timestamp 1679235063
transform 1 0 22448 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_239
timestamp 1679235063
transform 1 0 23092 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_251
timestamp 1679235063
transform 1 0 24196 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_5_278
timestamp 1679235063
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_281
timestamp 1679235063
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_304
timestamp 1679235063
transform 1 0 29072 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1679235063
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1679235063
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1679235063
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1679235063
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1679235063
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1679235063
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1679235063
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1679235063
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1679235063
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1679235063
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1679235063
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1679235063
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1679235063
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1679235063
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1679235063
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1679235063
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1679235063
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1679235063
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1679235063
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1679235063
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1679235063
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_517
timestamp 1679235063
transform 1 0 48668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1679235063
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1679235063
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1679235063
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_19
timestamp 1679235063
transform 1 0 2852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1679235063
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_31
timestamp 1679235063
transform 1 0 3956 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1679235063
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_48
timestamp 1679235063
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_58
timestamp 1679235063
transform 1 0 6440 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_70
timestamp 1679235063
transform 1 0 7544 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1679235063
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_85
timestamp 1679235063
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_90
timestamp 1679235063
transform 1 0 9384 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_102
timestamp 1679235063
transform 1 0 10488 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_114
timestamp 1679235063
transform 1 0 11592 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_126
timestamp 1679235063
transform 1 0 12696 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1679235063
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1679235063
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_164
timestamp 1679235063
transform 1 0 16192 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_168
timestamp 1679235063
transform 1 0 16560 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1679235063
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_209
timestamp 1679235063
transform 1 0 20332 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_216
timestamp 1679235063
transform 1 0 20976 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_230
timestamp 1679235063
transform 1 0 22264 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1679235063
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_244
timestamp 1679235063
transform 1 0 23552 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1679235063
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1679235063
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1679235063
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1679235063
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1679235063
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1679235063
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1679235063
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1679235063
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1679235063
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1679235063
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1679235063
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1679235063
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1679235063
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1679235063
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1679235063
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1679235063
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1679235063
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1679235063
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1679235063
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1679235063
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1679235063
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1679235063
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1679235063
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1679235063
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1679235063
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1679235063
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1679235063
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_501
timestamp 1679235063
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_513
timestamp 1679235063
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1679235063
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1679235063
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_15
timestamp 1679235063
transform 1 0 2484 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_22
timestamp 1679235063
transform 1 0 3128 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_30
timestamp 1679235063
transform 1 0 3864 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_42
timestamp 1679235063
transform 1 0 4968 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1679235063
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_62
timestamp 1679235063
transform 1 0 6808 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1679235063
transform 1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_86
timestamp 1679235063
transform 1 0 9016 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_98
timestamp 1679235063
transform 1 0 10120 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1679235063
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1679235063
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_116
timestamp 1679235063
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_126
timestamp 1679235063
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_132
timestamp 1679235063
transform 1 0 13248 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_142
timestamp 1679235063
transform 1 0 14168 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_154
timestamp 1679235063
transform 1 0 15272 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1679235063
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_169
timestamp 1679235063
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_179
timestamp 1679235063
transform 1 0 17572 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_191
timestamp 1679235063
transform 1 0 18676 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_203
timestamp 1679235063
transform 1 0 19780 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_215
timestamp 1679235063
transform 1 0 20884 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_222
timestamp 1679235063
transform 1 0 21528 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_225
timestamp 1679235063
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_230
timestamp 1679235063
transform 1 0 22264 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 1679235063
transform 1 0 22632 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_243
timestamp 1679235063
transform 1 0 23460 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_247
timestamp 1679235063
transform 1 0 23828 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_259
timestamp 1679235063
transform 1 0 24932 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_271
timestamp 1679235063
transform 1 0 26036 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1679235063
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1679235063
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1679235063
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1679235063
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1679235063
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1679235063
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1679235063
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1679235063
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1679235063
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1679235063
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1679235063
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1679235063
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1679235063
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1679235063
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1679235063
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1679235063
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1679235063
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1679235063
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1679235063
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1679235063
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1679235063
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1679235063
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1679235063
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1679235063
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1679235063
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1679235063
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1679235063
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1679235063
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1679235063
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_9
timestamp 1679235063
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_13
timestamp 1679235063
transform 1 0 2300 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_18
timestamp 1679235063
transform 1 0 2760 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1679235063
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1679235063
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_46
timestamp 1679235063
transform 1 0 5336 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_58
timestamp 1679235063
transform 1 0 6440 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_70
timestamp 1679235063
transform 1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1679235063
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 1679235063
transform 1 0 9384 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_96
timestamp 1679235063
transform 1 0 9936 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_107
timestamp 1679235063
transform 1 0 10948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_114
timestamp 1679235063
transform 1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_126
timestamp 1679235063
transform 1 0 12696 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1679235063
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_141
timestamp 1679235063
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_145
timestamp 1679235063
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_149
timestamp 1679235063
transform 1 0 14812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1679235063
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp 1679235063
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_178
timestamp 1679235063
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1679235063
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1679235063
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_208
timestamp 1679235063
transform 1 0 20240 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_220
timestamp 1679235063
transform 1 0 21344 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_224
timestamp 1679235063
transform 1 0 21712 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_233
timestamp 1679235063
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_241
timestamp 1679235063
transform 1 0 23276 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_8_249
timestamp 1679235063
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1679235063
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1679235063
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1679235063
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1679235063
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1679235063
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1679235063
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1679235063
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1679235063
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1679235063
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1679235063
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1679235063
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1679235063
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1679235063
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1679235063
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1679235063
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_401
timestamp 1679235063
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1679235063
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1679235063
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1679235063
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1679235063
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1679235063
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1679235063
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1679235063
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1679235063
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1679235063
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1679235063
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_501
timestamp 1679235063
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_513
timestamp 1679235063
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1679235063
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1679235063
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_6
timestamp 1679235063
transform 1 0 1656 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_16
timestamp 1679235063
transform 1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_28
timestamp 1679235063
transform 1 0 3680 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_40
timestamp 1679235063
transform 1 0 4784 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_44
timestamp 1679235063
transform 1 0 5152 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1679235063
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1679235063
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1679235063
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_81
timestamp 1679235063
transform 1 0 8556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_93
timestamp 1679235063
transform 1 0 9660 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1679235063
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1679235063
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1679235063
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_141
timestamp 1679235063
transform 1 0 14076 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_145
timestamp 1679235063
transform 1 0 14444 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_154
timestamp 1679235063
transform 1 0 15272 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1679235063
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_169
timestamp 1679235063
transform 1 0 16652 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_174
timestamp 1679235063
transform 1 0 17112 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_178
timestamp 1679235063
transform 1 0 17480 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_188
timestamp 1679235063
transform 1 0 18400 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_195
timestamp 1679235063
transform 1 0 19044 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_207
timestamp 1679235063
transform 1 0 20148 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_219
timestamp 1679235063
transform 1 0 21252 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1679235063
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 1679235063
transform 1 0 21804 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_247
timestamp 1679235063
transform 1 0 23828 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_255
timestamp 1679235063
transform 1 0 24564 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_259
timestamp 1679235063
transform 1 0 24932 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_271
timestamp 1679235063
transform 1 0 26036 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1679235063
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1679235063
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1679235063
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1679235063
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1679235063
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1679235063
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1679235063
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1679235063
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1679235063
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1679235063
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1679235063
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1679235063
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1679235063
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1679235063
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1679235063
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1679235063
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1679235063
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1679235063
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1679235063
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1679235063
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1679235063
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1679235063
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1679235063
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1679235063
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1679235063
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_505
timestamp 1679235063
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_517
timestamp 1679235063
transform 1 0 48668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1679235063
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1679235063
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_14
timestamp 1679235063
transform 1 0 2392 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1679235063
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 1679235063
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_40
timestamp 1679235063
transform 1 0 4784 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_52
timestamp 1679235063
transform 1 0 5888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_57
timestamp 1679235063
transform 1 0 6348 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_67
timestamp 1679235063
transform 1 0 7268 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_71
timestamp 1679235063
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1679235063
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_85
timestamp 1679235063
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_91
timestamp 1679235063
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_104
timestamp 1679235063
transform 1 0 10672 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1679235063
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_114
timestamp 1679235063
transform 1 0 11592 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_126
timestamp 1679235063
transform 1 0 12696 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1679235063
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1679235063
transform 1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_150
timestamp 1679235063
transform 1 0 14904 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1679235063
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_174
timestamp 1679235063
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1679235063
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1679235063
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1679235063
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_10_209
timestamp 1679235063
transform 1 0 20332 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1679235063
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_235
timestamp 1679235063
transform 1 0 22724 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_247
timestamp 1679235063
transform 1 0 23828 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1679235063
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 1679235063
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_259
timestamp 1679235063
transform 1 0 24932 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_263
timestamp 1679235063
transform 1 0 25300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_275
timestamp 1679235063
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_287
timestamp 1679235063
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_299
timestamp 1679235063
transform 1 0 28612 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1679235063
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1679235063
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1679235063
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1679235063
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1679235063
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1679235063
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1679235063
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1679235063
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1679235063
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1679235063
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1679235063
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1679235063
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1679235063
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1679235063
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1679235063
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1679235063
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1679235063
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1679235063
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1679235063
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1679235063
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1679235063
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_501
timestamp 1679235063
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_513
timestamp 1679235063
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1679235063
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1679235063
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_8
timestamp 1679235063
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_18
timestamp 1679235063
transform 1 0 2760 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1679235063
transform 1 0 3864 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_42
timestamp 1679235063
transform 1 0 4968 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1679235063
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 1679235063
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_67
timestamp 1679235063
transform 1 0 7268 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_79
timestamp 1679235063
transform 1 0 8372 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1679235063
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1679235063
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1679235063
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_115
timestamp 1679235063
transform 1 0 11684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1679235063
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1679235063
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_154
timestamp 1679235063
transform 1 0 15272 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1679235063
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_171
timestamp 1679235063
transform 1 0 16836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_185
timestamp 1679235063
transform 1 0 18124 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1679235063
transform 1 0 19596 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_213
timestamp 1679235063
transform 1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_220
timestamp 1679235063
transform 1 0 21344 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_225
timestamp 1679235063
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_235
timestamp 1679235063
transform 1 0 22724 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_247
timestamp 1679235063
transform 1 0 23828 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_253
timestamp 1679235063
transform 1 0 24380 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_259
timestamp 1679235063
transform 1 0 24932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_267
timestamp 1679235063
transform 1 0 25668 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_274
timestamp 1679235063
transform 1 0 26312 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1679235063
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1679235063
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1679235063
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1679235063
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1679235063
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1679235063
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1679235063
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1679235063
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1679235063
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1679235063
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1679235063
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1679235063
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1679235063
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1679235063
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1679235063
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1679235063
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1679235063
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1679235063
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1679235063
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1679235063
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_473
timestamp 1679235063
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_485
timestamp 1679235063
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1679235063
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1679235063
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_505
timestamp 1679235063
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_517
timestamp 1679235063
transform 1 0 48668 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1679235063
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_3
timestamp 1679235063
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_14
timestamp 1679235063
transform 1 0 2392 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1679235063
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_31
timestamp 1679235063
transform 1 0 3956 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_42
timestamp 1679235063
transform 1 0 4968 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_47
timestamp 1679235063
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1679235063
transform 1 0 6348 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_69
timestamp 1679235063
transform 1 0 7452 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_73
timestamp 1679235063
transform 1 0 7820 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1679235063
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1679235063
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_95
timestamp 1679235063
transform 1 0 9844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1679235063
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_123
timestamp 1679235063
transform 1 0 12420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_127
timestamp 1679235063
transform 1 0 12788 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1679235063
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_141
timestamp 1679235063
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_152
timestamp 1679235063
transform 1 0 15088 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_156
timestamp 1679235063
transform 1 0 15456 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_166
timestamp 1679235063
transform 1 0 16376 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_172
timestamp 1679235063
transform 1 0 16928 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_182
timestamp 1679235063
transform 1 0 17848 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1679235063
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1679235063
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_207
timestamp 1679235063
transform 1 0 20148 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_223
timestamp 1679235063
transform 1 0 21620 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_235
timestamp 1679235063
transform 1 0 22724 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_247
timestamp 1679235063
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1679235063
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 1679235063
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_263
timestamp 1679235063
transform 1 0 25300 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_275
timestamp 1679235063
transform 1 0 26404 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_290
timestamp 1679235063
transform 1 0 27784 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_296
timestamp 1679235063
transform 1 0 28336 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1679235063
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1679235063
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1679235063
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1679235063
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1679235063
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1679235063
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1679235063
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1679235063
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1679235063
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1679235063
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1679235063
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1679235063
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1679235063
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1679235063
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1679235063
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1679235063
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1679235063
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1679235063
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_477
timestamp 1679235063
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_489
timestamp 1679235063
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_501
timestamp 1679235063
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_513
timestamp 1679235063
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_525
timestamp 1679235063
transform 1 0 49404 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1679235063
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1679235063
transform 1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_18
timestamp 1679235063
transform 1 0 2760 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_30
timestamp 1679235063
transform 1 0 3864 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_42
timestamp 1679235063
transform 1 0 4968 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1679235063
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1679235063
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_62
timestamp 1679235063
transform 1 0 6808 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1679235063
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_79
timestamp 1679235063
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_100
timestamp 1679235063
transform 1 0 10304 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_108
timestamp 1679235063
transform 1 0 11040 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1679235063
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_135
timestamp 1679235063
transform 1 0 13524 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_143
timestamp 1679235063
transform 1 0 14260 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1679235063
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1679235063
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_191
timestamp 1679235063
transform 1 0 18676 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_208
timestamp 1679235063
transform 1 0 20240 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_220
timestamp 1679235063
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 1679235063
transform 1 0 21804 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_235
timestamp 1679235063
transform 1 0 22724 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_239
timestamp 1679235063
transform 1 0 23092 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_248
timestamp 1679235063
transform 1 0 23920 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_254
timestamp 1679235063
transform 1 0 24472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_263
timestamp 1679235063
transform 1 0 25300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_275
timestamp 1679235063
transform 1 0 26404 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1679235063
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_281
timestamp 1679235063
transform 1 0 26956 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_291
timestamp 1679235063
transform 1 0 27876 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_303
timestamp 1679235063
transform 1 0 28980 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_315
timestamp 1679235063
transform 1 0 30084 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_327
timestamp 1679235063
transform 1 0 31188 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1679235063
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1679235063
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1679235063
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1679235063
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1679235063
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1679235063
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1679235063
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1679235063
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1679235063
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1679235063
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1679235063
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1679235063
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1679235063
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1679235063
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1679235063
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1679235063
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_485
timestamp 1679235063
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1679235063
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1679235063
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_505
timestamp 1679235063
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_517
timestamp 1679235063
transform 1 0 48668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1679235063
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 1679235063
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1679235063
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1679235063
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_29
timestamp 1679235063
transform 1 0 3772 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 1679235063
transform 1 0 4048 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1679235063
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1679235063
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_55
timestamp 1679235063
transform 1 0 6164 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1679235063
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_71
timestamp 1679235063
transform 1 0 7636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1679235063
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_85
timestamp 1679235063
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1679235063
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1679235063
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_133
timestamp 1679235063
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1679235063
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_143
timestamp 1679235063
transform 1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1679235063
transform 1 0 16284 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1679235063
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_193
timestamp 1679235063
transform 1 0 18860 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1679235063
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_220
timestamp 1679235063
transform 1 0 21344 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_14_236
timestamp 1679235063
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1679235063
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_253
timestamp 1679235063
transform 1 0 24380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_260
timestamp 1679235063
transform 1 0 25024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_272
timestamp 1679235063
transform 1 0 26128 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_276
timestamp 1679235063
transform 1 0 26496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_279
timestamp 1679235063
transform 1 0 26772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_291
timestamp 1679235063
transform 1 0 27876 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_298
timestamp 1679235063
transform 1 0 28520 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_306
timestamp 1679235063
transform 1 0 29256 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1679235063
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1679235063
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1679235063
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1679235063
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1679235063
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1679235063
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1679235063
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1679235063
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1679235063
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1679235063
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1679235063
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1679235063
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1679235063
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1679235063
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1679235063
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1679235063
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1679235063
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1679235063
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1679235063
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1679235063
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_501
timestamp 1679235063
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_513
timestamp 1679235063
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1679235063
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_7
timestamp 1679235063
transform 1 0 1748 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_17
timestamp 1679235063
transform 1 0 2668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_29
timestamp 1679235063
transform 1 0 3772 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_41
timestamp 1679235063
transform 1 0 4876 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_45
timestamp 1679235063
transform 1 0 5244 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1679235063
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1679235063
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_68
timestamp 1679235063
transform 1 0 7360 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_95
timestamp 1679235063
transform 1 0 9844 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1679235063
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_119
timestamp 1679235063
transform 1 0 12052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_141
timestamp 1679235063
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_147
timestamp 1679235063
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_161
timestamp 1679235063
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1679235063
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1679235063
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_174
timestamp 1679235063
transform 1 0 17112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_198
timestamp 1679235063
transform 1 0 19320 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 1679235063
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_225
timestamp 1679235063
transform 1 0 21804 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_236
timestamp 1679235063
transform 1 0 22816 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_240
timestamp 1679235063
transform 1 0 23184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_251
timestamp 1679235063
transform 1 0 24196 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_263
timestamp 1679235063
transform 1 0 25300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_275
timestamp 1679235063
transform 1 0 26404 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1679235063
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_281
timestamp 1679235063
transform 1 0 26956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_287
timestamp 1679235063
transform 1 0 27508 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_291
timestamp 1679235063
transform 1 0 27876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_299
timestamp 1679235063
transform 1 0 28612 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_309
timestamp 1679235063
transform 1 0 29532 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_321
timestamp 1679235063
transform 1 0 30636 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1679235063
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1679235063
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1679235063
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1679235063
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1679235063
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1679235063
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1679235063
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1679235063
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1679235063
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1679235063
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1679235063
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1679235063
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1679235063
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1679235063
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1679235063
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1679235063
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1679235063
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1679235063
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1679235063
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_505
timestamp 1679235063
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_517
timestamp 1679235063
transform 1 0 48668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1679235063
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1679235063
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_14
timestamp 1679235063
transform 1 0 2392 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1679235063
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_29
timestamp 1679235063
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_35
timestamp 1679235063
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_39
timestamp 1679235063
transform 1 0 4692 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_60
timestamp 1679235063
transform 1 0 6624 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1679235063
transform 1 0 7360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1679235063
transform 1 0 7728 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1679235063
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_89
timestamp 1679235063
transform 1 0 9292 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_100
timestamp 1679235063
transform 1 0 10304 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1679235063
transform 1 0 10672 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_109
timestamp 1679235063
transform 1 0 11132 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1679235063
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1679235063
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1679235063
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_167
timestamp 1679235063
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_171
timestamp 1679235063
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1679235063
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_197
timestamp 1679235063
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_210
timestamp 1679235063
transform 1 0 20424 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_214
timestamp 1679235063
transform 1 0 20792 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_236
timestamp 1679235063
transform 1 0 22816 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_249
timestamp 1679235063
transform 1 0 24012 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 1679235063
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_263
timestamp 1679235063
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_275
timestamp 1679235063
transform 1 0 26404 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_287
timestamp 1679235063
transform 1 0 27508 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_295
timestamp 1679235063
transform 1 0 28244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_303
timestamp 1679235063
transform 1 0 28980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1679235063
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_309
timestamp 1679235063
transform 1 0 29532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_334
timestamp 1679235063
transform 1 0 31832 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_338
timestamp 1679235063
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_350
timestamp 1679235063
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1679235063
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1679235063
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1679235063
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1679235063
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1679235063
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1679235063
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1679235063
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1679235063
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1679235063
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1679235063
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1679235063
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1679235063
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1679235063
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1679235063
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_489
timestamp 1679235063
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_501
timestamp 1679235063
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_513
timestamp 1679235063
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1679235063
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1679235063
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_17
timestamp 1679235063
transform 1 0 2668 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_29
timestamp 1679235063
transform 1 0 3772 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_41
timestamp 1679235063
transform 1 0 4876 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1679235063
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_62
timestamp 1679235063
transform 1 0 6808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_86
timestamp 1679235063
transform 1 0 9016 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_101
timestamp 1679235063
transform 1 0 10396 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1679235063
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1679235063
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1679235063
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1679235063
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_127
timestamp 1679235063
transform 1 0 12788 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1679235063
transform 1 0 14996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_155
timestamp 1679235063
transform 1 0 15364 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1679235063
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1679235063
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1679235063
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1679235063
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_206
timestamp 1679235063
transform 1 0 20056 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_220
timestamp 1679235063
transform 1 0 21344 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_229
timestamp 1679235063
transform 1 0 22172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_252
timestamp 1679235063
transform 1 0 24288 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_256
timestamp 1679235063
transform 1 0 24656 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_264
timestamp 1679235063
transform 1 0 25392 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_275
timestamp 1679235063
transform 1 0 26404 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1679235063
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_281
timestamp 1679235063
transform 1 0 26956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_291
timestamp 1679235063
transform 1 0 27876 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_298
timestamp 1679235063
transform 1 0 28520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_310
timestamp 1679235063
transform 1 0 29624 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_322
timestamp 1679235063
transform 1 0 30728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_334
timestamp 1679235063
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1679235063
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1679235063
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1679235063
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1679235063
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1679235063
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1679235063
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1679235063
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1679235063
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1679235063
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1679235063
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1679235063
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1679235063
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1679235063
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1679235063
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_473
timestamp 1679235063
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_485
timestamp 1679235063
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1679235063
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1679235063
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1679235063
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1679235063
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1679235063
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1679235063
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1679235063
transform 1 0 1840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_14
timestamp 1679235063
transform 1 0 2392 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1679235063
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_33
timestamp 1679235063
transform 1 0 4140 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_43
timestamp 1679235063
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_70
timestamp 1679235063
transform 1 0 7544 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1679235063
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1679235063
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1679235063
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_99
timestamp 1679235063
transform 1 0 10212 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_112
timestamp 1679235063
transform 1 0 11408 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_125
timestamp 1679235063
transform 1 0 12604 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1679235063
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_143
timestamp 1679235063
transform 1 0 14260 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_146
timestamp 1679235063
transform 1 0 14536 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_159
timestamp 1679235063
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_183
timestamp 1679235063
transform 1 0 17940 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1679235063
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1679235063
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1679235063
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_226
timestamp 1679235063
transform 1 0 21896 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_250
timestamp 1679235063
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_255
timestamp 1679235063
transform 1 0 24564 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_259
timestamp 1679235063
transform 1 0 24932 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_268
timestamp 1679235063
transform 1 0 25760 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_280
timestamp 1679235063
transform 1 0 26864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_291
timestamp 1679235063
transform 1 0 27876 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_299
timestamp 1679235063
transform 1 0 28612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_303
timestamp 1679235063
transform 1 0 28980 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1679235063
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1679235063
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1679235063
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1679235063
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1679235063
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1679235063
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1679235063
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1679235063
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1679235063
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1679235063
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1679235063
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1679235063
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1679235063
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1679235063
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1679235063
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1679235063
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_457
timestamp 1679235063
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1679235063
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1679235063
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1679235063
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1679235063
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_501
timestamp 1679235063
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_513
timestamp 1679235063
transform 1 0 48300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1679235063
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1679235063
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_15
timestamp 1679235063
transform 1 0 2484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_19
timestamp 1679235063
transform 1 0 2852 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_29
timestamp 1679235063
transform 1 0 3772 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1679235063
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_67
timestamp 1679235063
transform 1 0 7268 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_94
timestamp 1679235063
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_98
timestamp 1679235063
transform 1 0 10120 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1679235063
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1679235063
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_116
timestamp 1679235063
transform 1 0 11776 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_127
timestamp 1679235063
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_140
timestamp 1679235063
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_153
timestamp 1679235063
transform 1 0 15180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1679235063
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_173
timestamp 1679235063
transform 1 0 17020 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_184
timestamp 1679235063
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_198
timestamp 1679235063
transform 1 0 19320 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 1679235063
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1679235063
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_231
timestamp 1679235063
transform 1 0 22356 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_235
timestamp 1679235063
transform 1 0 22724 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_257
timestamp 1679235063
transform 1 0 24748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_272
timestamp 1679235063
transform 1 0 26128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_278
timestamp 1679235063
transform 1 0 26680 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1679235063
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_291
timestamp 1679235063
transform 1 0 27876 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_303
timestamp 1679235063
transform 1 0 28980 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_315
timestamp 1679235063
transform 1 0 30084 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_327
timestamp 1679235063
transform 1 0 31188 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1679235063
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1679235063
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1679235063
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1679235063
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1679235063
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1679235063
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1679235063
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1679235063
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1679235063
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1679235063
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1679235063
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1679235063
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1679235063
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1679235063
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_461
timestamp 1679235063
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_473
timestamp 1679235063
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_485
timestamp 1679235063
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1679235063
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1679235063
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_505
timestamp 1679235063
transform 1 0 47564 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_517
timestamp 1679235063
transform 1 0 48668 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1679235063
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1679235063
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_21
timestamp 1679235063
transform 1 0 3036 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1679235063
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_34
timestamp 1679235063
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_45
timestamp 1679235063
transform 1 0 5244 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_58
timestamp 1679235063
transform 1 0 6440 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1679235063
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1679235063
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1679235063
transform 1 0 9936 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1679235063
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1679235063
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1679235063
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1679235063
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_163
timestamp 1679235063
transform 1 0 16100 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_169
timestamp 1679235063
transform 1 0 16652 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_181
timestamp 1679235063
transform 1 0 17756 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1679235063
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_199
timestamp 1679235063
transform 1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_204
timestamp 1679235063
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_228
timestamp 1679235063
transform 1 0 22080 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_243
timestamp 1679235063
transform 1 0 23460 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 1679235063
transform 1 0 24104 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 1679235063
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_264
timestamp 1679235063
transform 1 0 25392 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_276
timestamp 1679235063
transform 1 0 26496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_280
timestamp 1679235063
transform 1 0 26864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_291
timestamp 1679235063
transform 1 0 27876 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_303
timestamp 1679235063
transform 1 0 28980 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1679235063
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_311
timestamp 1679235063
transform 1 0 29716 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_323
timestamp 1679235063
transform 1 0 30820 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_335
timestamp 1679235063
transform 1 0 31924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_347
timestamp 1679235063
transform 1 0 33028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_359
timestamp 1679235063
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1679235063
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1679235063
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1679235063
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1679235063
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_401
timestamp 1679235063
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1679235063
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1679235063
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_421
timestamp 1679235063
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_433
timestamp 1679235063
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_445
timestamp 1679235063
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_457
timestamp 1679235063
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1679235063
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1679235063
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1679235063
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1679235063
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_501
timestamp 1679235063
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_513
timestamp 1679235063
transform 1 0 48300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1679235063
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1679235063
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_21
timestamp 1679235063
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1679235063
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1679235063
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_61
timestamp 1679235063
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1679235063
transform 1 0 7728 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_85
timestamp 1679235063
transform 1 0 8924 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1679235063
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_115
timestamp 1679235063
transform 1 0 11684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1679235063
transform 1 0 11960 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1679235063
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_148
timestamp 1679235063
transform 1 0 14720 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_152
timestamp 1679235063
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1679235063
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_171
timestamp 1679235063
transform 1 0 16836 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_194
timestamp 1679235063
transform 1 0 18952 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_198
timestamp 1679235063
transform 1 0 19320 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_209
timestamp 1679235063
transform 1 0 20332 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_222
timestamp 1679235063
transform 1 0 21528 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 1679235063
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_232
timestamp 1679235063
transform 1 0 22448 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_243
timestamp 1679235063
transform 1 0 23460 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_256
timestamp 1679235063
transform 1 0 24656 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_260
timestamp 1679235063
transform 1 0 25024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_270
timestamp 1679235063
transform 1 0 25944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1679235063
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_281
timestamp 1679235063
transform 1 0 26956 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_291
timestamp 1679235063
transform 1 0 27876 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_297
timestamp 1679235063
transform 1 0 28428 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_306
timestamp 1679235063
transform 1 0 29256 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_313
timestamp 1679235063
transform 1 0 29900 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_320
timestamp 1679235063
transform 1 0 30544 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_324
timestamp 1679235063
transform 1 0 30912 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1679235063
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1679235063
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1679235063
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1679235063
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1679235063
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1679235063
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1679235063
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_405
timestamp 1679235063
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_417
timestamp 1679235063
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_429
timestamp 1679235063
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1679235063
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1679235063
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1679235063
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1679235063
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1679235063
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1679235063
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1679235063
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1679235063
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_505
timestamp 1679235063
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_517
timestamp 1679235063
transform 1 0 48668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1679235063
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_3
timestamp 1679235063
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_21
timestamp 1679235063
transform 1 0 3036 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1679235063
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_47
timestamp 1679235063
transform 1 0 5428 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_74
timestamp 1679235063
transform 1 0 7912 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1679235063
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_97
timestamp 1679235063
transform 1 0 10028 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_110
timestamp 1679235063
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1679235063
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_136
timestamp 1679235063
transform 1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_141
timestamp 1679235063
transform 1 0 14076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_144
timestamp 1679235063
transform 1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_167
timestamp 1679235063
transform 1 0 16468 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_171
timestamp 1679235063
transform 1 0 16836 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1679235063
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1679235063
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_210
timestamp 1679235063
transform 1 0 20424 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 1679235063
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_229
timestamp 1679235063
transform 1 0 22172 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_244
timestamp 1679235063
transform 1 0 23552 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_255
timestamp 1679235063
transform 1 0 24564 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_260
timestamp 1679235063
transform 1 0 25024 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_271
timestamp 1679235063
transform 1 0 26036 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_279
timestamp 1679235063
transform 1 0 26772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_291
timestamp 1679235063
transform 1 0 27876 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_303
timestamp 1679235063
transform 1 0 28980 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_309
timestamp 1679235063
transform 1 0 29532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_319
timestamp 1679235063
transform 1 0 30452 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1679235063
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1679235063
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1679235063
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1679235063
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1679235063
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1679235063
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1679235063
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_401
timestamp 1679235063
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1679235063
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1679235063
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_421
timestamp 1679235063
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_433
timestamp 1679235063
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_445
timestamp 1679235063
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_457
timestamp 1679235063
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1679235063
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1679235063
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1679235063
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1679235063
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1679235063
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1679235063
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1679235063
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 1679235063
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_21
timestamp 1679235063
transform 1 0 3036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_28
timestamp 1679235063
transform 1 0 3680 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_41
timestamp 1679235063
transform 1 0 4876 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1679235063
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1679235063
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_63
timestamp 1679235063
transform 1 0 6900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_68
timestamp 1679235063
transform 1 0 7360 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_79
timestamp 1679235063
transform 1 0 8372 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_86
timestamp 1679235063
transform 1 0 9016 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_97
timestamp 1679235063
transform 1 0 10028 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1679235063
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_119
timestamp 1679235063
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 1679235063
transform 1 0 13064 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1679235063
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_142
timestamp 1679235063
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_153
timestamp 1679235063
transform 1 0 15180 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1679235063
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_173
timestamp 1679235063
transform 1 0 17020 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1679235063
transform 1 0 19044 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_199
timestamp 1679235063
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1679235063
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_227
timestamp 1679235063
transform 1 0 21988 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_250
timestamp 1679235063
transform 1 0 24104 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_256
timestamp 1679235063
transform 1 0 24656 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1679235063
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_285
timestamp 1679235063
transform 1 0 27324 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_296
timestamp 1679235063
transform 1 0 28336 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1679235063
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_320
timestamp 1679235063
transform 1 0 30544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_332
timestamp 1679235063
transform 1 0 31648 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1679235063
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1679235063
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1679235063
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1679235063
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1679235063
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1679235063
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1679235063
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_405
timestamp 1679235063
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_417
timestamp 1679235063
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_429
timestamp 1679235063
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1679235063
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1679235063
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1679235063
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1679235063
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1679235063
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1679235063
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1679235063
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1679235063
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_505
timestamp 1679235063
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_517
timestamp 1679235063
transform 1 0 48668 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1679235063
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1679235063
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1679235063
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1679235063
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1679235063
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_38
timestamp 1679235063
transform 1 0 4600 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_65
timestamp 1679235063
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_69
timestamp 1679235063
transform 1 0 7452 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_79
timestamp 1679235063
transform 1 0 8372 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 1679235063
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1679235063
transform 1 0 9936 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1679235063
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_110
timestamp 1679235063
transform 1 0 11224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_134
timestamp 1679235063
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_143
timestamp 1679235063
transform 1 0 14260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_146
timestamp 1679235063
transform 1 0 14536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_168
timestamp 1679235063
transform 1 0 16560 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1679235063
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1679235063
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1679235063
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_213
timestamp 1679235063
transform 1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_236
timestamp 1679235063
transform 1 0 22816 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_240
timestamp 1679235063
transform 1 0 23184 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_250
timestamp 1679235063
transform 1 0 24104 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1679235063
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_265
timestamp 1679235063
transform 1 0 25484 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_272
timestamp 1679235063
transform 1 0 26128 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_284
timestamp 1679235063
transform 1 0 27232 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_294
timestamp 1679235063
transform 1 0 28152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1679235063
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1679235063
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_321
timestamp 1679235063
transform 1 0 30636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_325
timestamp 1679235063
transform 1 0 31004 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_331
timestamp 1679235063
transform 1 0 31556 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_338
timestamp 1679235063
transform 1 0 32200 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_346
timestamp 1679235063
transform 1 0 32936 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_358
timestamp 1679235063
transform 1 0 34040 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1679235063
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1679235063
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1679235063
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_401
timestamp 1679235063
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1679235063
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1679235063
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1679235063
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1679235063
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1679235063
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1679235063
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1679235063
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1679235063
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1679235063
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1679235063
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_501
timestamp 1679235063
transform 1 0 47196 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_513
timestamp 1679235063
transform 1 0 48300 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1679235063
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1679235063
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_21
timestamp 1679235063
transform 1 0 3036 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_41
timestamp 1679235063
transform 1 0 4876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1679235063
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1679235063
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_60
timestamp 1679235063
transform 1 0 6624 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_66
timestamp 1679235063
transform 1 0 7176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_79
timestamp 1679235063
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 1679235063
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1679235063
transform 1 0 9936 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1679235063
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 1679235063
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1679235063
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1679235063
transform 1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_141
timestamp 1679235063
transform 1 0 14076 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_154
timestamp 1679235063
transform 1 0 15272 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1679235063
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_169
timestamp 1679235063
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_191
timestamp 1679235063
transform 1 0 18676 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_196
timestamp 1679235063
transform 1 0 19136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1679235063
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_220
timestamp 1679235063
transform 1 0 21344 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_225
timestamp 1679235063
transform 1 0 21804 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_236
timestamp 1679235063
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_244
timestamp 1679235063
transform 1 0 23552 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_254
timestamp 1679235063
transform 1 0 24472 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1679235063
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1679235063
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_291
timestamp 1679235063
transform 1 0 27876 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_303
timestamp 1679235063
transform 1 0 28980 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1679235063
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_327
timestamp 1679235063
transform 1 0 31188 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1679235063
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_337
timestamp 1679235063
transform 1 0 32108 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_349
timestamp 1679235063
transform 1 0 33212 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_356
timestamp 1679235063
transform 1 0 33856 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_360
timestamp 1679235063
transform 1 0 34224 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_372
timestamp 1679235063
transform 1 0 35328 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_384
timestamp 1679235063
transform 1 0 36432 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1679235063
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_405
timestamp 1679235063
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_417
timestamp 1679235063
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_429
timestamp 1679235063
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1679235063
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1679235063
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1679235063
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1679235063
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1679235063
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1679235063
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1679235063
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1679235063
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_505
timestamp 1679235063
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_517
timestamp 1679235063
transform 1 0 48668 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1679235063
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1679235063
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 1679235063
transform 1 0 3036 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_29
timestamp 1679235063
transform 1 0 3772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_47
timestamp 1679235063
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_51
timestamp 1679235063
transform 1 0 5796 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_56
timestamp 1679235063
transform 1 0 6256 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_69
timestamp 1679235063
transform 1 0 7452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1679235063
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1679235063
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_97
timestamp 1679235063
transform 1 0 10028 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1679235063
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_114
timestamp 1679235063
transform 1 0 11592 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_125
timestamp 1679235063
transform 1 0 12604 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1679235063
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 1679235063
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1679235063
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_170
timestamp 1679235063
transform 1 0 16744 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1679235063
transform 1 0 17940 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_191
timestamp 1679235063
transform 1 0 18676 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1679235063
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1679235063
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_222
timestamp 1679235063
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_226
timestamp 1679235063
transform 1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_237
timestamp 1679235063
transform 1 0 22908 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_250
timestamp 1679235063
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_255
timestamp 1679235063
transform 1 0 24564 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_266
timestamp 1679235063
transform 1 0 25576 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_279
timestamp 1679235063
transform 1 0 26772 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_283
timestamp 1679235063
transform 1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_295
timestamp 1679235063
transform 1 0 28244 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_302
timestamp 1679235063
transform 1 0 28888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 1679235063
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_312
timestamp 1679235063
transform 1 0 29808 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_317
timestamp 1679235063
transform 1 0 30268 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_331
timestamp 1679235063
transform 1 0 31556 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_345
timestamp 1679235063
transform 1 0 32844 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_359
timestamp 1679235063
transform 1 0 34132 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1679235063
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1679235063
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_371
timestamp 1679235063
transform 1 0 35236 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_375
timestamp 1679235063
transform 1 0 35604 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_387
timestamp 1679235063
transform 1 0 36708 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_399
timestamp 1679235063
transform 1 0 37812 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_411
timestamp 1679235063
transform 1 0 38916 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1679235063
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1679235063
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1679235063
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1679235063
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1679235063
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1679235063
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1679235063
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1679235063
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1679235063
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_501
timestamp 1679235063
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_513
timestamp 1679235063
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1679235063
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1679235063
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_21
timestamp 1679235063
transform 1 0 3036 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_41
timestamp 1679235063
transform 1 0 4876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1679235063
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1679235063
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_67
timestamp 1679235063
transform 1 0 7268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_80
timestamp 1679235063
transform 1 0 8464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_93
timestamp 1679235063
transform 1 0 9660 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1679235063
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1679235063
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_113
timestamp 1679235063
transform 1 0 11500 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_135
timestamp 1679235063
transform 1 0 13524 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 1679235063
transform 1 0 15180 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1679235063
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1679235063
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1679235063
transform 1 0 17204 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_179
timestamp 1679235063
transform 1 0 17572 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_202
timestamp 1679235063
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_215
timestamp 1679235063
transform 1 0 20884 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1679235063
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 1679235063
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_237
timestamp 1679235063
transform 1 0 22908 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_241
timestamp 1679235063
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_252
timestamp 1679235063
transform 1 0 24288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_276
timestamp 1679235063
transform 1 0 26496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1679235063
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_287
timestamp 1679235063
transform 1 0 27508 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_311
timestamp 1679235063
transform 1 0 29716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_323
timestamp 1679235063
transform 1 0 30820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_327
timestamp 1679235063
transform 1 0 31188 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1679235063
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1679235063
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_347
timestamp 1679235063
transform 1 0 33028 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_359
timestamp 1679235063
transform 1 0 34132 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_367
timestamp 1679235063
transform 1 0 34868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_27_374
timestamp 1679235063
transform 1 0 35512 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_379
timestamp 1679235063
transform 1 0 35972 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1679235063
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1679235063
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_405
timestamp 1679235063
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_417
timestamp 1679235063
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_429
timestamp 1679235063
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1679235063
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1679235063
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1679235063
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_461
timestamp 1679235063
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_473
timestamp 1679235063
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_485
timestamp 1679235063
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1679235063
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1679235063
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1679235063
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1679235063
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1679235063
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_3
timestamp 1679235063
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_21
timestamp 1679235063
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_31
timestamp 1679235063
transform 1 0 3956 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_36
timestamp 1679235063
transform 1 0 4416 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_60
timestamp 1679235063
transform 1 0 6624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_64
timestamp 1679235063
transform 1 0 6992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_69
timestamp 1679235063
transform 1 0 7452 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1679235063
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_85
timestamp 1679235063
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_98
timestamp 1679235063
transform 1 0 10120 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1679235063
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_126
timestamp 1679235063
transform 1 0 12696 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1679235063
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1679235063
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_146
timestamp 1679235063
transform 1 0 14536 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_156
timestamp 1679235063
transform 1 0 15456 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_181
timestamp 1679235063
transform 1 0 17756 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_185
timestamp 1679235063
transform 1 0 18124 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1679235063
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1679235063
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1679235063
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_207
timestamp 1679235063
transform 1 0 20148 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_217
timestamp 1679235063
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_224
timestamp 1679235063
transform 1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_248
timestamp 1679235063
transform 1 0 23920 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_255
timestamp 1679235063
transform 1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_278
timestamp 1679235063
transform 1 0 26680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_302
timestamp 1679235063
transform 1 0 28888 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1679235063
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_320
timestamp 1679235063
transform 1 0 30544 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_332
timestamp 1679235063
transform 1 0 31648 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_344
timestamp 1679235063
transform 1 0 32752 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_356
timestamp 1679235063
transform 1 0 33856 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_365
timestamp 1679235063
transform 1 0 34684 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_375
timestamp 1679235063
transform 1 0 35604 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_382
timestamp 1679235063
transform 1 0 36248 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_390
timestamp 1679235063
transform 1 0 36984 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_397
timestamp 1679235063
transform 1 0 37628 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_401
timestamp 1679235063
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1679235063
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1679235063
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1679235063
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1679235063
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_445
timestamp 1679235063
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_457
timestamp 1679235063
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1679235063
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1679235063
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1679235063
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1679235063
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_501
timestamp 1679235063
transform 1 0 47196 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_513
timestamp 1679235063
transform 1 0 48300 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1679235063
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1679235063
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_21
timestamp 1679235063
transform 1 0 3036 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_41
timestamp 1679235063
transform 1 0 4876 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1679235063
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_57
timestamp 1679235063
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_75
timestamp 1679235063
transform 1 0 8004 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1679235063
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_96
timestamp 1679235063
transform 1 0 9936 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_109
timestamp 1679235063
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_119
timestamp 1679235063
transform 1 0 12052 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_130
timestamp 1679235063
transform 1 0 13064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_145
timestamp 1679235063
transform 1 0 14444 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_158
timestamp 1679235063
transform 1 0 15640 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1679235063
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1679235063
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1679235063
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_192
timestamp 1679235063
transform 1 0 18768 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1679235063
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_209
timestamp 1679235063
transform 1 0 20332 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_212
timestamp 1679235063
transform 1 0 20608 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1679235063
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_225
timestamp 1679235063
transform 1 0 21804 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_235
timestamp 1679235063
transform 1 0 22724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_259
timestamp 1679235063
transform 1 0 24932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_274
timestamp 1679235063
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1679235063
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_286
timestamp 1679235063
transform 1 0 27416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_290
timestamp 1679235063
transform 1 0 27784 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_313
timestamp 1679235063
transform 1 0 29900 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_325
timestamp 1679235063
transform 1 0 31004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_329
timestamp 1679235063
transform 1 0 31372 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_334
timestamp 1679235063
transform 1 0 31832 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_345
timestamp 1679235063
transform 1 0 32844 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_359
timestamp 1679235063
transform 1 0 34132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_373
timestamp 1679235063
transform 1 0 35420 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_385
timestamp 1679235063
transform 1 0 36524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_389
timestamp 1679235063
transform 1 0 36892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1679235063
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_399
timestamp 1679235063
transform 1 0 37812 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_407
timestamp 1679235063
transform 1 0 38548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_414
timestamp 1679235063
transform 1 0 39192 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_418
timestamp 1679235063
transform 1 0 39560 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_430
timestamp 1679235063
transform 1 0 40664 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_442
timestamp 1679235063
transform 1 0 41768 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1679235063
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1679235063
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1679235063
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1679235063
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1679235063
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1679235063
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_505
timestamp 1679235063
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_517
timestamp 1679235063
transform 1 0 48668 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1679235063
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 1679235063
transform 1 0 1380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_21
timestamp 1679235063
transform 1 0 3036 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1679235063
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_47
timestamp 1679235063
transform 1 0 5428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_67
timestamp 1679235063
transform 1 0 7268 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_80
timestamp 1679235063
transform 1 0 8464 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1679235063
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_96
timestamp 1679235063
transform 1 0 9936 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1679235063
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_126
timestamp 1679235063
transform 1 0 12696 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1679235063
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1679235063
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1679235063
transform 1 0 14536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1679235063
transform 1 0 16560 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_175
timestamp 1679235063
transform 1 0 17204 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1679235063
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_199
timestamp 1679235063
transform 1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_212
timestamp 1679235063
transform 1 0 20608 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_216
timestamp 1679235063
transform 1 0 20976 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_237
timestamp 1679235063
transform 1 0 22908 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1679235063
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1679235063
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_259
timestamp 1679235063
transform 1 0 24932 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_263
timestamp 1679235063
transform 1 0 25300 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_285
timestamp 1679235063
transform 1 0 27324 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_292
timestamp 1679235063
transform 1 0 27968 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_296
timestamp 1679235063
transform 1 0 28336 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1679235063
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_309
timestamp 1679235063
transform 1 0 29532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_319
timestamp 1679235063
transform 1 0 30452 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_331
timestamp 1679235063
transform 1 0 31556 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_337
timestamp 1679235063
transform 1 0 32108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_347
timestamp 1679235063
transform 1 0 33028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_354
timestamp 1679235063
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_362
timestamp 1679235063
transform 1 0 34408 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_377
timestamp 1679235063
transform 1 0 35788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_389
timestamp 1679235063
transform 1 0 36892 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_393
timestamp 1679235063
transform 1 0 37260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1679235063
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_411
timestamp 1679235063
transform 1 0 38916 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_418
timestamp 1679235063
transform 1 0 39560 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_427
timestamp 1679235063
transform 1 0 40388 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_439
timestamp 1679235063
transform 1 0 41492 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_451
timestamp 1679235063
transform 1 0 42596 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_463
timestamp 1679235063
transform 1 0 43700 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1679235063
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1679235063
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1679235063
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_501
timestamp 1679235063
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_513
timestamp 1679235063
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1679235063
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_3
timestamp 1679235063
transform 1 0 1380 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_21
timestamp 1679235063
transform 1 0 3036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1679235063
transform 1 0 4876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1679235063
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1679235063
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_79
timestamp 1679235063
transform 1 0 8372 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1679235063
transform 1 0 9016 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_97
timestamp 1679235063
transform 1 0 10028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1679235063
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1679235063
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1679235063
transform 1 0 12420 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_138
timestamp 1679235063
transform 1 0 13800 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_142
timestamp 1679235063
transform 1 0 14168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_152
timestamp 1679235063
transform 1 0 15088 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1679235063
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_169
timestamp 1679235063
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_180
timestamp 1679235063
transform 1 0 17664 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_193
timestamp 1679235063
transform 1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_200
timestamp 1679235063
transform 1 0 19504 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_222
timestamp 1679235063
transform 1 0 21528 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1679235063
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_236
timestamp 1679235063
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_244
timestamp 1679235063
transform 1 0 23552 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_255
timestamp 1679235063
transform 1 0 24564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_270
timestamp 1679235063
transform 1 0 25944 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1679235063
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1679235063
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_292
timestamp 1679235063
transform 1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_316
timestamp 1679235063
transform 1 0 30176 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_328
timestamp 1679235063
transform 1 0 31280 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1679235063
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_347
timestamp 1679235063
transform 1 0 33028 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_359
timestamp 1679235063
transform 1 0 34132 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_365
timestamp 1679235063
transform 1 0 34684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_375
timestamp 1679235063
transform 1 0 35604 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_387
timestamp 1679235063
transform 1 0 36708 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1679235063
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_405
timestamp 1679235063
transform 1 0 38364 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_413
timestamp 1679235063
transform 1 0 39100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_420
timestamp 1679235063
transform 1 0 39744 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_426
timestamp 1679235063
transform 1 0 40296 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_433
timestamp 1679235063
transform 1 0 40940 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1679235063
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1679235063
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1679235063
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1679235063
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1679235063
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1679235063
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1679235063
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1679235063
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_505
timestamp 1679235063
transform 1 0 47564 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_517
timestamp 1679235063
transform 1 0 48668 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1679235063
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1679235063
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_21
timestamp 1679235063
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_34
timestamp 1679235063
transform 1 0 4232 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_58
timestamp 1679235063
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1679235063
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_87
timestamp 1679235063
transform 1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_93
timestamp 1679235063
transform 1 0 9660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_117
timestamp 1679235063
transform 1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_124
timestamp 1679235063
transform 1 0 12512 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_135
timestamp 1679235063
transform 1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_141
timestamp 1679235063
transform 1 0 14076 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_165
timestamp 1679235063
transform 1 0 16284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_170
timestamp 1679235063
transform 1 0 16744 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_181
timestamp 1679235063
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1679235063
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1679235063
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_204
timestamp 1679235063
transform 1 0 19872 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_228
timestamp 1679235063
transform 1 0 22080 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_234
timestamp 1679235063
transform 1 0 22632 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_245
timestamp 1679235063
transform 1 0 23644 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_32_253
timestamp 1679235063
transform 1 0 24380 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_265
timestamp 1679235063
transform 1 0 25484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_289
timestamp 1679235063
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_301
timestamp 1679235063
transform 1 0 28796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_305
timestamp 1679235063
transform 1 0 29164 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1679235063
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_320
timestamp 1679235063
transform 1 0 30544 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_332
timestamp 1679235063
transform 1 0 31648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_336
timestamp 1679235063
transform 1 0 32016 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_347
timestamp 1679235063
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_32_359
timestamp 1679235063
transform 1 0 34132 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1679235063
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_375
timestamp 1679235063
transform 1 0 35604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_387
timestamp 1679235063
transform 1 0 36708 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_399
timestamp 1679235063
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_411
timestamp 1679235063
transform 1 0 38916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_418
timestamp 1679235063
transform 1 0 39560 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_421
timestamp 1679235063
transform 1 0 39836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_427
timestamp 1679235063
transform 1 0 40388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_435
timestamp 1679235063
transform 1 0 41124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_442
timestamp 1679235063
transform 1 0 41768 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_452
timestamp 1679235063
transform 1 0 42688 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_464
timestamp 1679235063
transform 1 0 43792 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1679235063
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1679235063
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1679235063
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1679235063
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1679235063
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1679235063
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_21
timestamp 1679235063
transform 1 0 3036 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_29
timestamp 1679235063
transform 1 0 3772 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_33
timestamp 1679235063
transform 1 0 4140 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1679235063
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1679235063
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_75
timestamp 1679235063
transform 1 0 8004 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_102
timestamp 1679235063
transform 1 0 10488 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1679235063
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_113
timestamp 1679235063
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_118
timestamp 1679235063
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_131
timestamp 1679235063
transform 1 0 13156 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_155
timestamp 1679235063
transform 1 0 15364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_159
timestamp 1679235063
transform 1 0 15732 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1679235063
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_33_169
timestamp 1679235063
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1679235063
transform 1 0 16928 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_183
timestamp 1679235063
transform 1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_187
timestamp 1679235063
transform 1 0 18308 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_198
timestamp 1679235063
transform 1 0 19320 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1679235063
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_225
timestamp 1679235063
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_238
timestamp 1679235063
transform 1 0 23000 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_246
timestamp 1679235063
transform 1 0 23736 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_251
timestamp 1679235063
transform 1 0 24196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_273
timestamp 1679235063
transform 1 0 26220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_281
timestamp 1679235063
transform 1 0 26956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_292
timestamp 1679235063
transform 1 0 27968 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_296
timestamp 1679235063
transform 1 0 28336 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_317
timestamp 1679235063
transform 1 0 30268 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_330
timestamp 1679235063
transform 1 0 31464 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1679235063
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_347
timestamp 1679235063
transform 1 0 33028 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_359
timestamp 1679235063
transform 1 0 34132 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_365
timestamp 1679235063
transform 1 0 34684 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_375
timestamp 1679235063
transform 1 0 35604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_387
timestamp 1679235063
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_393
timestamp 1679235063
transform 1 0 37260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_405
timestamp 1679235063
transform 1 0 38364 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_419
timestamp 1679235063
transform 1 0 39652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_429
timestamp 1679235063
transform 1 0 40572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_433
timestamp 1679235063
transform 1 0 40940 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_446
timestamp 1679235063
transform 1 0 42136 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_449
timestamp 1679235063
transform 1 0 42412 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_454
timestamp 1679235063
transform 1 0 42872 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_464
timestamp 1679235063
transform 1 0 43792 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_476
timestamp 1679235063
transform 1 0 44896 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_488
timestamp 1679235063
transform 1 0 46000 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_500
timestamp 1679235063
transform 1 0 47104 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_505
timestamp 1679235063
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_517
timestamp 1679235063
transform 1 0 48668 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1679235063
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_21
timestamp 1679235063
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_29
timestamp 1679235063
transform 1 0 3772 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_47
timestamp 1679235063
transform 1 0 5428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_53
timestamp 1679235063
transform 1 0 5980 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_75
timestamp 1679235063
transform 1 0 8004 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_82
timestamp 1679235063
transform 1 0 8648 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1679235063
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_103
timestamp 1679235063
transform 1 0 10580 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_116
timestamp 1679235063
transform 1 0 11776 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1679235063
transform 1 0 13432 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_141
timestamp 1679235063
transform 1 0 14076 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_144
timestamp 1679235063
transform 1 0 14352 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_155
timestamp 1679235063
transform 1 0 15364 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_168
timestamp 1679235063
transform 1 0 16560 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_181
timestamp 1679235063
transform 1 0 17756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_194
timestamp 1679235063
transform 1 0 18952 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_197
timestamp 1679235063
transform 1 0 19228 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_219
timestamp 1679235063
transform 1 0 21252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_234
timestamp 1679235063
transform 1 0 22632 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_34_247
timestamp 1679235063
transform 1 0 23828 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_34_253
timestamp 1679235063
transform 1 0 24380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_265
timestamp 1679235063
transform 1 0 25484 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_269
timestamp 1679235063
transform 1 0 25852 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_290
timestamp 1679235063
transform 1 0 27784 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_302
timestamp 1679235063
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_34_309
timestamp 1679235063
transform 1 0 29532 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_323
timestamp 1679235063
transform 1 0 30820 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1679235063
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_348
timestamp 1679235063
transform 1 0 33120 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_360
timestamp 1679235063
transform 1 0 34224 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1679235063
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_371
timestamp 1679235063
transform 1 0 35236 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_375
timestamp 1679235063
transform 1 0 35604 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_387
timestamp 1679235063
transform 1 0 36708 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_399
timestamp 1679235063
transform 1 0 37812 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_411
timestamp 1679235063
transform 1 0 38916 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_418
timestamp 1679235063
transform 1 0 39560 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_421
timestamp 1679235063
transform 1 0 39836 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_431
timestamp 1679235063
transform 1 0 40756 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_439
timestamp 1679235063
transform 1 0 41492 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_447
timestamp 1679235063
transform 1 0 42228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_455
timestamp 1679235063
transform 1 0 42964 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_462
timestamp 1679235063
transform 1 0 43608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_469
timestamp 1679235063
transform 1 0 44252 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1679235063
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1679235063
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1679235063
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_501
timestamp 1679235063
transform 1 0 47196 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_509
timestamp 1679235063
transform 1 0 47932 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_515
timestamp 1679235063
transform 1 0 48484 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1679235063
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_3
timestamp 1679235063
transform 1 0 1380 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_21
timestamp 1679235063
transform 1 0 3036 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_41
timestamp 1679235063
transform 1 0 4876 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_54
timestamp 1679235063
transform 1 0 6072 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_68
timestamp 1679235063
transform 1 0 7360 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_92
timestamp 1679235063
transform 1 0 9568 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_97
timestamp 1679235063
transform 1 0 10028 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_110
timestamp 1679235063
transform 1 0 11224 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_113
timestamp 1679235063
transform 1 0 11500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_124
timestamp 1679235063
transform 1 0 12512 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_149
timestamp 1679235063
transform 1 0 14812 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1679235063
transform 1 0 15364 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1679235063
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_169
timestamp 1679235063
transform 1 0 16652 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1679235063
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_211
timestamp 1679235063
transform 1 0 20516 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_215
timestamp 1679235063
transform 1 0 20884 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1679235063
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1679235063
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_238
timestamp 1679235063
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1679235063
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_275
timestamp 1679235063
transform 1 0 26404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1679235063
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_281
timestamp 1679235063
transform 1 0 26956 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_293
timestamp 1679235063
transform 1 0 28060 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_317
timestamp 1679235063
transform 1 0 30268 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_330
timestamp 1679235063
transform 1 0 31464 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1679235063
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_347
timestamp 1679235063
transform 1 0 33028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_359
timestamp 1679235063
transform 1 0 34132 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_365
timestamp 1679235063
transform 1 0 34684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_375
timestamp 1679235063
transform 1 0 35604 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_35_387
timestamp 1679235063
transform 1 0 36708 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_393
timestamp 1679235063
transform 1 0 37260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_405
timestamp 1679235063
transform 1 0 38364 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_417
timestamp 1679235063
transform 1 0 39468 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_429
timestamp 1679235063
transform 1 0 40572 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_441
timestamp 1679235063
transform 1 0 41676 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1679235063
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_449
timestamp 1679235063
transform 1 0 42412 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_455
timestamp 1679235063
transform 1 0 42964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_463
timestamp 1679235063
transform 1 0 43700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_470
timestamp 1679235063
transform 1 0 44344 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_477
timestamp 1679235063
transform 1 0 44988 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_487
timestamp 1679235063
transform 1 0 45908 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_502
timestamp 1679235063
transform 1 0 47288 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_507
timestamp 1679235063
transform 1 0 47748 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1679235063
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1679235063
transform 1 0 1380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_21
timestamp 1679235063
transform 1 0 3036 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_29
timestamp 1679235063
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_47
timestamp 1679235063
transform 1 0 5428 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1679235063
transform 1 0 5888 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_58
timestamp 1679235063
transform 1 0 6440 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_78
timestamp 1679235063
transform 1 0 8280 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_87
timestamp 1679235063
transform 1 0 9108 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_98
timestamp 1679235063
transform 1 0 10120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_118
timestamp 1679235063
transform 1 0 11960 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1679235063
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_143
timestamp 1679235063
transform 1 0 14260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_149
timestamp 1679235063
transform 1 0 14812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_169
timestamp 1679235063
transform 1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_173
timestamp 1679235063
transform 1 0 17020 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_194
timestamp 1679235063
transform 1 0 18952 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1679235063
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1679235063
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_225
timestamp 1679235063
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1679235063
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1679235063
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_253
timestamp 1679235063
transform 1 0 24380 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_264
timestamp 1679235063
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_288
timestamp 1679235063
transform 1 0 27600 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_300
timestamp 1679235063
transform 1 0 28704 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1679235063
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_320
timestamp 1679235063
transform 1 0 30544 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_332
timestamp 1679235063
transform 1 0 31648 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_336
timestamp 1679235063
transform 1 0 32016 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_347
timestamp 1679235063
transform 1 0 33028 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_359
timestamp 1679235063
transform 1 0 34132 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1679235063
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_365
timestamp 1679235063
transform 1 0 34684 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1679235063
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_387
timestamp 1679235063
transform 1 0 36708 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_393
timestamp 1679235063
transform 1 0 37260 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1679235063
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_415
timestamp 1679235063
transform 1 0 39284 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_419
timestamp 1679235063
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_421
timestamp 1679235063
transform 1 0 39836 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_433
timestamp 1679235063
transform 1 0 40940 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_447
timestamp 1679235063
transform 1 0 42228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_459
timestamp 1679235063
transform 1 0 43332 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_471
timestamp 1679235063
transform 1 0 44436 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1679235063
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_477
timestamp 1679235063
transform 1 0 44988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_483
timestamp 1679235063
transform 1 0 45540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_491
timestamp 1679235063
transform 1 0 46276 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_499
timestamp 1679235063
transform 1 0 47012 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_505
timestamp 1679235063
transform 1 0 47564 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_513
timestamp 1679235063
transform 1 0 48300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1679235063
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1679235063
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_21
timestamp 1679235063
transform 1 0 3036 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_36
timestamp 1679235063
transform 1 0 4416 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1679235063
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1679235063
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_63
timestamp 1679235063
transform 1 0 6900 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_67
timestamp 1679235063
transform 1 0 7268 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_84
timestamp 1679235063
transform 1 0 8832 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_108
timestamp 1679235063
transform 1 0 11040 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_119
timestamp 1679235063
transform 1 0 12052 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_142
timestamp 1679235063
transform 1 0 14168 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_148
timestamp 1679235063
transform 1 0 14720 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_166
timestamp 1679235063
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_169
timestamp 1679235063
transform 1 0 16652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_191
timestamp 1679235063
transform 1 0 18676 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1679235063
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1679235063
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_225
timestamp 1679235063
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_235
timestamp 1679235063
transform 1 0 22724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_259
timestamp 1679235063
transform 1 0 24932 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_272
timestamp 1679235063
transform 1 0 26128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_281
timestamp 1679235063
transform 1 0 26956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_293
timestamp 1679235063
transform 1 0 28060 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_317
timestamp 1679235063
transform 1 0 30268 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_330
timestamp 1679235063
transform 1 0 31464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1679235063
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_347
timestamp 1679235063
transform 1 0 33028 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_359
timestamp 1679235063
transform 1 0 34132 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_365
timestamp 1679235063
transform 1 0 34684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_375
timestamp 1679235063
transform 1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_387
timestamp 1679235063
transform 1 0 36708 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1679235063
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1679235063
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1679235063
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_415
timestamp 1679235063
transform 1 0 39284 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_427
timestamp 1679235063
transform 1 0 40388 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_439
timestamp 1679235063
transform 1 0 41492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_446
timestamp 1679235063
transform 1 0 42136 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_449
timestamp 1679235063
transform 1 0 42412 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_461
timestamp 1679235063
transform 1 0 43516 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_473
timestamp 1679235063
transform 1 0 44620 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_481
timestamp 1679235063
transform 1 0 45356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_489
timestamp 1679235063
transform 1 0 46092 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_497
timestamp 1679235063
transform 1 0 46828 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1679235063
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_505
timestamp 1679235063
transform 1 0 47564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_511
timestamp 1679235063
transform 1 0 48116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_515
timestamp 1679235063
transform 1 0 48484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1679235063
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1679235063
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_21
timestamp 1679235063
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_29
timestamp 1679235063
transform 1 0 3772 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_41
timestamp 1679235063
transform 1 0 4876 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1679235063
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_62
timestamp 1679235063
transform 1 0 6808 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1679235063
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_87
timestamp 1679235063
transform 1 0 9108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_105
timestamp 1679235063
transform 1 0 10764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_132
timestamp 1679235063
transform 1 0 13248 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_141
timestamp 1679235063
transform 1 0 14076 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_144
timestamp 1679235063
transform 1 0 14352 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_150
timestamp 1679235063
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_170
timestamp 1679235063
transform 1 0 16744 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1679235063
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1679235063
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_202
timestamp 1679235063
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_226
timestamp 1679235063
transform 1 0 21896 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1679235063
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1679235063
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1679235063
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_277
timestamp 1679235063
transform 1 0 26588 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_283
timestamp 1679235063
transform 1 0 27140 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_305
timestamp 1679235063
transform 1 0 29164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1679235063
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_331
timestamp 1679235063
transform 1 0 31556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_337
timestamp 1679235063
transform 1 0 32108 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_347
timestamp 1679235063
transform 1 0 33028 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_359
timestamp 1679235063
transform 1 0 34132 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1679235063
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1679235063
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_375
timestamp 1679235063
transform 1 0 35604 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_387
timestamp 1679235063
transform 1 0 36708 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_394
timestamp 1679235063
transform 1 0 37352 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_418
timestamp 1679235063
transform 1 0 39560 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1679235063
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_431
timestamp 1679235063
transform 1 0 40756 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_443
timestamp 1679235063
transform 1 0 41860 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_455
timestamp 1679235063
transform 1 0 42964 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_467
timestamp 1679235063
transform 1 0 44068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_474
timestamp 1679235063
transform 1 0 44712 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_477
timestamp 1679235063
transform 1 0 44988 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_487
timestamp 1679235063
transform 1 0 45908 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_491
timestamp 1679235063
transform 1 0 46276 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_501
timestamp 1679235063
transform 1 0 47196 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_513
timestamp 1679235063
transform 1 0 48300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1679235063
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_3
timestamp 1679235063
transform 1 0 1380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_14
timestamp 1679235063
transform 1 0 2392 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_34
timestamp 1679235063
transform 1 0 4232 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_54
timestamp 1679235063
transform 1 0 6072 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_57
timestamp 1679235063
transform 1 0 6348 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_69
timestamp 1679235063
transform 1 0 7452 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_73
timestamp 1679235063
transform 1 0 7820 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_90
timestamp 1679235063
transform 1 0 9384 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_110
timestamp 1679235063
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_126
timestamp 1679235063
transform 1 0 12696 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_146
timestamp 1679235063
transform 1 0 14536 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_166
timestamp 1679235063
transform 1 0 16376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_169
timestamp 1679235063
transform 1 0 16652 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_188
timestamp 1679235063
transform 1 0 18400 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_213
timestamp 1679235063
transform 1 0 20700 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1679235063
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_247
timestamp 1679235063
transform 1 0 23828 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_254
timestamp 1679235063
transform 1 0 24472 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1679235063
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_281
timestamp 1679235063
transform 1 0 26956 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_303
timestamp 1679235063
transform 1 0 28980 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_317
timestamp 1679235063
transform 1 0 30268 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_321
timestamp 1679235063
transform 1 0 30636 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_334
timestamp 1679235063
transform 1 0 31832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1679235063
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_347
timestamp 1679235063
transform 1 0 33028 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_359
timestamp 1679235063
transform 1 0 34132 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_365
timestamp 1679235063
transform 1 0 34684 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_375
timestamp 1679235063
transform 1 0 35604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_387
timestamp 1679235063
transform 1 0 36708 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1679235063
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1679235063
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_415
timestamp 1679235063
transform 1 0 39284 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_427
timestamp 1679235063
transform 1 0 40388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_439
timestamp 1679235063
transform 1 0 41492 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_446
timestamp 1679235063
transform 1 0 42136 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_449
timestamp 1679235063
transform 1 0 42412 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_455
timestamp 1679235063
transform 1 0 42964 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_459
timestamp 1679235063
transform 1 0 43332 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_471
timestamp 1679235063
transform 1 0 44436 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_483
timestamp 1679235063
transform 1 0 45540 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_497
timestamp 1679235063
transform 1 0 46828 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1679235063
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_505
timestamp 1679235063
transform 1 0 47564 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_515
timestamp 1679235063
transform 1 0 48484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_523
timestamp 1679235063
transform 1 0 49220 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_3
timestamp 1679235063
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_8
timestamp 1679235063
transform 1 0 1840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_26
timestamp 1679235063
transform 1 0 3496 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_29
timestamp 1679235063
transform 1 0 3772 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_34
timestamp 1679235063
transform 1 0 4232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_54
timestamp 1679235063
transform 1 0 6072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_57
timestamp 1679235063
transform 1 0 6348 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_62
timestamp 1679235063
transform 1 0 6808 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_82
timestamp 1679235063
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_90
timestamp 1679235063
transform 1 0 9384 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_110
timestamp 1679235063
transform 1 0 11224 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1679235063
transform 1 0 11960 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_138
timestamp 1679235063
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_141
timestamp 1679235063
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_146
timestamp 1679235063
transform 1 0 14536 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_166
timestamp 1679235063
transform 1 0 16376 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_169
timestamp 1679235063
transform 1 0 16652 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_192
timestamp 1679235063
transform 1 0 18768 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1679235063
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_202
timestamp 1679235063
transform 1 0 19688 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_222
timestamp 1679235063
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_225
timestamp 1679235063
transform 1 0 21804 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_243
timestamp 1679235063
transform 1 0 23460 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1679235063
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1679235063
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_264
timestamp 1679235063
transform 1 0 25392 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_277
timestamp 1679235063
transform 1 0 26588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_281
timestamp 1679235063
transform 1 0 26956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_292
timestamp 1679235063
transform 1 0 27968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_304
timestamp 1679235063
transform 1 0 29072 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1679235063
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_321
timestamp 1679235063
transform 1 0 30636 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_333
timestamp 1679235063
transform 1 0 31740 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_337
timestamp 1679235063
transform 1 0 32108 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_347
timestamp 1679235063
transform 1 0 33028 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_359
timestamp 1679235063
transform 1 0 34132 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1679235063
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1679235063
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_375
timestamp 1679235063
transform 1 0 35604 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_387
timestamp 1679235063
transform 1 0 36708 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_393
timestamp 1679235063
transform 1 0 37260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1679235063
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_415
timestamp 1679235063
transform 1 0 39284 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1679235063
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1679235063
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_431
timestamp 1679235063
transform 1 0 40756 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_435
timestamp 1679235063
transform 1 0 41124 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_446
timestamp 1679235063
transform 1 0 42136 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_449
timestamp 1679235063
transform 1 0 42412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_461
timestamp 1679235063
transform 1 0 43516 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_473
timestamp 1679235063
transform 1 0 44620 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_477
timestamp 1679235063
transform 1 0 44988 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_487
timestamp 1679235063
transform 1 0 45908 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_491
timestamp 1679235063
transform 1 0 46276 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_502
timestamp 1679235063
transform 1 0 47288 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1679235063
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_515
timestamp 1679235063
transform 1 0 48484 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_523
timestamp 1679235063
transform 1 0 49220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1679235063
transform 1 0 45172 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1679235063
transform 1 0 1656 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1679235063
transform 1 0 6532 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1679235063
transform 1 0 37444 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1679235063
transform 1 0 30912 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold7 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1679235063
transform 1 0 28152 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1679235063
transform 1 0 35972 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1679235063
transform 1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1679235063
transform 1 0 20608 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1679235063
transform 1 0 38180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1679235063
transform 1 0 23092 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1679235063
transform 1 0 37076 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1679235063
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1679235063
transform 1 0 6532 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1679235063
transform 1 0 7912 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1679235063
transform 1 0 30912 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold19
timestamp 1679235063
transform 1 0 27140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold20
timestamp 1679235063
transform 1 0 8740 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1679235063
transform 1 0 43332 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1679235063
transform 1 0 8280 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1679235063
transform 1 0 28704 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1679235063
transform 1 0 4232 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1679235063
transform 1 0 14536 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1679235063
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1679235063
transform 1 0 18216 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1679235063
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1679235063
transform 1 0 11960 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold30
timestamp 1679235063
transform 1 0 13524 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1679235063
transform 1 0 40020 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold32
timestamp 1679235063
transform 1 0 10856 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1679235063
transform 1 0 25024 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1679235063
transform 1 0 37444 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 29348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1679235063
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold37
timestamp 1679235063
transform 1 0 5428 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold38
timestamp 1679235063
transform 1 0 24564 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold39
timestamp 1679235063
transform 1 0 37444 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1679235063
transform 1 0 17940 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1679235063
transform 1 0 34868 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1679235063
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1679235063
transform 1 0 33396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1679235063
transform 1 0 40020 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1679235063
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold46
timestamp 1679235063
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1679235063
transform 1 0 8924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold48
timestamp 1679235063
transform 1 0 17112 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold49
timestamp 1679235063
transform 1 0 18032 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1679235063
transform 1 0 25760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1679235063
transform 1 0 8280 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1679235063
transform 1 0 12420 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold53
timestamp 1679235063
transform 1 0 37076 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold54
timestamp 1679235063
transform 1 0 9108 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1679235063
transform 1 0 38548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1679235063
transform 1 0 30268 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold57
timestamp 1679235063
transform 1 0 9292 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1679235063
transform 1 0 33396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold59
timestamp 1679235063
transform 1 0 6716 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1679235063
transform 1 0 32292 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1679235063
transform 1 0 34868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold62
timestamp 1679235063
transform 1 0 14628 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1679235063
transform 1 0 9476 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1679235063
transform 1 0 32292 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1679235063
transform 1 0 34868 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1679235063
transform 1 0 32292 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1679235063
transform 1 0 32292 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1679235063
transform 1 0 19964 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1679235063
transform 1 0 14536 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1679235063
transform 1 0 11684 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold71
timestamp 1679235063
transform 1 0 6808 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1679235063
transform 1 0 4600 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold73
timestamp 1679235063
transform 1 0 28336 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1679235063
transform 1 0 43884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold75
timestamp 1679235063
transform 1 0 5612 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1679235063
transform 1 0 33396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1679235063
transform 1 0 33396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1679235063
transform 1 0 45172 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold79
timestamp 1679235063
transform 1 0 21988 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold80
timestamp 1679235063
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1679235063
transform 1 0 32016 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1679235063
transform 1 0 41124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1679235063
transform 1 0 35972 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1679235063
transform 1 0 27140 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1679235063
transform 1 0 32292 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1679235063
transform 1 0 35972 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold87
timestamp 1679235063
transform 1 0 28520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold88
timestamp 1679235063
transform 1 0 14720 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold89
timestamp 1679235063
transform 1 0 38732 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold90
timestamp 1679235063
transform 1 0 13340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1679235063
transform 1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1679235063
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold93
timestamp 1679235063
transform 1 0 27140 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1679235063
transform 1 0 21988 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold95
timestamp 1679235063
transform 1 0 6532 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1679235063
transform 1 0 7912 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1679235063
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1679235063
transform 1 0 24564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1679235063
transform 1 0 5336 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1679235063
transform 1 0 21988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1679235063
transform 1 0 20516 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold102
timestamp 1679235063
transform 1 0 19044 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1679235063
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold104
timestamp 1679235063
transform 1 0 27140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold105
timestamp 1679235063
transform 1 0 32292 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold106
timestamp 1679235063
transform 1 0 25668 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold107
timestamp 1679235063
transform 1 0 26772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold108
timestamp 1679235063
transform 1 0 25668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold109
timestamp 1679235063
transform 1 0 34868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold110
timestamp 1679235063
transform 1 0 42596 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1679235063
transform 1 0 4048 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold112
timestamp 1679235063
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold113
timestamp 1679235063
transform 1 0 14536 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold114
timestamp 1679235063
transform 1 0 4232 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold115
timestamp 1679235063
transform 1 0 1656 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold116
timestamp 1679235063
transform 1 0 3128 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1679235063
transform 1 0 48668 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold118
timestamp 1679235063
transform 1 0 47564 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold119
timestamp 1679235063
transform 1 0 47748 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1679235063
transform 1 0 42596 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold121
timestamp 1679235063
transform 1 0 3956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold122
timestamp 1679235063
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold123
timestamp 1679235063
transform 1 0 4600 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1679235063
transform 1 0 7728 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold125
timestamp 1679235063
transform 1 0 38548 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold126
timestamp 1679235063
transform 1 0 35972 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold127
timestamp 1679235063
transform 1 0 32292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold128
timestamp 1679235063
transform 1 0 32292 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold129
timestamp 1679235063
transform 1 0 4232 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold130
timestamp 1679235063
transform 1 0 1932 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold131
timestamp 1679235063
transform 1 0 32384 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold132
timestamp 1679235063
transform 1 0 27968 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold133
timestamp 1679235063
transform 1 0 20148 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold134
timestamp 1679235063
transform 1 0 21804 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold135
timestamp 1679235063
transform 1 0 21988 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold136
timestamp 1679235063
transform 1 0 23092 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold137
timestamp 1679235063
transform 1 0 33120 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold138
timestamp 1679235063
transform 1 0 33212 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold139
timestamp 1679235063
transform 1 0 35972 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold140
timestamp 1679235063
transform 1 0 37444 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold141
timestamp 1679235063
transform 1 0 16836 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold142
timestamp 1679235063
transform 1 0 23092 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold143
timestamp 1679235063
transform 1 0 13340 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold144
timestamp 1679235063
transform 1 0 14260 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold145
timestamp 1679235063
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold146
timestamp 1679235063
transform 1 0 4324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold147
timestamp 1679235063
transform 1 0 38732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold148
timestamp 1679235063
transform 1 0 40020 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold149
timestamp 1679235063
transform 1 0 21988 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold150
timestamp 1679235063
transform 1 0 23184 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold151
timestamp 1679235063
transform 1 0 2024 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold152
timestamp 1679235063
transform 1 0 7176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold153
timestamp 1679235063
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold154
timestamp 1679235063
transform 1 0 28244 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold155
timestamp 1679235063
transform 1 0 7820 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold156
timestamp 1679235063
transform 1 0 2760 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold157
timestamp 1679235063
transform 1 0 44804 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold158
timestamp 1679235063
transform 1 0 41860 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold159
timestamp 1679235063
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold160
timestamp 1679235063
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold161
timestamp 1679235063
transform 1 0 29716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1679235063
transform 1 0 28244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold163
timestamp 1679235063
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold164
timestamp 1679235063
transform 1 0 16744 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold165
timestamp 1679235063
transform 1 0 5704 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold166
timestamp 1679235063
transform 1 0 1840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold167
timestamp 1679235063
transform 1 0 30636 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold168
timestamp 1679235063
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold169
timestamp 1679235063
transform 1 0 2760 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold170
timestamp 1679235063
transform 1 0 13064 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold171
timestamp 1679235063
transform 1 0 3036 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold172
timestamp 1679235063
transform 1 0 12144 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold173
timestamp 1679235063
transform 1 0 18860 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold174
timestamp 1679235063
transform 1 0 19412 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold175
timestamp 1679235063
transform 1 0 6532 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold176
timestamp 1679235063
transform 1 0 39652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold177
timestamp 1679235063
transform 1 0 11684 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold178
timestamp 1679235063
transform 1 0 43516 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold179
timestamp 1679235063
transform 1 0 23736 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold180
timestamp 1679235063
transform 1 0 27600 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold181
timestamp 1679235063
transform 1 0 39652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold182
timestamp 1679235063
transform 1 0 35788 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold183
timestamp 1679235063
transform 1 0 11960 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold184
timestamp 1679235063
transform 1 0 11960 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold185
timestamp 1679235063
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold186
timestamp 1679235063
transform 1 0 29808 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold187
timestamp 1679235063
transform 1 0 15180 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold188
timestamp 1679235063
transform 1 0 34500 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold189
timestamp 1679235063
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold190
timestamp 1679235063
transform 1 0 30452 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold191
timestamp 1679235063
transform 1 0 24564 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold192
timestamp 1679235063
transform 1 0 16836 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold193
timestamp 1679235063
transform 1 0 12328 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold194
timestamp 1679235063
transform 1 0 17940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold195
timestamp 1679235063
transform 1 0 9108 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold196
timestamp 1679235063
transform 1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold197
timestamp 1679235063
transform 1 0 4232 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold198
timestamp 1679235063
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold199
timestamp 1679235063
transform 1 0 15272 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold200
timestamp 1679235063
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold201
timestamp 1679235063
transform 1 0 6532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold202
timestamp 1679235063
transform 1 0 10856 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold203
timestamp 1679235063
transform 1 0 32292 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold204
timestamp 1679235063
transform 1 0 16008 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold205
timestamp 1679235063
transform 1 0 4140 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold206
timestamp 1679235063
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold207
timestamp 1679235063
transform 1 0 34868 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold208
timestamp 1679235063
transform 1 0 35972 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold209
timestamp 1679235063
transform 1 0 27140 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold210
timestamp 1679235063
transform 1 0 27140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold211
timestamp 1679235063
transform 1 0 38180 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold212
timestamp 1679235063
transform 1 0 41308 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold213
timestamp 1679235063
transform 1 0 4232 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold214
timestamp 1679235063
transform 1 0 1656 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold215
timestamp 1679235063
transform 1 0 20792 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold216
timestamp 1679235063
transform 1 0 22172 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold217
timestamp 1679235063
transform 1 0 34868 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold218
timestamp 1679235063
transform 1 0 33212 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold219
timestamp 1679235063
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold220
timestamp 1679235063
transform 1 0 7176 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold221
timestamp 1679235063
transform 1 0 31924 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold222
timestamp 1679235063
transform 1 0 16376 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold223
timestamp 1679235063
transform 1 0 33396 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold224
timestamp 1679235063
transform 1 0 32292 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold225
timestamp 1679235063
transform 1 0 9384 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold226
timestamp 1679235063
transform 1 0 2760 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold227
timestamp 1679235063
transform 1 0 7636 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold228
timestamp 1679235063
transform 1 0 5336 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold229
timestamp 1679235063
transform 1 0 35972 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold230
timestamp 1679235063
transform 1 0 35972 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold231
timestamp 1679235063
transform 1 0 19412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold232
timestamp 1679235063
transform 1 0 20608 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold233
timestamp 1679235063
transform 1 0 33396 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold234
timestamp 1679235063
transform 1 0 32292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold235
timestamp 1679235063
transform 1 0 9568 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold236
timestamp 1679235063
transform 1 0 10580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold237
timestamp 1679235063
transform 1 0 33396 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold238
timestamp 1679235063
transform 1 0 33396 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold239
timestamp 1679235063
transform 1 0 30544 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold240
timestamp 1679235063
transform 1 0 30912 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold241
timestamp 1679235063
transform 1 0 40020 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold242
timestamp 1679235063
transform 1 0 38548 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold243
timestamp 1679235063
transform 1 0 13432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold244
timestamp 1679235063
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold245
timestamp 1679235063
transform 1 0 27140 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold246
timestamp 1679235063
transform 1 0 25668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold247
timestamp 1679235063
transform 1 0 32292 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold248
timestamp 1679235063
transform 1 0 31004 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold249
timestamp 1679235063
transform 1 0 6808 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold250
timestamp 1679235063
transform 1 0 3128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold251
timestamp 1679235063
transform 1 0 30820 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold252
timestamp 1679235063
transform 1 0 28060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold253
timestamp 1679235063
transform 1 0 40756 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold254
timestamp 1679235063
transform 1 0 42228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold255
timestamp 1679235063
transform 1 0 37444 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold256
timestamp 1679235063
transform 1 0 37444 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold257
timestamp 1679235063
transform 1 0 34868 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold258
timestamp 1679235063
transform 1 0 33488 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold259
timestamp 1679235063
transform 1 0 6532 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold260
timestamp 1679235063
transform 1 0 1656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold261
timestamp 1679235063
transform 1 0 22172 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold262
timestamp 1679235063
transform 1 0 21988 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold263
timestamp 1679235063
transform 1 0 9384 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold264
timestamp 1679235063
transform 1 0 9752 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold265
timestamp 1679235063
transform 1 0 3404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold266
timestamp 1679235063
transform 1 0 40756 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold267
timestamp 1679235063
transform 1 0 36156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold268
timestamp 1679235063
transform 1 0 28244 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold269
timestamp 1679235063
transform 1 0 16928 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold270
timestamp 1679235063
transform 1 0 6532 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold271
timestamp 1679235063
transform 1 0 40940 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold272
timestamp 1679235063
transform 1 0 42596 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold273
timestamp 1679235063
transform 1 0 34868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold274
timestamp 1679235063
transform 1 0 34868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold275
timestamp 1679235063
transform 1 0 33396 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold276
timestamp 1679235063
transform 1 0 35972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold277
timestamp 1679235063
transform 1 0 30084 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold278
timestamp 1679235063
transform 1 0 28244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold279
timestamp 1679235063
transform 1 0 25668 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold280
timestamp 1679235063
transform 1 0 28796 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold281
timestamp 1679235063
transform 1 0 18216 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold282
timestamp 1679235063
transform 1 0 29716 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold283
timestamp 1679235063
transform 1 0 34868 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold284
timestamp 1679235063
transform 1 0 33396 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold285
timestamp 1679235063
transform 1 0 2024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold286
timestamp 1679235063
transform 1 0 38548 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold287
timestamp 1679235063
transform 1 0 23184 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold288
timestamp 1679235063
transform 1 0 43884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold289
timestamp 1679235063
transform 1 0 33396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold290
timestamp 1679235063
transform 1 0 29716 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold291
timestamp 1679235063
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold292
timestamp 1679235063
transform 1 0 4600 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold293
timestamp 1679235063
transform 1 0 31464 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold294
timestamp 1679235063
transform 1 0 22080 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold295
timestamp 1679235063
transform 1 0 6808 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold296
timestamp 1679235063
transform 1 0 24564 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold297
timestamp 1679235063
transform 1 0 25668 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold298
timestamp 1679235063
transform 1 0 19504 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold299
timestamp 1679235063
transform 1 0 4232 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold300
timestamp 1679235063
transform 1 0 3036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold301
timestamp 1679235063
transform 1 0 25392 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold302
timestamp 1679235063
transform 1 0 27140 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold303
timestamp 1679235063
transform 1 0 17848 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold304
timestamp 1679235063
transform 1 0 30912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold305
timestamp 1679235063
transform 1 0 35788 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold306
timestamp 1679235063
transform 1 0 15640 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold307
timestamp 1679235063
transform 1 0 23460 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold308
timestamp 1679235063
transform 1 0 20884 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold309
timestamp 1679235063
transform 1 0 43700 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold310
timestamp 1679235063
transform 1 0 1656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold311
timestamp 1679235063
transform 1 0 5152 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold312
timestamp 1679235063
transform 1 0 1932 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold313
timestamp 1679235063
transform 1 0 39836 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold314
timestamp 1679235063
transform 1 0 6716 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold315
timestamp 1679235063
transform 1 0 5704 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  hold316
timestamp 1679235063
transform 1 0 31280 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold317
timestamp 1679235063
transform 1 0 4600 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold318
timestamp 1679235063
transform 1 0 3956 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold319
timestamp 1679235063
transform 1 0 1656 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold320
timestamp 1679235063
transform 1 0 3496 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold321
timestamp 1679235063
transform 1 0 2760 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold322
timestamp 1679235063
transform 1 0 48668 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold323
timestamp 1679235063
transform 1 0 46552 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold324
timestamp 1679235063
transform 1 0 48668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold325
timestamp 1679235063
transform 1 0 46460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold326
timestamp 1679235063
transform 1 0 47748 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1679235063
transform 1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1679235063
transform 1 0 47012 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1679235063
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1679235063
transform 1 0 1564 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1679235063
transform 1 0 1564 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1679235063
transform 1 0 13340 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1679235063
transform 1 0 21988 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1679235063
transform 1 0 21344 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1679235063
transform 1 0 17572 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1679235063
transform 1 0 15456 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1679235063
transform 1 0 18400 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1679235063
transform 1 0 20700 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1679235063
transform 1 0 20976 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1679235063
transform 1 0 19412 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1679235063
transform 1 0 19688 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1679235063
transform 1 0 16284 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1679235063
transform 1 0 26956 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1679235063
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1679235063
transform 1 0 19412 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1679235063
transform 1 0 28612 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1679235063
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1679235063
transform 1 0 16928 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1679235063
transform 1 0 16008 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1679235063
transform 1 0 1564 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1679235063
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1679235063
transform 1 0 1564 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1679235063
transform 1 0 18216 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1679235063
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1679235063
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1679235063
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1679235063
transform 1 0 1564 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1679235063
transform 1 0 1564 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1679235063
transform 1 0 2760 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1679235063
transform 1 0 42596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1679235063
transform 1 0 29716 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1679235063
transform 1 0 34868 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1679235063
transform 1 0 33580 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1679235063
transform 1 0 44436 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1679235063
transform 1 0 43976 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1679235063
transform 1 0 44712 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1679235063
transform 1 0 31464 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1679235063
transform 1 0 48852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1679235063
transform 1 0 38548 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1679235063
transform 1 0 29992 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input45
timestamp 1679235063
transform 1 0 44988 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1679235063
transform 1 0 39284 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1679235063
transform 1 0 44068 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1679235063
transform 1 0 38916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1679235063
transform 1 0 39468 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1679235063
transform 1 0 38732 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1679235063
transform 1 0 40572 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1679235063
transform 1 0 41216 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1679235063
transform 1 0 41492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1679235063
transform 1 0 43332 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1679235063
transform 1 0 30268 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1679235063
transform 1 0 37444 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1679235063
transform 1 0 31924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1679235063
transform 1 0 14260 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1679235063
transform 1 0 31556 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1679235063
transform 1 0 37076 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1679235063
transform 1 0 37352 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1679235063
transform 1 0 45908 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1679235063
transform 1 0 25484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1679235063
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1679235063
transform 1 0 30820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1679235063
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1679235063
transform 1 0 36064 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1679235063
transform 1 0 41216 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1679235063
transform 1 0 45724 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input70
timestamp 1679235063
transform 1 0 46460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1679235063
transform 1 0 47196 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1679235063
transform 1 0 48852 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1679235063
transform 1 0 47748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input74
timestamp 1679235063
transform 1 0 47932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input75
timestamp 1679235063
transform 1 0 45908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1679235063
transform 1 0 45172 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  output77 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1679235063
transform 1 0 6532 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1679235063
transform 1 0 1564 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1679235063
transform 1 0 1564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1679235063
transform 1 0 1564 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1679235063
transform 1 0 1564 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1679235063
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1679235063
transform 1 0 1564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1679235063
transform 1 0 1564 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1679235063
transform 1 0 1564 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1679235063
transform 1 0 3956 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1679235063
transform 1 0 1564 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1679235063
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1679235063
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1679235063
transform 1 0 3956 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1679235063
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1679235063
transform 1 0 3956 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1679235063
transform 1 0 3404 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1679235063
transform 1 0 5796 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1679235063
transform 1 0 3404 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1679235063
transform 1 0 3956 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1679235063
transform 1 0 6532 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1679235063
transform 1 0 3404 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1679235063
transform 1 0 9108 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1679235063
transform 1 0 1564 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1679235063
transform 1 0 1564 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output103
timestamp 1679235063
transform 1 0 1564 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output104
timestamp 1679235063
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output105
timestamp 1679235063
transform 1 0 1564 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output106
timestamp 1679235063
transform 1 0 1564 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output107
timestamp 1679235063
transform 1 0 1564 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output108
timestamp 1679235063
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output109
timestamp 1679235063
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output110
timestamp 1679235063
transform 1 0 7176 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output111
timestamp 1679235063
transform 1 0 7912 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output112
timestamp 1679235063
transform 1 0 9292 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output113
timestamp 1679235063
transform 1 0 10488 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output114
timestamp 1679235063
transform 1 0 11960 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output115
timestamp 1679235063
transform 1 0 9752 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output116
timestamp 1679235063
transform 1 0 12328 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output117
timestamp 1679235063
transform 1 0 9752 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output118
timestamp 1679235063
transform 1 0 12328 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output119
timestamp 1679235063
transform 1 0 15180 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1679235063
transform 1 0 2024 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1679235063
transform 1 0 13064 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1679235063
transform 1 0 14904 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1679235063
transform 1 0 16836 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1679235063
transform 1 0 15272 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1679235063
transform 1 0 14904 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1679235063
transform 1 0 14904 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1679235063
transform 1 0 16928 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1679235063
transform 1 0 20332 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1679235063
transform 1 0 20056 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1679235063
transform 1 0 21988 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1679235063
transform 1 0 2760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1679235063
transform 1 0 4600 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1679235063
transform 1 0 4600 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1679235063
transform 1 0 5336 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1679235063
transform 1 0 6808 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1679235063
transform 1 0 4600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1679235063
transform 1 0 7176 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1679235063
transform 1 0 7360 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1679235063
transform 1 0 4140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1679235063
transform 1 0 6808 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1679235063
transform 1 0 9476 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1679235063
transform 1 0 12144 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1679235063
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1679235063
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1679235063
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1679235063
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1679235063
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1679235063
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1679235063
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1679235063
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1679235063
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1679235063
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1679235063
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1679235063
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1679235063
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1679235063
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1679235063
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1679235063
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1679235063
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1679235063
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1679235063
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1679235063
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1679235063
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1679235063
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1679235063
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1679235063
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1679235063
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1679235063
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1679235063
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1679235063
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1679235063
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1679235063
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1679235063
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1679235063
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1679235063
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1679235063
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1679235063
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1679235063
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1679235063
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1679235063
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1679235063
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1679235063
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1679235063
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1679235063
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1679235063
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1679235063
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1679235063
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1679235063
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1679235063
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1679235063
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1679235063
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1679235063
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1679235063
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1679235063
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1679235063
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1679235063
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1679235063
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1679235063
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1679235063
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1679235063
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1679235063
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1679235063
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1679235063
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1679235063
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1679235063
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1679235063
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1679235063
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1679235063
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1679235063
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1679235063
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1679235063
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1679235063
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1679235063
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1679235063
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1679235063
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1679235063
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1679235063
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1679235063
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1679235063
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1679235063
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1679235063
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1679235063
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1679235063
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1679235063
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22080 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 18676 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19412 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20240 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 21068 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_9.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_left_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16836 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_left_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 18768 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 19688 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_15.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20056 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 21988 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_17.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22264 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 23092 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_19.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 23368 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24380 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25484 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25852 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_31.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 25944 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 25760 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_33.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24840 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27140 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_35.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27324 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28428 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28428 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_47.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28428 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 28336 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_49.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 28060 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 27048 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_left_track_51.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 24656 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 37720 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 27876 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 24840 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 24840 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22448 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19504 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20976 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 19688 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 18216 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 20240 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20976 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 22908 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 19688 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 22264 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 20056 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1679235063
transform 1 0 17112 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17480 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16652 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14444 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14444 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14628 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16100 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17112 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 17112 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 16928 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 16836 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14720 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14628 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14260 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 13156 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12236 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11500 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11684 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11500 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11776 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 11592 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11684 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 10856 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 10028 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 8648 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 6808 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6532 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 4600 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 6164 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 7728 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_42.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 9200 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 11132 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 12236 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 12880 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 13524 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 14352 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 14720 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1679235063
transform 1 0 15824 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_8__0_.mem_top_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1679235063
transform 1 0 17848 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_0_
timestamp 1679235063
transform 1 0 31188 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l1_in_1_
timestamp 1679235063
transform 1 0 27416 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_1.mux_l1_in_1__196
timestamp 1679235063
transform 1 0 27232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_1.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l1_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_3.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_3.mux_l2_in_0__155
timestamp 1679235063
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5704 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_5.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17112 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_5.mux_l2_in_0__162
timestamp 1679235063
transform 1 0 23276 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24564 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_7.mux_l1_in_1__164
timestamp 1679235063
transform 1 0 16928 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_7.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15732 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_9.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_9.mux_l2_in_0__165
timestamp 1679235063
transform 1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 27876 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_11.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11868 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_11.mux_l2_in_0__197
timestamp 1679235063
transform 1 0 41860 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 10672 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_13.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14536 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_13.mux_l2_in_0__198
timestamp 1679235063
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28336 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_15.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_15.mux_l2_in_0__199
timestamp 1679235063
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25760 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_17.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18492 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_17.mux_l2_in_0__200
timestamp 1679235063
transform 1 0 8372 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29348 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l1_in_0_
timestamp 1679235063
transform 1 0 25300 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_19.mux_l2_in_0__153
timestamp 1679235063
transform 1 0 19412 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_19.mux_l2_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_29.mux_l2_in_0__154
timestamp 1679235063
transform 1 0 19044 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_29.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22816 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27232 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_31.mux_l2_in_0__156
timestamp 1679235063
transform 1 0 6532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_31.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23000 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l1_in_0_
timestamp 1679235063
transform 1 0 27232 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_33.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21804 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_33.mux_l2_in_0__157
timestamp 1679235063
transform 1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 34868 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_35.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_35.mux_l2_in_0__158
timestamp 1679235063
transform 1 0 23828 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_45.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_45.mux_l2_in_0__159
timestamp 1679235063
transform 1 0 24196 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  sb_8__0_.mux_left_track_45.mux_l2_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 25576 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_47.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24656 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_47.mux_l2_in_0__160
timestamp 1679235063
transform 1 0 27692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l1_in_0_
timestamp 1679235063
transform 1 0 30636 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_49.mux_l2_in_0__161
timestamp 1679235063
transform 1 0 27140 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_49.mux_l2_in_0_
timestamp 1679235063
transform 1 0 25944 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 16836 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l1_in_0_
timestamp 1679235063
transform 1 0 29716 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_left_track_51.mux_l2_in_0__163
timestamp 1679235063
transform 1 0 21436 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_left_track_51.mux_l2_in_0_
timestamp 1679235063
transform 1 0 22080 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_0_
timestamp 1679235063
transform 1 0 28428 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l1_in_1_
timestamp 1679235063
transform 1 0 29716 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_0_
timestamp 1679235063
transform 1 0 27140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l2_in_1_
timestamp 1679235063
transform 1 0 20056 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_0.mux_l2_in_1__166
timestamp 1679235063
transform 1 0 19596 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_0.mux_l3_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 23828 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_0_
timestamp 1679235063
transform 1 0 26404 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25116 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_0_
timestamp 1679235063
transform 1 0 24564 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l2_in_1_
timestamp 1679235063
transform 1 0 13156 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_2.mux_l2_in_1__172
timestamp 1679235063
transform 1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_2.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19412 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_0_
timestamp 1679235063
transform 1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l1_in_1_
timestamp 1679235063
transform 1 0 21344 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l2_in_1_
timestamp 1679235063
transform 1 0 11960 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_4.mux_l2_in_1__183
timestamp 1679235063
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_4.mux_l3_in_0_
timestamp 1679235063
transform 1 0 16928 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 9108 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23736 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23460 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_0_
timestamp 1679235063
transform 1 0 21988 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15456 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_6.mux_l2_in_1__190
timestamp 1679235063
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_6.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19320 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_0_
timestamp 1679235063
transform 1 0 24748 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l1_in_1_
timestamp 1679235063
transform 1 0 25208 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_0_
timestamp 1679235063
transform 1 0 20700 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l2_in_1_
timestamp 1679235063
transform 1 0 15548 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_8.mux_l2_in_1__191
timestamp 1679235063
transform 1 0 14628 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_8.mux_l3_in_0_
timestamp 1679235063
transform 1 0 19504 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 19412 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_0_
timestamp 1679235063
transform 1 0 23276 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l1_in_1_
timestamp 1679235063
transform 1 0 23828 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_0_
timestamp 1679235063
transform 1 0 23184 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l2_in_1_
timestamp 1679235063
transform 1 0 14260 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_10.mux_l2_in_1__167
timestamp 1679235063
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_10.mux_l3_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 14352 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19504 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l1_in_1_
timestamp 1679235063
transform 1 0 14352 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_12.mux_l1_in_1__168
timestamp 1679235063
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_12.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17204 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_14.mux_l1_in_1__169
timestamp 1679235063
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_14.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12972 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 3956 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18124 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_16.mux_l1_in_1__170
timestamp 1679235063
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_16.mux_l2_in_0_
timestamp 1679235063
transform 1 0 13156 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 29624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20516 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l1_in_1_
timestamp 1679235063
transform 1 0 13892 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_18.mux_l1_in_1__171
timestamp 1679235063
transform 1 0 6532 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_18.mux_l2_in_0_
timestamp 1679235063
transform 1 0 17112 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_20.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15548 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_20.mux_l2_in_0__173
timestamp 1679235063
transform 1 0 26312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 18400 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l1_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_22.mux_l2_in_0__174
timestamp 1679235063
transform 1 0 3956 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_22.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14352 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 28612 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l1_in_0_
timestamp 1679235063
transform 1 0 15180 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_24.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14444 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_24.mux_l2_in_0__175
timestamp 1679235063
transform 1 0 3956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 24748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_26.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11776 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_26.mux_l2_in_0__176
timestamp 1679235063
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l1_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_28.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10580 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_28.mux_l2_in_0__177
timestamp 1679235063
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 5704 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_30.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11960 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_30.mux_l2_in_0__178
timestamp 1679235063
transform 1 0 9108 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_32.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  sb_8__0_.mux_top_track_32.mux_l2_in_0_
timestamp 1679235063
transform 1 0 11684 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_32.mux_l2_in_0__179
timestamp 1679235063
transform 1 0 13524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 39284 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12236 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_34.mux_l2_in_0_
timestamp 1679235063
transform 1 0 10396 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_34.mux_l2_in_0__180
timestamp 1679235063
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l1_in_0_
timestamp 1679235063
transform 1 0 12880 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_36.mux_l2_in_0_
timestamp 1679235063
transform 1 0 9292 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_36.mux_l2_in_0__181
timestamp 1679235063
transform 1 0 6532 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_38.mux_l2_in_0_
timestamp 1679235063
transform 1 0 5244 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_38.mux_l2_in_0__182
timestamp 1679235063
transform 1 0 20700 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21988 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l1_in_0_
timestamp 1679235063
transform 1 0 7636 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_40.mux_l2_in_0_
timestamp 1679235063
transform 1 0 15456 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_40.mux_l2_in_0__184
timestamp 1679235063
transform 1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l1_in_0_
timestamp 1679235063
transform 1 0 11684 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_42.mux_l2_in_0_
timestamp 1679235063
transform 1 0 6532 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_42.mux_l2_in_0__185
timestamp 1679235063
transform 1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_0_
timestamp 1679235063
transform 1 0 17572 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l1_in_1_
timestamp 1679235063
transform 1 0 9200 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_44.mux_l1_in_1__186
timestamp 1679235063
transform 1 0 20700 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_44.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14260 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 35972 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_0_
timestamp 1679235063
transform 1 0 18032 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l1_in_1_
timestamp 1679235063
transform 1 0 10304 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_46.mux_l1_in_1__187
timestamp 1679235063
transform 1 0 28244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_46.mux_l2_in_0_
timestamp 1679235063
transform 1 0 12328 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 37444 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_0_
timestamp 1679235063
transform 1 0 19136 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l1_in_1_
timestamp 1679235063
transform 1 0 11776 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_48.mux_l1_in_1__188
timestamp 1679235063
transform 1 0 3956 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_48.mux_l2_in_0_
timestamp 1679235063
transform 1 0 14812 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 41860 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_0_
timestamp 1679235063
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l1_in_1_
timestamp 1679235063
transform 1 0 12972 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_8__0_.mux_top_track_50.mux_l1_in_1__189
timestamp 1679235063
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_8__0_.mux_top_track_50.mux_l2_in_0_
timestamp 1679235063
transform 1 0 16836 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1679235063
transform 1 0 42596 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1679235063
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1679235063
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1679235063
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1679235063
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1679235063
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1679235063
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1679235063
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1679235063
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1679235063
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1679235063
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1679235063
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1679235063
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1679235063
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1679235063
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1679235063
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1679235063
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1679235063
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1679235063
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1679235063
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1679235063
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1679235063
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1679235063
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1679235063
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1679235063
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1679235063
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1679235063
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1679235063
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1679235063
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1679235063
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1679235063
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1679235063
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1679235063
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1679235063
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1679235063
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1679235063
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1679235063
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1679235063
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1679235063
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1679235063
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1679235063
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1679235063
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1679235063
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1679235063
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1679235063
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1679235063
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1679235063
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1679235063
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1679235063
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1679235063
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1679235063
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1679235063
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1679235063
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1679235063
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1679235063
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1679235063
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1679235063
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1679235063
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1679235063
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1679235063
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1679235063
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1679235063
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1679235063
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1679235063
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1679235063
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1679235063
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1679235063
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1679235063
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1679235063
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1679235063
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1679235063
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1679235063
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1679235063
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1679235063
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1679235063
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1679235063
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1679235063
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1679235063
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1679235063
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1679235063
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1679235063
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1679235063
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1679235063
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1679235063
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1679235063
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1679235063
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1679235063
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1679235063
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1679235063
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1679235063
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1679235063
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1679235063
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1679235063
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1679235063
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1679235063
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1679235063
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1679235063
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1679235063
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1679235063
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1679235063
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1679235063
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1679235063
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1679235063
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1679235063
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1679235063
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1679235063
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1679235063
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1679235063
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1679235063
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1679235063
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1679235063
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1679235063
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1679235063
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1679235063
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1679235063
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1679235063
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1679235063
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1679235063
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1679235063
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1679235063
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1679235063
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1679235063
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1679235063
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1679235063
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1679235063
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1679235063
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1679235063
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1679235063
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1679235063
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1679235063
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1679235063
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1679235063
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1679235063
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1679235063
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1679235063
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1679235063
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1679235063
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1679235063
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1679235063
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1679235063
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1679235063
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1679235063
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1679235063
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1679235063
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1679235063
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1679235063
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1679235063
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1679235063
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1679235063
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1679235063
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1679235063
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1679235063
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1679235063
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1679235063
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1679235063
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1679235063
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1679235063
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1679235063
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1679235063
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1679235063
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1679235063
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1679235063
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1679235063
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1679235063
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1679235063
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1679235063
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1679235063
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1679235063
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1679235063
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1679235063
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1679235063
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1679235063
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1679235063
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1679235063
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1679235063
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1679235063
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1679235063
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1679235063
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1679235063
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1679235063
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1679235063
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1679235063
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1679235063
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1679235063
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1679235063
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1679235063
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1679235063
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1679235063
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1679235063
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1679235063
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1679235063
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1679235063
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1679235063
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1679235063
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1679235063
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1679235063
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1679235063
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1679235063
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1679235063
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1679235063
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1679235063
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1679235063
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1679235063
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1679235063
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1679235063
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1679235063
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1679235063
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1679235063
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1679235063
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1679235063
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1679235063
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1679235063
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1679235063
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1679235063
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1679235063
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1679235063
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1679235063
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1679235063
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1679235063
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1679235063
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1679235063
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1679235063
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1679235063
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1679235063
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1679235063
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1679235063
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1679235063
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1679235063
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1679235063
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1679235063
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1679235063
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1679235063
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1679235063
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1679235063
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1679235063
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1679235063
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1679235063
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1679235063
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1679235063
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1679235063
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1679235063
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1679235063
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1679235063
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1679235063
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1679235063
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1679235063
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1679235063
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1679235063
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1679235063
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1679235063
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1679235063
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1679235063
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1679235063
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1679235063
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1679235063
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1679235063
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1679235063
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1679235063
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1679235063
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1679235063
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1679235063
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1679235063
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1679235063
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1679235063
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1679235063
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1679235063
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1679235063
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1679235063
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1679235063
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1679235063
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1679235063
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1679235063
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1679235063
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1679235063
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1679235063
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1679235063
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1679235063
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1679235063
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1679235063
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1679235063
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1679235063
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1679235063
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1679235063
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1679235063
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1679235063
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1679235063
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1679235063
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1679235063
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1679235063
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1679235063
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1679235063
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1679235063
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1679235063
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1679235063
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1679235063
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1679235063
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1679235063
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1679235063
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1679235063
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1679235063
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1679235063
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1679235063
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1679235063
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1679235063
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1679235063
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1679235063
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1679235063
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1679235063
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1679235063
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1679235063
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1679235063
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1679235063
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1679235063
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1679235063
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1679235063
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1679235063
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1679235063
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1679235063
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1679235063
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1679235063
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1679235063
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1679235063
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1679235063
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1679235063
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1679235063
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1679235063
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1679235063
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1679235063
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1679235063
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1679235063
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1679235063
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1679235063
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1679235063
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1679235063
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1679235063
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1679235063
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1679235063
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1679235063
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1679235063
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1679235063
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1679235063
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1679235063
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1679235063
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1679235063
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1679235063
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1679235063
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1679235063
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1679235063
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1679235063
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1679235063
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1679235063
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1679235063
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1679235063
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1679235063
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1679235063
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1679235063
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1679235063
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1679235063
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1679235063
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1679235063
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1679235063
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1679235063
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1679235063
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1679235063
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1679235063
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1679235063
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1679235063
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1679235063
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1679235063
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1679235063
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1679235063
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1679235063
transform 1 0 6256 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1679235063
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1679235063
transform 1 0 11408 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1679235063
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1679235063
transform 1 0 16560 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1679235063
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1679235063
transform 1 0 21712 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1679235063
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1679235063
transform 1 0 26864 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1679235063
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1679235063
transform 1 0 32016 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1679235063
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1679235063
transform 1 0 37168 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1679235063
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1679235063
transform 1 0 42320 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1679235063
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1679235063
transform 1 0 47472 0 1 23936
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 24528 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 24528 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 1398 0 1454 800 0 FreeSans 224 90 0 0 ccff_head
port 2 nsew signal input
flabel metal2 s 48594 26200 48650 27000 0 FreeSans 224 90 0 0 ccff_head_1
port 3 nsew signal input
flabel metal3 s 50200 20952 51000 21072 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 2226 26200 2282 27000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 0 1504 800 1624 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 6 nsew signal input
flabel metal3 s 0 5584 800 5704 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 7 nsew signal input
flabel metal3 s 0 5992 800 6112 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 8 nsew signal input
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 9 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 10 nsew signal input
flabel metal3 s 0 7216 800 7336 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 11 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 12 nsew signal input
flabel metal3 s 0 8032 800 8152 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 13 nsew signal input
flabel metal3 s 0 8440 800 8560 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 14 nsew signal input
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 15 nsew signal input
flabel metal3 s 0 9256 800 9376 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 16 nsew signal input
flabel metal3 s 0 1912 800 2032 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 17 nsew signal input
flabel metal3 s 0 9664 800 9784 0 FreeSans 480 0 0 0 chanx_left_in[20]
port 18 nsew signal input
flabel metal3 s 0 10072 800 10192 0 FreeSans 480 0 0 0 chanx_left_in[21]
port 19 nsew signal input
flabel metal3 s 0 10480 800 10600 0 FreeSans 480 0 0 0 chanx_left_in[22]
port 20 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 chanx_left_in[23]
port 21 nsew signal input
flabel metal3 s 0 11296 800 11416 0 FreeSans 480 0 0 0 chanx_left_in[24]
port 22 nsew signal input
flabel metal3 s 0 11704 800 11824 0 FreeSans 480 0 0 0 chanx_left_in[25]
port 23 nsew signal input
flabel metal3 s 0 12112 800 12232 0 FreeSans 480 0 0 0 chanx_left_in[26]
port 24 nsew signal input
flabel metal3 s 0 12520 800 12640 0 FreeSans 480 0 0 0 chanx_left_in[27]
port 25 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 chanx_left_in[28]
port 26 nsew signal input
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 chanx_left_in[29]
port 27 nsew signal input
flabel metal3 s 0 2320 800 2440 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 28 nsew signal input
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 29 nsew signal input
flabel metal3 s 0 3136 800 3256 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 30 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 31 nsew signal input
flabel metal3 s 0 3952 800 4072 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 32 nsew signal input
flabel metal3 s 0 4360 800 4480 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 33 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 34 nsew signal input
flabel metal3 s 0 5176 800 5296 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 35 nsew signal input
flabel metal3 s 0 13744 800 13864 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 36 nsew signal tristate
flabel metal3 s 0 17824 800 17944 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 37 nsew signal tristate
flabel metal3 s 0 18232 800 18352 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 38 nsew signal tristate
flabel metal3 s 0 18640 800 18760 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 39 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 40 nsew signal tristate
flabel metal3 s 0 19456 800 19576 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 41 nsew signal tristate
flabel metal3 s 0 19864 800 19984 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 42 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 43 nsew signal tristate
flabel metal3 s 0 20680 800 20800 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 44 nsew signal tristate
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 45 nsew signal tristate
flabel metal3 s 0 21496 800 21616 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 46 nsew signal tristate
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 47 nsew signal tristate
flabel metal3 s 0 21904 800 22024 0 FreeSans 480 0 0 0 chanx_left_out[20]
port 48 nsew signal tristate
flabel metal3 s 0 22312 800 22432 0 FreeSans 480 0 0 0 chanx_left_out[21]
port 49 nsew signal tristate
flabel metal3 s 0 22720 800 22840 0 FreeSans 480 0 0 0 chanx_left_out[22]
port 50 nsew signal tristate
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 chanx_left_out[23]
port 51 nsew signal tristate
flabel metal3 s 0 23536 800 23656 0 FreeSans 480 0 0 0 chanx_left_out[24]
port 52 nsew signal tristate
flabel metal3 s 0 23944 800 24064 0 FreeSans 480 0 0 0 chanx_left_out[25]
port 53 nsew signal tristate
flabel metal3 s 0 24352 800 24472 0 FreeSans 480 0 0 0 chanx_left_out[26]
port 54 nsew signal tristate
flabel metal3 s 0 24760 800 24880 0 FreeSans 480 0 0 0 chanx_left_out[27]
port 55 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 chanx_left_out[28]
port 56 nsew signal tristate
flabel metal3 s 0 25576 800 25696 0 FreeSans 480 0 0 0 chanx_left_out[29]
port 57 nsew signal tristate
flabel metal3 s 0 14560 800 14680 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 58 nsew signal tristate
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 59 nsew signal tristate
flabel metal3 s 0 15376 800 15496 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 60 nsew signal tristate
flabel metal3 s 0 15784 800 15904 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 61 nsew signal tristate
flabel metal3 s 0 16192 800 16312 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 62 nsew signal tristate
flabel metal3 s 0 16600 800 16720 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 63 nsew signal tristate
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 64 nsew signal tristate
flabel metal3 s 0 17416 800 17536 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 65 nsew signal tristate
flabel metal2 s 22190 26200 22246 27000 0 FreeSans 224 90 0 0 chany_top_in[0]
port 66 nsew signal input
flabel metal2 s 28630 26200 28686 27000 0 FreeSans 224 90 0 0 chany_top_in[10]
port 67 nsew signal input
flabel metal2 s 29274 26200 29330 27000 0 FreeSans 224 90 0 0 chany_top_in[11]
port 68 nsew signal input
flabel metal2 s 29918 26200 29974 27000 0 FreeSans 224 90 0 0 chany_top_in[12]
port 69 nsew signal input
flabel metal2 s 30562 26200 30618 27000 0 FreeSans 224 90 0 0 chany_top_in[13]
port 70 nsew signal input
flabel metal2 s 31206 26200 31262 27000 0 FreeSans 224 90 0 0 chany_top_in[14]
port 71 nsew signal input
flabel metal2 s 31850 26200 31906 27000 0 FreeSans 224 90 0 0 chany_top_in[15]
port 72 nsew signal input
flabel metal2 s 32494 26200 32550 27000 0 FreeSans 224 90 0 0 chany_top_in[16]
port 73 nsew signal input
flabel metal2 s 33138 26200 33194 27000 0 FreeSans 224 90 0 0 chany_top_in[17]
port 74 nsew signal input
flabel metal2 s 33782 26200 33838 27000 0 FreeSans 224 90 0 0 chany_top_in[18]
port 75 nsew signal input
flabel metal2 s 34426 26200 34482 27000 0 FreeSans 224 90 0 0 chany_top_in[19]
port 76 nsew signal input
flabel metal2 s 22834 26200 22890 27000 0 FreeSans 224 90 0 0 chany_top_in[1]
port 77 nsew signal input
flabel metal2 s 35070 26200 35126 27000 0 FreeSans 224 90 0 0 chany_top_in[20]
port 78 nsew signal input
flabel metal2 s 35714 26200 35770 27000 0 FreeSans 224 90 0 0 chany_top_in[21]
port 79 nsew signal input
flabel metal2 s 36358 26200 36414 27000 0 FreeSans 224 90 0 0 chany_top_in[22]
port 80 nsew signal input
flabel metal2 s 37002 26200 37058 27000 0 FreeSans 224 90 0 0 chany_top_in[23]
port 81 nsew signal input
flabel metal2 s 37646 26200 37702 27000 0 FreeSans 224 90 0 0 chany_top_in[24]
port 82 nsew signal input
flabel metal2 s 38290 26200 38346 27000 0 FreeSans 224 90 0 0 chany_top_in[25]
port 83 nsew signal input
flabel metal2 s 38934 26200 38990 27000 0 FreeSans 224 90 0 0 chany_top_in[26]
port 84 nsew signal input
flabel metal2 s 39578 26200 39634 27000 0 FreeSans 224 90 0 0 chany_top_in[27]
port 85 nsew signal input
flabel metal2 s 40222 26200 40278 27000 0 FreeSans 224 90 0 0 chany_top_in[28]
port 86 nsew signal input
flabel metal2 s 40866 26200 40922 27000 0 FreeSans 224 90 0 0 chany_top_in[29]
port 87 nsew signal input
flabel metal2 s 23478 26200 23534 27000 0 FreeSans 224 90 0 0 chany_top_in[2]
port 88 nsew signal input
flabel metal2 s 24122 26200 24178 27000 0 FreeSans 224 90 0 0 chany_top_in[3]
port 89 nsew signal input
flabel metal2 s 24766 26200 24822 27000 0 FreeSans 224 90 0 0 chany_top_in[4]
port 90 nsew signal input
flabel metal2 s 25410 26200 25466 27000 0 FreeSans 224 90 0 0 chany_top_in[5]
port 91 nsew signal input
flabel metal2 s 26054 26200 26110 27000 0 FreeSans 224 90 0 0 chany_top_in[6]
port 92 nsew signal input
flabel metal2 s 26698 26200 26754 27000 0 FreeSans 224 90 0 0 chany_top_in[7]
port 93 nsew signal input
flabel metal2 s 27342 26200 27398 27000 0 FreeSans 224 90 0 0 chany_top_in[8]
port 94 nsew signal input
flabel metal2 s 27986 26200 28042 27000 0 FreeSans 224 90 0 0 chany_top_in[9]
port 95 nsew signal input
flabel metal2 s 2870 26200 2926 27000 0 FreeSans 224 90 0 0 chany_top_out[0]
port 96 nsew signal tristate
flabel metal2 s 9310 26200 9366 27000 0 FreeSans 224 90 0 0 chany_top_out[10]
port 97 nsew signal tristate
flabel metal2 s 9954 26200 10010 27000 0 FreeSans 224 90 0 0 chany_top_out[11]
port 98 nsew signal tristate
flabel metal2 s 10598 26200 10654 27000 0 FreeSans 224 90 0 0 chany_top_out[12]
port 99 nsew signal tristate
flabel metal2 s 11242 26200 11298 27000 0 FreeSans 224 90 0 0 chany_top_out[13]
port 100 nsew signal tristate
flabel metal2 s 11886 26200 11942 27000 0 FreeSans 224 90 0 0 chany_top_out[14]
port 101 nsew signal tristate
flabel metal2 s 12530 26200 12586 27000 0 FreeSans 224 90 0 0 chany_top_out[15]
port 102 nsew signal tristate
flabel metal2 s 13174 26200 13230 27000 0 FreeSans 224 90 0 0 chany_top_out[16]
port 103 nsew signal tristate
flabel metal2 s 13818 26200 13874 27000 0 FreeSans 224 90 0 0 chany_top_out[17]
port 104 nsew signal tristate
flabel metal2 s 14462 26200 14518 27000 0 FreeSans 224 90 0 0 chany_top_out[18]
port 105 nsew signal tristate
flabel metal2 s 15106 26200 15162 27000 0 FreeSans 224 90 0 0 chany_top_out[19]
port 106 nsew signal tristate
flabel metal2 s 3514 26200 3570 27000 0 FreeSans 224 90 0 0 chany_top_out[1]
port 107 nsew signal tristate
flabel metal2 s 15750 26200 15806 27000 0 FreeSans 224 90 0 0 chany_top_out[20]
port 108 nsew signal tristate
flabel metal2 s 16394 26200 16450 27000 0 FreeSans 224 90 0 0 chany_top_out[21]
port 109 nsew signal tristate
flabel metal2 s 17038 26200 17094 27000 0 FreeSans 224 90 0 0 chany_top_out[22]
port 110 nsew signal tristate
flabel metal2 s 17682 26200 17738 27000 0 FreeSans 224 90 0 0 chany_top_out[23]
port 111 nsew signal tristate
flabel metal2 s 18326 26200 18382 27000 0 FreeSans 224 90 0 0 chany_top_out[24]
port 112 nsew signal tristate
flabel metal2 s 18970 26200 19026 27000 0 FreeSans 224 90 0 0 chany_top_out[25]
port 113 nsew signal tristate
flabel metal2 s 19614 26200 19670 27000 0 FreeSans 224 90 0 0 chany_top_out[26]
port 114 nsew signal tristate
flabel metal2 s 20258 26200 20314 27000 0 FreeSans 224 90 0 0 chany_top_out[27]
port 115 nsew signal tristate
flabel metal2 s 20902 26200 20958 27000 0 FreeSans 224 90 0 0 chany_top_out[28]
port 116 nsew signal tristate
flabel metal2 s 21546 26200 21602 27000 0 FreeSans 224 90 0 0 chany_top_out[29]
port 117 nsew signal tristate
flabel metal2 s 4158 26200 4214 27000 0 FreeSans 224 90 0 0 chany_top_out[2]
port 118 nsew signal tristate
flabel metal2 s 4802 26200 4858 27000 0 FreeSans 224 90 0 0 chany_top_out[3]
port 119 nsew signal tristate
flabel metal2 s 5446 26200 5502 27000 0 FreeSans 224 90 0 0 chany_top_out[4]
port 120 nsew signal tristate
flabel metal2 s 6090 26200 6146 27000 0 FreeSans 224 90 0 0 chany_top_out[5]
port 121 nsew signal tristate
flabel metal2 s 6734 26200 6790 27000 0 FreeSans 224 90 0 0 chany_top_out[6]
port 122 nsew signal tristate
flabel metal2 s 7378 26200 7434 27000 0 FreeSans 224 90 0 0 chany_top_out[7]
port 123 nsew signal tristate
flabel metal2 s 8022 26200 8078 27000 0 FreeSans 224 90 0 0 chany_top_out[8]
port 124 nsew signal tristate
flabel metal2 s 8666 26200 8722 27000 0 FreeSans 224 90 0 0 chany_top_out[9]
port 125 nsew signal tristate
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[0]
port 126 nsew signal tristate
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[1]
port 127 nsew signal tristate
flabel metal2 s 9402 0 9458 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[2]
port 128 nsew signal tristate
flabel metal2 s 12070 0 12126 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_dir[3]
port 129 nsew signal tristate
flabel metal2 s 25410 0 25466 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[0]
port 130 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[1]
port 131 nsew signal input
flabel metal2 s 30746 0 30802 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[2]
port 132 nsew signal input
flabel metal2 s 33414 0 33470 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_in[3]
port 133 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[0]
port 134 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[1]
port 135 nsew signal tristate
flabel metal2 s 20074 0 20130 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[2]
port 136 nsew signal tristate
flabel metal2 s 22742 0 22798 800 0 FreeSans 224 90 0 0 gfpga_pad_io_soc_out[3]
port 137 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 isol_n
port 138 nsew signal input
flabel metal2 s 38750 0 38806 800 0 FreeSans 224 90 0 0 prog_clk
port 139 nsew signal input
flabel metal2 s 41510 26200 41566 27000 0 FreeSans 224 90 0 0 prog_reset
port 140 nsew signal input
flabel metal2 s 42154 26200 42210 27000 0 FreeSans 224 90 0 0 reset
port 141 nsew signal input
flabel metal2 s 42798 26200 42854 27000 0 FreeSans 224 90 0 0 test_enable
port 142 nsew signal input
flabel metal2 s 44730 26200 44786 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
port 143 nsew signal input
flabel metal2 s 45374 26200 45430 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
port 144 nsew signal input
flabel metal2 s 46018 26200 46074 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
port 145 nsew signal input
flabel metal2 s 46662 26200 46718 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
port 146 nsew signal input
flabel metal2 s 47306 26200 47362 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
port 147 nsew signal input
flabel metal2 s 47950 26200 48006 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
port 148 nsew signal input
flabel metal2 s 43442 26200 43498 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
port 149 nsew signal input
flabel metal2 s 44086 26200 44142 27000 0 FreeSans 224 90 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
port 150 nsew signal input
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
port 151 nsew signal input
flabel metal3 s 50200 22856 51000 22976 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
port 152 nsew signal input
flabel metal3 s 50200 23808 51000 23928 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
port 153 nsew signal input
flabel metal3 s 50200 24760 51000 24880 0 FreeSans 480 0 0 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
port 154 nsew signal input
flabel metal2 s 41418 0 41474 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_0__pin_inpad_0_
port 155 nsew signal tristate
flabel metal2 s 44086 0 44142 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_1__pin_inpad_0_
port 156 nsew signal tristate
flabel metal2 s 46754 0 46810 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_2__pin_inpad_0_
port 157 nsew signal tristate
flabel metal2 s 49422 0 49478 800 0 FreeSans 224 90 0 0 top_width_0_height_0_subtile_3__pin_inpad_0_
port 158 nsew signal tristate
rlabel metal1 25484 23936 25484 23936 0 VGND
rlabel metal1 25484 24480 25484 24480 0 VPWR
rlabel metal1 14490 3672 14490 3672 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal1 9200 3638 9200 3638 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 15686 4862 15686 4862 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal1 19918 4250 19918 4250 0 cbx_8__0_.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 26450 17000 26450 17000 0 cbx_8__0_.cbx_8__0_.ccff_head
rlabel metal1 10212 9350 10212 9350 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.ccff_tail
rlabel metal1 21528 16558 21528 16558 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[0\]
rlabel metal2 9246 12988 9246 12988 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[1\]
rlabel metal1 10442 7854 10442 7854 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_0.mem_out\[2\]
rlabel metal2 7222 9792 7222 9792 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.ccff_tail
rlabel metal2 4048 20604 4048 20604 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[0\]
rlabel metal3 5980 9452 5980 9452 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[1\]
rlabel metal1 5842 12954 5842 12954 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_1.mem_out\[2\]
rlabel metal1 8418 11152 8418 11152 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.ccff_tail
rlabel metal2 7084 19924 7084 19924 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[0\]
rlabel metal1 4508 8942 4508 8942 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[1\]
rlabel metal1 6302 13430 6302 13430 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_2.mem_out\[2\]
rlabel metal1 2346 23630 2346 23630 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[0\]
rlabel metal2 5750 20502 5750 20502 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[1\]
rlabel metal1 2484 2618 2484 2618 0 cbx_8__0_.cbx_8__0_.mem_top_ipin_3.mem_out\[2\]
rlabel metal1 9844 13294 9844 13294 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9890 8279 9890 8279 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal2 11914 6154 11914 6154 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 9476 13158 9476 13158 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9246 15130 9246 15130 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 10028 15062 10028 15062 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9798 14008 9798 14008 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 9982 11271 9982 11271 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 9982 11118 9982 11118 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 10304 7718 10304 7718 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 10396 12614 10396 12614 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 10810 9690 10810 9690 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 4508 15130 4508 15130 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 6946 11152 6946 11152 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 7084 3502 7084 3502 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 3358 12954 3358 12954 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 9062 16048 9062 16048 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 7176 16218 7176 16218 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9568 14518 9568 14518 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 5106 14620 5106 14620 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 5014 15096 5014 15096 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 6486 9350 6486 9350 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 5658 12206 5658 12206 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 5428 13396 5428 13396 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 5750 15215 5750 15215 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9430 11560 9430 11560 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 6026 4080 6026 4080 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 7314 15062 7314 15062 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 7176 14042 7176 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6992 13974 6992 13974 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 10120 12070 10120 12070 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 5704 13362 5704 13362 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 6348 13226 6348 13226 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 9522 13260 9522 13260 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 11132 13294 11132 13294 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 6716 13158 6716 13158 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 7314 17034 7314 17034 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8556 17578 8556 17578 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal4 13524 13452 13524 13452 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal2 2622 22168 2622 22168 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6716 17306 6716 17306 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 6992 15674 6992 15674 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 9154 14042 9154 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 10810 17714 10810 17714 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 5290 17272 5290 17272 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 8280 14042 8280 14042 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 9476 18666 9476 18666 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 9430 17510 9430 17510 0 cbx_8__0_.cbx_8__0_.mux_top_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 19550 3740 19550 3740 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 17296 3094 17296 3094 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 27209 4726 27209 4726 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 20608 6290 20608 6290 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 17112 4046 17112 4046 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal1 25231 4794 25231 4794 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 24748 7514 24748 7514 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal1 16468 4522 16468 4522 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal1 24242 4658 24242 4658 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 17618 5542 17618 5542 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 24978 5440 24978 5440 0 cbx_8__0_.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 8740 2618 8740 2618 0 ccff_head
rlabel metal1 48530 21114 48530 21114 0 ccff_head_1
rlabel metal2 49174 21233 49174 21233 0 ccff_tail
rlabel metal2 2530 23851 2530 23851 0 ccff_tail_0
rlabel metal3 2062 1564 2062 1564 0 chanx_left_in[0]
rlabel metal1 1472 5678 1472 5678 0 chanx_left_in[10]
rlabel metal1 1794 6290 1794 6290 0 chanx_left_in[11]
rlabel metal1 13708 2618 13708 2618 0 chanx_left_in[12]
rlabel metal2 22218 6579 22218 6579 0 chanx_left_in[13]
rlabel metal2 21206 6222 21206 6222 0 chanx_left_in[14]
rlabel metal1 11316 918 11316 918 0 chanx_left_in[15]
rlabel metal2 3404 2380 3404 2380 0 chanx_left_in[16]
rlabel metal3 8303 1156 8303 1156 0 chanx_left_in[17]
rlabel metal1 12604 986 12604 986 0 chanx_left_in[18]
rlabel metal1 11408 578 11408 578 0 chanx_left_in[19]
rlabel metal3 2108 1972 2108 1972 0 chanx_left_in[1]
rlabel metal3 7820 9656 7820 9656 0 chanx_left_in[20]
rlabel metal2 15778 5117 15778 5117 0 chanx_left_in[21]
rlabel metal3 16215 1020 16215 1020 0 chanx_left_in[22]
rlabel metal2 14214 1853 14214 1853 0 chanx_left_in[23]
rlabel metal1 19366 4658 19366 4658 0 chanx_left_in[24]
rlabel metal2 11730 1632 11730 1632 0 chanx_left_in[25]
rlabel metal1 2438 11152 2438 11152 0 chanx_left_in[26]
rlabel metal2 15962 4709 15962 4709 0 chanx_left_in[27]
rlabel metal1 8878 442 8878 442 0 chanx_left_in[28]
rlabel metal1 1380 12750 1380 12750 0 chanx_left_in[29]
rlabel metal1 1610 2380 1610 2380 0 chanx_left_in[2]
rlabel metal2 11178 1938 11178 1938 0 chanx_left_in[3]
rlabel metal1 17434 2482 17434 2482 0 chanx_left_in[4]
rlabel metal1 8027 1802 8027 1802 0 chanx_left_in[5]
rlabel metal1 11362 238 11362 238 0 chanx_left_in[6]
rlabel metal1 11224 1054 11224 1054 0 chanx_left_in[7]
rlabel metal2 11546 2176 11546 2176 0 chanx_left_in[8]
rlabel metal1 2852 2414 2852 2414 0 chanx_left_in[9]
rlabel metal3 1372 13804 1372 13804 0 chanx_left_out[0]
rlabel metal3 1050 17884 1050 17884 0 chanx_left_out[10]
rlabel metal3 1372 18292 1372 18292 0 chanx_left_out[11]
rlabel metal3 1096 18700 1096 18700 0 chanx_left_out[12]
rlabel metal3 1050 19108 1050 19108 0 chanx_left_out[13]
rlabel metal3 1372 19516 1372 19516 0 chanx_left_out[14]
rlabel metal2 2806 20689 2806 20689 0 chanx_left_out[15]
rlabel metal3 1096 20332 1096 20332 0 chanx_left_out[16]
rlabel metal2 3818 20859 3818 20859 0 chanx_left_out[17]
rlabel metal3 1464 21148 1464 21148 0 chanx_left_out[18]
rlabel metal3 1694 21556 1694 21556 0 chanx_left_out[19]
rlabel metal3 1004 14212 1004 14212 0 chanx_left_out[1]
rlabel metal2 3358 22015 3358 22015 0 chanx_left_out[20]
rlabel metal3 1487 22372 1487 22372 0 chanx_left_out[21]
rlabel metal1 3726 21114 3726 21114 0 chanx_left_out[22]
rlabel metal3 1717 23188 1717 23188 0 chanx_left_out[23]
rlabel metal1 5382 21590 5382 21590 0 chanx_left_out[24]
rlabel metal1 3956 19754 3956 19754 0 chanx_left_out[25]
rlabel metal2 2806 24021 2806 24021 0 chanx_left_out[26]
rlabel metal2 4002 24599 4002 24599 0 chanx_left_out[27]
rlabel metal2 4784 19924 4784 19924 0 chanx_left_out[28]
rlabel metal2 4094 25347 4094 25347 0 chanx_left_out[29]
rlabel metal3 1004 14620 1004 14620 0 chanx_left_out[2]
rlabel metal3 1004 15028 1004 15028 0 chanx_left_out[3]
rlabel metal3 1004 15436 1004 15436 0 chanx_left_out[4]
rlabel metal3 1004 15844 1004 15844 0 chanx_left_out[5]
rlabel metal3 1004 16252 1004 16252 0 chanx_left_out[6]
rlabel metal3 1004 16660 1004 16660 0 chanx_left_out[7]
rlabel metal3 958 17068 958 17068 0 chanx_left_out[8]
rlabel metal3 1372 17476 1372 17476 0 chanx_left_out[9]
rlabel metal2 13754 4114 13754 4114 0 chany_top_in[0]
rlabel metal1 43010 20298 43010 20298 0 chany_top_in[10]
rlabel metal1 29532 24242 29532 24242 0 chany_top_in[11]
rlabel metal1 34546 20842 34546 20842 0 chany_top_in[12]
rlabel metal1 33810 16116 33810 16116 0 chany_top_in[13]
rlabel metal2 44666 22882 44666 22882 0 chany_top_in[14]
rlabel metal1 44206 20944 44206 20944 0 chany_top_in[15]
rlabel metal1 44942 21556 44942 21556 0 chany_top_in[16]
rlabel metal1 33212 18394 33212 18394 0 chany_top_in[17]
rlabel metal1 49082 24174 49082 24174 0 chany_top_in[18]
rlabel metal1 37996 18666 37996 18666 0 chany_top_in[19]
rlabel metal3 28290 21556 28290 21556 0 chany_top_in[1]
rlabel metal2 45034 22372 45034 22372 0 chany_top_in[20]
rlabel metal1 39514 18836 39514 18836 0 chany_top_in[21]
rlabel metal1 44160 21522 44160 21522 0 chany_top_in[22]
rlabel metal1 39146 18326 39146 18326 0 chany_top_in[23]
rlabel metal1 39146 19346 39146 19346 0 chany_top_in[24]
rlabel metal1 38640 19414 38640 19414 0 chany_top_in[25]
rlabel metal1 40618 19414 40618 19414 0 chany_top_in[26]
rlabel metal2 41262 20230 41262 20230 0 chany_top_in[27]
rlabel metal2 41722 21012 41722 21012 0 chany_top_in[28]
rlabel metal1 43516 20910 43516 20910 0 chany_top_in[29]
rlabel metal2 30498 15232 30498 15232 0 chany_top_in[2]
rlabel metal1 36800 21318 36800 21318 0 chany_top_in[3]
rlabel metal1 32108 15470 32108 15470 0 chany_top_in[4]
rlabel metal2 1794 23936 1794 23936 0 chany_top_in[5]
rlabel metal2 31786 15878 31786 15878 0 chany_top_in[6]
rlabel metal1 36892 22746 36892 22746 0 chany_top_in[7]
rlabel metal1 37536 17646 37536 17646 0 chany_top_in[8]
rlabel metal2 45954 24990 45954 24990 0 chany_top_in[9]
rlabel metal1 3542 23290 3542 23290 0 chany_top_out[0]
rlabel metal1 8786 24242 8786 24242 0 chany_top_out[10]
rlabel metal1 9568 23630 9568 23630 0 chany_top_out[11]
rlabel metal2 10534 24735 10534 24735 0 chany_top_out[12]
rlabel metal2 11270 24184 11270 24184 0 chany_top_out[13]
rlabel metal2 12834 22066 12834 22066 0 chany_top_out[14]
rlabel metal2 12466 24157 12466 24157 0 chany_top_out[15]
rlabel metal2 13478 24191 13478 24191 0 chany_top_out[16]
rlabel metal2 13846 25204 13846 25204 0 chany_top_out[17]
rlabel metal1 13570 24276 13570 24276 0 chany_top_out[18]
rlabel metal1 15410 22066 15410 22066 0 chany_top_out[19]
rlabel metal1 3404 24242 3404 24242 0 chany_top_out[1]
rlabel metal1 15042 23766 15042 23766 0 chany_top_out[20]
rlabel metal2 16146 24497 16146 24497 0 chany_top_out[21]
rlabel metal2 17211 26588 17211 26588 0 chany_top_out[22]
rlabel metal1 16698 23086 16698 23086 0 chany_top_out[23]
rlabel metal1 17250 23630 17250 23630 0 chany_top_out[24]
rlabel metal1 17572 24242 17572 24242 0 chany_top_out[25]
rlabel metal1 18676 23766 18676 23766 0 chany_top_out[26]
rlabel metal1 20792 22066 20792 22066 0 chany_top_out[27]
rlabel metal2 20930 25272 20930 25272 0 chany_top_out[28]
rlabel metal2 21574 25272 21574 25272 0 chany_top_out[29]
rlabel metal1 4094 23698 4094 23698 0 chany_top_out[2]
rlabel metal2 5106 24429 5106 24429 0 chany_top_out[3]
rlabel metal2 5474 24966 5474 24966 0 chany_top_out[4]
rlabel metal2 6118 24728 6118 24728 0 chany_top_out[5]
rlabel metal1 7176 22066 7176 22066 0 chany_top_out[6]
rlabel metal1 6624 24242 6624 24242 0 chany_top_out[7]
rlabel metal2 7866 24735 7866 24735 0 chany_top_out[8]
rlabel metal2 8602 24497 8602 24497 0 chany_top_out[9]
rlabel metal1 12650 19346 12650 19346 0 clknet_0_prog_clk
rlabel metal2 8510 6256 8510 6256 0 clknet_4_0_0_prog_clk
rlabel metal2 21942 9282 21942 9282 0 clknet_4_10_0_prog_clk
rlabel metal1 19596 16626 19596 16626 0 clknet_4_11_0_prog_clk
rlabel metal2 15870 19278 15870 19278 0 clknet_4_12_0_prog_clk
rlabel metal1 21022 18802 21022 18802 0 clknet_4_13_0_prog_clk
rlabel metal2 25806 18496 25806 18496 0 clknet_4_14_0_prog_clk
rlabel metal1 20332 23834 20332 23834 0 clknet_4_15_0_prog_clk
rlabel metal2 4186 13056 4186 13056 0 clknet_4_1_0_prog_clk
rlabel metal2 16882 7616 16882 7616 0 clknet_4_2_0_prog_clk
rlabel metal2 14674 14178 14674 14178 0 clknet_4_3_0_prog_clk
rlabel metal1 5566 17714 5566 17714 0 clknet_4_4_0_prog_clk
rlabel metal1 9844 19822 9844 19822 0 clknet_4_5_0_prog_clk
rlabel metal1 14352 18326 14352 18326 0 clknet_4_6_0_prog_clk
rlabel metal2 13570 19890 13570 19890 0 clknet_4_7_0_prog_clk
rlabel metal1 17296 11186 17296 11186 0 clknet_4_8_0_prog_clk
rlabel metal2 19734 14688 19734 14688 0 clknet_4_9_0_prog_clk
rlabel metal2 4094 1622 4094 1622 0 gfpga_pad_io_soc_dir[0]
rlabel metal2 6762 1622 6762 1622 0 gfpga_pad_io_soc_dir[1]
rlabel metal2 9430 1622 9430 1622 0 gfpga_pad_io_soc_dir[2]
rlabel metal2 12098 1622 12098 1622 0 gfpga_pad_io_soc_dir[3]
rlabel metal1 25576 2414 25576 2414 0 gfpga_pad_io_soc_in[0]
rlabel metal2 28382 1581 28382 1581 0 gfpga_pad_io_soc_in[1]
rlabel metal1 30912 2414 30912 2414 0 gfpga_pad_io_soc_in[2]
rlabel metal1 33580 2414 33580 2414 0 gfpga_pad_io_soc_in[3]
rlabel metal1 15042 4114 15042 4114 0 gfpga_pad_io_soc_out[0]
rlabel metal1 17480 4522 17480 4522 0 gfpga_pad_io_soc_out[1]
rlabel metal1 19412 4046 19412 4046 0 gfpga_pad_io_soc_out[2]
rlabel metal1 21574 3094 21574 3094 0 gfpga_pad_io_soc_out[3]
rlabel metal2 36110 1588 36110 1588 0 isol_n
rlabel metal2 17618 2567 17618 2567 0 net1
rlabel metal2 15778 1768 15778 1768 0 net10
rlabel metal1 9338 20876 9338 20876 0 net100
rlabel metal2 3634 14892 3634 14892 0 net101
rlabel metal1 2254 14994 2254 14994 0 net102
rlabel metal1 1840 15470 1840 15470 0 net103
rlabel metal2 1794 15470 1794 15470 0 net104
rlabel metal1 1794 16660 1794 16660 0 net105
rlabel metal2 1794 16865 1794 16865 0 net106
rlabel metal1 2277 17646 2277 17646 0 net107
rlabel metal2 3358 15759 3358 15759 0 net108
rlabel metal4 13524 8908 13524 8908 0 net109
rlabel metal1 14306 15470 14306 15470 0 net11
rlabel metal2 22126 1241 22126 1241 0 net110
rlabel metal1 12558 7480 12558 7480 0 net111
rlabel metal2 40986 15657 40986 15657 0 net112
rlabel metal2 38410 12461 38410 12461 0 net113
rlabel via2 36938 17765 36938 17765 0 net114
rlabel metal2 35098 15793 35098 15793 0 net115
rlabel metal1 40664 19958 40664 19958 0 net116
rlabel metal2 34730 10846 34730 10846 0 net117
rlabel metal2 42826 17646 42826 17646 0 net118
rlabel metal2 18446 20825 18446 20825 0 net119
rlabel metal2 23874 7735 23874 7735 0 net12
rlabel metal2 2254 24225 2254 24225 0 net120
rlabel metal2 43562 20128 43562 20128 0 net121
rlabel metal3 17572 20468 17572 20468 0 net122
rlabel metal1 17112 21522 17112 21522 0 net123
rlabel metal2 41998 23443 41998 23443 0 net124
rlabel metal3 16077 21148 16077 21148 0 net125
rlabel metal3 18354 20332 18354 20332 0 net126
rlabel metal2 21068 16796 21068 16796 0 net127
rlabel metal3 18492 21964 18492 21964 0 net128
rlabel metal2 20102 25194 20102 25194 0 net129
rlabel metal1 12604 850 12604 850 0 net13
rlabel metal3 30130 20740 30130 20740 0 net130
rlabel metal3 14605 16932 14605 16932 0 net131
rlabel metal1 1288 22542 1288 22542 0 net132
rlabel via2 3933 884 3933 884 0 net133
rlabel via2 5382 4131 5382 4131 0 net134
rlabel metal4 1012 18786 1012 18786 0 net135
rlabel via2 34362 20349 34362 20349 0 net136
rlabel metal2 12696 19346 12696 19346 0 net137
rlabel metal2 34362 21777 34362 21777 0 net138
rlabel metal2 4370 2040 4370 2040 0 net139
rlabel metal1 18814 2380 18814 2380 0 net14
rlabel metal1 7038 2380 7038 2380 0 net140
rlabel metal1 10718 2414 10718 2414 0 net141
rlabel metal2 15226 2516 15226 2516 0 net142
rlabel metal2 6210 12512 6210 12512 0 net143
rlabel metal1 17611 5610 17611 5610 0 net144
rlabel metal1 6433 14314 6433 14314 0 net145
rlabel metal1 12841 23018 12841 23018 0 net146
rlabel metal2 21022 19584 21022 19584 0 net147
rlabel metal1 22264 21454 22264 21454 0 net148
rlabel metal1 6118 21964 6118 21964 0 net149
rlabel via2 20010 5219 20010 5219 0 net15
rlabel metal2 26450 18700 26450 18700 0 net150
rlabel metal1 24242 14246 24242 14246 0 net151
rlabel metal2 42826 23358 42826 23358 0 net152
rlabel metal1 18768 20910 18768 20910 0 net153
rlabel metal1 23230 19856 23230 19856 0 net154
rlabel metal1 18492 12274 18492 12274 0 net155
rlabel metal2 21390 24276 21390 24276 0 net156
rlabel metal2 24012 17884 24012 17884 0 net157
rlabel metal1 24426 24106 24426 24106 0 net158
rlabel metal1 26036 21590 26036 21590 0 net159
rlabel via2 16698 14059 16698 14059 0 net16
rlabel metal1 27002 18802 27002 18802 0 net160
rlabel metal1 26772 16558 26772 16558 0 net161
rlabel metal2 18630 18292 18630 18292 0 net162
rlabel metal2 22494 17408 22494 17408 0 net163
rlabel metal1 21206 18836 21206 18836 0 net164
rlabel metal1 16238 21522 16238 21522 0 net165
rlabel metal2 19642 15266 19642 15266 0 net166
rlabel metal1 16974 7446 16974 7446 0 net167
rlabel metal3 15617 2652 15617 2652 0 net168
rlabel metal1 12926 3400 12926 3400 0 net169
rlabel metal2 20654 13005 20654 13005 0 net17
rlabel metal1 7544 3094 7544 3094 0 net170
rlabel metal1 13708 13702 13708 13702 0 net171
rlabel metal2 14582 7650 14582 7650 0 net172
rlabel metal1 16560 17238 16560 17238 0 net173
rlabel metal2 14214 17731 14214 17731 0 net174
rlabel metal2 14306 15776 14306 15776 0 net175
rlabel metal1 3312 2482 3312 2482 0 net176
rlabel metal1 18630 7956 18630 7956 0 net177
rlabel via2 9062 6749 9062 6749 0 net178
rlabel metal1 17572 1190 17572 1190 0 net179
rlabel metal1 14490 2618 14490 2618 0 net18
rlabel metal2 20838 3383 20838 3383 0 net180
rlabel metal3 10327 20740 10327 20740 0 net181
rlabel metal2 10994 1751 10994 1751 0 net182
rlabel metal1 8832 3366 8832 3366 0 net183
rlabel via2 21942 4675 21942 4675 0 net184
rlabel metal2 34822 15997 34822 15997 0 net185
rlabel metal1 20930 3570 20930 3570 0 net186
rlabel metal4 20884 15640 20884 15640 0 net187
rlabel metal4 1932 14336 1932 14336 0 net188
rlabel metal1 9430 7922 9430 7922 0 net189
rlabel metal1 20332 9894 20332 9894 0 net19
rlabel metal2 15870 10982 15870 10982 0 net190
rlabel metal1 15318 7922 15318 7922 0 net191
rlabel metal1 9246 5746 9246 5746 0 net192
rlabel metal2 13800 2652 13800 2652 0 net193
rlabel metal2 14122 15997 14122 15997 0 net194
rlabel metal1 15824 10574 15824 10574 0 net195
rlabel metal1 27554 16558 27554 16558 0 net196
rlabel metal2 41906 16541 41906 16541 0 net197
rlabel metal1 17848 17850 17848 17850 0 net198
rlabel metal1 19458 12342 19458 12342 0 net199
rlabel metal2 47058 22678 47058 22678 0 net2
rlabel metal2 10994 11577 10994 11577 0 net20
rlabel metal2 7912 23052 7912 23052 0 net200
rlabel metal2 48714 22202 48714 22202 0 net201
rlabel metal1 42642 22032 42642 22032 0 net202
rlabel metal2 1702 4250 1702 4250 0 net203
rlabel metal1 7498 3026 7498 3026 0 net204
rlabel metal1 37766 22746 37766 22746 0 net205
rlabel metal1 31970 21998 31970 21998 0 net206
rlabel metal2 1978 11271 1978 11271 0 net207
rlabel metal2 28842 21522 28842 21522 0 net208
rlabel metal2 36662 19924 36662 19924 0 net209
rlabel metal1 1978 23596 1978 23596 0 net21
rlabel metal1 22908 8942 22908 8942 0 net210
rlabel metal1 21574 6766 21574 6766 0 net211
rlabel metal2 38870 21556 38870 21556 0 net212
rlabel metal1 23598 8058 23598 8058 0 net213
rlabel metal1 33258 18292 33258 18292 0 net214
rlabel metal1 14306 4624 14306 4624 0 net215
rlabel metal1 5796 10166 5796 10166 0 net216
rlabel metal1 8418 4794 8418 4794 0 net217
rlabel metal1 29992 12818 29992 12818 0 net218
rlabel metal1 23874 9554 23874 9554 0 net219
rlabel metal2 35282 17221 35282 17221 0 net22
rlabel metal1 12006 6800 12006 6800 0 net220
rlabel metal1 43746 23290 43746 23290 0 net221
rlabel metal1 3174 11118 3174 11118 0 net222
rlabel metal1 28842 14382 28842 14382 0 net223
rlabel metal2 1886 6460 1886 6460 0 net224
rlabel metal1 16008 6426 16008 6426 0 net225
rlabel metal1 11684 5202 11684 5202 0 net226
rlabel metal1 19182 8942 19182 8942 0 net227
rlabel metal1 12926 18734 12926 18734 0 net228
rlabel metal1 12880 7854 12880 7854 0 net229
rlabel via3 19205 21148 19205 21148 0 net23
rlabel metal1 16054 4250 16054 4250 0 net230
rlabel metal2 39698 23868 39698 23868 0 net231
rlabel metal1 43470 23698 43470 23698 0 net232
rlabel metal1 26680 12410 26680 12410 0 net233
rlabel metal1 35834 21012 35834 21012 0 net234
rlabel metal1 16100 16558 16100 16558 0 net235
rlabel metal2 15686 6732 15686 6732 0 net236
rlabel metal1 12006 5712 12006 5712 0 net237
rlabel metal1 26956 13294 26956 13294 0 net238
rlabel metal1 33258 16660 33258 16660 0 net239
rlabel metal1 20148 17102 20148 17102 0 net24
rlabel metal1 16882 6256 16882 6256 0 net240
rlabel metal1 35742 20570 35742 20570 0 net241
rlabel metal2 16422 8058 16422 8058 0 net242
rlabel metal1 34316 17306 34316 17306 0 net243
rlabel metal2 40710 21556 40710 21556 0 net244
rlabel metal2 2438 8500 2438 8500 0 net245
rlabel metal1 9614 1360 9614 1360 0 net246
rlabel metal1 8096 7514 8096 7514 0 net247
rlabel via2 17894 8891 17894 8891 0 net248
rlabel metal1 19412 18054 19412 18054 0 net249
rlabel metal1 1288 2482 1288 2482 0 net25
rlabel metal1 26358 13158 26358 13158 0 net250
rlabel metal2 8970 5780 8970 5780 0 net251
rlabel metal1 12765 4794 12765 4794 0 net252
rlabel metal2 37582 16490 37582 16490 0 net253
rlabel metal4 17756 12648 17756 12648 0 net254
rlabel metal2 38594 23052 38594 23052 0 net255
rlabel metal1 30544 18326 30544 18326 0 net256
rlabel metal2 9982 4947 9982 4947 0 net257
rlabel metal1 33718 22066 33718 22066 0 net258
rlabel metal2 8418 8126 8418 8126 0 net259
rlabel metal2 8786 6035 8786 6035 0 net26
rlabel metal2 32338 18938 32338 18938 0 net260
rlabel metal2 36018 20876 36018 20876 0 net261
rlabel metal2 15318 3757 15318 3757 0 net262
rlabel metal1 10396 3502 10396 3502 0 net263
rlabel metal1 33212 19822 33212 19822 0 net264
rlabel metal1 37490 23664 37490 23664 0 net265
rlabel metal2 31050 24004 31050 24004 0 net266
rlabel metal2 32246 20026 32246 20026 0 net267
rlabel metal2 20654 9078 20654 9078 0 net268
rlabel metal2 15226 5984 15226 5984 0 net269
rlabel metal2 7590 9503 7590 9503 0 net27
rlabel metal2 6578 17476 6578 17476 0 net270
rlabel metal1 7452 5882 7452 5882 0 net271
rlabel metal2 2254 6562 2254 6562 0 net272
rlabel metal1 22034 22576 22034 22576 0 net273
rlabel metal1 42274 23120 42274 23120 0 net274
rlabel metal2 9798 7378 9798 7378 0 net275
rlabel metal1 34500 22610 34500 22610 0 net276
rlabel metal2 33534 21114 33534 21114 0 net277
rlabel metal1 44252 24242 44252 24242 0 net278
rlabel metal2 22678 18496 22678 18496 0 net279
rlabel metal1 18906 2618 18906 2618 0 net28
rlabel metal1 4094 14042 4094 14042 0 net280
rlabel metal2 31878 15912 31878 15912 0 net281
rlabel metal2 41814 23494 41814 23494 0 net282
rlabel metal2 36018 23290 36018 23290 0 net283
rlabel metal1 28336 9690 28336 9690 0 net284
rlabel metal1 33212 24174 33212 24174 0 net285
rlabel metal1 36294 22746 36294 22746 0 net286
rlabel metal2 21942 14739 21942 14739 0 net287
rlabel metal1 15870 17850 15870 17850 0 net288
rlabel via2 39054 20451 39054 20451 0 net289
rlabel metal1 19964 3366 19964 3366 0 net29
rlabel metal1 20010 15096 20010 15096 0 net290
rlabel metal1 3910 7514 3910 7514 0 net291
rlabel metal1 6578 7310 6578 7310 0 net292
rlabel metal2 16974 11203 16974 11203 0 net293
rlabel metal1 22586 8602 22586 8602 0 net294
rlabel metal3 15364 13192 15364 13192 0 net295
rlabel metal2 8602 7616 8602 7616 0 net296
rlabel metal1 8924 9962 8924 9962 0 net297
rlabel metal2 21666 10778 21666 10778 0 net298
rlabel metal1 7084 13226 7084 13226 0 net299
rlabel metal1 16054 4794 16054 4794 0 net3
rlabel metal1 14858 1462 14858 1462 0 net30
rlabel metal1 21206 12750 21206 12750 0 net300
rlabel metal1 20240 7446 20240 7446 0 net301
rlabel metal1 19044 6426 19044 6426 0 net302
rlabel metal1 18170 11866 18170 11866 0 net303
rlabel metal1 26496 16014 26496 16014 0 net304
rlabel metal1 13984 20502 13984 20502 0 net305
rlabel metal2 24242 10302 24242 10302 0 net306
rlabel metal2 14950 11135 14950 11135 0 net307
rlabel via2 14766 9605 14766 9605 0 net308
rlabel metal2 35558 18343 35558 18343 0 net309
rlabel metal2 9062 15096 9062 15096 0 net31
rlabel metal2 12558 23188 12558 23188 0 net310
rlabel metal1 4600 7514 4600 7514 0 net311
rlabel metal1 4784 8058 4784 8058 0 net312
rlabel metal1 15272 7514 15272 7514 0 net313
rlabel metal2 5612 12716 5612 12716 0 net314
rlabel metal2 2346 13430 2346 13430 0 net315
rlabel metal1 4130 13702 4130 13702 0 net316
rlabel metal2 49358 23698 49358 23698 0 net317
rlabel metal1 46506 23120 46506 23120 0 net318
rlabel metal1 46414 23154 46414 23154 0 net319
rlabel metal1 15962 14926 15962 14926 0 net32
rlabel metal2 43286 21760 43286 21760 0 net320
rlabel metal2 4646 4352 4646 4352 0 net321
rlabel metal2 3542 3468 3542 3468 0 net322
rlabel metal1 5934 3026 5934 3026 0 net323
rlabel metal1 8786 2958 8786 2958 0 net324
rlabel metal2 37490 23324 37490 23324 0 net325
rlabel metal2 36662 24752 36662 24752 0 net326
rlabel metal2 30958 21828 30958 21828 0 net327
rlabel metal1 27554 21896 27554 21896 0 net328
rlabel metal1 7406 7854 7406 7854 0 net329
rlabel via2 17434 20757 17434 20757 0 net33
rlabel metal2 2622 15827 2622 15827 0 net330
rlabel metal1 31510 20876 31510 20876 0 net331
rlabel metal1 26673 18938 26673 18938 0 net332
rlabel metal2 20838 6596 20838 6596 0 net333
rlabel metal1 22402 6970 22402 6970 0 net334
rlabel metal2 20930 8500 20930 8500 0 net335
rlabel metal2 21390 10098 21390 10098 0 net336
rlabel metal1 35052 17714 35052 17714 0 net337
rlabel metal2 21804 13362 21804 13362 0 net338
rlabel metal2 36018 19516 36018 19516 0 net339
rlabel metal1 43424 20842 43424 20842 0 net34
rlabel metal1 18952 21590 18952 21590 0 net340
rlabel metal1 17940 5338 17940 5338 0 net341
rlabel metal1 19642 9452 19642 9452 0 net342
rlabel metal2 10994 5780 10994 5780 0 net343
rlabel metal1 14674 4794 14674 4794 0 net344
rlabel metal2 11086 9622 11086 9622 0 net345
rlabel metal1 5014 12376 5014 12376 0 net346
rlabel metal2 38226 21114 38226 21114 0 net347
rlabel metal1 40388 22066 40388 22066 0 net348
rlabel metal1 24748 9350 24748 9350 0 net349
rlabel metal2 19734 25381 19734 25381 0 net35
rlabel metal1 23874 9656 23874 9656 0 net350
rlabel metal1 7498 4590 7498 4590 0 net351
rlabel metal3 6739 20876 6739 20876 0 net352
rlabel metal2 16330 15453 16330 15453 0 net353
rlabel metal1 25760 14586 25760 14586 0 net354
rlabel metal2 8326 6732 8326 6732 0 net355
rlabel metal1 3496 11322 3496 11322 0 net356
rlabel metal1 43792 23086 43792 23086 0 net357
rlabel metal2 41906 24718 41906 24718 0 net358
rlabel metal2 8786 8636 8786 8636 0 net359
rlabel metal1 6164 2482 6164 2482 0 net36
rlabel metal1 12489 13158 12489 13158 0 net360
rlabel metal1 30682 14586 30682 14586 0 net361
rlabel metal3 16836 13940 16836 13940 0 net362
rlabel metal2 13754 6086 13754 6086 0 net363
rlabel metal1 17020 6834 17020 6834 0 net364
rlabel metal1 4784 5678 4784 5678 0 net365
rlabel metal2 2530 12546 2530 12546 0 net366
rlabel via2 13846 10149 13846 10149 0 net367
rlabel metal2 17986 24718 17986 24718 0 net368
rlabel metal1 12098 7854 12098 7854 0 net369
rlabel metal2 31694 15776 31694 15776 0 net37
rlabel via2 13731 14484 13731 14484 0 net370
rlabel metal1 10534 5236 10534 5236 0 net371
rlabel metal2 12834 5474 12834 5474 0 net372
rlabel metal1 19182 8602 19182 8602 0 net373
rlabel metal1 20194 9146 20194 9146 0 net374
rlabel metal2 37030 25058 37030 25058 0 net375
rlabel metal1 20332 23018 20332 23018 0 net376
rlabel metal1 11684 4182 11684 4182 0 net377
rlabel metal1 43838 23562 43838 23562 0 net378
rlabel metal1 24748 12206 24748 12206 0 net379
rlabel metal1 44436 23290 44436 23290 0 net38
rlabel metal1 26726 14926 26726 14926 0 net380
rlabel metal1 38916 21930 38916 21930 0 net381
rlabel metal1 19872 20842 19872 20842 0 net382
rlabel metal1 10166 6392 10166 6392 0 net383
rlabel metal1 12742 5882 12742 5882 0 net384
rlabel metal1 17664 8058 17664 8058 0 net385
rlabel metal1 18676 9146 18676 9146 0 net386
rlabel metal1 33764 17170 33764 17170 0 net387
rlabel metal3 18952 12852 18952 12852 0 net388
rlabel via2 18078 8381 18078 8381 0 net389
rlabel metal1 33856 21046 33856 21046 0 net39
rlabel metal2 17158 15725 17158 15725 0 net390
rlabel metal1 18998 6256 18998 6256 0 net391
rlabel metal1 17664 6426 17664 6426 0 net392
rlabel metal1 13294 3706 13294 3706 0 net393
rlabel metal2 18630 5270 18630 5270 0 net394
rlabel metal1 8188 9690 8188 9690 0 net395
rlabel metal2 12926 7429 12926 7429 0 net396
rlabel metal1 5198 9894 5198 9894 0 net397
rlabel metal1 7406 8534 7406 8534 0 net398
rlabel metal2 15686 7548 15686 7548 0 net399
rlabel metal1 14490 14994 14490 14994 0 net4
rlabel metal2 44758 20553 44758 20553 0 net40
rlabel metal1 14628 13226 14628 13226 0 net400
rlabel metal1 12466 4522 12466 4522 0 net401
rlabel metal1 11592 5882 11592 5882 0 net402
rlabel metal2 32430 16456 32430 16456 0 net403
rlabel metal1 18206 16762 18206 16762 0 net404
rlabel metal1 6348 8942 6348 8942 0 net405
rlabel metal1 13340 7446 13340 7446 0 net406
rlabel metal2 35558 20230 35558 20230 0 net407
rlabel metal1 20286 20366 20286 20366 0 net408
rlabel metal2 27784 13260 27784 13260 0 net409
rlabel via1 16974 17187 16974 17187 0 net41
rlabel metal1 23276 12886 23276 12886 0 net410
rlabel metal1 39468 20026 39468 20026 0 net411
rlabel metal2 41630 24276 41630 24276 0 net412
rlabel metal2 4922 7106 4922 7106 0 net413
rlabel metal1 4278 9112 4278 9112 0 net414
rlabel metal1 18078 18292 18078 18292 0 net415
rlabel metal1 23092 16558 23092 16558 0 net416
rlabel metal1 36524 17850 36524 17850 0 net417
rlabel metal1 33718 16626 33718 16626 0 net418
rlabel metal2 8326 5372 8326 5372 0 net419
rlabel metal1 49036 24038 49036 24038 0 net42
rlabel metal3 5635 16116 5635 16116 0 net420
rlabel metal1 32292 16626 32292 16626 0 net421
rlabel metal1 15088 15402 15088 15402 0 net422
rlabel metal1 33764 23222 33764 23222 0 net423
rlabel metal2 29762 22712 29762 22712 0 net424
rlabel metal2 9338 4794 9338 4794 0 net425
rlabel metal1 5750 10234 5750 10234 0 net426
rlabel metal1 12834 3468 12834 3468 0 net427
rlabel metal1 8418 10744 8418 10744 0 net428
rlabel metal1 35282 21522 35282 21522 0 net429
rlabel metal1 36340 15470 36340 15470 0 net43
rlabel metal1 31050 20332 31050 20332 0 net430
rlabel metal1 20056 7514 20056 7514 0 net431
rlabel metal1 20930 9350 20930 9350 0 net432
rlabel metal1 32844 19346 32844 19346 0 net433
rlabel metal2 32982 18394 32982 18394 0 net434
rlabel metal2 9522 3706 9522 3706 0 net435
rlabel metal1 12466 4148 12466 4148 0 net436
rlabel metal1 32338 19856 32338 19856 0 net437
rlabel metal1 28796 19414 28796 19414 0 net438
rlabel metal2 32338 19958 32338 19958 0 net439
rlabel metal1 30038 16456 30038 16456 0 net44
rlabel metal1 30406 19958 30406 19958 0 net440
rlabel metal1 40618 23290 40618 23290 0 net441
rlabel metal2 39238 23834 39238 23834 0 net442
rlabel metal2 14582 5644 14582 5644 0 net443
rlabel metal1 13616 6834 13616 6834 0 net444
rlabel metal1 25806 13328 25806 13328 0 net445
rlabel metal1 24564 11662 24564 11662 0 net446
rlabel metal1 32660 23290 32660 23290 0 net447
rlabel metal1 25162 23800 25162 23800 0 net448
rlabel metal2 7498 5236 7498 5236 0 net449
rlabel metal2 45218 15929 45218 15929 0 net45
rlabel metal2 506 14178 506 14178 0 net450
rlabel metal1 30452 18258 30452 18258 0 net451
rlabel metal1 27416 17578 27416 17578 0 net452
rlabel metal1 42688 22746 42688 22746 0 net453
rlabel metal1 43286 23222 43286 23222 0 net454
rlabel metal1 35282 23698 35282 23698 0 net455
rlabel metal1 34914 23596 34914 23596 0 net456
rlabel metal1 33948 21522 33948 21522 0 net457
rlabel metal2 34178 20672 34178 20672 0 net458
rlabel metal2 7222 4386 7222 4386 0 net459
rlabel metal1 35558 18734 35558 18734 0 net46
rlabel via2 2346 8075 2346 8075 0 net460
rlabel metal1 22816 22066 22816 22066 0 net461
rlabel metal1 24370 22202 24370 22202 0 net462
rlabel metal1 7866 6426 7866 6426 0 net463
rlabel metal1 7222 20502 7222 20502 0 net464
rlabel via2 46138 23205 46138 23205 0 net465
rlabel metal1 35282 23834 35282 23834 0 net466
rlabel metal1 36984 18938 36984 18938 0 net467
rlabel via2 28934 13243 28934 13243 0 net468
rlabel metal1 11730 19414 11730 19414 0 net469
rlabel metal2 44114 21607 44114 21607 0 net47
rlabel metal2 7222 17391 7222 17391 0 net470
rlabel metal1 43056 21454 43056 21454 0 net471
rlabel metal2 42918 26299 42918 26299 0 net472
rlabel metal1 33718 22610 33718 22610 0 net473
rlabel metal1 35512 22746 35512 22746 0 net474
rlabel metal1 36018 23732 36018 23732 0 net475
rlabel metal1 32338 23188 32338 23188 0 net476
rlabel metal2 32062 17476 32062 17476 0 net477
rlabel metal1 27554 15946 27554 15946 0 net478
rlabel metal2 26358 9350 26358 9350 0 net479
rlabel metal1 32246 17204 32246 17204 0 net48
rlabel metal1 29762 10778 29762 10778 0 net480
rlabel metal1 19688 17714 19688 17714 0 net481
rlabel metal2 30406 18224 30406 18224 0 net482
rlabel metal1 32338 24208 32338 24208 0 net483
rlabel metal2 27462 23868 27462 23868 0 net484
rlabel via1 2622 6987 2622 6987 0 net485
rlabel metal1 38226 22066 38226 22066 0 net486
rlabel metal2 23874 10302 23874 10302 0 net487
rlabel metal1 41630 20536 41630 20536 0 net488
rlabel metal1 14444 17850 14444 17850 0 net489
rlabel metal2 39514 19754 39514 19754 0 net49
rlabel metal3 18492 16184 18492 16184 0 net490
rlabel metal1 5060 7378 5060 7378 0 net491
rlabel metal2 5290 7038 5290 7038 0 net492
rlabel metal2 31970 15283 31970 15283 0 net493
rlabel metal2 22770 9180 22770 9180 0 net494
rlabel metal1 7728 6766 7728 6766 0 net495
rlabel metal1 24932 9554 24932 9554 0 net496
rlabel metal1 26772 11322 26772 11322 0 net497
rlabel metal1 20378 6970 20378 6970 0 net498
rlabel metal1 5152 8466 5152 8466 0 net499
rlabel metal2 2714 5457 2714 5457 0 net5
rlabel metal1 15502 16762 15502 16762 0 net50
rlabel metal1 4968 9554 4968 9554 0 net500
rlabel metal1 19090 6324 19090 6324 0 net501
rlabel metal1 28106 12614 28106 12614 0 net502
rlabel metal2 18538 7106 18538 7106 0 net503
rlabel metal2 31234 16864 31234 16864 0 net504
rlabel metal1 34408 16014 34408 16014 0 net505
rlabel metal2 16330 4862 16330 4862 0 net506
rlabel metal1 25714 10608 25714 10608 0 net507
rlabel metal2 25346 8772 25346 8772 0 net508
rlabel metal2 44390 22236 44390 22236 0 net509
rlabel metal2 40802 19193 40802 19193 0 net51
rlabel metal2 2346 9112 2346 9112 0 net510
rlabel metal1 4094 7888 4094 7888 0 net511
rlabel metal2 2622 9486 2622 9486 0 net512
rlabel metal1 34914 19380 34914 19380 0 net513
rlabel metal2 2162 9282 2162 9282 0 net514
rlabel metal2 6394 7684 6394 7684 0 net515
rlabel metal1 16468 6834 16468 6834 0 net516
rlabel metal1 4646 3706 4646 3706 0 net517
rlabel metal1 4600 4794 4600 4794 0 net518
rlabel metal2 2346 3910 2346 3910 0 net519
rlabel metal1 41492 20366 41492 20366 0 net52
rlabel metal2 17802 2176 17802 2176 0 net520
rlabel metal1 4278 3026 4278 3026 0 net521
rlabel metal2 49358 22100 49358 22100 0 net522
rlabel metal1 48530 22610 48530 22610 0 net523
rlabel metal1 48944 22066 48944 22066 0 net524
rlabel metal2 47242 22236 47242 22236 0 net525
rlabel metal2 48438 24004 48438 24004 0 net526
rlabel metal2 41630 18496 41630 18496 0 net53
rlabel metal2 43378 20825 43378 20825 0 net54
rlabel metal1 30130 14042 30130 14042 0 net55
rlabel metal2 37766 22559 37766 22559 0 net56
rlabel metal1 32108 15606 32108 15606 0 net57
rlabel metal2 14306 24089 14306 24089 0 net58
rlabel metal2 31602 15929 31602 15929 0 net59
rlabel metal2 12374 10727 12374 10727 0 net6
rlabel metal2 37122 23001 37122 23001 0 net60
rlabel metal4 32844 16116 32844 16116 0 net61
rlabel metal2 44942 23970 44942 23970 0 net62
rlabel metal1 25162 5066 25162 5066 0 net63
rlabel metal1 28014 2618 28014 2618 0 net64
rlabel metal1 29026 4998 29026 4998 0 net65
rlabel metal2 33534 3842 33534 3842 0 net66
rlabel metal2 36386 5542 36386 5542 0 net67
rlabel metal2 41538 21828 41538 21828 0 net68
rlabel metal2 44850 18666 44850 18666 0 net69
rlabel metal1 17250 6120 17250 6120 0 net7
rlabel metal2 46690 21148 46690 21148 0 net70
rlabel metal2 47426 19550 47426 19550 0 net71
rlabel metal2 49082 15742 49082 15742 0 net72
rlabel metal2 46874 19431 46874 19431 0 net73
rlabel metal1 48024 21862 48024 21862 0 net74
rlabel metal2 45494 20570 45494 20570 0 net75
rlabel metal2 45402 19856 45402 19856 0 net76
rlabel metal1 47886 21522 47886 21522 0 net77
rlabel metal1 6854 20434 6854 20434 0 net78
rlabel via2 1610 13277 1610 13277 0 net79
rlabel metal1 19504 5678 19504 5678 0 net8
rlabel metal1 2668 18734 2668 18734 0 net80
rlabel metal1 1978 19346 1978 19346 0 net81
rlabel metal1 1334 19822 1334 19822 0 net82
rlabel metal1 1380 20434 1380 20434 0 net83
rlabel metal1 2024 20910 2024 20910 0 net84
rlabel via3 1725 20876 1725 20876 0 net85
rlabel metal2 1564 18598 1564 18598 0 net86
rlabel metal3 16031 748 16031 748 0 net87
rlabel metal1 1932 22610 1932 22610 0 net88
rlabel metal1 1840 23086 1840 23086 0 net89
rlabel metal1 17802 3502 17802 3502 0 net9
rlabel metal1 1472 17850 1472 17850 0 net90
rlabel metal3 3795 21556 3795 21556 0 net91
rlabel metal2 14766 22576 14766 22576 0 net92
rlabel metal2 9982 19584 9982 19584 0 net93
rlabel via2 13662 15045 13662 15045 0 net94
rlabel metal1 15870 20434 15870 20434 0 net95
rlabel metal1 3956 17170 3956 17170 0 net96
rlabel metal1 4186 16524 4186 16524 0 net97
rlabel metal1 7452 18258 7452 18258 0 net98
rlabel metal1 5106 16082 5106 16082 0 net99
rlabel metal2 38778 4240 38778 4240 0 prog_clk
rlabel metal2 41446 24004 41446 24004 0 prog_reset
rlabel metal1 19412 17034 19412 17034 0 sb_8__0_.mem_left_track_1.ccff_head
rlabel metal1 20838 18224 20838 18224 0 sb_8__0_.mem_left_track_1.ccff_tail
rlabel metal2 27830 17051 27830 17051 0 sb_8__0_.mem_left_track_1.mem_out\[0\]
rlabel metal1 19044 21862 19044 21862 0 sb_8__0_.mem_left_track_11.ccff_head
rlabel metal1 41722 19278 41722 19278 0 sb_8__0_.mem_left_track_11.ccff_tail
rlabel metal1 43838 22610 43838 22610 0 sb_8__0_.mem_left_track_11.mem_out\[0\]
rlabel metal2 44850 23919 44850 23919 0 sb_8__0_.mem_left_track_13.ccff_tail
rlabel metal1 38594 22474 38594 22474 0 sb_8__0_.mem_left_track_13.mem_out\[0\]
rlabel metal1 3772 20434 3772 20434 0 sb_8__0_.mem_left_track_15.ccff_tail
rlabel via2 31786 19125 31786 19125 0 sb_8__0_.mem_left_track_15.mem_out\[0\]
rlabel metal2 19090 20910 19090 20910 0 sb_8__0_.mem_left_track_17.ccff_tail
rlabel metal1 38594 24276 38594 24276 0 sb_8__0_.mem_left_track_17.mem_out\[0\]
rlabel metal1 18814 21012 18814 21012 0 sb_8__0_.mem_left_track_19.ccff_tail
rlabel metal2 33166 22797 33166 22797 0 sb_8__0_.mem_left_track_19.mem_out\[0\]
rlabel metal1 27232 18598 27232 18598 0 sb_8__0_.mem_left_track_29.ccff_tail
rlabel metal2 27830 20604 27830 20604 0 sb_8__0_.mem_left_track_29.mem_out\[0\]
rlabel metal2 21482 19771 21482 19771 0 sb_8__0_.mem_left_track_3.ccff_tail
rlabel metal1 17296 19346 17296 19346 0 sb_8__0_.mem_left_track_3.mem_out\[0\]
rlabel metal1 22908 21998 22908 21998 0 sb_8__0_.mem_left_track_31.ccff_tail
rlabel metal1 29026 21624 29026 21624 0 sb_8__0_.mem_left_track_31.mem_out\[0\]
rlabel metal1 34914 24242 34914 24242 0 sb_8__0_.mem_left_track_33.ccff_tail
rlabel metal1 29072 22542 29072 22542 0 sb_8__0_.mem_left_track_33.mem_out\[0\]
rlabel metal2 32246 24004 32246 24004 0 sb_8__0_.mem_left_track_35.ccff_tail
rlabel metal2 37490 24378 37490 24378 0 sb_8__0_.mem_left_track_35.mem_out\[0\]
rlabel metal2 27922 21522 27922 21522 0 sb_8__0_.mem_left_track_45.ccff_tail
rlabel metal2 40066 22814 40066 22814 0 sb_8__0_.mem_left_track_45.mem_out\[0\]
rlabel metal1 25346 22678 25346 22678 0 sb_8__0_.mem_left_track_47.ccff_tail
rlabel metal2 35006 21726 35006 21726 0 sb_8__0_.mem_left_track_47.mem_out\[0\]
rlabel metal1 29026 18054 29026 18054 0 sb_8__0_.mem_left_track_49.ccff_tail
rlabel metal1 33442 19380 33442 19380 0 sb_8__0_.mem_left_track_49.mem_out\[0\]
rlabel metal1 20976 20774 20976 20774 0 sb_8__0_.mem_left_track_5.ccff_tail
rlabel metal2 39698 22406 39698 22406 0 sb_8__0_.mem_left_track_5.mem_out\[0\]
rlabel metal1 30222 17170 30222 17170 0 sb_8__0_.mem_left_track_51.mem_out\[0\]
rlabel metal2 34454 18445 34454 18445 0 sb_8__0_.mem_left_track_7.ccff_tail
rlabel metal1 24334 18802 24334 18802 0 sb_8__0_.mem_left_track_7.mem_out\[0\]
rlabel metal2 16330 21148 16330 21148 0 sb_8__0_.mem_left_track_9.mem_out\[0\]
rlabel metal1 23782 16150 23782 16150 0 sb_8__0_.mem_top_track_0.ccff_tail
rlabel metal2 39882 19856 39882 19856 0 sb_8__0_.mem_top_track_0.mem_out\[0\]
rlabel metal1 21114 17102 21114 17102 0 sb_8__0_.mem_top_track_0.mem_out\[1\]
rlabel metal1 20838 12614 20838 12614 0 sb_8__0_.mem_top_track_10.ccff_head
rlabel metal1 18860 9622 18860 9622 0 sb_8__0_.mem_top_track_10.ccff_tail
rlabel metal1 24196 13838 24196 13838 0 sb_8__0_.mem_top_track_10.mem_out\[0\]
rlabel metal2 21850 10574 21850 10574 0 sb_8__0_.mem_top_track_10.mem_out\[1\]
rlabel metal2 19458 7684 19458 7684 0 sb_8__0_.mem_top_track_12.ccff_tail
rlabel metal1 15548 12750 15548 12750 0 sb_8__0_.mem_top_track_12.mem_out\[0\]
rlabel metal1 8234 8534 8234 8534 0 sb_8__0_.mem_top_track_14.ccff_tail
rlabel metal1 20378 7854 20378 7854 0 sb_8__0_.mem_top_track_14.mem_out\[0\]
rlabel metal1 14214 12750 14214 12750 0 sb_8__0_.mem_top_track_16.ccff_tail
rlabel metal1 15778 5202 15778 5202 0 sb_8__0_.mem_top_track_16.mem_out\[0\]
rlabel metal1 18952 8466 18952 8466 0 sb_8__0_.mem_top_track_18.ccff_tail
rlabel metal2 21114 13124 21114 13124 0 sb_8__0_.mem_top_track_18.mem_out\[0\]
rlabel metal2 21298 8874 21298 8874 0 sb_8__0_.mem_top_track_2.ccff_tail
rlabel metal1 26726 13906 26726 13906 0 sb_8__0_.mem_top_track_2.mem_out\[0\]
rlabel metal1 13754 8364 13754 8364 0 sb_8__0_.mem_top_track_2.mem_out\[1\]
rlabel via2 18722 15317 18722 15317 0 sb_8__0_.mem_top_track_20.ccff_tail
rlabel metal1 18860 14586 18860 14586 0 sb_8__0_.mem_top_track_20.mem_out\[0\]
rlabel metal2 13432 9418 13432 9418 0 sb_8__0_.mem_top_track_22.ccff_tail
rlabel metal1 19320 15878 19320 15878 0 sb_8__0_.mem_top_track_22.mem_out\[0\]
rlabel metal1 14858 6358 14858 6358 0 sb_8__0_.mem_top_track_24.ccff_tail
rlabel metal1 15548 7854 15548 7854 0 sb_8__0_.mem_top_track_24.mem_out\[0\]
rlabel metal1 12098 10472 12098 10472 0 sb_8__0_.mem_top_track_26.ccff_tail
rlabel metal1 13294 11662 13294 11662 0 sb_8__0_.mem_top_track_26.mem_out\[0\]
rlabel metal1 10810 12274 10810 12274 0 sb_8__0_.mem_top_track_28.ccff_tail
rlabel metal1 6578 7922 6578 7922 0 sb_8__0_.mem_top_track_28.mem_out\[0\]
rlabel metal2 6854 11220 6854 11220 0 sb_8__0_.mem_top_track_30.ccff_tail
rlabel metal1 7958 8908 7958 8908 0 sb_8__0_.mem_top_track_30.mem_out\[0\]
rlabel metal2 12558 15249 12558 15249 0 sb_8__0_.mem_top_track_32.ccff_tail
rlabel metal1 8050 12240 8050 12240 0 sb_8__0_.mem_top_track_32.mem_out\[0\]
rlabel metal2 12650 19091 12650 19091 0 sb_8__0_.mem_top_track_34.ccff_tail
rlabel metal2 13340 9350 13340 9350 0 sb_8__0_.mem_top_track_34.mem_out\[0\]
rlabel metal1 10074 20230 10074 20230 0 sb_8__0_.mem_top_track_36.ccff_tail
rlabel metal1 11960 19686 11960 19686 0 sb_8__0_.mem_top_track_36.mem_out\[0\]
rlabel metal2 5566 5933 5566 5933 0 sb_8__0_.mem_top_track_38.ccff_tail
rlabel metal1 8142 15980 8142 15980 0 sb_8__0_.mem_top_track_38.mem_out\[0\]
rlabel metal1 19918 11526 19918 11526 0 sb_8__0_.mem_top_track_4.ccff_tail
rlabel metal1 23230 13804 23230 13804 0 sb_8__0_.mem_top_track_4.mem_out\[0\]
rlabel metal1 19458 6766 19458 6766 0 sb_8__0_.mem_top_track_4.mem_out\[1\]
rlabel metal1 2484 2550 2484 2550 0 sb_8__0_.mem_top_track_40.ccff_tail
rlabel via2 8234 17085 8234 17085 0 sb_8__0_.mem_top_track_40.mem_out\[0\]
rlabel metal1 13892 9350 13892 9350 0 sb_8__0_.mem_top_track_42.ccff_tail
rlabel metal2 13846 11543 13846 11543 0 sb_8__0_.mem_top_track_42.mem_out\[0\]
rlabel metal3 14444 20196 14444 20196 0 sb_8__0_.mem_top_track_44.ccff_tail
rlabel metal1 43746 21964 43746 21964 0 sb_8__0_.mem_top_track_44.mem_out\[0\]
rlabel metal1 15916 20366 15916 20366 0 sb_8__0_.mem_top_track_46.ccff_tail
rlabel metal1 14812 21318 14812 21318 0 sb_8__0_.mem_top_track_46.mem_out\[0\]
rlabel via2 15410 18173 15410 18173 0 sb_8__0_.mem_top_track_48.ccff_tail
rlabel metal1 19872 18190 19872 18190 0 sb_8__0_.mem_top_track_48.mem_out\[0\]
rlabel metal1 19412 18598 19412 18598 0 sb_8__0_.mem_top_track_50.mem_out\[0\]
rlabel metal1 21068 15130 21068 15130 0 sb_8__0_.mem_top_track_6.ccff_tail
rlabel metal1 22080 13362 22080 13362 0 sb_8__0_.mem_top_track_6.mem_out\[0\]
rlabel metal1 17066 11050 17066 11050 0 sb_8__0_.mem_top_track_6.mem_out\[1\]
rlabel metal1 25898 14416 25898 14416 0 sb_8__0_.mem_top_track_8.mem_out\[0\]
rlabel metal1 16238 9044 16238 9044 0 sb_8__0_.mem_top_track_8.mem_out\[1\]
rlabel metal1 14122 17272 14122 17272 0 sb_8__0_.mux_left_track_1.out
rlabel metal1 25254 19822 25254 19822 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 26266 16762 26266 16762 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 21298 18496 21298 18496 0 sb_8__0_.mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 12834 20502 12834 20502 0 sb_8__0_.mux_left_track_11.out
rlabel metal2 12374 24208 12374 24208 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 11638 4794 11638 4794 0 sb_8__0_.mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 28658 15300 28658 15300 0 sb_8__0_.mux_left_track_13.out
rlabel via2 27186 24293 27186 24293 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 15134 21063 15134 21063 0 sb_8__0_.mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21022 17306 21022 17306 0 sb_8__0_.mux_left_track_15.out
rlabel metal1 19918 19686 19918 19686 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 21022 17170 21022 17170 0 sb_8__0_.mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 14674 23137 14674 23137 0 sb_8__0_.mux_left_track_17.out
rlabel via2 18998 20451 18998 20451 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 29026 24191 29026 24191 0 sb_8__0_.mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 9062 2142 9062 2142 0 sb_8__0_.mux_left_track_19.out
rlabel metal2 18630 21862 18630 21862 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22034 13039 22034 13039 0 sb_8__0_.mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 8694 6800 8694 6800 0 sb_8__0_.mux_left_track_29.out
rlabel metal1 23322 19924 23322 19924 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11730 5865 11730 5865 0 sb_8__0_.mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16514 24905 16514 24905 0 sb_8__0_.mux_left_track_3.out
rlabel metal2 17434 20060 17434 20060 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 10994 2652 10994 2652 0 sb_8__0_.mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2208 12138 2208 12138 0 sb_8__0_.mux_left_track_31.out
rlabel metal1 23552 20910 23552 20910 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 19458 7956 19458 7956 0 sb_8__0_.mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal3 23943 1972 23943 1972 0 sb_8__0_.mux_left_track_33.out
rlabel metal1 22356 20978 22356 20978 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34868 18598 34868 18598 0 sb_8__0_.mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 12742 3910 12742 3910 0 sb_8__0_.mux_left_track_35.out
rlabel metal2 27278 23800 27278 23800 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 13110 3111 13110 3111 0 sb_8__0_.mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 22034 2635 22034 2635 0 sb_8__0_.mux_left_track_45.out
rlabel metal1 26634 22202 26634 22202 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23000 2618 23000 2618 0 sb_8__0_.mux_left_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6532 9622 6532 9622 0 sb_8__0_.mux_left_track_47.out
rlabel metal1 26358 20774 26358 20774 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19366 5100 19366 5100 0 sb_8__0_.mux_left_track_47.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 16836 7514 16836 7514 0 sb_8__0_.mux_left_track_49.out
rlabel metal1 26542 16422 26542 16422 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17112 7378 17112 7378 0 sb_8__0_.mux_left_track_49.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 16146 18615 16146 18615 0 sb_8__0_.mux_left_track_5.out
rlabel metal2 17618 21216 17618 21216 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22264 15674 22264 15674 0 sb_8__0_.mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4186 13362 4186 13362 0 sb_8__0_.mux_left_track_51.out
rlabel metal1 22908 17306 22908 17306 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 3634 14960 3634 14960 0 sb_8__0_.mux_left_track_51.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 2714 23630 2714 23630 0 sb_8__0_.mux_left_track_7.out
rlabel metal1 22908 19482 22908 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22862 18938 22862 18938 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21988 19482 21988 19482 0 sb_8__0_.mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 19228 1870 19228 1870 0 sb_8__0_.mux_left_track_9.out
rlabel metal2 15778 21284 15778 21284 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal3 18561 14620 18561 14620 0 sb_8__0_.mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27370 13498 27370 13498 0 sb_8__0_.mux_top_track_0.out
rlabel metal1 28060 18938 28060 18938 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28612 19482 28612 19482 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23782 16660 23782 16660 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 21390 17000 21390 17000 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23598 13294 23598 13294 0 sb_8__0_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33948 18666 33948 18666 0 sb_8__0_.mux_top_track_10.out
rlabel metal1 23368 15334 23368 15334 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23736 14042 23736 14042 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17802 11543 17802 11543 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15088 9146 15088 9146 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 14904 8398 14904 8398 0 sb_8__0_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 41308 20842 41308 20842 0 sb_8__0_.mux_top_track_12.out
rlabel metal2 17986 13855 17986 13855 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 17020 11866 17020 11866 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15502 7208 15502 7208 0 sb_8__0_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 3726 6222 3726 6222 0 sb_8__0_.mux_top_track_14.out
rlabel metal1 17112 12614 17112 12614 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13524 12070 13524 12070 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 4232 6766 4232 6766 0 sb_8__0_.mux_top_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 29486 14042 29486 14042 0 sb_8__0_.mux_top_track_16.out
rlabel metal1 18170 13362 18170 13362 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10534 7514 10534 7514 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 13202 12699 13202 12699 0 sb_8__0_.mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43562 21522 43562 21522 0 sb_8__0_.mux_top_track_18.out
rlabel metal1 19918 15946 19918 15946 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13938 13804 13938 13804 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 17342 4556 17342 4556 0 sb_8__0_.mux_top_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 11408 20570 11408 20570 0 sb_8__0_.mux_top_track_2.out
rlabel metal1 25622 13158 25622 13158 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24978 13498 24978 13498 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24334 13158 24334 13158 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 15824 8602 15824 8602 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal3 15732 13328 15732 13328 0 sb_8__0_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36892 18054 36892 18054 0 sb_8__0_.mux_top_track_20.out
rlabel metal1 15824 15130 15824 15130 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 16790 16150 16790 16150 0 sb_8__0_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 42642 21522 42642 21522 0 sb_8__0_.mux_top_track_22.out
rlabel metal1 14628 15130 14628 15130 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 24610 15028 24610 15028 0 sb_8__0_.mux_top_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34592 17170 34592 17170 0 sb_8__0_.mux_top_track_24.out
rlabel metal1 15226 13838 15226 13838 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 14490 15963 14490 15963 0 sb_8__0_.mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32798 6001 32798 6001 0 sb_8__0_.mux_top_track_26.out
rlabel metal2 12006 12036 12006 12036 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 8418 4182 8418 4182 0 sb_8__0_.mux_top_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20700 714 20700 714 0 sb_8__0_.mux_top_track_28.out
rlabel metal1 10580 8330 10580 8330 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 7130 5270 7130 5270 0 sb_8__0_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38042 17578 38042 17578 0 sb_8__0_.mux_top_track_30.out
rlabel metal2 12006 13600 12006 13600 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39376 20910 39376 20910 0 sb_8__0_.mux_top_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38456 18258 38456 18258 0 sb_8__0_.mux_top_track_32.out
rlabel metal2 12282 16320 12282 16320 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 12742 17816 12742 17816 0 sb_8__0_.mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40894 20026 40894 20026 0 sb_8__0_.mux_top_track_34.out
rlabel metal1 11914 18394 11914 18394 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 42964 20434 42964 20434 0 sb_8__0_.mux_top_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 15134 3298 15134 3298 0 sb_8__0_.mux_top_track_36.out
rlabel metal1 12880 17850 12880 17850 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 9338 21777 9338 21777 0 sb_8__0_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 13386 170 13386 170 0 sb_8__0_.mux_top_track_38.out
rlabel metal2 7590 17272 7590 17272 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 690 17238 690 17238 0 sb_8__0_.mux_top_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 6578 23732 6578 23732 0 sb_8__0_.mux_top_track_4.out
rlabel metal1 22586 10778 22586 10778 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21344 11594 21344 11594 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 21620 10506 21620 10506 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 12006 8687 12006 8687 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal3 15111 19380 15111 19380 0 sb_8__0_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 23046 6562 23046 6562 0 sb_8__0_.mux_top_track_40.out
rlabel metal2 9982 17306 9982 17306 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 21482 7531 21482 7531 0 sb_8__0_.mux_top_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 14858 3077 14858 3077 0 sb_8__0_.mux_top_track_42.out
rlabel metal1 10074 21658 10074 21658 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_0_X
rlabel via2 12742 6069 12742 6069 0 sb_8__0_.mux_top_track_42.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35995 10642 35995 10642 0 sb_8__0_.mux_top_track_44.out
rlabel metal1 17480 18938 17480 18938 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 9246 19448 9246 19448 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35926 17595 35926 17595 0 sb_8__0_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38134 19346 38134 19346 0 sb_8__0_.mux_top_track_46.out
rlabel metal2 16422 19431 16422 19431 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 10626 18394 10626 18394 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36846 19142 36846 19142 0 sb_8__0_.mux_top_track_46.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 5980 2618 5980 2618 0 sb_8__0_.mux_top_track_48.out
rlabel metal1 17250 18394 17250 18394 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 11822 16881 11822 16881 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 42044 20910 42044 20910 0 sb_8__0_.mux_top_track_48.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 43378 24038 43378 24038 0 sb_8__0_.mux_top_track_50.out
rlabel metal1 19550 17782 19550 17782 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 13018 16456 13018 16456 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel via2 42734 23749 42734 23749 0 sb_8__0_.mux_top_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20148 11730 20148 11730 0 sb_8__0_.mux_top_track_6.out
rlabel metal1 22954 16150 22954 16150 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 22954 16218 22954 16218 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20930 16218 20930 16218 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 15502 11951 15502 11951 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19412 16218 19412 16218 0 sb_8__0_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 24656 15980 24656 15980 0 sb_8__0_.mux_top_track_8.out
rlabel metal1 21344 13906 21344 13906 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 21114 13855 21114 13855 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20792 14042 20792 14042 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20194 15334 20194 15334 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 19458 15674 19458 15674 0 sb_8__0_.mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 45126 24463 45126 24463 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_
rlabel metal2 45402 24490 45402 24490 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_
rlabel metal1 46460 22134 46460 22134 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_
rlabel metal2 48898 23494 48898 23494 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_
rlabel metal1 47610 22678 47610 22678 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_
rlabel metal1 47932 21998 47932 21998 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_
rlabel metal2 43562 22967 43562 22967 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_
rlabel metal1 45218 21964 45218 21964 0 top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_
rlabel metal3 48446 21964 48446 21964 0 top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 46782 21301 46782 21301 0 top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 47449 23732 47449 23732 0 top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 48262 24820 48262 24820 0 top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal2 41446 2778 41446 2778 0 top_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal2 44114 2132 44114 2132 0 top_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal2 46782 2098 46782 2098 0 top_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal2 49450 2880 49450 2880 0 top_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 27000
<< end >>
