magic
tech sky130A
magscale 1 2
timestamp 1679321912
<< obsli1 >>
rect 1104 2159 49864 54417
<< obsm1 >>
rect 382 1640 49864 55752
<< metal2 >>
rect 386 56200 442 57000
rect 1122 56200 1178 57000
rect 1858 56200 1914 57000
rect 2594 56200 2650 57000
rect 3330 56200 3386 57000
rect 4066 56200 4122 57000
rect 4802 56200 4858 57000
rect 5538 56200 5594 57000
rect 6274 56200 6330 57000
rect 7010 56200 7066 57000
rect 7746 56200 7802 57000
rect 8482 56200 8538 57000
rect 9218 56200 9274 57000
rect 9954 56200 10010 57000
rect 10690 56200 10746 57000
rect 11426 56200 11482 57000
rect 12162 56200 12218 57000
rect 12898 56200 12954 57000
rect 13634 56200 13690 57000
rect 14370 56200 14426 57000
rect 15106 56200 15162 57000
rect 15842 56200 15898 57000
rect 16578 56200 16634 57000
rect 17314 56200 17370 57000
rect 18050 56200 18106 57000
rect 18786 56200 18842 57000
rect 19522 56200 19578 57000
rect 20258 56200 20314 57000
rect 20994 56200 21050 57000
rect 21730 56200 21786 57000
rect 22466 56200 22522 57000
rect 23202 56200 23258 57000
rect 23938 56200 23994 57000
rect 24674 56200 24730 57000
rect 25410 56200 25466 57000
rect 26146 56200 26202 57000
rect 26882 56200 26938 57000
rect 27618 56200 27674 57000
rect 28354 56200 28410 57000
rect 29090 56200 29146 57000
rect 29826 56200 29882 57000
rect 30562 56200 30618 57000
rect 31298 56200 31354 57000
rect 32034 56200 32090 57000
rect 32770 56200 32826 57000
rect 33506 56200 33562 57000
rect 34242 56200 34298 57000
rect 34978 56200 35034 57000
rect 35714 56200 35770 57000
rect 36450 56200 36506 57000
rect 37186 56200 37242 57000
rect 37922 56200 37978 57000
rect 38658 56200 38714 57000
rect 39394 56200 39450 57000
rect 40130 56200 40186 57000
rect 40866 56200 40922 57000
rect 41602 56200 41658 57000
rect 42338 56200 42394 57000
rect 43074 56200 43130 57000
rect 43810 56200 43866 57000
rect 44546 56200 44602 57000
rect 46754 56200 46810 57000
rect 47490 56200 47546 57000
rect 48226 56200 48282 57000
rect 48962 56200 49018 57000
rect 49698 56200 49754 57000
rect 50434 56200 50490 57000
rect 754 0 810 800
rect 1490 0 1546 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22098 0 22154 800
rect 22834 0 22890 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
rect 49330 0 49386 800
<< obsm2 >>
rect 498 56144 1066 56250
rect 1234 56144 1802 56250
rect 1970 56144 2538 56250
rect 2706 56144 3274 56250
rect 3442 56144 4010 56250
rect 4178 56144 4746 56250
rect 4914 56144 5482 56250
rect 5650 56144 6218 56250
rect 6386 56144 6954 56250
rect 7122 56144 7690 56250
rect 7858 56144 8426 56250
rect 8594 56144 9162 56250
rect 9330 56144 9898 56250
rect 10066 56144 10634 56250
rect 10802 56144 11370 56250
rect 11538 56144 12106 56250
rect 12274 56144 12842 56250
rect 13010 56144 13578 56250
rect 13746 56144 14314 56250
rect 14482 56144 15050 56250
rect 15218 56144 15786 56250
rect 15954 56144 16522 56250
rect 16690 56144 17258 56250
rect 17426 56144 17994 56250
rect 18162 56144 18730 56250
rect 18898 56144 19466 56250
rect 19634 56144 20202 56250
rect 20370 56144 20938 56250
rect 21106 56144 21674 56250
rect 21842 56144 22410 56250
rect 22578 56144 23146 56250
rect 23314 56144 23882 56250
rect 24050 56144 24618 56250
rect 24786 56144 25354 56250
rect 25522 56144 26090 56250
rect 26258 56144 26826 56250
rect 26994 56144 27562 56250
rect 27730 56144 28298 56250
rect 28466 56144 29034 56250
rect 29202 56144 29770 56250
rect 29938 56144 30506 56250
rect 30674 56144 31242 56250
rect 31410 56144 31978 56250
rect 32146 56144 32714 56250
rect 32882 56144 33450 56250
rect 33618 56144 34186 56250
rect 34354 56144 34922 56250
rect 35090 56144 35658 56250
rect 35826 56144 36394 56250
rect 36562 56144 37130 56250
rect 37298 56144 37866 56250
rect 38034 56144 38602 56250
rect 38770 56144 39338 56250
rect 39506 56144 40074 56250
rect 40242 56144 40810 56250
rect 40978 56144 41546 56250
rect 41714 56144 42282 56250
rect 42450 56144 43018 56250
rect 43186 56144 43754 56250
rect 43922 56144 44490 56250
rect 44658 56144 46698 56250
rect 46866 56144 47434 56250
rect 47602 56144 48170 56250
rect 48338 56144 48906 56250
rect 49074 56144 49642 56250
rect 388 856 49752 56144
rect 388 734 698 856
rect 866 734 1434 856
rect 1602 734 2170 856
rect 2338 734 2906 856
rect 3074 734 3642 856
rect 3810 734 4378 856
rect 4546 734 5114 856
rect 5282 734 5850 856
rect 6018 734 6586 856
rect 6754 734 7322 856
rect 7490 734 8058 856
rect 8226 734 8794 856
rect 8962 734 9530 856
rect 9698 734 10266 856
rect 10434 734 11002 856
rect 11170 734 11738 856
rect 11906 734 12474 856
rect 12642 734 13210 856
rect 13378 734 13946 856
rect 14114 734 14682 856
rect 14850 734 15418 856
rect 15586 734 16154 856
rect 16322 734 16890 856
rect 17058 734 17626 856
rect 17794 734 18362 856
rect 18530 734 19098 856
rect 19266 734 19834 856
rect 20002 734 20570 856
rect 20738 734 21306 856
rect 21474 734 22042 856
rect 22210 734 22778 856
rect 22946 734 23514 856
rect 23682 734 24250 856
rect 24418 734 24986 856
rect 25154 734 25722 856
rect 25890 734 26458 856
rect 26626 734 27194 856
rect 27362 734 27930 856
rect 28098 734 28666 856
rect 28834 734 29402 856
rect 29570 734 30138 856
rect 30306 734 30874 856
rect 31042 734 31610 856
rect 31778 734 32346 856
rect 32514 734 33082 856
rect 33250 734 33818 856
rect 33986 734 34554 856
rect 34722 734 35290 856
rect 35458 734 36026 856
rect 36194 734 36762 856
rect 36930 734 37498 856
rect 37666 734 38234 856
rect 38402 734 38970 856
rect 39138 734 39706 856
rect 39874 734 40442 856
rect 40610 734 41178 856
rect 41346 734 41914 856
rect 42082 734 42650 856
rect 42818 734 43386 856
rect 43554 734 44122 856
rect 44290 734 44858 856
rect 45026 734 45594 856
rect 45762 734 46330 856
rect 46498 734 47066 856
rect 47234 734 47802 856
rect 47970 734 48538 856
rect 48706 734 49274 856
rect 49442 734 49752 856
<< metal3 >>
rect 0 54952 800 55072
rect 0 52640 800 52760
rect 50200 52504 51000 52624
rect 50200 51824 51000 51944
rect 50200 51144 51000 51264
rect 0 50328 800 50448
rect 50200 50464 51000 50584
rect 50200 49784 51000 49904
rect 50200 49104 51000 49224
rect 50200 48424 51000 48544
rect 0 48016 800 48136
rect 50200 47744 51000 47864
rect 50200 47064 51000 47184
rect 50200 46384 51000 46504
rect 0 45704 800 45824
rect 50200 45704 51000 45824
rect 50200 45024 51000 45144
rect 50200 44344 51000 44464
rect 50200 43664 51000 43784
rect 0 43392 800 43512
rect 50200 42984 51000 43104
rect 50200 42304 51000 42424
rect 50200 41624 51000 41744
rect 0 41080 800 41200
rect 50200 40944 51000 41064
rect 50200 40264 51000 40384
rect 50200 39584 51000 39704
rect 0 38768 800 38888
rect 50200 38904 51000 39024
rect 50200 38224 51000 38344
rect 50200 37544 51000 37664
rect 50200 36864 51000 36984
rect 0 36456 800 36576
rect 50200 36184 51000 36304
rect 50200 35504 51000 35624
rect 50200 34824 51000 34944
rect 0 34144 800 34264
rect 50200 34144 51000 34264
rect 50200 33464 51000 33584
rect 50200 32784 51000 32904
rect 50200 32104 51000 32224
rect 0 31832 800 31952
rect 50200 31424 51000 31544
rect 50200 30744 51000 30864
rect 50200 30064 51000 30184
rect 0 29520 800 29640
rect 50200 29384 51000 29504
rect 50200 28704 51000 28824
rect 50200 28024 51000 28144
rect 0 27208 800 27328
rect 50200 27344 51000 27464
rect 50200 26664 51000 26784
rect 50200 25984 51000 26104
rect 50200 25304 51000 25424
rect 0 24896 800 25016
rect 50200 24624 51000 24744
rect 50200 23944 51000 24064
rect 50200 23264 51000 23384
rect 0 22584 800 22704
rect 50200 22584 51000 22704
rect 50200 21904 51000 22024
rect 50200 21224 51000 21344
rect 50200 20544 51000 20664
rect 0 20272 800 20392
rect 50200 19864 51000 19984
rect 50200 19184 51000 19304
rect 50200 18504 51000 18624
rect 0 17960 800 18080
rect 50200 17824 51000 17944
rect 50200 17144 51000 17264
rect 50200 16464 51000 16584
rect 0 15648 800 15768
rect 50200 15784 51000 15904
rect 50200 15104 51000 15224
rect 50200 14424 51000 14544
rect 50200 13744 51000 13864
rect 0 13336 800 13456
rect 50200 13064 51000 13184
rect 50200 12384 51000 12504
rect 50200 11704 51000 11824
rect 0 11024 800 11144
rect 50200 11024 51000 11144
rect 50200 10344 51000 10464
rect 50200 9664 51000 9784
rect 50200 8984 51000 9104
rect 0 8712 800 8832
rect 50200 8304 51000 8424
rect 50200 7624 51000 7744
rect 50200 6944 51000 7064
rect 0 6400 800 6520
rect 50200 6264 51000 6384
rect 50200 5584 51000 5704
rect 50200 4904 51000 5024
rect 0 4088 800 4208
rect 50200 4224 51000 4344
rect 0 1776 800 1896
<< obsm3 >>
rect 880 54872 50200 55045
rect 800 52840 50200 54872
rect 880 52704 50200 52840
rect 880 52560 50120 52704
rect 800 52424 50120 52560
rect 800 52024 50200 52424
rect 800 51744 50120 52024
rect 800 51344 50200 51744
rect 800 51064 50120 51344
rect 800 50664 50200 51064
rect 800 50528 50120 50664
rect 880 50384 50120 50528
rect 880 50248 50200 50384
rect 800 49984 50200 50248
rect 800 49704 50120 49984
rect 800 49304 50200 49704
rect 800 49024 50120 49304
rect 800 48624 50200 49024
rect 800 48344 50120 48624
rect 800 48216 50200 48344
rect 880 47944 50200 48216
rect 880 47936 50120 47944
rect 800 47664 50120 47936
rect 800 47264 50200 47664
rect 800 46984 50120 47264
rect 800 46584 50200 46984
rect 800 46304 50120 46584
rect 800 45904 50200 46304
rect 880 45624 50120 45904
rect 800 45224 50200 45624
rect 800 44944 50120 45224
rect 800 44544 50200 44944
rect 800 44264 50120 44544
rect 800 43864 50200 44264
rect 800 43592 50120 43864
rect 880 43584 50120 43592
rect 880 43312 50200 43584
rect 800 43184 50200 43312
rect 800 42904 50120 43184
rect 800 42504 50200 42904
rect 800 42224 50120 42504
rect 800 41824 50200 42224
rect 800 41544 50120 41824
rect 800 41280 50200 41544
rect 880 41144 50200 41280
rect 880 41000 50120 41144
rect 800 40864 50120 41000
rect 800 40464 50200 40864
rect 800 40184 50120 40464
rect 800 39784 50200 40184
rect 800 39504 50120 39784
rect 800 39104 50200 39504
rect 800 38968 50120 39104
rect 880 38824 50120 38968
rect 880 38688 50200 38824
rect 800 38424 50200 38688
rect 800 38144 50120 38424
rect 800 37744 50200 38144
rect 800 37464 50120 37744
rect 800 37064 50200 37464
rect 800 36784 50120 37064
rect 800 36656 50200 36784
rect 880 36384 50200 36656
rect 880 36376 50120 36384
rect 800 36104 50120 36376
rect 800 35704 50200 36104
rect 800 35424 50120 35704
rect 800 35024 50200 35424
rect 800 34744 50120 35024
rect 800 34344 50200 34744
rect 880 34064 50120 34344
rect 800 33664 50200 34064
rect 800 33384 50120 33664
rect 800 32984 50200 33384
rect 800 32704 50120 32984
rect 800 32304 50200 32704
rect 800 32032 50120 32304
rect 880 32024 50120 32032
rect 880 31752 50200 32024
rect 800 31624 50200 31752
rect 800 31344 50120 31624
rect 800 30944 50200 31344
rect 800 30664 50120 30944
rect 800 30264 50200 30664
rect 800 29984 50120 30264
rect 800 29720 50200 29984
rect 880 29584 50200 29720
rect 880 29440 50120 29584
rect 800 29304 50120 29440
rect 800 28904 50200 29304
rect 800 28624 50120 28904
rect 800 28224 50200 28624
rect 800 27944 50120 28224
rect 800 27544 50200 27944
rect 800 27408 50120 27544
rect 880 27264 50120 27408
rect 880 27128 50200 27264
rect 800 26864 50200 27128
rect 800 26584 50120 26864
rect 800 26184 50200 26584
rect 800 25904 50120 26184
rect 800 25504 50200 25904
rect 800 25224 50120 25504
rect 800 25096 50200 25224
rect 880 24824 50200 25096
rect 880 24816 50120 24824
rect 800 24544 50120 24816
rect 800 24144 50200 24544
rect 800 23864 50120 24144
rect 800 23464 50200 23864
rect 800 23184 50120 23464
rect 800 22784 50200 23184
rect 880 22504 50120 22784
rect 800 22104 50200 22504
rect 800 21824 50120 22104
rect 800 21424 50200 21824
rect 800 21144 50120 21424
rect 800 20744 50200 21144
rect 800 20472 50120 20744
rect 880 20464 50120 20472
rect 880 20192 50200 20464
rect 800 20064 50200 20192
rect 800 19784 50120 20064
rect 800 19384 50200 19784
rect 800 19104 50120 19384
rect 800 18704 50200 19104
rect 800 18424 50120 18704
rect 800 18160 50200 18424
rect 880 18024 50200 18160
rect 880 17880 50120 18024
rect 800 17744 50120 17880
rect 800 17344 50200 17744
rect 800 17064 50120 17344
rect 800 16664 50200 17064
rect 800 16384 50120 16664
rect 800 15984 50200 16384
rect 800 15848 50120 15984
rect 880 15704 50120 15848
rect 880 15568 50200 15704
rect 800 15304 50200 15568
rect 800 15024 50120 15304
rect 800 14624 50200 15024
rect 800 14344 50120 14624
rect 800 13944 50200 14344
rect 800 13664 50120 13944
rect 800 13536 50200 13664
rect 880 13264 50200 13536
rect 880 13256 50120 13264
rect 800 12984 50120 13256
rect 800 12584 50200 12984
rect 800 12304 50120 12584
rect 800 11904 50200 12304
rect 800 11624 50120 11904
rect 800 11224 50200 11624
rect 880 10944 50120 11224
rect 800 10544 50200 10944
rect 800 10264 50120 10544
rect 800 9864 50200 10264
rect 800 9584 50120 9864
rect 800 9184 50200 9584
rect 800 8912 50120 9184
rect 880 8904 50120 8912
rect 880 8632 50200 8904
rect 800 8504 50200 8632
rect 800 8224 50120 8504
rect 800 7824 50200 8224
rect 800 7544 50120 7824
rect 800 7144 50200 7544
rect 800 6864 50120 7144
rect 800 6600 50200 6864
rect 880 6464 50200 6600
rect 880 6320 50120 6464
rect 800 6184 50120 6320
rect 800 5784 50200 6184
rect 800 5504 50120 5784
rect 800 5104 50200 5504
rect 800 4824 50120 5104
rect 800 4424 50200 4824
rect 800 4288 50120 4424
rect 880 4144 50120 4288
rect 880 4008 50200 4144
rect 800 1976 50200 4008
rect 880 1803 50200 1976
<< metal4 >>
rect 2944 2128 3264 54448
rect 7944 2128 8264 54448
rect 12944 2128 13264 54448
rect 17944 2128 18264 54448
rect 22944 2128 23264 54448
rect 27944 2128 28264 54448
rect 32944 2128 33264 54448
rect 37944 2128 38264 54448
rect 42944 2128 43264 54448
rect 47944 2128 48264 54448
<< obsm4 >>
rect 22691 2048 22864 44709
rect 23344 2048 27864 44709
rect 28344 2048 32864 44709
rect 33344 2048 37864 44709
rect 38344 2048 40605 44709
rect 22691 1803 40605 2048
<< labels >>
rlabel metal4 s 7944 2128 8264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 17944 2128 18264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 27944 2128 28264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 37944 2128 38264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 47944 2128 48264 54448 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2944 2128 3264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 12944 2128 13264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 22944 2128 23264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 32944 2128 33264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 42944 2128 43264 54448 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 54952 800 55072 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 ccff_head_0
port 4 nsew signal input
rlabel metal3 s 50200 4224 51000 4344 6 ccff_tail
port 5 nsew signal output
rlabel metal2 s 386 56200 442 57000 6 ccff_tail_0
port 6 nsew signal output
rlabel metal3 s 50200 25304 51000 25424 6 chanx_right_in[0]
port 7 nsew signal input
rlabel metal3 s 50200 32104 51000 32224 6 chanx_right_in[10]
port 8 nsew signal input
rlabel metal3 s 50200 32784 51000 32904 6 chanx_right_in[11]
port 9 nsew signal input
rlabel metal3 s 50200 33464 51000 33584 6 chanx_right_in[12]
port 10 nsew signal input
rlabel metal3 s 50200 34144 51000 34264 6 chanx_right_in[13]
port 11 nsew signal input
rlabel metal3 s 50200 34824 51000 34944 6 chanx_right_in[14]
port 12 nsew signal input
rlabel metal3 s 50200 35504 51000 35624 6 chanx_right_in[15]
port 13 nsew signal input
rlabel metal3 s 50200 36184 51000 36304 6 chanx_right_in[16]
port 14 nsew signal input
rlabel metal3 s 50200 36864 51000 36984 6 chanx_right_in[17]
port 15 nsew signal input
rlabel metal3 s 50200 37544 51000 37664 6 chanx_right_in[18]
port 16 nsew signal input
rlabel metal3 s 50200 38224 51000 38344 6 chanx_right_in[19]
port 17 nsew signal input
rlabel metal3 s 50200 25984 51000 26104 6 chanx_right_in[1]
port 18 nsew signal input
rlabel metal3 s 50200 38904 51000 39024 6 chanx_right_in[20]
port 19 nsew signal input
rlabel metal3 s 50200 39584 51000 39704 6 chanx_right_in[21]
port 20 nsew signal input
rlabel metal3 s 50200 40264 51000 40384 6 chanx_right_in[22]
port 21 nsew signal input
rlabel metal3 s 50200 40944 51000 41064 6 chanx_right_in[23]
port 22 nsew signal input
rlabel metal3 s 50200 41624 51000 41744 6 chanx_right_in[24]
port 23 nsew signal input
rlabel metal3 s 50200 42304 51000 42424 6 chanx_right_in[25]
port 24 nsew signal input
rlabel metal3 s 50200 42984 51000 43104 6 chanx_right_in[26]
port 25 nsew signal input
rlabel metal3 s 50200 43664 51000 43784 6 chanx_right_in[27]
port 26 nsew signal input
rlabel metal3 s 50200 44344 51000 44464 6 chanx_right_in[28]
port 27 nsew signal input
rlabel metal3 s 50200 45024 51000 45144 6 chanx_right_in[29]
port 28 nsew signal input
rlabel metal3 s 50200 26664 51000 26784 6 chanx_right_in[2]
port 29 nsew signal input
rlabel metal3 s 50200 27344 51000 27464 6 chanx_right_in[3]
port 30 nsew signal input
rlabel metal3 s 50200 28024 51000 28144 6 chanx_right_in[4]
port 31 nsew signal input
rlabel metal3 s 50200 28704 51000 28824 6 chanx_right_in[5]
port 32 nsew signal input
rlabel metal3 s 50200 29384 51000 29504 6 chanx_right_in[6]
port 33 nsew signal input
rlabel metal3 s 50200 30064 51000 30184 6 chanx_right_in[7]
port 34 nsew signal input
rlabel metal3 s 50200 30744 51000 30864 6 chanx_right_in[8]
port 35 nsew signal input
rlabel metal3 s 50200 31424 51000 31544 6 chanx_right_in[9]
port 36 nsew signal input
rlabel metal3 s 50200 4904 51000 5024 6 chanx_right_out[0]
port 37 nsew signal output
rlabel metal3 s 50200 11704 51000 11824 6 chanx_right_out[10]
port 38 nsew signal output
rlabel metal3 s 50200 12384 51000 12504 6 chanx_right_out[11]
port 39 nsew signal output
rlabel metal3 s 50200 13064 51000 13184 6 chanx_right_out[12]
port 40 nsew signal output
rlabel metal3 s 50200 13744 51000 13864 6 chanx_right_out[13]
port 41 nsew signal output
rlabel metal3 s 50200 14424 51000 14544 6 chanx_right_out[14]
port 42 nsew signal output
rlabel metal3 s 50200 15104 51000 15224 6 chanx_right_out[15]
port 43 nsew signal output
rlabel metal3 s 50200 15784 51000 15904 6 chanx_right_out[16]
port 44 nsew signal output
rlabel metal3 s 50200 16464 51000 16584 6 chanx_right_out[17]
port 45 nsew signal output
rlabel metal3 s 50200 17144 51000 17264 6 chanx_right_out[18]
port 46 nsew signal output
rlabel metal3 s 50200 17824 51000 17944 6 chanx_right_out[19]
port 47 nsew signal output
rlabel metal3 s 50200 5584 51000 5704 6 chanx_right_out[1]
port 48 nsew signal output
rlabel metal3 s 50200 18504 51000 18624 6 chanx_right_out[20]
port 49 nsew signal output
rlabel metal3 s 50200 19184 51000 19304 6 chanx_right_out[21]
port 50 nsew signal output
rlabel metal3 s 50200 19864 51000 19984 6 chanx_right_out[22]
port 51 nsew signal output
rlabel metal3 s 50200 20544 51000 20664 6 chanx_right_out[23]
port 52 nsew signal output
rlabel metal3 s 50200 21224 51000 21344 6 chanx_right_out[24]
port 53 nsew signal output
rlabel metal3 s 50200 21904 51000 22024 6 chanx_right_out[25]
port 54 nsew signal output
rlabel metal3 s 50200 22584 51000 22704 6 chanx_right_out[26]
port 55 nsew signal output
rlabel metal3 s 50200 23264 51000 23384 6 chanx_right_out[27]
port 56 nsew signal output
rlabel metal3 s 50200 23944 51000 24064 6 chanx_right_out[28]
port 57 nsew signal output
rlabel metal3 s 50200 24624 51000 24744 6 chanx_right_out[29]
port 58 nsew signal output
rlabel metal3 s 50200 6264 51000 6384 6 chanx_right_out[2]
port 59 nsew signal output
rlabel metal3 s 50200 6944 51000 7064 6 chanx_right_out[3]
port 60 nsew signal output
rlabel metal3 s 50200 7624 51000 7744 6 chanx_right_out[4]
port 61 nsew signal output
rlabel metal3 s 50200 8304 51000 8424 6 chanx_right_out[5]
port 62 nsew signal output
rlabel metal3 s 50200 8984 51000 9104 6 chanx_right_out[6]
port 63 nsew signal output
rlabel metal3 s 50200 9664 51000 9784 6 chanx_right_out[7]
port 64 nsew signal output
rlabel metal3 s 50200 10344 51000 10464 6 chanx_right_out[8]
port 65 nsew signal output
rlabel metal3 s 50200 11024 51000 11144 6 chanx_right_out[9]
port 66 nsew signal output
rlabel metal2 s 754 0 810 800 6 chany_bottom_in[0]
port 67 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[10]
port 68 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 chany_bottom_in[11]
port 69 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 70 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[13]
port 71 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[14]
port 72 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[15]
port 73 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_in[16]
port 74 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_in[17]
port 75 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_in[18]
port 76 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in[19]
port 77 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_in[1]
port 78 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_in[20]
port 79 nsew signal input
rlabel metal2 s 16210 0 16266 800 6 chany_bottom_in[21]
port 80 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in[22]
port 81 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_in[23]
port 82 nsew signal input
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_in[24]
port 83 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_in[25]
port 84 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_in[26]
port 85 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_in[27]
port 86 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_in[28]
port 87 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_in[29]
port 88 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_in[2]
port 89 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 chany_bottom_in[3]
port 90 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[4]
port 91 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_in[5]
port 92 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[6]
port 93 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[7]
port 94 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_in[8]
port 95 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[9]
port 96 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 chany_bottom_out[0]
port 97 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 chany_bottom_out[10]
port 98 nsew signal output
rlabel metal2 s 30930 0 30986 800 6 chany_bottom_out[11]
port 99 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 chany_bottom_out[12]
port 100 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 chany_bottom_out[13]
port 101 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 chany_bottom_out[14]
port 102 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 chany_bottom_out[15]
port 103 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 chany_bottom_out[16]
port 104 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 chany_bottom_out[17]
port 105 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 chany_bottom_out[18]
port 106 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 chany_bottom_out[19]
port 107 nsew signal output
rlabel metal2 s 23570 0 23626 800 6 chany_bottom_out[1]
port 108 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 chany_bottom_out[20]
port 109 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 chany_bottom_out[21]
port 110 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 chany_bottom_out[22]
port 111 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 chany_bottom_out[23]
port 112 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 chany_bottom_out[24]
port 113 nsew signal output
rlabel metal2 s 41234 0 41290 800 6 chany_bottom_out[25]
port 114 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 chany_bottom_out[26]
port 115 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 chany_bottom_out[27]
port 116 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 chany_bottom_out[28]
port 117 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 chany_bottom_out[29]
port 118 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 chany_bottom_out[2]
port 119 nsew signal output
rlabel metal2 s 25042 0 25098 800 6 chany_bottom_out[3]
port 120 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 chany_bottom_out[4]
port 121 nsew signal output
rlabel metal2 s 26514 0 26570 800 6 chany_bottom_out[5]
port 122 nsew signal output
rlabel metal2 s 27250 0 27306 800 6 chany_bottom_out[6]
port 123 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 chany_bottom_out[7]
port 124 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 chany_bottom_out[8]
port 125 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 chany_bottom_out[9]
port 126 nsew signal output
rlabel metal2 s 23202 56200 23258 57000 6 chany_top_in_0[0]
port 127 nsew signal input
rlabel metal2 s 30562 56200 30618 57000 6 chany_top_in_0[10]
port 128 nsew signal input
rlabel metal2 s 31298 56200 31354 57000 6 chany_top_in_0[11]
port 129 nsew signal input
rlabel metal2 s 32034 56200 32090 57000 6 chany_top_in_0[12]
port 130 nsew signal input
rlabel metal2 s 32770 56200 32826 57000 6 chany_top_in_0[13]
port 131 nsew signal input
rlabel metal2 s 33506 56200 33562 57000 6 chany_top_in_0[14]
port 132 nsew signal input
rlabel metal2 s 34242 56200 34298 57000 6 chany_top_in_0[15]
port 133 nsew signal input
rlabel metal2 s 34978 56200 35034 57000 6 chany_top_in_0[16]
port 134 nsew signal input
rlabel metal2 s 35714 56200 35770 57000 6 chany_top_in_0[17]
port 135 nsew signal input
rlabel metal2 s 36450 56200 36506 57000 6 chany_top_in_0[18]
port 136 nsew signal input
rlabel metal2 s 37186 56200 37242 57000 6 chany_top_in_0[19]
port 137 nsew signal input
rlabel metal2 s 23938 56200 23994 57000 6 chany_top_in_0[1]
port 138 nsew signal input
rlabel metal2 s 37922 56200 37978 57000 6 chany_top_in_0[20]
port 139 nsew signal input
rlabel metal2 s 38658 56200 38714 57000 6 chany_top_in_0[21]
port 140 nsew signal input
rlabel metal2 s 39394 56200 39450 57000 6 chany_top_in_0[22]
port 141 nsew signal input
rlabel metal2 s 40130 56200 40186 57000 6 chany_top_in_0[23]
port 142 nsew signal input
rlabel metal2 s 40866 56200 40922 57000 6 chany_top_in_0[24]
port 143 nsew signal input
rlabel metal2 s 41602 56200 41658 57000 6 chany_top_in_0[25]
port 144 nsew signal input
rlabel metal2 s 42338 56200 42394 57000 6 chany_top_in_0[26]
port 145 nsew signal input
rlabel metal2 s 43074 56200 43130 57000 6 chany_top_in_0[27]
port 146 nsew signal input
rlabel metal2 s 43810 56200 43866 57000 6 chany_top_in_0[28]
port 147 nsew signal input
rlabel metal2 s 44546 56200 44602 57000 6 chany_top_in_0[29]
port 148 nsew signal input
rlabel metal2 s 24674 56200 24730 57000 6 chany_top_in_0[2]
port 149 nsew signal input
rlabel metal2 s 25410 56200 25466 57000 6 chany_top_in_0[3]
port 150 nsew signal input
rlabel metal2 s 26146 56200 26202 57000 6 chany_top_in_0[4]
port 151 nsew signal input
rlabel metal2 s 26882 56200 26938 57000 6 chany_top_in_0[5]
port 152 nsew signal input
rlabel metal2 s 27618 56200 27674 57000 6 chany_top_in_0[6]
port 153 nsew signal input
rlabel metal2 s 28354 56200 28410 57000 6 chany_top_in_0[7]
port 154 nsew signal input
rlabel metal2 s 29090 56200 29146 57000 6 chany_top_in_0[8]
port 155 nsew signal input
rlabel metal2 s 29826 56200 29882 57000 6 chany_top_in_0[9]
port 156 nsew signal input
rlabel metal2 s 1122 56200 1178 57000 6 chany_top_out_0[0]
port 157 nsew signal output
rlabel metal2 s 8482 56200 8538 57000 6 chany_top_out_0[10]
port 158 nsew signal output
rlabel metal2 s 9218 56200 9274 57000 6 chany_top_out_0[11]
port 159 nsew signal output
rlabel metal2 s 9954 56200 10010 57000 6 chany_top_out_0[12]
port 160 nsew signal output
rlabel metal2 s 10690 56200 10746 57000 6 chany_top_out_0[13]
port 161 nsew signal output
rlabel metal2 s 11426 56200 11482 57000 6 chany_top_out_0[14]
port 162 nsew signal output
rlabel metal2 s 12162 56200 12218 57000 6 chany_top_out_0[15]
port 163 nsew signal output
rlabel metal2 s 12898 56200 12954 57000 6 chany_top_out_0[16]
port 164 nsew signal output
rlabel metal2 s 13634 56200 13690 57000 6 chany_top_out_0[17]
port 165 nsew signal output
rlabel metal2 s 14370 56200 14426 57000 6 chany_top_out_0[18]
port 166 nsew signal output
rlabel metal2 s 15106 56200 15162 57000 6 chany_top_out_0[19]
port 167 nsew signal output
rlabel metal2 s 1858 56200 1914 57000 6 chany_top_out_0[1]
port 168 nsew signal output
rlabel metal2 s 15842 56200 15898 57000 6 chany_top_out_0[20]
port 169 nsew signal output
rlabel metal2 s 16578 56200 16634 57000 6 chany_top_out_0[21]
port 170 nsew signal output
rlabel metal2 s 17314 56200 17370 57000 6 chany_top_out_0[22]
port 171 nsew signal output
rlabel metal2 s 18050 56200 18106 57000 6 chany_top_out_0[23]
port 172 nsew signal output
rlabel metal2 s 18786 56200 18842 57000 6 chany_top_out_0[24]
port 173 nsew signal output
rlabel metal2 s 19522 56200 19578 57000 6 chany_top_out_0[25]
port 174 nsew signal output
rlabel metal2 s 20258 56200 20314 57000 6 chany_top_out_0[26]
port 175 nsew signal output
rlabel metal2 s 20994 56200 21050 57000 6 chany_top_out_0[27]
port 176 nsew signal output
rlabel metal2 s 21730 56200 21786 57000 6 chany_top_out_0[28]
port 177 nsew signal output
rlabel metal2 s 22466 56200 22522 57000 6 chany_top_out_0[29]
port 178 nsew signal output
rlabel metal2 s 2594 56200 2650 57000 6 chany_top_out_0[2]
port 179 nsew signal output
rlabel metal2 s 3330 56200 3386 57000 6 chany_top_out_0[3]
port 180 nsew signal output
rlabel metal2 s 4066 56200 4122 57000 6 chany_top_out_0[4]
port 181 nsew signal output
rlabel metal2 s 4802 56200 4858 57000 6 chany_top_out_0[5]
port 182 nsew signal output
rlabel metal2 s 5538 56200 5594 57000 6 chany_top_out_0[6]
port 183 nsew signal output
rlabel metal2 s 6274 56200 6330 57000 6 chany_top_out_0[7]
port 184 nsew signal output
rlabel metal2 s 7010 56200 7066 57000 6 chany_top_out_0[8]
port 185 nsew signal output
rlabel metal2 s 7746 56200 7802 57000 6 chany_top_out_0[9]
port 186 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 gfpga_pad_io_soc_dir[0]
port 187 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 gfpga_pad_io_soc_dir[1]
port 188 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 gfpga_pad_io_soc_dir[2]
port 189 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 gfpga_pad_io_soc_dir[3]
port 190 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 gfpga_pad_io_soc_in[0]
port 191 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 gfpga_pad_io_soc_in[1]
port 192 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 gfpga_pad_io_soc_in[2]
port 193 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 gfpga_pad_io_soc_in[3]
port 194 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 gfpga_pad_io_soc_out[0]
port 195 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 gfpga_pad_io_soc_out[1]
port 196 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 gfpga_pad_io_soc_out[2]
port 197 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 gfpga_pad_io_soc_out[3]
port 198 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 isol_n
port 199 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 prog_clk
port 200 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 prog_reset_bottom_in
port 201 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 prog_reset_bottom_out
port 202 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 prog_reset_left_in
port 203 nsew signal input
rlabel metal3 s 50200 45704 51000 45824 6 prog_reset_right_out
port 204 nsew signal output
rlabel metal2 s 47490 56200 47546 57000 6 prog_reset_top_in
port 205 nsew signal input
rlabel metal2 s 46754 56200 46810 57000 6 prog_reset_top_out
port 206 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 reset_bottom_in
port 207 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 reset_bottom_out
port 208 nsew signal output
rlabel metal3 s 50200 46384 51000 46504 6 reset_right_in
port 209 nsew signal input
rlabel metal2 s 48962 56200 49018 57000 6 reset_top_in
port 210 nsew signal input
rlabel metal2 s 48226 56200 48282 57000 6 reset_top_out
port 211 nsew signal output
rlabel metal3 s 50200 47064 51000 47184 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 212 nsew signal input
rlabel metal3 s 50200 47744 51000 47864 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 213 nsew signal input
rlabel metal3 s 50200 48424 51000 48544 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 214 nsew signal input
rlabel metal3 s 50200 49104 51000 49224 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 215 nsew signal input
rlabel metal3 s 50200 49784 51000 49904 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 216 nsew signal input
rlabel metal3 s 50200 50464 51000 50584 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 217 nsew signal input
rlabel metal3 s 50200 51144 51000 51264 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 218 nsew signal input
rlabel metal3 s 50200 51824 51000 51944 6 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 219 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 right_width_0_height_0_subtile_0__pin_inpad_0_
port 220 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 right_width_0_height_0_subtile_1__pin_inpad_0_
port 221 nsew signal output
rlabel metal3 s 0 8712 800 8832 6 right_width_0_height_0_subtile_2__pin_inpad_0_
port 222 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 right_width_0_height_0_subtile_3__pin_inpad_0_
port 223 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 test_enable_bottom_in
port 224 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 test_enable_bottom_out
port 225 nsew signal output
rlabel metal3 s 50200 52504 51000 52624 6 test_enable_right_in
port 226 nsew signal input
rlabel metal2 s 50434 56200 50490 57000 6 test_enable_top_in
port 227 nsew signal input
rlabel metal2 s 49698 56200 49754 57000 6 test_enable_top_out
port 228 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 229 nsew signal input
rlabel metal3 s 0 48016 800 48136 6 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 230 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 231 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 232 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 51000 57000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3101854
string GDS_FILE /home/hosni/OpenFPGA/clear/openlane/left_tile/runs/23_03_20_07_16/results/signoff/left_tile.magic.gds
string GDS_START 175900
<< end >>

