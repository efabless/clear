magic
tech sky130A
magscale 1 2
timestamp 1625783863
<< locali >>
rect 11989 20315 12023 20417
rect 12449 20383 12483 20485
rect 12541 20315 12575 20417
rect 15301 20315 15335 20553
rect 15485 19703 15519 19873
rect 7113 19159 7147 19397
rect 13369 19295 13403 19465
rect 9873 19159 9907 19261
rect 11805 19159 11839 19261
rect 13461 19159 13495 19261
rect 15025 19159 15059 19329
rect 11805 18819 11839 18921
rect 17509 18819 17543 18921
rect 17785 18207 17819 18309
rect 9137 16983 9171 17153
rect 9229 17119 9263 17289
rect 12633 16983 12667 17221
rect 9781 16643 9815 16745
rect 14473 16575 14507 16745
rect 8677 16031 8711 16201
rect 18153 14943 18187 15113
rect 10517 14807 10551 14909
rect 14197 14467 14231 14569
rect 14197 14433 14289 14467
rect 11437 12631 11471 12937
rect 14289 12631 14323 12937
rect 8493 11067 8527 11237
rect 16497 10999 16531 11101
rect 9229 9911 9263 10217
rect 10701 10047 10735 10217
rect 12265 10047 12299 10149
rect 16129 9979 16163 10217
rect 17693 9911 17727 10149
rect 11805 9367 11839 9469
rect 13921 9435 13955 9537
rect 16129 8891 16163 9129
rect 19625 8483 19659 8585
rect 13645 8279 13679 8449
rect 10149 7803 10183 8041
rect 12449 7327 12483 7497
rect 11989 7191 12023 7293
rect 11437 6715 11471 6885
rect 9137 6103 9171 6409
rect 11989 6103 12023 6273
rect 9965 5015 9999 5117
rect 10425 5015 10459 5321
rect 10517 5151 10551 5253
rect 11253 4539 11287 4709
rect 19717 4675 19751 4777
rect 9505 4063 9539 4233
rect 11805 3927 11839 4029
rect 7941 3383 7975 3689
rect 9689 3587 9723 3689
rect 8861 3383 8895 3553
rect 7849 2839 7883 3009
rect 10609 2975 10643 3145
rect 15025 2839 15059 3009
rect 16773 2907 16807 3077
rect 19625 2907 19659 3009
rect 11897 2363 11931 2601
rect 22017 1411 22051 2533
rect 22109 1479 22143 2465
<< viali >>
rect 1593 20553 1627 20587
rect 15301 20553 15335 20587
rect 16221 20553 16255 20587
rect 4353 20485 4387 20519
rect 12081 20485 12115 20519
rect 12449 20485 12483 20519
rect 12633 20485 12667 20519
rect 13185 20485 13219 20519
rect 13737 20485 13771 20519
rect 2237 20417 2271 20451
rect 3341 20417 3375 20451
rect 5549 20417 5583 20451
rect 11989 20417 12023 20451
rect 2513 20349 2547 20383
rect 3157 20349 3191 20383
rect 4169 20349 4203 20383
rect 5365 20349 5399 20383
rect 6009 20349 6043 20383
rect 6837 20349 6871 20383
rect 7665 20349 7699 20383
rect 8217 20349 8251 20383
rect 8677 20349 8711 20383
rect 9597 20349 9631 20383
rect 10701 20349 10735 20383
rect 12265 20349 12299 20383
rect 12449 20349 12483 20383
rect 12541 20417 12575 20451
rect 14565 20417 14599 20451
rect 2053 20281 2087 20315
rect 4721 20281 4755 20315
rect 4905 20281 4939 20315
rect 7021 20281 7055 20315
rect 7849 20281 7883 20315
rect 10057 20281 10091 20315
rect 10241 20281 10275 20315
rect 10517 20281 10551 20315
rect 11253 20281 11287 20315
rect 11989 20281 12023 20315
rect 15025 20349 15059 20383
rect 16865 20485 16899 20519
rect 17877 20485 17911 20519
rect 18429 20485 18463 20519
rect 18981 20485 19015 20519
rect 19533 20485 19567 20519
rect 15761 20417 15795 20451
rect 20085 20349 20119 20383
rect 12541 20281 12575 20315
rect 12817 20281 12851 20315
rect 13369 20281 13403 20315
rect 13921 20281 13955 20315
rect 15209 20281 15243 20315
rect 15301 20281 15335 20315
rect 15577 20281 15611 20315
rect 16129 20281 16163 20315
rect 16681 20281 16715 20315
rect 17693 20281 17727 20315
rect 18245 20281 18279 20315
rect 18797 20281 18831 20315
rect 19349 20281 19383 20315
rect 20637 20281 20671 20315
rect 20821 20281 20855 20315
rect 21189 20281 21223 20315
rect 21373 20281 21407 20315
rect 2697 20213 2731 20247
rect 5917 20213 5951 20247
rect 8309 20213 8343 20247
rect 8861 20213 8895 20247
rect 9505 20213 9539 20247
rect 11161 20213 11195 20247
rect 17233 20213 17267 20247
rect 20269 20213 20303 20247
rect 2329 20009 2363 20043
rect 3433 20009 3467 20043
rect 3893 20009 3927 20043
rect 4353 20009 4387 20043
rect 4905 20009 4939 20043
rect 5825 20009 5859 20043
rect 7849 20009 7883 20043
rect 8309 20009 8343 20043
rect 8769 20009 8803 20043
rect 9597 20009 9631 20043
rect 13829 20009 13863 20043
rect 18153 20009 18187 20043
rect 19165 20009 19199 20043
rect 10149 19941 10183 19975
rect 10241 19941 10275 19975
rect 13093 19941 13127 19975
rect 14565 19941 14599 19975
rect 15117 19941 15151 19975
rect 15301 19941 15335 19975
rect 15669 19941 15703 19975
rect 16221 19941 16255 19975
rect 16405 19941 16439 19975
rect 16773 19941 16807 19975
rect 17325 19941 17359 19975
rect 19809 19941 19843 19975
rect 20361 19941 20395 19975
rect 1685 19873 1719 19907
rect 2145 19873 2179 19907
rect 2605 19873 2639 19907
rect 4721 19873 4755 19907
rect 6101 19873 6135 19907
rect 6561 19873 6595 19907
rect 7021 19873 7055 19907
rect 7665 19873 7699 19907
rect 8125 19873 8159 19907
rect 8585 19873 8619 19907
rect 9413 19873 9447 19907
rect 11233 19873 11267 19907
rect 13185 19873 13219 19907
rect 14013 19873 14047 19907
rect 14749 19873 14783 19907
rect 15485 19873 15519 19907
rect 15853 19873 15887 19907
rect 16957 19873 16991 19907
rect 17509 19873 17543 19907
rect 17969 19873 18003 19907
rect 18521 19873 18555 19907
rect 19073 19873 19107 19907
rect 19993 19873 20027 19907
rect 20545 19873 20579 19907
rect 21189 19873 21223 19907
rect 3065 19805 3099 19839
rect 5457 19805 5491 19839
rect 10057 19805 10091 19839
rect 10977 19805 11011 19839
rect 13001 19805 13035 19839
rect 2789 19737 2823 19771
rect 7205 19737 7239 19771
rect 21373 19737 21407 19771
rect 1777 19669 1811 19703
rect 6285 19669 6319 19703
rect 6745 19669 6779 19703
rect 10609 19669 10643 19703
rect 12357 19669 12391 19703
rect 13553 19669 13587 19703
rect 15485 19669 15519 19703
rect 18613 19669 18647 19703
rect 1961 19465 1995 19499
rect 2513 19465 2547 19499
rect 4997 19465 5031 19499
rect 6561 19465 6595 19499
rect 13277 19465 13311 19499
rect 13369 19465 13403 19499
rect 18613 19465 18647 19499
rect 7113 19397 7147 19431
rect 9689 19397 9723 19431
rect 1409 19261 1443 19295
rect 5641 19261 5675 19295
rect 4353 19193 4387 19227
rect 6101 19193 6135 19227
rect 15025 19329 15059 19363
rect 15301 19329 15335 19363
rect 7205 19261 7239 19295
rect 7665 19261 7699 19295
rect 8125 19261 8159 19295
rect 8585 19261 8619 19295
rect 9045 19261 9079 19295
rect 9505 19261 9539 19295
rect 9873 19261 9907 19295
rect 9965 19261 9999 19295
rect 11805 19261 11839 19295
rect 11897 19261 11931 19295
rect 13369 19261 13403 19295
rect 13461 19261 13495 19295
rect 13553 19261 13587 19295
rect 13809 19261 13843 19295
rect 10232 19193 10266 19227
rect 12164 19193 12198 19227
rect 4721 19125 4755 19159
rect 7113 19125 7147 19159
rect 7389 19125 7423 19159
rect 7849 19125 7883 19159
rect 8309 19125 8343 19159
rect 8769 19125 8803 19159
rect 9229 19125 9263 19159
rect 9873 19125 9907 19159
rect 11345 19125 11379 19159
rect 11805 19125 11839 19159
rect 16957 19261 16991 19295
rect 17509 19261 17543 19295
rect 17969 19261 18003 19295
rect 18429 19261 18463 19295
rect 18889 19261 18923 19295
rect 19349 19261 19383 19295
rect 20637 19261 20671 19295
rect 21189 19261 21223 19295
rect 15485 19193 15519 19227
rect 15577 19193 15611 19227
rect 16221 19193 16255 19227
rect 19993 19193 20027 19227
rect 21373 19193 21407 19227
rect 13461 19125 13495 19159
rect 14933 19125 14967 19159
rect 15025 19125 15059 19159
rect 15945 19125 15979 19159
rect 17693 19125 17727 19159
rect 18153 19125 18187 19159
rect 19073 19125 19107 19159
rect 19533 19125 19567 19159
rect 6009 18921 6043 18955
rect 7297 18921 7331 18955
rect 8309 18921 8343 18955
rect 10701 18921 10735 18955
rect 11253 18921 11287 18955
rect 11713 18921 11747 18955
rect 11805 18921 11839 18955
rect 12449 18921 12483 18955
rect 13461 18921 13495 18955
rect 13921 18921 13955 18955
rect 16589 18921 16623 18955
rect 17509 18921 17543 18955
rect 17693 18921 17727 18955
rect 19717 18921 19751 18955
rect 20177 18921 20211 18955
rect 4997 18853 5031 18887
rect 6929 18853 6963 18887
rect 9566 18853 9600 18887
rect 14810 18853 14844 18887
rect 20637 18853 20671 18887
rect 20821 18853 20855 18887
rect 7665 18785 7699 18819
rect 8125 18785 8159 18819
rect 8585 18785 8619 18819
rect 11345 18785 11379 18819
rect 11805 18785 11839 18819
rect 12357 18785 12391 18819
rect 13001 18785 13035 18819
rect 13645 18785 13679 18819
rect 14565 18785 14599 18819
rect 17417 18785 17451 18819
rect 17509 18785 17543 18819
rect 17877 18785 17911 18819
rect 18153 18785 18187 18819
rect 18613 18785 18647 18819
rect 19073 18785 19107 18819
rect 20085 18785 20119 18819
rect 21189 18785 21223 18819
rect 5733 18717 5767 18751
rect 6469 18717 6503 18751
rect 9321 18717 9355 18751
rect 11161 18717 11195 18751
rect 12541 18717 12575 18751
rect 16681 18717 16715 18751
rect 16773 18717 16807 18751
rect 4629 18649 4663 18683
rect 5365 18649 5399 18683
rect 7849 18649 7883 18683
rect 15945 18649 15979 18683
rect 17233 18649 17267 18683
rect 18797 18649 18831 18683
rect 21373 18649 21407 18683
rect 4261 18581 4295 18615
rect 8769 18581 8803 18615
rect 11989 18581 12023 18615
rect 16221 18581 16255 18615
rect 18337 18581 18371 18615
rect 19257 18581 19291 18615
rect 6653 18377 6687 18411
rect 14841 18377 14875 18411
rect 17601 18377 17635 18411
rect 9045 18309 9079 18343
rect 10885 18309 10919 18343
rect 17785 18309 17819 18343
rect 5365 18241 5399 18275
rect 9965 18241 9999 18275
rect 12357 18241 12391 18275
rect 12449 18241 12483 18275
rect 13737 18241 13771 18275
rect 14197 18241 14231 18275
rect 14381 18241 14415 18275
rect 17877 18241 17911 18275
rect 19625 18241 19659 18275
rect 19809 18241 19843 18275
rect 7665 18173 7699 18207
rect 10701 18173 10735 18207
rect 11161 18173 11195 18207
rect 13553 18173 13587 18207
rect 15209 18173 15243 18207
rect 15476 18173 15510 18207
rect 17049 18173 17083 18207
rect 17417 18173 17451 18207
rect 17785 18173 17819 18207
rect 20637 18173 20671 18207
rect 4997 18105 5031 18139
rect 7932 18105 7966 18139
rect 13461 18105 13495 18139
rect 18144 18105 18178 18139
rect 21189 18105 21223 18139
rect 21373 18105 21407 18139
rect 5641 18037 5675 18071
rect 6101 18037 6135 18071
rect 7021 18037 7055 18071
rect 7389 18037 7423 18071
rect 9413 18037 9447 18071
rect 9781 18037 9815 18071
rect 9873 18037 9907 18071
rect 11345 18037 11379 18071
rect 11897 18037 11931 18071
rect 12265 18037 12299 18071
rect 13093 18037 13127 18071
rect 14473 18037 14507 18071
rect 16589 18037 16623 18071
rect 19257 18037 19291 18071
rect 19901 18037 19935 18071
rect 20269 18037 20303 18071
rect 20729 18037 20763 18071
rect 6009 17833 6043 17867
rect 6837 17833 6871 17867
rect 7849 17833 7883 17867
rect 8769 17833 8803 17867
rect 9321 17833 9355 17867
rect 12357 17833 12391 17867
rect 13277 17833 13311 17867
rect 13737 17833 13771 17867
rect 15025 17833 15059 17867
rect 18981 17833 19015 17867
rect 20177 17833 20211 17867
rect 13369 17765 13403 17799
rect 15577 17765 15611 17799
rect 17846 17765 17880 17799
rect 8585 17697 8619 17731
rect 10434 17697 10468 17731
rect 11069 17697 11103 17731
rect 11529 17697 11563 17731
rect 14933 17697 14967 17731
rect 17058 17697 17092 17731
rect 17325 17697 17359 17731
rect 17601 17697 17635 17731
rect 21189 17697 21223 17731
rect 6469 17629 6503 17663
rect 7573 17629 7607 17663
rect 7757 17629 7791 17663
rect 10701 17629 10735 17663
rect 12449 17629 12483 17663
rect 12541 17629 12575 17663
rect 13185 17629 13219 17663
rect 15117 17629 15151 17663
rect 20269 17629 20303 17663
rect 20361 17629 20395 17663
rect 11713 17561 11747 17595
rect 11989 17561 12023 17595
rect 14565 17561 14599 17595
rect 15945 17561 15979 17595
rect 21373 17561 21407 17595
rect 5733 17493 5767 17527
rect 7113 17493 7147 17527
rect 8217 17493 8251 17527
rect 11253 17493 11287 17527
rect 19809 17493 19843 17527
rect 6101 17289 6135 17323
rect 6653 17289 6687 17323
rect 6929 17289 6963 17323
rect 9229 17289 9263 17323
rect 10057 17289 10091 17323
rect 12449 17289 12483 17323
rect 14105 17289 14139 17323
rect 14473 17289 14507 17323
rect 14749 17289 14783 17323
rect 20545 17289 20579 17323
rect 1593 17221 1627 17255
rect 8309 17153 8343 17187
rect 9137 17153 9171 17187
rect 8861 17085 8895 17119
rect 1777 17017 1811 17051
rect 8042 17017 8076 17051
rect 10333 17221 10367 17255
rect 12633 17221 12667 17255
rect 15853 17221 15887 17255
rect 9505 17153 9539 17187
rect 9597 17153 9631 17187
rect 10885 17153 10919 17187
rect 11713 17153 11747 17187
rect 9229 17085 9263 17119
rect 10701 17085 10735 17119
rect 12265 17085 12299 17119
rect 12725 17153 12759 17187
rect 15301 17153 15335 17187
rect 16497 17153 16531 17187
rect 17693 17153 17727 17187
rect 18153 17153 18187 17187
rect 19901 17153 19935 17187
rect 20085 17153 20119 17187
rect 12992 17085 13026 17119
rect 17601 17085 17635 17119
rect 18420 17085 18454 17119
rect 21189 17085 21223 17119
rect 15209 17017 15243 17051
rect 16221 17017 16255 17051
rect 2237 16949 2271 16983
rect 5365 16949 5399 16983
rect 5733 16949 5767 16983
rect 9045 16949 9079 16983
rect 9137 16949 9171 16983
rect 9689 16949 9723 16983
rect 10793 16949 10827 16983
rect 12633 16949 12667 16983
rect 15117 16949 15151 16983
rect 16313 16949 16347 16983
rect 17141 16949 17175 16983
rect 17509 16949 17543 16983
rect 19533 16949 19567 16983
rect 20177 16949 20211 16983
rect 21281 16949 21315 16983
rect 5733 16745 5767 16779
rect 6285 16745 6319 16779
rect 8309 16745 8343 16779
rect 8769 16745 8803 16779
rect 9137 16745 9171 16779
rect 9689 16745 9723 16779
rect 9781 16745 9815 16779
rect 10149 16745 10183 16779
rect 13829 16745 13863 16779
rect 14473 16745 14507 16779
rect 14933 16745 14967 16779
rect 15301 16745 15335 16779
rect 15577 16745 15611 16779
rect 16221 16745 16255 16779
rect 16497 16745 16531 16779
rect 16957 16745 16991 16779
rect 17509 16745 17543 16779
rect 18337 16745 18371 16779
rect 19809 16745 19843 16779
rect 5457 16609 5491 16643
rect 6101 16609 6135 16643
rect 7685 16609 7719 16643
rect 8585 16609 8619 16643
rect 9505 16609 9539 16643
rect 9781 16609 9815 16643
rect 11630 16609 11664 16643
rect 11897 16609 11931 16643
rect 12173 16609 12207 16643
rect 12429 16609 12463 16643
rect 14013 16609 14047 16643
rect 17969 16677 18003 16711
rect 18797 16677 18831 16711
rect 21189 16677 21223 16711
rect 14841 16609 14875 16643
rect 16037 16609 16071 16643
rect 16865 16609 16899 16643
rect 18705 16609 18739 16643
rect 20637 16609 20671 16643
rect 21373 16609 21407 16643
rect 7941 16541 7975 16575
rect 14473 16541 14507 16575
rect 14749 16541 14783 16575
rect 17049 16541 17083 16575
rect 18981 16541 19015 16575
rect 6561 16473 6595 16507
rect 13553 16473 13587 16507
rect 10517 16405 10551 16439
rect 20269 16405 20303 16439
rect 20821 16405 20855 16439
rect 6009 16201 6043 16235
rect 8677 16201 8711 16235
rect 13093 16201 13127 16235
rect 15761 16201 15795 16235
rect 17049 16201 17083 16235
rect 11345 16133 11379 16167
rect 17325 16133 17359 16167
rect 19717 16133 19751 16167
rect 9321 16065 9355 16099
rect 10241 16065 10275 16099
rect 10333 16065 10367 16099
rect 12449 16065 12483 16099
rect 14473 16065 14507 16099
rect 14841 16065 14875 16099
rect 16313 16065 16347 16099
rect 17877 16065 17911 16099
rect 20545 16065 20579 16099
rect 20637 16065 20671 16099
rect 5365 15997 5399 16031
rect 8226 15997 8260 16031
rect 8493 15997 8527 16031
rect 8677 15997 8711 16031
rect 9137 15997 9171 16031
rect 10425 15997 10459 16031
rect 11161 15997 11195 16031
rect 16221 15997 16255 16031
rect 17693 15997 17727 16031
rect 18337 15997 18371 16031
rect 18593 15997 18627 16031
rect 21189 15997 21223 16031
rect 5733 15929 5767 15963
rect 9229 15929 9263 15963
rect 12357 15929 12391 15963
rect 14206 15929 14240 15963
rect 20453 15929 20487 15963
rect 21373 15929 21407 15963
rect 4997 15861 5031 15895
rect 6745 15861 6779 15895
rect 7113 15861 7147 15895
rect 8769 15861 8803 15895
rect 10793 15861 10827 15895
rect 11897 15861 11931 15895
rect 12265 15861 12299 15895
rect 15025 15861 15059 15895
rect 15117 15861 15151 15895
rect 15485 15861 15519 15895
rect 16129 15861 16163 15895
rect 17785 15861 17819 15895
rect 20085 15861 20119 15895
rect 5733 15657 5767 15691
rect 6101 15657 6135 15691
rect 6653 15657 6687 15691
rect 7113 15657 7147 15691
rect 11345 15657 11379 15691
rect 11989 15657 12023 15691
rect 12725 15657 12759 15691
rect 13553 15657 13587 15691
rect 14013 15657 14047 15691
rect 15301 15657 15335 15691
rect 16129 15657 16163 15691
rect 16957 15657 16991 15691
rect 17325 15657 17359 15691
rect 18981 15657 19015 15691
rect 19809 15657 19843 15691
rect 6745 15589 6779 15623
rect 9321 15589 9355 15623
rect 18460 15589 18494 15623
rect 21189 15589 21223 15623
rect 8513 15521 8547 15555
rect 10232 15521 10266 15555
rect 11805 15521 11839 15555
rect 12633 15521 12667 15555
rect 13645 15521 13679 15555
rect 14933 15521 14967 15555
rect 16221 15521 16255 15555
rect 16773 15521 16807 15555
rect 20177 15521 20211 15555
rect 6561 15453 6595 15487
rect 8769 15453 8803 15487
rect 9965 15453 9999 15487
rect 12909 15453 12943 15487
rect 13369 15453 13403 15487
rect 14657 15453 14691 15487
rect 14841 15453 14875 15487
rect 16405 15453 16439 15487
rect 18705 15453 18739 15487
rect 20269 15453 20303 15487
rect 20361 15453 20395 15487
rect 7389 15317 7423 15351
rect 12265 15317 12299 15351
rect 15761 15317 15795 15351
rect 21281 15317 21315 15351
rect 7389 15113 7423 15147
rect 11345 15113 11379 15147
rect 18153 15113 18187 15147
rect 18521 15113 18555 15147
rect 7849 15045 7883 15079
rect 9321 15045 9355 15079
rect 10333 15045 10367 15079
rect 14933 15045 14967 15079
rect 16589 15045 16623 15079
rect 8585 14977 8619 15011
rect 8677 14977 8711 15011
rect 9689 14977 9723 15011
rect 9873 14977 9907 15011
rect 10793 14977 10827 15011
rect 12449 14977 12483 15011
rect 12909 14977 12943 15011
rect 18981 14977 19015 15011
rect 7665 14909 7699 14943
rect 9137 14909 9171 14943
rect 10517 14909 10551 14943
rect 10885 14909 10919 14943
rect 12265 14909 12299 14943
rect 13553 14909 13587 14943
rect 13820 14909 13854 14943
rect 15209 14909 15243 14943
rect 15465 14909 15499 14943
rect 17877 14909 17911 14943
rect 18153 14909 18187 14943
rect 18337 14909 18371 14943
rect 20370 14909 20404 14943
rect 20637 14909 20671 14943
rect 21189 14909 21223 14943
rect 6653 14841 6687 14875
rect 9965 14841 9999 14875
rect 17141 14841 17175 14875
rect 21373 14841 21407 14875
rect 7021 14773 7055 14807
rect 8125 14773 8159 14807
rect 8493 14773 8527 14807
rect 10517 14773 10551 14807
rect 10977 14773 11011 14807
rect 11897 14773 11931 14807
rect 12357 14773 12391 14807
rect 18061 14773 18095 14807
rect 19257 14773 19291 14807
rect 5641 14569 5675 14603
rect 6009 14569 6043 14603
rect 6469 14569 6503 14603
rect 7481 14569 7515 14603
rect 7941 14569 7975 14603
rect 8401 14569 8435 14603
rect 12909 14569 12943 14603
rect 13369 14569 13403 14603
rect 14197 14569 14231 14603
rect 14381 14569 14415 14603
rect 14933 14569 14967 14603
rect 18337 14569 18371 14603
rect 11529 14501 11563 14535
rect 15577 14501 15611 14535
rect 21189 14501 21223 14535
rect 7665 14433 7699 14467
rect 8309 14433 8343 14467
rect 9505 14433 9539 14467
rect 9772 14433 9806 14467
rect 12173 14433 12207 14467
rect 13001 14433 13035 14467
rect 13829 14433 13863 14467
rect 14289 14433 14323 14467
rect 14749 14433 14783 14467
rect 17610 14433 17644 14467
rect 18153 14433 18187 14467
rect 18613 14433 18647 14467
rect 19073 14433 19107 14467
rect 20453 14433 20487 14467
rect 8493 14365 8527 14399
rect 11621 14365 11655 14399
rect 11713 14365 11747 14399
rect 12817 14365 12851 14399
rect 15669 14365 15703 14399
rect 15853 14365 15887 14399
rect 17877 14365 17911 14399
rect 20545 14365 20579 14399
rect 20637 14365 20671 14399
rect 7205 14297 7239 14331
rect 12357 14297 12391 14331
rect 14013 14297 14047 14331
rect 15209 14297 15243 14331
rect 16497 14297 16531 14331
rect 19257 14297 19291 14331
rect 21373 14297 21407 14331
rect 6837 14229 6871 14263
rect 9229 14229 9263 14263
rect 10885 14229 10919 14263
rect 11161 14229 11195 14263
rect 18797 14229 18831 14263
rect 19625 14229 19659 14263
rect 20085 14229 20119 14263
rect 7113 14025 7147 14059
rect 7573 14025 7607 14059
rect 8401 14025 8435 14059
rect 9321 14025 9355 14059
rect 12173 14025 12207 14059
rect 13829 14025 13863 14059
rect 14105 14025 14139 14059
rect 19901 14025 19935 14059
rect 7849 13957 7883 13991
rect 9597 13957 9631 13991
rect 11345 13957 11379 13991
rect 17141 13957 17175 13991
rect 6837 13889 6871 13923
rect 14749 13889 14783 13923
rect 16405 13889 16439 13923
rect 18521 13889 18555 13923
rect 19533 13889 19567 13923
rect 20361 13889 20395 13923
rect 20453 13889 20487 13923
rect 8217 13821 8251 13855
rect 8861 13821 8895 13855
rect 9137 13821 9171 13855
rect 10977 13821 11011 13855
rect 11989 13821 12023 13855
rect 12449 13821 12483 13855
rect 16313 13821 16347 13855
rect 21189 13821 21223 13855
rect 21373 13821 21407 13855
rect 10710 13753 10744 13787
rect 12716 13753 12750 13787
rect 14565 13753 14599 13787
rect 16221 13753 16255 13787
rect 18254 13753 18288 13787
rect 20269 13753 20303 13787
rect 8677 13685 8711 13719
rect 14473 13685 14507 13719
rect 15117 13685 15151 13719
rect 15853 13685 15887 13719
rect 18889 13685 18923 13719
rect 19257 13685 19291 13719
rect 19349 13685 19383 13719
rect 6745 13481 6779 13515
rect 8769 13481 8803 13515
rect 14565 13481 14599 13515
rect 15393 13481 15427 13515
rect 15761 13481 15795 13515
rect 16405 13481 16439 13515
rect 18429 13481 18463 13515
rect 20085 13481 20119 13515
rect 7481 13413 7515 13447
rect 9137 13413 9171 13447
rect 11354 13413 11388 13447
rect 12265 13413 12299 13447
rect 21189 13413 21223 13447
rect 8309 13345 8343 13379
rect 8585 13345 8619 13379
rect 9505 13345 9539 13379
rect 11621 13345 11655 13379
rect 13645 13345 13679 13379
rect 14933 13345 14967 13379
rect 15853 13345 15887 13379
rect 17518 13345 17552 13379
rect 19257 13345 19291 13379
rect 20453 13345 20487 13379
rect 20545 13345 20579 13379
rect 7849 13277 7883 13311
rect 12357 13277 12391 13311
rect 12449 13277 12483 13311
rect 13737 13277 13771 13311
rect 13921 13277 13955 13311
rect 16037 13277 16071 13311
rect 17785 13277 17819 13311
rect 18521 13277 18555 13311
rect 18613 13277 18647 13311
rect 19809 13277 19843 13311
rect 20729 13277 20763 13311
rect 9689 13209 9723 13243
rect 21373 13209 21407 13243
rect 7113 13141 7147 13175
rect 8125 13141 8159 13175
rect 10241 13141 10275 13175
rect 11897 13141 11931 13175
rect 12909 13141 12943 13175
rect 13277 13141 13311 13175
rect 15117 13141 15151 13175
rect 18061 13141 18095 13175
rect 7021 12937 7055 12971
rect 7849 12937 7883 12971
rect 11345 12937 11379 12971
rect 11437 12937 11471 12971
rect 7297 12869 7331 12903
rect 9873 12869 9907 12903
rect 10149 12869 10183 12903
rect 10793 12801 10827 12835
rect 10885 12801 10919 12835
rect 7665 12733 7699 12767
rect 9249 12733 9283 12767
rect 9505 12733 9539 12767
rect 10333 12733 10367 12767
rect 14289 12937 14323 12971
rect 15209 12937 15243 12971
rect 20453 12937 20487 12971
rect 13093 12801 13127 12835
rect 14105 12801 14139 12835
rect 12817 12733 12851 12767
rect 13829 12665 13863 12699
rect 18521 12869 18555 12903
rect 14565 12801 14599 12835
rect 16313 12801 16347 12835
rect 17509 12801 17543 12835
rect 21005 12801 21039 12835
rect 14841 12733 14875 12767
rect 16957 12733 16991 12767
rect 17693 12733 17727 12767
rect 19634 12733 19668 12767
rect 19901 12733 19935 12767
rect 16221 12665 16255 12699
rect 8125 12597 8159 12631
rect 10977 12597 11011 12631
rect 11437 12597 11471 12631
rect 11897 12597 11931 12631
rect 12449 12597 12483 12631
rect 12909 12597 12943 12631
rect 13461 12597 13495 12631
rect 13921 12597 13955 12631
rect 14289 12597 14323 12631
rect 14749 12597 14783 12631
rect 15761 12597 15795 12631
rect 16129 12597 16163 12631
rect 17785 12597 17819 12631
rect 18153 12597 18187 12631
rect 20821 12597 20855 12631
rect 20913 12597 20947 12631
rect 6929 12393 6963 12427
rect 7849 12393 7883 12427
rect 11713 12393 11747 12427
rect 14565 12393 14599 12427
rect 16497 12393 16531 12427
rect 16957 12393 16991 12427
rect 17509 12393 17543 12427
rect 17877 12393 17911 12427
rect 18981 12393 19015 12427
rect 19901 12393 19935 12427
rect 11345 12325 11379 12359
rect 7665 12257 7699 12291
rect 8125 12257 8159 12291
rect 8585 12257 8619 12291
rect 9597 12257 9631 12291
rect 9689 12257 9723 12291
rect 10517 12257 10551 12291
rect 12541 12257 12575 12291
rect 12808 12257 12842 12291
rect 15678 12257 15712 12291
rect 15945 12257 15979 12291
rect 16865 12257 16899 12291
rect 18889 12257 18923 12291
rect 21014 12257 21048 12291
rect 21281 12257 21315 12291
rect 7389 12189 7423 12223
rect 9413 12189 9447 12223
rect 11069 12189 11103 12223
rect 11253 12189 11287 12223
rect 12265 12189 12299 12223
rect 17141 12189 17175 12223
rect 17969 12189 18003 12223
rect 18061 12189 18095 12223
rect 19073 12189 19107 12223
rect 8769 12121 8803 12155
rect 8309 12053 8343 12087
rect 10057 12053 10091 12087
rect 10701 12053 10735 12087
rect 13921 12053 13955 12087
rect 18521 12053 18555 12087
rect 7757 11849 7791 11883
rect 10057 11849 10091 11883
rect 13277 11849 13311 11883
rect 13553 11849 13587 11883
rect 16129 11849 16163 11883
rect 17325 11849 17359 11883
rect 19993 11849 20027 11883
rect 9781 11781 9815 11815
rect 8401 11713 8435 11747
rect 10517 11713 10551 11747
rect 10609 11713 10643 11747
rect 11897 11713 11931 11747
rect 14105 11713 14139 11747
rect 8657 11645 8691 11679
rect 14749 11645 14783 11679
rect 15005 11645 15039 11679
rect 17141 11645 17175 11679
rect 18990 11645 19024 11679
rect 19257 11645 19291 11679
rect 19717 11645 19751 11679
rect 21373 11645 21407 11679
rect 10425 11577 10459 11611
rect 11069 11577 11103 11611
rect 12164 11577 12198 11611
rect 16405 11577 16439 11611
rect 21128 11577 21162 11611
rect 8125 11509 8159 11543
rect 13921 11509 13955 11543
rect 14013 11509 14047 11543
rect 17877 11509 17911 11543
rect 19533 11509 19567 11543
rect 7113 11305 7147 11339
rect 11713 11305 11747 11339
rect 12449 11305 12483 11339
rect 13737 11305 13771 11339
rect 18521 11305 18555 11339
rect 21189 11305 21223 11339
rect 8493 11237 8527 11271
rect 9588 11237 9622 11271
rect 13369 11237 13403 11271
rect 16834 11237 16868 11271
rect 20054 11237 20088 11271
rect 8125 11169 8159 11203
rect 7849 11101 7883 11135
rect 8585 11169 8619 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 12357 11169 12391 11203
rect 14565 11169 14599 11203
rect 16313 11169 16347 11203
rect 18889 11169 18923 11203
rect 18981 11169 19015 11203
rect 9321 11101 9355 11135
rect 11069 11101 11103 11135
rect 12633 11101 12667 11135
rect 13093 11101 13127 11135
rect 13277 11101 13311 11135
rect 16497 11101 16531 11135
rect 16589 11101 16623 11135
rect 19073 11101 19107 11135
rect 19809 11101 19843 11135
rect 7481 11033 7515 11067
rect 8309 11033 8343 11067
rect 8493 11033 8527 11067
rect 8769 11033 8803 11067
rect 11989 11033 12023 11067
rect 10701 10965 10735 10999
rect 16497 10965 16531 10999
rect 17969 10965 18003 10999
rect 7389 10761 7423 10795
rect 8677 10761 8711 10795
rect 13185 10761 13219 10795
rect 14749 10761 14783 10795
rect 18889 10761 18923 10795
rect 20545 10761 20579 10795
rect 16589 10693 16623 10727
rect 12081 10625 12115 10659
rect 12633 10625 12667 10659
rect 13553 10625 13587 10659
rect 15301 10625 15335 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 17233 10625 17267 10659
rect 17417 10625 17451 10659
rect 18613 10625 18647 10659
rect 21189 10625 21223 10659
rect 8493 10557 8527 10591
rect 8953 10557 8987 10591
rect 9413 10557 9447 10591
rect 9873 10557 9907 10591
rect 10140 10557 10174 10591
rect 13737 10557 13771 10591
rect 15209 10557 15243 10591
rect 16221 10557 16255 10591
rect 20269 10557 20303 10591
rect 8217 10489 8251 10523
rect 20024 10489 20058 10523
rect 7757 10421 7791 10455
rect 9137 10421 9171 10455
rect 9597 10421 9631 10455
rect 11253 10421 11287 10455
rect 12725 10421 12759 10455
rect 12817 10421 12851 10455
rect 13829 10421 13863 10455
rect 14197 10421 14231 10455
rect 15117 10421 15151 10455
rect 17509 10421 17543 10455
rect 17877 10421 17911 10455
rect 20913 10421 20947 10455
rect 21005 10421 21039 10455
rect 9229 10217 9263 10251
rect 10057 10217 10091 10251
rect 10149 10217 10183 10251
rect 10517 10217 10551 10251
rect 10701 10217 10735 10251
rect 12173 10217 12207 10251
rect 13829 10217 13863 10251
rect 14933 10217 14967 10251
rect 15945 10217 15979 10251
rect 16129 10217 16163 10251
rect 18245 10217 18279 10251
rect 18889 10217 18923 10251
rect 19809 10217 19843 10251
rect 21005 10217 21039 10251
rect 8769 10081 8803 10115
rect 9321 10081 9355 10115
rect 12265 10149 12299 10183
rect 12694 10149 12728 10183
rect 11060 10081 11094 10115
rect 15761 10081 15795 10115
rect 9873 10013 9907 10047
rect 10701 10013 10735 10047
rect 10793 10013 10827 10047
rect 12265 10013 12299 10047
rect 12449 10013 12483 10047
rect 15025 10013 15059 10047
rect 15117 10013 15151 10047
rect 17693 10149 17727 10183
rect 20177 10149 20211 10183
rect 16488 10081 16522 10115
rect 16221 10013 16255 10047
rect 14565 9945 14599 9979
rect 16129 9945 16163 9979
rect 19073 10081 19107 10115
rect 20821 10081 20855 10115
rect 18337 10013 18371 10047
rect 18521 10013 18555 10047
rect 20269 10013 20303 10047
rect 20361 10013 20395 10047
rect 8309 9877 8343 9911
rect 9229 9877 9263 9911
rect 9505 9877 9539 9911
rect 17601 9877 17635 9911
rect 17693 9877 17727 9911
rect 17877 9877 17911 9911
rect 21281 9877 21315 9911
rect 8033 9673 8067 9707
rect 18521 9673 18555 9707
rect 20177 9673 20211 9707
rect 9689 9605 9723 9639
rect 10149 9605 10183 9639
rect 11897 9605 11931 9639
rect 13737 9605 13771 9639
rect 10517 9537 10551 9571
rect 12541 9537 12575 9571
rect 13093 9537 13127 9571
rect 13921 9537 13955 9571
rect 14565 9537 14599 9571
rect 15577 9537 15611 9571
rect 16589 9537 16623 9571
rect 17141 9537 17175 9571
rect 21005 9537 21039 9571
rect 9229 9469 9263 9503
rect 9505 9469 9539 9503
rect 9965 9469 9999 9503
rect 11805 9469 11839 9503
rect 12265 9469 12299 9503
rect 18797 9469 18831 9503
rect 19053 9469 19087 9503
rect 20913 9469 20947 9503
rect 13921 9401 13955 9435
rect 14381 9401 14415 9435
rect 15485 9401 15519 9435
rect 17408 9401 17442 9435
rect 8401 9333 8435 9367
rect 8861 9333 8895 9367
rect 10701 9333 10735 9367
rect 10793 9333 10827 9367
rect 11161 9333 11195 9367
rect 11805 9333 11839 9367
rect 12357 9333 12391 9367
rect 13277 9333 13311 9367
rect 13369 9333 13403 9367
rect 14013 9333 14047 9367
rect 14473 9333 14507 9367
rect 15025 9333 15059 9367
rect 15393 9333 15427 9367
rect 16129 9333 16163 9367
rect 20453 9333 20487 9367
rect 20821 9333 20855 9367
rect 11069 9129 11103 9163
rect 12081 9129 12115 9163
rect 13645 9129 13679 9163
rect 15945 9129 15979 9163
rect 16129 9129 16163 9163
rect 16221 9129 16255 9163
rect 16681 9129 16715 9163
rect 17509 9129 17543 9163
rect 17969 9129 18003 9163
rect 18245 9129 18279 9163
rect 21005 9129 21039 9163
rect 8309 9061 8343 9095
rect 12357 9061 12391 9095
rect 13553 9061 13587 9095
rect 8769 8993 8803 9027
rect 9945 8993 9979 9027
rect 11713 8993 11747 9027
rect 14565 8993 14599 9027
rect 14832 8993 14866 9027
rect 9689 8925 9723 8959
rect 11437 8925 11471 8959
rect 11621 8925 11655 8959
rect 13737 8925 13771 8959
rect 17601 9061 17635 9095
rect 18613 9061 18647 9095
rect 16589 8993 16623 9027
rect 20361 8993 20395 9027
rect 16773 8925 16807 8959
rect 17325 8925 17359 8959
rect 18705 8925 18739 8959
rect 18797 8925 18831 8959
rect 20453 8925 20487 8959
rect 20637 8925 20671 8959
rect 8585 8857 8619 8891
rect 13185 8857 13219 8891
rect 16129 8857 16163 8891
rect 7849 8789 7883 8823
rect 9137 8789 9171 8823
rect 12817 8789 12851 8823
rect 19625 8789 19659 8823
rect 19993 8789 20027 8823
rect 7205 8585 7239 8619
rect 8401 8585 8435 8619
rect 9597 8585 9631 8619
rect 13553 8585 13587 8619
rect 13829 8585 13863 8619
rect 14289 8585 14323 8619
rect 18337 8585 18371 8619
rect 19625 8585 19659 8619
rect 19809 8585 19843 8619
rect 8861 8517 8895 8551
rect 9321 8517 9355 8551
rect 18797 8517 18831 8551
rect 11253 8449 11287 8483
rect 13645 8449 13679 8483
rect 14841 8449 14875 8483
rect 15485 8449 15519 8483
rect 16405 8449 16439 8483
rect 17785 8449 17819 8483
rect 19257 8449 19291 8483
rect 19441 8449 19475 8483
rect 19625 8449 19659 8483
rect 8217 8381 8251 8415
rect 8677 8381 8711 8415
rect 9137 8381 9171 8415
rect 10977 8381 11011 8415
rect 12173 8381 12207 8415
rect 12440 8381 12474 8415
rect 7573 8313 7607 8347
rect 10732 8313 10766 8347
rect 14013 8381 14047 8415
rect 17141 8381 17175 8415
rect 17969 8381 18003 8415
rect 19165 8381 19199 8415
rect 21189 8381 21223 8415
rect 14657 8313 14691 8347
rect 14749 8313 14783 8347
rect 16221 8313 16255 8347
rect 16313 8313 16347 8347
rect 20944 8313 20978 8347
rect 7849 8245 7883 8279
rect 11713 8245 11747 8279
rect 13645 8245 13679 8279
rect 15853 8245 15887 8279
rect 17325 8245 17359 8279
rect 17877 8245 17911 8279
rect 7021 8041 7055 8075
rect 9321 8041 9355 8075
rect 10149 8041 10183 8075
rect 10701 8041 10735 8075
rect 11069 8041 11103 8075
rect 12081 8041 12115 8075
rect 14933 8041 14967 8075
rect 17693 8041 17727 8075
rect 18797 8041 18831 8075
rect 21189 8041 21223 8075
rect 7849 7973 7883 8007
rect 7481 7905 7515 7939
rect 8125 7905 8159 7939
rect 8585 7905 8619 7939
rect 9689 7905 9723 7939
rect 9781 7837 9815 7871
rect 9965 7837 9999 7871
rect 12808 7973 12842 8007
rect 14473 7973 14507 8007
rect 11713 7905 11747 7939
rect 16046 7905 16080 7939
rect 17785 7905 17819 7939
rect 18705 7905 18739 7939
rect 19809 7905 19843 7939
rect 20076 7905 20110 7939
rect 10517 7837 10551 7871
rect 10609 7837 10643 7871
rect 11437 7837 11471 7871
rect 11621 7837 11655 7871
rect 12541 7837 12575 7871
rect 16313 7837 16347 7871
rect 16865 7837 16899 7871
rect 17509 7837 17543 7871
rect 18521 7837 18555 7871
rect 10149 7769 10183 7803
rect 8309 7701 8343 7735
rect 8769 7701 8803 7735
rect 13921 7701 13955 7735
rect 18153 7701 18187 7735
rect 19165 7701 19199 7735
rect 7389 7497 7423 7531
rect 9505 7497 9539 7531
rect 11161 7497 11195 7531
rect 12357 7497 12391 7531
rect 12449 7497 12483 7531
rect 15117 7497 15151 7531
rect 17141 7497 17175 7531
rect 7021 7429 7055 7463
rect 13185 7361 13219 7395
rect 14197 7361 14231 7395
rect 16497 7361 16531 7395
rect 19257 7361 19291 7395
rect 19349 7361 19383 7395
rect 20453 7361 20487 7395
rect 7849 7293 7883 7327
rect 8125 7293 8159 7327
rect 9781 7293 9815 7327
rect 10048 7293 10082 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 12449 7293 12483 7327
rect 14013 7293 14047 7327
rect 14841 7293 14875 7327
rect 16241 7293 16275 7327
rect 18521 7293 18555 7327
rect 19165 7293 19199 7327
rect 8392 7225 8426 7259
rect 13001 7225 13035 7259
rect 14105 7225 14139 7259
rect 18254 7225 18288 7259
rect 7665 7157 7699 7191
rect 11897 7157 11931 7191
rect 11989 7157 12023 7191
rect 12633 7157 12667 7191
rect 13093 7157 13127 7191
rect 13645 7157 13679 7191
rect 14657 7157 14691 7191
rect 18797 7157 18831 7191
rect 19901 7157 19935 7191
rect 20269 7157 20303 7191
rect 20361 7157 20395 7191
rect 20913 7157 20947 7191
rect 10057 6953 10091 6987
rect 10885 6953 10919 6987
rect 11529 6953 11563 6987
rect 13645 6953 13679 6987
rect 16405 6953 16439 6987
rect 18889 6953 18923 6987
rect 11437 6885 11471 6919
rect 14933 6885 14967 6919
rect 17417 6885 17451 6919
rect 20076 6885 20110 6919
rect 6561 6817 6595 6851
rect 7021 6817 7055 6851
rect 7665 6817 7699 6851
rect 8125 6817 8159 6851
rect 8769 6817 8803 6851
rect 9689 6817 9723 6851
rect 10977 6817 11011 6851
rect 7389 6749 7423 6783
rect 9413 6749 9447 6783
rect 9597 6749 9631 6783
rect 11069 6749 11103 6783
rect 12642 6817 12676 6851
rect 12909 6817 12943 6851
rect 15577 6817 15611 6851
rect 17509 6817 17543 6851
rect 18245 6817 18279 6851
rect 13737 6749 13771 6783
rect 13921 6749 13955 6783
rect 15025 6749 15059 6783
rect 15117 6749 15151 6783
rect 16497 6749 16531 6783
rect 16589 6749 16623 6783
rect 17601 6749 17635 6783
rect 18613 6749 18647 6783
rect 18797 6749 18831 6783
rect 19809 6749 19843 6783
rect 11437 6681 11471 6715
rect 16037 6681 16071 6715
rect 17049 6681 17083 6715
rect 6285 6613 6319 6647
rect 7849 6613 7883 6647
rect 8309 6613 8343 6647
rect 10517 6613 10551 6647
rect 13277 6613 13311 6647
rect 14565 6613 14599 6647
rect 15761 6613 15795 6647
rect 18061 6613 18095 6647
rect 19257 6613 19291 6647
rect 21189 6613 21223 6647
rect 9137 6409 9171 6443
rect 9321 6409 9355 6443
rect 20637 6409 20671 6443
rect 7297 6341 7331 6375
rect 7665 6273 7699 6307
rect 6929 6205 6963 6239
rect 7932 6137 7966 6171
rect 12817 6341 12851 6375
rect 20361 6341 20395 6375
rect 9873 6273 9907 6307
rect 10885 6273 10919 6307
rect 11989 6273 12023 6307
rect 12173 6273 12207 6307
rect 12357 6273 12391 6307
rect 15301 6273 15335 6307
rect 21189 6273 21223 6307
rect 9781 6137 9815 6171
rect 10701 6137 10735 6171
rect 11805 6137 11839 6171
rect 14473 6205 14507 6239
rect 15577 6205 15611 6239
rect 16221 6205 16255 6239
rect 17325 6205 17359 6239
rect 18981 6205 19015 6239
rect 19248 6205 19282 6239
rect 21005 6205 21039 6239
rect 12449 6137 12483 6171
rect 14206 6137 14240 6171
rect 17570 6137 17604 6171
rect 6101 6069 6135 6103
rect 6653 6069 6687 6103
rect 9045 6069 9079 6103
rect 9137 6069 9171 6103
rect 9689 6069 9723 6103
rect 10333 6069 10367 6103
rect 10793 6069 10827 6103
rect 11989 6069 12023 6103
rect 13093 6069 13127 6103
rect 14749 6069 14783 6103
rect 15485 6069 15519 6103
rect 15945 6069 15979 6103
rect 16405 6069 16439 6103
rect 17049 6069 17083 6103
rect 18705 6069 18739 6103
rect 21097 6069 21131 6103
rect 1777 5865 1811 5899
rect 5825 5865 5859 5899
rect 6285 5865 6319 5899
rect 7941 5865 7975 5899
rect 8769 5865 8803 5899
rect 9597 5865 9631 5899
rect 9965 5865 9999 5899
rect 12909 5865 12943 5899
rect 13185 5865 13219 5899
rect 13553 5865 13587 5899
rect 15945 5865 15979 5899
rect 16681 5865 16715 5899
rect 17325 5865 17359 5899
rect 20177 5865 20211 5899
rect 20545 5865 20579 5899
rect 6806 5797 6840 5831
rect 10057 5797 10091 5831
rect 11814 5797 11848 5831
rect 16589 5797 16623 5831
rect 18460 5797 18494 5831
rect 21189 5797 21223 5831
rect 1593 5729 1627 5763
rect 2053 5729 2087 5763
rect 6561 5729 6595 5763
rect 8309 5729 8343 5763
rect 8585 5729 8619 5763
rect 12081 5729 12115 5763
rect 12725 5729 12759 5763
rect 13645 5729 13679 5763
rect 14565 5729 14599 5763
rect 15577 5729 15611 5763
rect 19165 5729 19199 5763
rect 10149 5661 10183 5695
rect 13737 5661 13771 5695
rect 15301 5661 15335 5695
rect 15485 5661 15519 5695
rect 16773 5661 16807 5695
rect 18705 5661 18739 5695
rect 19993 5661 20027 5695
rect 20085 5661 20119 5695
rect 12449 5593 12483 5627
rect 16221 5593 16255 5627
rect 21005 5593 21039 5627
rect 9321 5525 9355 5559
rect 10701 5525 10735 5559
rect 14749 5525 14783 5559
rect 18981 5525 19015 5559
rect 6653 5321 6687 5355
rect 10333 5321 10367 5355
rect 10425 5321 10459 5355
rect 6009 5253 6043 5287
rect 7389 5253 7423 5287
rect 7757 5253 7791 5287
rect 9873 5253 9907 5287
rect 8493 5185 8527 5219
rect 8769 5117 8803 5151
rect 9229 5117 9263 5151
rect 9689 5117 9723 5151
rect 9965 5117 9999 5151
rect 10149 5117 10183 5151
rect 7021 5049 7055 5083
rect 8125 5049 8159 5083
rect 8953 4981 8987 5015
rect 9413 4981 9447 5015
rect 9965 4981 9999 5015
rect 10517 5253 10551 5287
rect 16129 5253 16163 5287
rect 19625 5253 19659 5287
rect 10793 5185 10827 5219
rect 12541 5185 12575 5219
rect 17693 5185 17727 5219
rect 20085 5185 20119 5219
rect 20269 5185 20303 5219
rect 21189 5185 21223 5219
rect 10517 5117 10551 5151
rect 10885 5117 10919 5151
rect 12357 5117 12391 5151
rect 13093 5117 13127 5151
rect 14749 5117 14783 5151
rect 15016 5117 15050 5151
rect 19993 5117 20027 5151
rect 13360 5049 13394 5083
rect 16589 5049 16623 5083
rect 17509 5049 17543 5083
rect 17601 5049 17635 5083
rect 18245 5049 18279 5083
rect 19349 5049 19383 5083
rect 21005 5049 21039 5083
rect 10425 4981 10459 5015
rect 10977 4981 11011 5015
rect 11345 4981 11379 5015
rect 11897 4981 11931 5015
rect 12265 4981 12299 5015
rect 14473 4981 14507 5015
rect 17141 4981 17175 5015
rect 18705 4981 18739 5015
rect 20637 4981 20671 5015
rect 21097 4981 21131 5015
rect 6193 4777 6227 4811
rect 6561 4777 6595 4811
rect 7297 4777 7331 4811
rect 17325 4777 17359 4811
rect 19717 4777 19751 4811
rect 21189 4777 21223 4811
rect 6837 4709 6871 4743
rect 11253 4709 11287 4743
rect 11682 4709 11716 4743
rect 15025 4709 15059 4743
rect 16212 4709 16246 4743
rect 17785 4709 17819 4743
rect 18705 4709 18739 4743
rect 8769 4641 8803 4675
rect 9321 4641 9355 4675
rect 10048 4641 10082 4675
rect 9781 4573 9815 4607
rect 13369 4641 13403 4675
rect 13921 4641 13955 4675
rect 15577 4641 15611 4675
rect 18521 4641 18555 4675
rect 19073 4641 19107 4675
rect 19717 4641 19751 4675
rect 19809 4641 19843 4675
rect 20076 4641 20110 4675
rect 11437 4573 11471 4607
rect 15945 4573 15979 4607
rect 11161 4505 11195 4539
rect 11253 4505 11287 4539
rect 13185 4505 13219 4539
rect 13737 4505 13771 4539
rect 14841 4505 14875 4539
rect 15393 4505 15427 4539
rect 17601 4505 17635 4539
rect 7665 4437 7699 4471
rect 8033 4437 8067 4471
rect 8401 4437 8435 4471
rect 9505 4437 9539 4471
rect 12817 4437 12851 4471
rect 14565 4437 14599 4471
rect 19165 4437 19199 4471
rect 5733 4233 5767 4267
rect 9505 4233 9539 4267
rect 20729 4233 20763 4267
rect 6561 4097 6595 4131
rect 7665 4097 7699 4131
rect 12909 4165 12943 4199
rect 19717 4165 19751 4199
rect 10793 4097 10827 4131
rect 12357 4097 12391 4131
rect 12541 4097 12575 4131
rect 13461 4097 13495 4131
rect 14565 4097 14599 4131
rect 16221 4097 16255 4131
rect 16405 4097 16439 4131
rect 17693 4097 17727 4131
rect 18337 4097 18371 4131
rect 20085 4097 20119 4131
rect 6929 4029 6963 4063
rect 8309 4029 8343 4063
rect 8769 4029 8803 4063
rect 9229 4029 9263 4063
rect 9505 4029 9539 4063
rect 9713 4029 9747 4063
rect 10149 4029 10183 4063
rect 10977 4029 11011 4063
rect 11805 4029 11839 4063
rect 13277 4029 13311 4063
rect 14087 4029 14121 4063
rect 15025 4029 15059 4063
rect 16129 4029 16163 4063
rect 21281 4029 21315 4063
rect 7205 3961 7239 3995
rect 10885 3961 10919 3995
rect 13369 3961 13403 3995
rect 14657 3961 14691 3995
rect 15209 3961 15243 3995
rect 17325 3961 17359 3995
rect 17877 3961 17911 3995
rect 18604 3961 18638 3995
rect 21097 3961 21131 3995
rect 6101 3893 6135 3927
rect 8033 3893 8067 3927
rect 8493 3893 8527 3927
rect 8953 3893 8987 3927
rect 9413 3893 9447 3927
rect 9873 3893 9907 3927
rect 10333 3893 10367 3927
rect 11345 3893 11379 3927
rect 11805 3893 11839 3927
rect 11897 3893 11931 3927
rect 12265 3893 12299 3927
rect 14565 3893 14599 3927
rect 15761 3893 15795 3927
rect 17233 3893 17267 3927
rect 20269 3893 20303 3927
rect 20361 3893 20395 3927
rect 5365 3689 5399 3723
rect 7941 3689 7975 3723
rect 6653 3621 6687 3655
rect 4997 3553 5031 3587
rect 5641 3485 5675 3519
rect 1777 3417 1811 3451
rect 9689 3689 9723 3723
rect 10425 3689 10459 3723
rect 11529 3689 11563 3723
rect 12173 3689 12207 3723
rect 14013 3689 14047 3723
rect 16681 3689 16715 3723
rect 18889 3689 18923 3723
rect 14810 3621 14844 3655
rect 19993 3621 20027 3655
rect 20545 3621 20579 3655
rect 21281 3621 21315 3655
rect 8125 3553 8159 3587
rect 8585 3553 8619 3587
rect 8861 3553 8895 3587
rect 9321 3553 9355 3587
rect 9689 3553 9723 3587
rect 9781 3553 9815 3587
rect 10241 3553 10275 3587
rect 10701 3553 10735 3587
rect 12817 3553 12851 3587
rect 13645 3553 13679 3587
rect 14565 3553 14599 3587
rect 17776 3553 17810 3587
rect 20729 3553 20763 3587
rect 8309 3417 8343 3451
rect 11253 3485 11287 3519
rect 11437 3485 11471 3519
rect 13369 3485 13403 3519
rect 13553 3485 13587 3519
rect 16773 3485 16807 3519
rect 16957 3485 16991 3519
rect 17509 3485 17543 3519
rect 9505 3417 9539 3451
rect 9965 3417 9999 3451
rect 12633 3417 12667 3451
rect 19809 3417 19843 3451
rect 1409 3349 1443 3383
rect 6193 3349 6227 3383
rect 7021 3349 7055 3383
rect 7297 3349 7331 3383
rect 7757 3349 7791 3383
rect 7941 3349 7975 3383
rect 8769 3349 8803 3383
rect 8861 3349 8895 3383
rect 10885 3349 10919 3383
rect 11897 3349 11931 3383
rect 15945 3349 15979 3383
rect 16313 3349 16347 3383
rect 19165 3349 19199 3383
rect 21189 3349 21223 3383
rect 4905 3145 4939 3179
rect 10609 3145 10643 3179
rect 10885 3145 10919 3179
rect 13277 3145 13311 3179
rect 14933 3145 14967 3179
rect 18521 3145 18555 3179
rect 1593 3077 1627 3111
rect 4445 3077 4479 3111
rect 6101 3077 6135 3111
rect 7849 3009 7883 3043
rect 1409 2941 1443 2975
rect 1869 2941 1903 2975
rect 2789 2941 2823 2975
rect 4721 2941 4755 2975
rect 5549 2941 5583 2975
rect 7021 2941 7055 2975
rect 7481 2941 7515 2975
rect 2329 2873 2363 2907
rect 3065 2873 3099 2907
rect 16589 3077 16623 3111
rect 16773 3077 16807 3111
rect 11897 3009 11931 3043
rect 15025 3009 15059 3043
rect 7941 2941 7975 2975
rect 8401 2941 8435 2975
rect 8861 2941 8895 2975
rect 9321 2941 9355 2975
rect 9781 2941 9815 2975
rect 10241 2941 10275 2975
rect 10609 2941 10643 2975
rect 10701 2941 10735 2975
rect 11161 2941 11195 2975
rect 13553 2941 13587 2975
rect 13809 2941 13843 2975
rect 12142 2873 12176 2907
rect 15209 2941 15243 2975
rect 15476 2941 15510 2975
rect 19349 3009 19383 3043
rect 19625 3009 19659 3043
rect 20545 3009 20579 3043
rect 21097 3009 21131 3043
rect 17141 2941 17175 2975
rect 19165 2941 19199 2975
rect 19257 2941 19291 2975
rect 20729 2941 20763 2975
rect 21281 2941 21315 2975
rect 16773 2873 16807 2907
rect 17386 2873 17420 2907
rect 19625 2873 19659 2907
rect 19809 2873 19843 2907
rect 19993 2873 20027 2907
rect 2053 2805 2087 2839
rect 3433 2805 3467 2839
rect 3985 2805 4019 2839
rect 5181 2805 5215 2839
rect 6561 2805 6595 2839
rect 7205 2805 7239 2839
rect 7665 2805 7699 2839
rect 7849 2805 7883 2839
rect 8125 2805 8159 2839
rect 8585 2805 8619 2839
rect 9045 2805 9079 2839
rect 9505 2805 9539 2839
rect 9965 2805 9999 2839
rect 10425 2805 10459 2839
rect 11345 2805 11379 2839
rect 15025 2805 15059 2839
rect 18797 2805 18831 2839
rect 1593 2601 1627 2635
rect 4261 2601 4295 2635
rect 4813 2601 4847 2635
rect 6929 2601 6963 2635
rect 10701 2601 10735 2635
rect 11161 2601 11195 2635
rect 11897 2601 11931 2635
rect 14749 2601 14783 2635
rect 16037 2601 16071 2635
rect 16497 2601 16531 2635
rect 17325 2601 17359 2635
rect 20085 2601 20119 2635
rect 2237 2533 2271 2567
rect 4169 2533 4203 2567
rect 5549 2533 5583 2567
rect 7573 2533 7607 2567
rect 8401 2533 8435 2567
rect 10241 2533 10275 2567
rect 1409 2465 1443 2499
rect 2053 2465 2087 2499
rect 2513 2465 2547 2499
rect 3157 2465 3191 2499
rect 4721 2465 4755 2499
rect 5365 2465 5399 2499
rect 6009 2465 6043 2499
rect 6837 2465 6871 2499
rect 7757 2465 7791 2499
rect 8217 2465 8251 2499
rect 8677 2465 8711 2499
rect 9505 2465 9539 2499
rect 10057 2465 10091 2499
rect 10609 2465 10643 2499
rect 11253 2465 11287 2499
rect 9689 2397 9723 2431
rect 12265 2533 12299 2567
rect 12909 2533 12943 2567
rect 15301 2533 15335 2567
rect 18797 2533 18831 2567
rect 20545 2533 20579 2567
rect 20729 2533 20763 2567
rect 22017 2533 22051 2567
rect 13461 2465 13495 2499
rect 14013 2465 14047 2499
rect 16129 2465 16163 2499
rect 17969 2465 18003 2499
rect 19441 2465 19475 2499
rect 21281 2465 21315 2499
rect 15945 2397 15979 2431
rect 16773 2397 16807 2431
rect 17693 2397 17727 2431
rect 17877 2397 17911 2431
rect 19257 2397 19291 2431
rect 11897 2329 11931 2363
rect 12081 2329 12115 2363
rect 15485 2329 15519 2363
rect 18613 2329 18647 2363
rect 21097 2329 21131 2363
rect 2697 2261 2731 2295
rect 3249 2261 3283 2295
rect 5917 2261 5951 2295
rect 8861 2261 8895 2295
rect 13001 2261 13035 2295
rect 13553 2261 13587 2295
rect 14105 2261 14139 2295
rect 18337 2261 18371 2295
rect 22109 2465 22143 2499
rect 22109 1445 22143 1479
rect 22017 1377 22051 1411
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 4447 20698
rect 4499 20646 4511 20698
rect 4563 20646 4575 20698
rect 4627 20646 4639 20698
rect 4691 20646 11378 20698
rect 11430 20646 11442 20698
rect 11494 20646 11506 20698
rect 11558 20646 11570 20698
rect 11622 20646 18308 20698
rect 18360 20646 18372 20698
rect 18424 20646 18436 20698
rect 18488 20646 18500 20698
rect 18552 20646 21896 20698
rect 1104 20624 21896 20646
rect 842 20544 848 20596
rect 900 20584 906 20596
rect 1581 20587 1639 20593
rect 1581 20584 1593 20587
rect 900 20556 1593 20584
rect 900 20544 906 20556
rect 1581 20553 1593 20556
rect 1627 20553 1639 20587
rect 5074 20584 5080 20596
rect 1581 20547 1639 20553
rect 2746 20556 5080 20584
rect 1596 20380 1624 20547
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 2746 20448 2774 20556
rect 5074 20544 5080 20556
rect 5132 20544 5138 20596
rect 8938 20544 8944 20596
rect 8996 20584 9002 20596
rect 8996 20556 12204 20584
rect 8996 20544 9002 20556
rect 4341 20519 4399 20525
rect 4341 20485 4353 20519
rect 4387 20516 4399 20519
rect 5994 20516 6000 20528
rect 4387 20488 6000 20516
rect 4387 20485 4399 20488
rect 4341 20479 4399 20485
rect 5994 20476 6000 20488
rect 6052 20476 6058 20528
rect 7098 20476 7104 20528
rect 7156 20516 7162 20528
rect 7558 20516 7564 20528
rect 7156 20488 7564 20516
rect 7156 20476 7162 20488
rect 7558 20476 7564 20488
rect 7616 20476 7622 20528
rect 8202 20476 8208 20528
rect 8260 20516 8266 20528
rect 11422 20516 11428 20528
rect 8260 20488 11428 20516
rect 8260 20476 8266 20488
rect 11422 20476 11428 20488
rect 11480 20476 11486 20528
rect 12066 20516 12072 20528
rect 12027 20488 12072 20516
rect 12066 20476 12072 20488
rect 12124 20476 12130 20528
rect 12176 20516 12204 20556
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 12308 20556 14412 20584
rect 12308 20544 12314 20556
rect 12437 20519 12495 20525
rect 12437 20516 12449 20519
rect 12176 20488 12449 20516
rect 12437 20485 12449 20488
rect 12483 20485 12495 20519
rect 12618 20516 12624 20528
rect 12579 20488 12624 20516
rect 12437 20479 12495 20485
rect 12618 20476 12624 20488
rect 12676 20476 12682 20528
rect 13170 20516 13176 20528
rect 13131 20488 13176 20516
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 13722 20516 13728 20528
rect 13683 20488 13728 20516
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 14384 20516 14412 20556
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 14516 20556 15301 20584
rect 14516 20544 14522 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 15289 20547 15347 20553
rect 16209 20587 16267 20593
rect 16209 20553 16221 20587
rect 16255 20584 16267 20587
rect 18138 20584 18144 20596
rect 16255 20556 18144 20584
rect 16255 20553 16267 20556
rect 16209 20547 16267 20553
rect 18138 20544 18144 20556
rect 18196 20544 18202 20596
rect 16390 20516 16396 20528
rect 14384 20488 16396 20516
rect 16390 20476 16396 20488
rect 16448 20476 16454 20528
rect 16853 20519 16911 20525
rect 16853 20485 16865 20519
rect 16899 20516 16911 20519
rect 17678 20516 17684 20528
rect 16899 20488 17684 20516
rect 16899 20485 16911 20488
rect 16853 20479 16911 20485
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 17865 20519 17923 20525
rect 17865 20485 17877 20519
rect 17911 20516 17923 20519
rect 17954 20516 17960 20528
rect 17911 20488 17960 20516
rect 17911 20485 17923 20488
rect 17865 20479 17923 20485
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 18417 20519 18475 20525
rect 18417 20485 18429 20519
rect 18463 20516 18475 20519
rect 18598 20516 18604 20528
rect 18463 20488 18604 20516
rect 18463 20485 18475 20488
rect 18417 20479 18475 20485
rect 18598 20476 18604 20488
rect 18656 20476 18662 20528
rect 18966 20516 18972 20528
rect 18927 20488 18972 20516
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19518 20516 19524 20528
rect 19479 20488 19524 20516
rect 19518 20476 19524 20488
rect 19576 20476 19582 20528
rect 2271 20420 2774 20448
rect 3329 20451 3387 20457
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 3329 20417 3341 20451
rect 3375 20448 3387 20451
rect 5166 20448 5172 20460
rect 3375 20420 5172 20448
rect 3375 20417 3387 20420
rect 3329 20411 3387 20417
rect 5166 20408 5172 20420
rect 5224 20408 5230 20460
rect 5537 20451 5595 20457
rect 5537 20417 5549 20451
rect 5583 20448 5595 20451
rect 6914 20448 6920 20460
rect 5583 20420 6920 20448
rect 5583 20417 5595 20420
rect 5537 20411 5595 20417
rect 6914 20408 6920 20420
rect 6972 20408 6978 20460
rect 10042 20448 10048 20460
rect 7300 20420 10048 20448
rect 2501 20383 2559 20389
rect 2501 20380 2513 20383
rect 1596 20352 2513 20380
rect 2501 20349 2513 20352
rect 2547 20349 2559 20383
rect 2501 20343 2559 20349
rect 3050 20340 3056 20392
rect 3108 20380 3114 20392
rect 3145 20383 3203 20389
rect 3145 20380 3157 20383
rect 3108 20352 3157 20380
rect 3108 20340 3114 20352
rect 3145 20349 3157 20352
rect 3191 20349 3203 20383
rect 3145 20343 3203 20349
rect 3602 20340 3608 20392
rect 3660 20380 3666 20392
rect 4157 20383 4215 20389
rect 4157 20380 4169 20383
rect 3660 20352 4169 20380
rect 3660 20340 3666 20352
rect 4157 20349 4169 20352
rect 4203 20349 4215 20383
rect 4157 20343 4215 20349
rect 5258 20340 5264 20392
rect 5316 20380 5322 20392
rect 5353 20383 5411 20389
rect 5353 20380 5365 20383
rect 5316 20352 5365 20380
rect 5316 20340 5322 20352
rect 5353 20349 5365 20352
rect 5399 20349 5411 20383
rect 5353 20343 5411 20349
rect 5810 20340 5816 20392
rect 5868 20380 5874 20392
rect 5997 20383 6055 20389
rect 5997 20380 6009 20383
rect 5868 20352 6009 20380
rect 5868 20340 5874 20352
rect 5997 20349 6009 20352
rect 6043 20349 6055 20383
rect 5997 20343 6055 20349
rect 6454 20340 6460 20392
rect 6512 20380 6518 20392
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6512 20352 6837 20380
rect 6512 20340 6518 20352
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7300 20324 7328 20420
rect 10042 20408 10048 20420
rect 10100 20408 10106 20460
rect 11977 20451 12035 20457
rect 11977 20448 11989 20451
rect 10244 20420 11989 20448
rect 7558 20340 7564 20392
rect 7616 20380 7622 20392
rect 7653 20383 7711 20389
rect 7653 20380 7665 20383
rect 7616 20352 7665 20380
rect 7616 20340 7622 20352
rect 7653 20349 7665 20352
rect 7699 20349 7711 20383
rect 8110 20380 8116 20392
rect 7653 20343 7711 20349
rect 7760 20352 8116 20380
rect 1946 20272 1952 20324
rect 2004 20312 2010 20324
rect 2041 20315 2099 20321
rect 2041 20312 2053 20315
rect 2004 20284 2053 20312
rect 2004 20272 2010 20284
rect 2041 20281 2053 20284
rect 2087 20281 2099 20315
rect 4709 20315 4767 20321
rect 4709 20312 4721 20315
rect 2041 20275 2099 20281
rect 4172 20284 4721 20312
rect 4172 20256 4200 20284
rect 4709 20281 4721 20284
rect 4755 20281 4767 20315
rect 4890 20312 4896 20324
rect 4851 20284 4896 20312
rect 4709 20275 4767 20281
rect 4890 20272 4896 20284
rect 4948 20272 4954 20324
rect 7009 20315 7067 20321
rect 7009 20281 7021 20315
rect 7055 20312 7067 20315
rect 7282 20312 7288 20324
rect 7055 20284 7288 20312
rect 7055 20281 7067 20284
rect 7009 20275 7067 20281
rect 7282 20272 7288 20284
rect 7340 20272 7346 20324
rect 7466 20272 7472 20324
rect 7524 20312 7530 20324
rect 7760 20312 7788 20352
rect 8110 20340 8116 20352
rect 8168 20380 8174 20392
rect 8205 20383 8263 20389
rect 8205 20380 8217 20383
rect 8168 20352 8217 20380
rect 8168 20340 8174 20352
rect 8205 20349 8217 20352
rect 8251 20349 8263 20383
rect 8205 20343 8263 20349
rect 8665 20383 8723 20389
rect 8665 20349 8677 20383
rect 8711 20349 8723 20383
rect 8665 20343 8723 20349
rect 7524 20284 7788 20312
rect 7837 20315 7895 20321
rect 7524 20272 7530 20284
rect 7837 20281 7849 20315
rect 7883 20312 7895 20315
rect 8386 20312 8392 20324
rect 7883 20284 8392 20312
rect 7883 20281 7895 20284
rect 7837 20275 7895 20281
rect 2682 20244 2688 20256
rect 2643 20216 2688 20244
rect 2682 20204 2688 20216
rect 2740 20204 2746 20256
rect 4154 20204 4160 20256
rect 4212 20204 4218 20256
rect 5902 20244 5908 20256
rect 5863 20216 5908 20244
rect 5902 20204 5908 20216
rect 5960 20204 5966 20256
rect 7374 20204 7380 20256
rect 7432 20244 7438 20256
rect 7852 20244 7880 20275
rect 8386 20272 8392 20284
rect 8444 20272 8450 20324
rect 8680 20312 8708 20343
rect 8754 20340 8760 20392
rect 8812 20380 8818 20392
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 8812 20352 9597 20380
rect 8812 20340 8818 20352
rect 9585 20349 9597 20352
rect 9631 20380 9643 20383
rect 10244 20380 10272 20420
rect 11977 20417 11989 20420
rect 12023 20417 12035 20451
rect 11977 20411 12035 20417
rect 12529 20451 12587 20457
rect 12529 20417 12541 20451
rect 12575 20448 12587 20451
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 12575 20420 14565 20448
rect 12575 20417 12587 20420
rect 12529 20411 12587 20417
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 18782 20448 18788 20460
rect 15795 20420 18788 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 18782 20408 18788 20420
rect 18840 20408 18846 20460
rect 20438 20448 20444 20460
rect 18892 20420 20444 20448
rect 9631 20352 10272 20380
rect 9631 20349 9643 20352
rect 9585 20343 9643 20349
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10376 20352 10701 20380
rect 10376 20340 10382 20352
rect 10689 20349 10701 20352
rect 10735 20380 10747 20383
rect 10778 20380 10784 20392
rect 10735 20352 10784 20380
rect 10735 20349 10747 20352
rect 10689 20343 10747 20349
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 12253 20383 12311 20389
rect 12253 20380 12265 20383
rect 10928 20352 12265 20380
rect 10928 20340 10934 20352
rect 12253 20349 12265 20352
rect 12299 20349 12311 20383
rect 12253 20343 12311 20349
rect 12437 20383 12495 20389
rect 12437 20349 12449 20383
rect 12483 20380 12495 20383
rect 15013 20383 15071 20389
rect 15013 20380 15025 20383
rect 12483 20352 15025 20380
rect 12483 20349 12495 20352
rect 12437 20343 12495 20349
rect 15013 20349 15025 20352
rect 15059 20349 15071 20383
rect 18892 20380 18920 20420
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 15013 20343 15071 20349
rect 17512 20352 18920 20380
rect 20073 20383 20131 20389
rect 8680 20284 9812 20312
rect 7432 20216 7880 20244
rect 8297 20247 8355 20253
rect 7432 20204 7438 20216
rect 8297 20213 8309 20247
rect 8343 20244 8355 20247
rect 8662 20244 8668 20256
rect 8343 20216 8668 20244
rect 8343 20213 8355 20216
rect 8297 20207 8355 20213
rect 8662 20204 8668 20216
rect 8720 20204 8726 20256
rect 8846 20244 8852 20256
rect 8807 20216 8852 20244
rect 8846 20204 8852 20216
rect 8904 20204 8910 20256
rect 9490 20244 9496 20256
rect 9451 20216 9496 20244
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 9784 20244 9812 20284
rect 9858 20272 9864 20324
rect 9916 20312 9922 20324
rect 10045 20315 10103 20321
rect 10045 20312 10057 20315
rect 9916 20284 10057 20312
rect 9916 20272 9922 20284
rect 10045 20281 10057 20284
rect 10091 20281 10103 20315
rect 10045 20275 10103 20281
rect 10229 20315 10287 20321
rect 10229 20281 10241 20315
rect 10275 20312 10287 20315
rect 10410 20312 10416 20324
rect 10275 20284 10416 20312
rect 10275 20281 10287 20284
rect 10229 20275 10287 20281
rect 10410 20272 10416 20284
rect 10468 20272 10474 20324
rect 10502 20272 10508 20324
rect 10560 20312 10566 20324
rect 10560 20284 10605 20312
rect 10560 20272 10566 20284
rect 11054 20272 11060 20324
rect 11112 20312 11118 20324
rect 11241 20315 11299 20321
rect 11241 20312 11253 20315
rect 11112 20284 11253 20312
rect 11112 20272 11118 20284
rect 11241 20281 11253 20284
rect 11287 20312 11299 20315
rect 11698 20312 11704 20324
rect 11287 20284 11704 20312
rect 11287 20281 11299 20284
rect 11241 20275 11299 20281
rect 11698 20272 11704 20284
rect 11756 20272 11762 20324
rect 11977 20315 12035 20321
rect 11977 20281 11989 20315
rect 12023 20312 12035 20315
rect 12529 20315 12587 20321
rect 12529 20312 12541 20315
rect 12023 20284 12541 20312
rect 12023 20281 12035 20284
rect 11977 20275 12035 20281
rect 12529 20281 12541 20284
rect 12575 20281 12587 20315
rect 12802 20312 12808 20324
rect 12763 20284 12808 20312
rect 12529 20275 12587 20281
rect 12802 20272 12808 20284
rect 12860 20272 12866 20324
rect 13357 20315 13415 20321
rect 13357 20281 13369 20315
rect 13403 20312 13415 20315
rect 13722 20312 13728 20324
rect 13403 20284 13728 20312
rect 13403 20281 13415 20284
rect 13357 20275 13415 20281
rect 13722 20272 13728 20284
rect 13780 20272 13786 20324
rect 13906 20312 13912 20324
rect 13867 20284 13912 20312
rect 13906 20272 13912 20284
rect 13964 20272 13970 20324
rect 15197 20315 15255 20321
rect 15197 20281 15209 20315
rect 15243 20281 15255 20315
rect 15197 20275 15255 20281
rect 15289 20315 15347 20321
rect 15289 20281 15301 20315
rect 15335 20312 15347 20315
rect 15565 20315 15623 20321
rect 15565 20312 15577 20315
rect 15335 20284 15577 20312
rect 15335 20281 15347 20284
rect 15289 20275 15347 20281
rect 15565 20281 15577 20284
rect 15611 20281 15623 20315
rect 16114 20312 16120 20324
rect 16075 20284 16120 20312
rect 15565 20275 15623 20281
rect 9950 20244 9956 20256
rect 9784 20216 9956 20244
rect 9950 20204 9956 20216
rect 10008 20204 10014 20256
rect 11146 20244 11152 20256
rect 11107 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 15212 20244 15240 20275
rect 16114 20272 16120 20284
rect 16172 20272 16178 20324
rect 16666 20312 16672 20324
rect 16627 20284 16672 20312
rect 16666 20272 16672 20284
rect 16724 20272 16730 20324
rect 17512 20312 17540 20352
rect 20073 20349 20085 20383
rect 20119 20380 20131 20383
rect 20162 20380 20168 20392
rect 20119 20352 20168 20380
rect 20119 20349 20131 20352
rect 20073 20343 20131 20349
rect 20162 20340 20168 20352
rect 20220 20340 20226 20392
rect 17678 20312 17684 20324
rect 17144 20284 17540 20312
rect 17639 20284 17684 20312
rect 17144 20244 17172 20284
rect 17678 20272 17684 20284
rect 17736 20272 17742 20324
rect 17954 20272 17960 20324
rect 18012 20312 18018 20324
rect 18233 20315 18291 20321
rect 18233 20312 18245 20315
rect 18012 20284 18245 20312
rect 18012 20272 18018 20284
rect 18233 20281 18245 20284
rect 18279 20281 18291 20315
rect 18782 20312 18788 20324
rect 18743 20284 18788 20312
rect 18233 20275 18291 20281
rect 18782 20272 18788 20284
rect 18840 20272 18846 20324
rect 19337 20315 19395 20321
rect 19337 20281 19349 20315
rect 19383 20312 19395 20315
rect 19426 20312 19432 20324
rect 19383 20284 19432 20312
rect 19383 20281 19395 20284
rect 19337 20275 19395 20281
rect 19426 20272 19432 20284
rect 19484 20272 19490 20324
rect 20622 20312 20628 20324
rect 20583 20284 20628 20312
rect 20622 20272 20628 20284
rect 20680 20272 20686 20324
rect 20806 20312 20812 20324
rect 20767 20284 20812 20312
rect 20806 20272 20812 20284
rect 20864 20272 20870 20324
rect 21174 20312 21180 20324
rect 21135 20284 21180 20312
rect 21174 20272 21180 20284
rect 21232 20272 21238 20324
rect 21361 20315 21419 20321
rect 21361 20281 21373 20315
rect 21407 20312 21419 20315
rect 21450 20312 21456 20324
rect 21407 20284 21456 20312
rect 21407 20281 21419 20284
rect 21361 20275 21419 20281
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 15212 20216 17172 20244
rect 17218 20204 17224 20256
rect 17276 20244 17282 20256
rect 20257 20247 20315 20253
rect 17276 20216 17321 20244
rect 17276 20204 17282 20216
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 21082 20244 21088 20256
rect 20303 20216 21088 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 1104 20154 21896 20176
rect 1104 20102 7912 20154
rect 7964 20102 7976 20154
rect 8028 20102 8040 20154
rect 8092 20102 8104 20154
rect 8156 20102 14843 20154
rect 14895 20102 14907 20154
rect 14959 20102 14971 20154
rect 15023 20102 15035 20154
rect 15087 20102 21896 20154
rect 1104 20080 21896 20102
rect 2314 20040 2320 20052
rect 2275 20012 2320 20040
rect 2314 20000 2320 20012
rect 2372 20000 2378 20052
rect 3050 20000 3056 20052
rect 3108 20040 3114 20052
rect 3421 20043 3479 20049
rect 3421 20040 3433 20043
rect 3108 20012 3433 20040
rect 3108 20000 3114 20012
rect 3421 20009 3433 20012
rect 3467 20009 3479 20043
rect 3421 20003 3479 20009
rect 3602 20000 3608 20052
rect 3660 20040 3666 20052
rect 3881 20043 3939 20049
rect 3881 20040 3893 20043
rect 3660 20012 3893 20040
rect 3660 20000 3666 20012
rect 3881 20009 3893 20012
rect 3927 20009 3939 20043
rect 3881 20003 3939 20009
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4341 20043 4399 20049
rect 4341 20040 4353 20043
rect 4212 20012 4353 20040
rect 4212 20000 4218 20012
rect 4341 20009 4353 20012
rect 4387 20009 4399 20043
rect 4341 20003 4399 20009
rect 4893 20043 4951 20049
rect 4893 20009 4905 20043
rect 4939 20009 4951 20043
rect 4893 20003 4951 20009
rect 5813 20043 5871 20049
rect 5813 20009 5825 20043
rect 5859 20040 5871 20043
rect 7098 20040 7104 20052
rect 5859 20012 7104 20040
rect 5859 20009 5871 20012
rect 5813 20003 5871 20009
rect 1394 19932 1400 19984
rect 1452 19972 1458 19984
rect 1946 19972 1952 19984
rect 1452 19944 1952 19972
rect 1452 19932 1458 19944
rect 1946 19932 1952 19944
rect 2004 19972 2010 19984
rect 4908 19972 4936 20003
rect 7098 20000 7104 20012
rect 7156 20000 7162 20052
rect 7837 20043 7895 20049
rect 7837 20009 7849 20043
rect 7883 20040 7895 20043
rect 8202 20040 8208 20052
rect 7883 20012 8208 20040
rect 7883 20009 7895 20012
rect 7837 20003 7895 20009
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 8297 20043 8355 20049
rect 8297 20009 8309 20043
rect 8343 20009 8355 20043
rect 8297 20003 8355 20009
rect 8757 20043 8815 20049
rect 8757 20009 8769 20043
rect 8803 20040 8815 20043
rect 8938 20040 8944 20052
rect 8803 20012 8944 20040
rect 8803 20009 8815 20012
rect 8757 20003 8815 20009
rect 8312 19972 8340 20003
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 9585 20043 9643 20049
rect 9585 20009 9597 20043
rect 9631 20040 9643 20043
rect 9631 20012 11376 20040
rect 9631 20009 9643 20012
rect 9585 20003 9643 20009
rect 9766 19972 9772 19984
rect 2004 19944 2176 19972
rect 4908 19944 8248 19972
rect 8312 19944 9772 19972
rect 2004 19932 2010 19944
rect 1670 19904 1676 19916
rect 1631 19876 1676 19904
rect 1670 19864 1676 19876
rect 1728 19864 1734 19916
rect 2148 19913 2176 19944
rect 2133 19907 2191 19913
rect 2133 19873 2145 19907
rect 2179 19873 2191 19907
rect 2133 19867 2191 19873
rect 2498 19864 2504 19916
rect 2556 19904 2562 19916
rect 2593 19907 2651 19913
rect 2593 19904 2605 19907
rect 2556 19876 2605 19904
rect 2556 19864 2562 19876
rect 2593 19873 2605 19876
rect 2639 19873 2651 19907
rect 2593 19867 2651 19873
rect 4709 19907 4767 19913
rect 4709 19873 4721 19907
rect 4755 19904 4767 19907
rect 4798 19904 4804 19916
rect 4755 19876 4804 19904
rect 4755 19873 4767 19876
rect 4709 19867 4767 19873
rect 4798 19864 4804 19876
rect 4856 19864 4862 19916
rect 6086 19904 6092 19916
rect 6047 19876 6092 19904
rect 6086 19864 6092 19876
rect 6144 19864 6150 19916
rect 6546 19904 6552 19916
rect 6507 19876 6552 19904
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7006 19904 7012 19916
rect 6967 19876 7012 19904
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 7650 19904 7656 19916
rect 7611 19876 7656 19904
rect 7650 19864 7656 19876
rect 7708 19864 7714 19916
rect 8110 19904 8116 19916
rect 8071 19876 8116 19904
rect 8110 19864 8116 19876
rect 8168 19864 8174 19916
rect 8220 19904 8248 19944
rect 9766 19932 9772 19944
rect 9824 19932 9830 19984
rect 10042 19932 10048 19984
rect 10100 19972 10106 19984
rect 10137 19975 10195 19981
rect 10137 19972 10149 19975
rect 10100 19944 10149 19972
rect 10100 19932 10106 19944
rect 10137 19941 10149 19944
rect 10183 19941 10195 19975
rect 10137 19935 10195 19941
rect 10229 19975 10287 19981
rect 10229 19941 10241 19975
rect 10275 19972 10287 19975
rect 11348 19972 11376 20012
rect 11422 20000 11428 20052
rect 11480 20040 11486 20052
rect 11480 20012 13584 20040
rect 11480 20000 11486 20012
rect 10275 19944 10364 19972
rect 11348 19944 12020 19972
rect 10275 19941 10287 19944
rect 10229 19935 10287 19941
rect 10336 19916 10364 19944
rect 8386 19904 8392 19916
rect 8220 19876 8392 19904
rect 8386 19864 8392 19876
rect 8444 19864 8450 19916
rect 8570 19904 8576 19916
rect 8483 19876 8576 19904
rect 8570 19864 8576 19876
rect 8628 19904 8634 19916
rect 9306 19904 9312 19916
rect 8628 19876 9312 19904
rect 8628 19864 8634 19876
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 9401 19907 9459 19913
rect 9401 19873 9413 19907
rect 9447 19904 9459 19907
rect 9582 19904 9588 19916
rect 9447 19876 9588 19904
rect 9447 19873 9459 19876
rect 9401 19867 9459 19873
rect 9582 19864 9588 19876
rect 9640 19864 9646 19916
rect 10318 19864 10324 19916
rect 10376 19864 10382 19916
rect 11054 19864 11060 19916
rect 11112 19904 11118 19916
rect 11221 19907 11279 19913
rect 11221 19904 11233 19907
rect 11112 19876 11233 19904
rect 11112 19864 11118 19876
rect 11221 19873 11233 19876
rect 11267 19873 11279 19907
rect 11221 19867 11279 19873
rect 2038 19796 2044 19848
rect 2096 19836 2102 19848
rect 3053 19839 3111 19845
rect 3053 19836 3065 19839
rect 2096 19808 3065 19836
rect 2096 19796 2102 19808
rect 3053 19805 3065 19808
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 5445 19839 5503 19845
rect 5445 19805 5457 19839
rect 5491 19836 5503 19839
rect 6638 19836 6644 19848
rect 5491 19808 6644 19836
rect 5491 19805 5503 19808
rect 5445 19799 5503 19805
rect 6638 19796 6644 19808
rect 6696 19796 6702 19848
rect 6822 19796 6828 19848
rect 6880 19836 6886 19848
rect 9858 19836 9864 19848
rect 6880 19808 9864 19836
rect 6880 19796 6886 19808
rect 9858 19796 9864 19808
rect 9916 19796 9922 19848
rect 10042 19836 10048 19848
rect 10003 19808 10048 19836
rect 10042 19796 10048 19808
rect 10100 19796 10106 19848
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 2774 19728 2780 19780
rect 2832 19768 2838 19780
rect 7190 19768 7196 19780
rect 2832 19740 2877 19768
rect 7151 19740 7196 19768
rect 2832 19728 2838 19740
rect 7190 19728 7196 19740
rect 7248 19728 7254 19780
rect 8110 19728 8116 19780
rect 8168 19768 8174 19780
rect 10134 19768 10140 19780
rect 8168 19740 10140 19768
rect 8168 19728 8174 19740
rect 10134 19728 10140 19740
rect 10192 19728 10198 19780
rect 10226 19728 10232 19780
rect 10284 19768 10290 19780
rect 10980 19768 11008 19796
rect 10284 19740 11008 19768
rect 11992 19768 12020 19944
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 13081 19975 13139 19981
rect 13081 19972 13093 19975
rect 12124 19944 13093 19972
rect 12124 19932 12130 19944
rect 13081 19941 13093 19944
rect 13127 19941 13139 19975
rect 13081 19935 13139 19941
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 13173 19907 13231 19913
rect 13173 19904 13185 19907
rect 12952 19876 13185 19904
rect 12952 19864 12958 19876
rect 13173 19873 13185 19876
rect 13219 19873 13231 19907
rect 13173 19867 13231 19873
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19836 13047 19839
rect 13262 19836 13268 19848
rect 13035 19808 13268 19836
rect 13035 19805 13047 19808
rect 12989 19799 13047 19805
rect 13262 19796 13268 19808
rect 13320 19796 13326 19848
rect 13556 19836 13584 20012
rect 13722 20000 13728 20052
rect 13780 20040 13786 20052
rect 13817 20043 13875 20049
rect 13817 20040 13829 20043
rect 13780 20012 13829 20040
rect 13780 20000 13786 20012
rect 13817 20009 13829 20012
rect 13863 20009 13875 20043
rect 14458 20040 14464 20052
rect 13817 20003 13875 20009
rect 13924 20012 14464 20040
rect 13814 19864 13820 19916
rect 13872 19904 13878 19916
rect 13924 19904 13952 20012
rect 14458 20000 14464 20012
rect 14516 20000 14522 20052
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 14792 20012 15148 20040
rect 14792 20000 14798 20012
rect 14274 19932 14280 19984
rect 14332 19972 14338 19984
rect 15120 19981 15148 20012
rect 15194 20000 15200 20052
rect 15252 20000 15258 20052
rect 18141 20043 18199 20049
rect 18141 20009 18153 20043
rect 18187 20040 18199 20043
rect 18782 20040 18788 20052
rect 18187 20012 18788 20040
rect 18187 20009 18199 20012
rect 18141 20003 18199 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 19153 20043 19211 20049
rect 19153 20009 19165 20043
rect 19199 20040 19211 20043
rect 21542 20040 21548 20052
rect 19199 20012 21548 20040
rect 19199 20009 19211 20012
rect 19153 20003 19211 20009
rect 21542 20000 21548 20012
rect 21600 20000 21606 20052
rect 14553 19975 14611 19981
rect 14553 19972 14565 19975
rect 14332 19944 14565 19972
rect 14332 19932 14338 19944
rect 14553 19941 14565 19944
rect 14599 19941 14611 19975
rect 14553 19935 14611 19941
rect 15105 19975 15163 19981
rect 15105 19941 15117 19975
rect 15151 19941 15163 19975
rect 15212 19972 15240 20000
rect 15289 19975 15347 19981
rect 15289 19972 15301 19975
rect 15212 19944 15301 19972
rect 15105 19935 15163 19941
rect 15289 19941 15301 19944
rect 15335 19941 15347 19975
rect 15289 19935 15347 19941
rect 15378 19932 15384 19984
rect 15436 19972 15442 19984
rect 15657 19975 15715 19981
rect 15657 19972 15669 19975
rect 15436 19944 15669 19972
rect 15436 19932 15442 19944
rect 15657 19941 15669 19944
rect 15703 19941 15715 19975
rect 15657 19935 15715 19941
rect 15930 19932 15936 19984
rect 15988 19972 15994 19984
rect 16209 19975 16267 19981
rect 16209 19972 16221 19975
rect 15988 19944 16221 19972
rect 15988 19932 15994 19944
rect 16209 19941 16221 19944
rect 16255 19941 16267 19975
rect 16390 19972 16396 19984
rect 16351 19944 16396 19972
rect 16209 19935 16267 19941
rect 16390 19932 16396 19944
rect 16448 19932 16454 19984
rect 16574 19932 16580 19984
rect 16632 19972 16638 19984
rect 16761 19975 16819 19981
rect 16761 19972 16773 19975
rect 16632 19944 16773 19972
rect 16632 19932 16638 19944
rect 16761 19941 16773 19944
rect 16807 19941 16819 19975
rect 16761 19935 16819 19941
rect 17034 19932 17040 19984
rect 17092 19972 17098 19984
rect 17313 19975 17371 19981
rect 17313 19972 17325 19975
rect 17092 19944 17325 19972
rect 17092 19932 17098 19944
rect 17313 19941 17325 19944
rect 17359 19941 17371 19975
rect 17313 19935 17371 19941
rect 19334 19932 19340 19984
rect 19392 19972 19398 19984
rect 19797 19975 19855 19981
rect 19797 19972 19809 19975
rect 19392 19944 19809 19972
rect 19392 19932 19398 19944
rect 19797 19941 19809 19944
rect 19843 19941 19855 19975
rect 19797 19935 19855 19941
rect 19886 19932 19892 19984
rect 19944 19972 19950 19984
rect 20349 19975 20407 19981
rect 20349 19972 20361 19975
rect 19944 19944 20361 19972
rect 19944 19932 19950 19944
rect 20349 19941 20361 19944
rect 20395 19941 20407 19975
rect 20349 19935 20407 19941
rect 13872 19876 13952 19904
rect 14001 19907 14059 19913
rect 13872 19864 13878 19876
rect 14001 19873 14013 19907
rect 14047 19904 14059 19907
rect 14458 19904 14464 19916
rect 14047 19876 14464 19904
rect 14047 19873 14059 19876
rect 14001 19867 14059 19873
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 14737 19907 14795 19913
rect 14737 19873 14749 19907
rect 14783 19904 14795 19907
rect 15194 19904 15200 19916
rect 14783 19876 15200 19904
rect 14783 19873 14795 19876
rect 14737 19867 14795 19873
rect 15194 19864 15200 19876
rect 15252 19864 15258 19916
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19904 15531 19907
rect 15841 19907 15899 19913
rect 15841 19904 15853 19907
rect 15519 19876 15853 19904
rect 15519 19873 15531 19876
rect 15473 19867 15531 19873
rect 15841 19873 15853 19876
rect 15887 19873 15899 19907
rect 16942 19904 16948 19916
rect 16903 19876 16948 19904
rect 15841 19867 15899 19873
rect 16942 19864 16948 19876
rect 17000 19864 17006 19916
rect 17494 19904 17500 19916
rect 17455 19876 17500 19904
rect 17494 19864 17500 19876
rect 17552 19864 17558 19916
rect 17957 19907 18015 19913
rect 17957 19873 17969 19907
rect 18003 19873 18015 19907
rect 18506 19904 18512 19916
rect 18467 19876 18512 19904
rect 17957 19867 18015 19873
rect 17972 19836 18000 19867
rect 18506 19864 18512 19876
rect 18564 19864 18570 19916
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 19061 19907 19119 19913
rect 19061 19904 19073 19907
rect 18656 19876 19073 19904
rect 18656 19864 18662 19876
rect 19061 19873 19073 19876
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 19610 19864 19616 19916
rect 19668 19904 19674 19916
rect 19981 19907 20039 19913
rect 19981 19904 19993 19907
rect 19668 19876 19993 19904
rect 19668 19864 19674 19876
rect 19981 19873 19993 19876
rect 20027 19873 20039 19907
rect 20530 19904 20536 19916
rect 20491 19876 20536 19904
rect 19981 19867 20039 19873
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 21177 19907 21235 19913
rect 21177 19873 21189 19907
rect 21223 19873 21235 19907
rect 21177 19867 21235 19873
rect 13556 19808 18000 19836
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 21192 19836 21220 19867
rect 19392 19808 21220 19836
rect 19392 19796 19398 19808
rect 16666 19768 16672 19780
rect 11992 19740 16672 19768
rect 10284 19728 10290 19740
rect 16666 19728 16672 19740
rect 16724 19728 16730 19780
rect 21358 19768 21364 19780
rect 21319 19740 21364 19768
rect 21358 19728 21364 19740
rect 21416 19728 21422 19780
rect 1762 19700 1768 19712
rect 1723 19672 1768 19700
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 6273 19703 6331 19709
rect 6273 19669 6285 19703
rect 6319 19700 6331 19703
rect 6638 19700 6644 19712
rect 6319 19672 6644 19700
rect 6319 19669 6331 19672
rect 6273 19663 6331 19669
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 6733 19703 6791 19709
rect 6733 19669 6745 19703
rect 6779 19700 6791 19703
rect 6822 19700 6828 19712
rect 6779 19672 6828 19700
rect 6779 19669 6791 19672
rect 6733 19663 6791 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 7098 19660 7104 19712
rect 7156 19700 7162 19712
rect 10318 19700 10324 19712
rect 7156 19672 10324 19700
rect 7156 19660 7162 19672
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 10597 19703 10655 19709
rect 10597 19669 10609 19703
rect 10643 19700 10655 19703
rect 11238 19700 11244 19712
rect 10643 19672 11244 19700
rect 10643 19669 10655 19672
rect 10597 19663 10655 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 12342 19700 12348 19712
rect 12303 19672 12348 19700
rect 12342 19660 12348 19672
rect 12400 19660 12406 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 14366 19700 14372 19712
rect 13587 19672 14372 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 14550 19660 14556 19712
rect 14608 19700 14614 19712
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 14608 19672 15485 19700
rect 14608 19660 14614 19672
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15473 19663 15531 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 22094 19700 22100 19712
rect 18647 19672 22100 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 1104 19610 21896 19632
rect 1104 19558 4447 19610
rect 4499 19558 4511 19610
rect 4563 19558 4575 19610
rect 4627 19558 4639 19610
rect 4691 19558 11378 19610
rect 11430 19558 11442 19610
rect 11494 19558 11506 19610
rect 11558 19558 11570 19610
rect 11622 19558 18308 19610
rect 18360 19558 18372 19610
rect 18424 19558 18436 19610
rect 18488 19558 18500 19610
rect 18552 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19496 1952 19508
rect 1907 19468 1952 19496
rect 1946 19456 1952 19468
rect 2004 19456 2010 19508
rect 2498 19496 2504 19508
rect 2459 19468 2504 19496
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 4798 19456 4804 19508
rect 4856 19496 4862 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 4856 19468 4997 19496
rect 4856 19456 4862 19468
rect 4985 19465 4997 19468
rect 5031 19465 5043 19499
rect 4985 19459 5043 19465
rect 6454 19456 6460 19508
rect 6512 19496 6518 19508
rect 6549 19499 6607 19505
rect 6549 19496 6561 19499
rect 6512 19468 6561 19496
rect 6512 19456 6518 19468
rect 6549 19465 6561 19468
rect 6595 19465 6607 19499
rect 6549 19459 6607 19465
rect 6638 19456 6644 19508
rect 6696 19496 6702 19508
rect 12894 19496 12900 19508
rect 6696 19468 12900 19496
rect 6696 19456 6702 19468
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 13262 19496 13268 19508
rect 13223 19468 13268 19496
rect 13262 19456 13268 19468
rect 13320 19456 13326 19508
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 13403 19468 14504 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 7101 19431 7159 19437
rect 7101 19397 7113 19431
rect 7147 19428 7159 19431
rect 9677 19431 9735 19437
rect 7147 19400 8248 19428
rect 7147 19397 7159 19400
rect 7101 19391 7159 19397
rect 7282 19360 7288 19372
rect 6932 19332 7288 19360
rect 290 19252 296 19304
rect 348 19292 354 19304
rect 1397 19295 1455 19301
rect 1397 19292 1409 19295
rect 348 19264 1409 19292
rect 348 19252 354 19264
rect 1397 19261 1409 19264
rect 1443 19292 1455 19295
rect 1670 19292 1676 19304
rect 1443 19264 1676 19292
rect 1443 19261 1455 19264
rect 1397 19255 1455 19261
rect 1670 19252 1676 19264
rect 1728 19252 1734 19304
rect 5258 19252 5264 19304
rect 5316 19292 5322 19304
rect 5629 19295 5687 19301
rect 5629 19292 5641 19295
rect 5316 19264 5641 19292
rect 5316 19252 5322 19264
rect 5629 19261 5641 19264
rect 5675 19261 5687 19295
rect 6932 19292 6960 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7558 19320 7564 19372
rect 7616 19360 7622 19372
rect 7616 19332 7788 19360
rect 7616 19320 7622 19332
rect 5629 19255 5687 19261
rect 5736 19264 6960 19292
rect 4341 19227 4399 19233
rect 4341 19193 4353 19227
rect 4387 19224 4399 19227
rect 5736 19224 5764 19264
rect 7098 19252 7104 19304
rect 7156 19292 7162 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7156 19264 7205 19292
rect 7156 19252 7162 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 7432 19264 7665 19292
rect 7432 19252 7438 19264
rect 7653 19261 7665 19264
rect 7699 19261 7711 19295
rect 7760 19292 7788 19332
rect 8113 19295 8171 19301
rect 8113 19292 8125 19295
rect 7760 19264 8125 19292
rect 7653 19255 7711 19261
rect 8113 19261 8125 19264
rect 8159 19261 8171 19295
rect 8220 19292 8248 19400
rect 9677 19397 9689 19431
rect 9723 19397 9735 19431
rect 9677 19391 9735 19397
rect 9692 19360 9720 19391
rect 9692 19332 10088 19360
rect 8573 19295 8631 19301
rect 8573 19292 8585 19295
rect 8220 19264 8585 19292
rect 8113 19255 8171 19261
rect 8573 19261 8585 19264
rect 8619 19292 8631 19295
rect 8846 19292 8852 19304
rect 8619 19264 8852 19292
rect 8619 19261 8631 19264
rect 8573 19255 8631 19261
rect 8846 19252 8852 19264
rect 8904 19252 8910 19304
rect 9030 19292 9036 19304
rect 8991 19264 9036 19292
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 9214 19292 9220 19304
rect 9140 19264 9220 19292
rect 4387 19196 5764 19224
rect 6089 19227 6147 19233
rect 4387 19193 4399 19196
rect 4341 19187 4399 19193
rect 6089 19193 6101 19227
rect 6135 19224 6147 19227
rect 6546 19224 6552 19236
rect 6135 19196 6552 19224
rect 6135 19193 6147 19196
rect 6089 19187 6147 19193
rect 6546 19184 6552 19196
rect 6604 19224 6610 19236
rect 9140 19224 9168 19264
rect 9214 19252 9220 19264
rect 9272 19252 9278 19304
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 9674 19292 9680 19304
rect 9539 19264 9680 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19292 9919 19295
rect 9953 19295 10011 19301
rect 9953 19292 9965 19295
rect 9907 19264 9965 19292
rect 9907 19261 9919 19264
rect 9861 19255 9919 19261
rect 9953 19261 9965 19264
rect 9999 19261 10011 19295
rect 10060 19292 10088 19332
rect 10962 19320 10968 19372
rect 11020 19360 11026 19372
rect 13280 19360 13308 19456
rect 14476 19428 14504 19468
rect 14734 19456 14740 19508
rect 14792 19496 14798 19508
rect 17218 19496 17224 19508
rect 14792 19468 17224 19496
rect 14792 19456 14798 19468
rect 17218 19456 17224 19468
rect 17276 19456 17282 19508
rect 18601 19499 18659 19505
rect 18601 19465 18613 19499
rect 18647 19496 18659 19499
rect 20622 19496 20628 19508
rect 18647 19468 20628 19496
rect 18647 19465 18659 19468
rect 18601 19459 18659 19465
rect 20622 19456 20628 19468
rect 20680 19456 20686 19508
rect 16114 19428 16120 19440
rect 14476 19400 16120 19428
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 19426 19428 19432 19440
rect 19168 19400 19432 19428
rect 15013 19363 15071 19369
rect 11020 19332 11652 19360
rect 13280 19332 13676 19360
rect 11020 19320 11026 19332
rect 10594 19292 10600 19304
rect 10060 19264 10600 19292
rect 9953 19255 10011 19261
rect 10594 19252 10600 19264
rect 10652 19252 10658 19304
rect 11624 19292 11652 19332
rect 11793 19295 11851 19301
rect 11793 19292 11805 19295
rect 11624 19264 11805 19292
rect 11793 19261 11805 19264
rect 11839 19292 11851 19295
rect 11885 19295 11943 19301
rect 11885 19292 11897 19295
rect 11839 19264 11897 19292
rect 11839 19261 11851 19264
rect 11793 19255 11851 19261
rect 11885 19261 11897 19264
rect 11931 19261 11943 19295
rect 13357 19295 13415 19301
rect 13357 19292 13369 19295
rect 11885 19255 11943 19261
rect 11992 19264 13369 19292
rect 10220 19227 10278 19233
rect 6604 19196 9168 19224
rect 9232 19196 10180 19224
rect 6604 19184 6610 19196
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 6178 19156 6184 19168
rect 4755 19128 6184 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 6270 19116 6276 19168
rect 6328 19156 6334 19168
rect 7101 19159 7159 19165
rect 7101 19156 7113 19159
rect 6328 19128 7113 19156
rect 6328 19116 6334 19128
rect 7101 19125 7113 19128
rect 7147 19125 7159 19159
rect 7374 19156 7380 19168
rect 7335 19128 7380 19156
rect 7101 19119 7159 19125
rect 7374 19116 7380 19128
rect 7432 19116 7438 19168
rect 7742 19116 7748 19168
rect 7800 19156 7806 19168
rect 7837 19159 7895 19165
rect 7837 19156 7849 19159
rect 7800 19128 7849 19156
rect 7800 19116 7806 19128
rect 7837 19125 7849 19128
rect 7883 19125 7895 19159
rect 8294 19156 8300 19168
rect 8255 19128 8300 19156
rect 7837 19119 7895 19125
rect 8294 19116 8300 19128
rect 8352 19116 8358 19168
rect 8754 19156 8760 19168
rect 8715 19128 8760 19156
rect 8754 19116 8760 19128
rect 8812 19116 8818 19168
rect 9232 19165 9260 19196
rect 9217 19159 9275 19165
rect 9217 19125 9229 19159
rect 9263 19125 9275 19159
rect 9217 19119 9275 19125
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9861 19159 9919 19165
rect 9861 19156 9873 19159
rect 9364 19128 9873 19156
rect 9364 19116 9370 19128
rect 9861 19125 9873 19128
rect 9907 19156 9919 19159
rect 10042 19156 10048 19168
rect 9907 19128 10048 19156
rect 9907 19125 9919 19128
rect 9861 19119 9919 19125
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 10152 19156 10180 19196
rect 10220 19193 10232 19227
rect 10266 19224 10278 19227
rect 10686 19224 10692 19236
rect 10266 19196 10692 19224
rect 10266 19193 10278 19196
rect 10220 19187 10278 19193
rect 10686 19184 10692 19196
rect 10744 19184 10750 19236
rect 11992 19224 12020 19264
rect 13357 19261 13369 19264
rect 13403 19261 13415 19295
rect 13357 19255 13415 19261
rect 13449 19295 13507 19301
rect 13449 19261 13461 19295
rect 13495 19292 13507 19295
rect 13541 19295 13599 19301
rect 13541 19292 13553 19295
rect 13495 19264 13553 19292
rect 13495 19261 13507 19264
rect 13449 19255 13507 19261
rect 13541 19261 13553 19264
rect 13587 19261 13599 19295
rect 13648 19292 13676 19332
rect 15013 19329 15025 19363
rect 15059 19360 15071 19363
rect 15289 19363 15347 19369
rect 15289 19360 15301 19363
rect 15059 19332 15301 19360
rect 15059 19329 15071 19332
rect 15013 19323 15071 19329
rect 15289 19329 15301 19332
rect 15335 19329 15347 19363
rect 18598 19360 18604 19372
rect 15289 19323 15347 19329
rect 15396 19332 18604 19360
rect 13797 19295 13855 19301
rect 13797 19292 13809 19295
rect 13648 19264 13809 19292
rect 13541 19255 13599 19261
rect 13797 19261 13809 19264
rect 13843 19261 13855 19295
rect 13797 19255 13855 19261
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 15396 19292 15424 19332
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 16945 19295 17003 19301
rect 16945 19292 16957 19295
rect 14332 19264 15424 19292
rect 15488 19264 16957 19292
rect 14332 19252 14338 19264
rect 12158 19233 12164 19236
rect 12152 19224 12164 19233
rect 11256 19196 12020 19224
rect 12071 19196 12164 19224
rect 11256 19156 11284 19196
rect 12152 19187 12164 19196
rect 12216 19224 12222 19236
rect 12342 19224 12348 19236
rect 12216 19196 12348 19224
rect 12158 19184 12164 19187
rect 12216 19184 12222 19196
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 12434 19184 12440 19236
rect 12492 19224 12498 19236
rect 15488 19233 15516 19264
rect 16945 19261 16957 19264
rect 16991 19261 17003 19295
rect 16945 19255 17003 19261
rect 17034 19252 17040 19304
rect 17092 19292 17098 19304
rect 17497 19295 17555 19301
rect 17497 19292 17509 19295
rect 17092 19264 17509 19292
rect 17092 19252 17098 19264
rect 17497 19261 17509 19264
rect 17543 19261 17555 19295
rect 17497 19255 17555 19261
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 17957 19295 18015 19301
rect 17957 19292 17969 19295
rect 17644 19264 17969 19292
rect 17644 19252 17650 19264
rect 17957 19261 17969 19264
rect 18003 19261 18015 19295
rect 18414 19292 18420 19304
rect 18375 19264 18420 19292
rect 17957 19255 18015 19261
rect 18414 19252 18420 19264
rect 18472 19252 18478 19304
rect 18877 19295 18935 19301
rect 18877 19261 18889 19295
rect 18923 19292 18935 19295
rect 19058 19292 19064 19304
rect 18923 19264 19064 19292
rect 18923 19261 18935 19264
rect 18877 19255 18935 19261
rect 19058 19252 19064 19264
rect 19116 19252 19122 19304
rect 15473 19227 15531 19233
rect 15473 19224 15485 19227
rect 12492 19196 15485 19224
rect 12492 19184 12498 19196
rect 15473 19193 15485 19196
rect 15519 19193 15531 19227
rect 15473 19187 15531 19193
rect 15565 19227 15623 19233
rect 15565 19193 15577 19227
rect 15611 19224 15623 19227
rect 16209 19227 16267 19233
rect 16209 19224 16221 19227
rect 15611 19196 16221 19224
rect 15611 19193 15623 19196
rect 15565 19187 15623 19193
rect 16209 19193 16221 19196
rect 16255 19193 16267 19227
rect 19168 19224 19196 19400
rect 19426 19388 19432 19400
rect 19484 19388 19490 19440
rect 19260 19332 19564 19360
rect 19260 19304 19288 19332
rect 19242 19252 19248 19304
rect 19300 19252 19306 19304
rect 19337 19295 19395 19301
rect 19337 19261 19349 19295
rect 19383 19261 19395 19295
rect 19536 19292 19564 19332
rect 20625 19295 20683 19301
rect 20625 19292 20637 19295
rect 19536 19264 20637 19292
rect 19337 19255 19395 19261
rect 20625 19261 20637 19264
rect 20671 19261 20683 19295
rect 20625 19255 20683 19261
rect 16209 19187 16267 19193
rect 18156 19196 19196 19224
rect 19352 19224 19380 19255
rect 21082 19252 21088 19304
rect 21140 19292 21146 19304
rect 21177 19295 21235 19301
rect 21177 19292 21189 19295
rect 21140 19264 21189 19292
rect 21140 19252 21146 19264
rect 21177 19261 21189 19264
rect 21223 19261 21235 19295
rect 21177 19255 21235 19261
rect 19702 19224 19708 19236
rect 19352 19196 19708 19224
rect 10152 19128 11284 19156
rect 11333 19159 11391 19165
rect 11333 19125 11345 19159
rect 11379 19156 11391 19159
rect 11422 19156 11428 19168
rect 11379 19128 11428 19156
rect 11379 19125 11391 19128
rect 11333 19119 11391 19125
rect 11422 19116 11428 19128
rect 11480 19116 11486 19168
rect 11793 19159 11851 19165
rect 11793 19125 11805 19159
rect 11839 19156 11851 19159
rect 12710 19156 12716 19168
rect 11839 19128 12716 19156
rect 11839 19125 11851 19128
rect 11793 19119 11851 19125
rect 12710 19116 12716 19128
rect 12768 19156 12774 19168
rect 13449 19159 13507 19165
rect 13449 19156 13461 19159
rect 12768 19128 13461 19156
rect 12768 19116 12774 19128
rect 13449 19125 13461 19128
rect 13495 19125 13507 19159
rect 13449 19119 13507 19125
rect 14182 19116 14188 19168
rect 14240 19156 14246 19168
rect 14921 19159 14979 19165
rect 14921 19156 14933 19159
rect 14240 19128 14933 19156
rect 14240 19116 14246 19128
rect 14921 19125 14933 19128
rect 14967 19156 14979 19159
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14967 19128 15025 19156
rect 14967 19125 14979 19128
rect 14921 19119 14979 19125
rect 15013 19125 15025 19128
rect 15059 19125 15071 19159
rect 15013 19119 15071 19125
rect 15933 19159 15991 19165
rect 15933 19125 15945 19159
rect 15979 19156 15991 19159
rect 16574 19156 16580 19168
rect 15979 19128 16580 19156
rect 15979 19125 15991 19128
rect 15933 19119 15991 19125
rect 16574 19116 16580 19128
rect 16632 19116 16638 19168
rect 17681 19159 17739 19165
rect 17681 19125 17693 19159
rect 17727 19156 17739 19159
rect 17954 19156 17960 19168
rect 17727 19128 17960 19156
rect 17727 19125 17739 19128
rect 17681 19119 17739 19125
rect 17954 19116 17960 19128
rect 18012 19116 18018 19168
rect 18156 19165 18184 19196
rect 19702 19184 19708 19196
rect 19760 19184 19766 19236
rect 19978 19224 19984 19236
rect 19939 19196 19984 19224
rect 19978 19184 19984 19196
rect 20036 19184 20042 19236
rect 21358 19224 21364 19236
rect 21319 19196 21364 19224
rect 21358 19184 21364 19196
rect 21416 19184 21422 19236
rect 18141 19159 18199 19165
rect 18141 19125 18153 19159
rect 18187 19125 18199 19159
rect 18141 19119 18199 19125
rect 19061 19159 19119 19165
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19334 19156 19340 19168
rect 19107 19128 19340 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 19521 19159 19579 19165
rect 19521 19125 19533 19159
rect 19567 19156 19579 19159
rect 21082 19156 21088 19168
rect 19567 19128 21088 19156
rect 19567 19125 19579 19128
rect 19521 19119 19579 19125
rect 21082 19116 21088 19128
rect 21140 19116 21146 19168
rect 1104 19066 21896 19088
rect 1104 19014 7912 19066
rect 7964 19014 7976 19066
rect 8028 19014 8040 19066
rect 8092 19014 8104 19066
rect 8156 19014 14843 19066
rect 14895 19014 14907 19066
rect 14959 19014 14971 19066
rect 15023 19014 15035 19066
rect 15087 19014 21896 19066
rect 1104 18992 21896 19014
rect 5810 18912 5816 18964
rect 5868 18952 5874 18964
rect 5997 18955 6055 18961
rect 5997 18952 6009 18955
rect 5868 18924 6009 18952
rect 5868 18912 5874 18924
rect 5997 18921 6009 18924
rect 6043 18921 6055 18955
rect 5997 18915 6055 18921
rect 7006 18912 7012 18964
rect 7064 18952 7070 18964
rect 7285 18955 7343 18961
rect 7285 18952 7297 18955
rect 7064 18924 7297 18952
rect 7064 18912 7070 18924
rect 7285 18921 7297 18924
rect 7331 18921 7343 18955
rect 7466 18952 7472 18964
rect 7285 18915 7343 18921
rect 7392 18924 7472 18952
rect 4985 18887 5043 18893
rect 4985 18853 4997 18887
rect 5031 18884 5043 18887
rect 6178 18884 6184 18896
rect 5031 18856 6184 18884
rect 5031 18853 5043 18856
rect 4985 18847 5043 18853
rect 6178 18844 6184 18856
rect 6236 18844 6242 18896
rect 6917 18887 6975 18893
rect 6917 18853 6929 18887
rect 6963 18884 6975 18887
rect 7392 18884 7420 18924
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 8297 18955 8355 18961
rect 8297 18921 8309 18955
rect 8343 18952 8355 18955
rect 10686 18952 10692 18964
rect 8343 18924 9674 18952
rect 10647 18924 10692 18952
rect 8343 18921 8355 18924
rect 8297 18915 8355 18921
rect 6963 18856 7420 18884
rect 7576 18856 8688 18884
rect 6963 18853 6975 18856
rect 6917 18847 6975 18853
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6144 18788 6500 18816
rect 6144 18776 6150 18788
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 6270 18748 6276 18760
rect 5767 18720 6276 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 6270 18708 6276 18720
rect 6328 18708 6334 18760
rect 6472 18757 6500 18788
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18748 6515 18751
rect 7576 18748 7604 18856
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18785 7711 18819
rect 7653 18779 7711 18785
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 6503 18720 7604 18748
rect 6503 18717 6515 18720
rect 6457 18711 6515 18717
rect 4617 18683 4675 18689
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 5258 18680 5264 18692
rect 4663 18652 5264 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 5353 18683 5411 18689
rect 5353 18649 5365 18683
rect 5399 18680 5411 18683
rect 5399 18652 6040 18680
rect 5399 18649 5411 18652
rect 5353 18643 5411 18649
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 5534 18612 5540 18624
rect 4295 18584 5540 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 5534 18572 5540 18584
rect 5592 18572 5598 18624
rect 6012 18612 6040 18652
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 7668 18680 7696 18779
rect 7926 18708 7932 18760
rect 7984 18748 7990 18760
rect 8128 18748 8156 18779
rect 8478 18776 8484 18828
rect 8536 18816 8542 18828
rect 8573 18819 8631 18825
rect 8573 18816 8585 18819
rect 8536 18788 8585 18816
rect 8536 18776 8542 18788
rect 8573 18785 8585 18788
rect 8619 18785 8631 18819
rect 8660 18816 8688 18856
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 9554 18887 9612 18893
rect 9554 18884 9566 18887
rect 9364 18856 9566 18884
rect 9364 18844 9370 18856
rect 9554 18853 9566 18856
rect 9600 18853 9612 18887
rect 9646 18884 9674 18924
rect 10686 18912 10692 18924
rect 10744 18912 10750 18964
rect 11238 18952 11244 18964
rect 11199 18924 11244 18952
rect 11238 18912 11244 18924
rect 11296 18912 11302 18964
rect 11701 18955 11759 18961
rect 11701 18921 11713 18955
rect 11747 18952 11759 18955
rect 11793 18955 11851 18961
rect 11793 18952 11805 18955
rect 11747 18924 11805 18952
rect 11747 18921 11759 18924
rect 11701 18915 11759 18921
rect 11793 18921 11805 18924
rect 11839 18921 11851 18955
rect 11793 18915 11851 18921
rect 12250 18912 12256 18964
rect 12308 18952 12314 18964
rect 12437 18955 12495 18961
rect 12437 18952 12449 18955
rect 12308 18924 12449 18952
rect 12308 18912 12314 18924
rect 12437 18921 12449 18924
rect 12483 18921 12495 18955
rect 12437 18915 12495 18921
rect 12802 18912 12808 18964
rect 12860 18952 12866 18964
rect 13449 18955 13507 18961
rect 13449 18952 13461 18955
rect 12860 18924 13461 18952
rect 12860 18912 12866 18924
rect 13449 18921 13461 18924
rect 13495 18921 13507 18955
rect 13449 18915 13507 18921
rect 13538 18912 13544 18964
rect 13596 18952 13602 18964
rect 13909 18955 13967 18961
rect 13909 18952 13921 18955
rect 13596 18924 13921 18952
rect 13596 18912 13602 18924
rect 13909 18921 13921 18924
rect 13955 18921 13967 18955
rect 13909 18915 13967 18921
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 16574 18952 16580 18964
rect 14240 18924 14688 18952
rect 16535 18924 16580 18952
rect 14240 18912 14246 18924
rect 13998 18884 14004 18896
rect 9646 18856 14004 18884
rect 9554 18847 9612 18853
rect 13998 18844 14004 18856
rect 14056 18844 14062 18896
rect 14660 18884 14688 18924
rect 16574 18912 16580 18924
rect 16632 18912 16638 18964
rect 16666 18912 16672 18964
rect 16724 18952 16730 18964
rect 17497 18955 17555 18961
rect 17497 18952 17509 18955
rect 16724 18924 17509 18952
rect 16724 18912 16730 18924
rect 17497 18921 17509 18924
rect 17543 18921 17555 18955
rect 17678 18952 17684 18964
rect 17639 18924 17684 18952
rect 17497 18915 17555 18921
rect 17678 18912 17684 18924
rect 17736 18912 17742 18964
rect 19242 18912 19248 18964
rect 19300 18952 19306 18964
rect 19705 18955 19763 18961
rect 19705 18952 19717 18955
rect 19300 18924 19717 18952
rect 19300 18912 19306 18924
rect 19705 18921 19717 18924
rect 19751 18921 19763 18955
rect 19705 18915 19763 18921
rect 20165 18955 20223 18961
rect 20165 18921 20177 18955
rect 20211 18952 20223 18955
rect 22646 18952 22652 18964
rect 20211 18924 22652 18952
rect 20211 18921 20223 18924
rect 20165 18915 20223 18921
rect 22646 18912 22652 18924
rect 22704 18912 22710 18964
rect 14798 18887 14856 18893
rect 14798 18884 14810 18887
rect 14660 18856 14810 18884
rect 14798 18853 14810 18856
rect 14844 18853 14856 18887
rect 15378 18884 15384 18896
rect 14798 18847 14856 18853
rect 15120 18856 15384 18884
rect 11238 18816 11244 18828
rect 8660 18788 11244 18816
rect 8573 18779 8631 18785
rect 11238 18776 11244 18788
rect 11296 18776 11302 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 11793 18819 11851 18825
rect 11388 18788 11433 18816
rect 11388 18776 11394 18788
rect 11793 18785 11805 18819
rect 11839 18816 11851 18819
rect 12066 18816 12072 18828
rect 11839 18788 12072 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 12345 18819 12403 18825
rect 12345 18785 12357 18819
rect 12391 18816 12403 18819
rect 12989 18819 13047 18825
rect 12989 18816 13001 18819
rect 12391 18788 13001 18816
rect 12391 18785 12403 18788
rect 12345 18779 12403 18785
rect 12989 18785 13001 18788
rect 13035 18785 13047 18819
rect 12989 18779 13047 18785
rect 13446 18776 13452 18828
rect 13504 18816 13510 18828
rect 13633 18819 13691 18825
rect 13633 18816 13645 18819
rect 13504 18788 13645 18816
rect 13504 18776 13510 18788
rect 13633 18785 13645 18788
rect 13679 18785 13691 18819
rect 13633 18779 13691 18785
rect 14553 18819 14611 18825
rect 14553 18785 14565 18819
rect 14599 18816 14611 18819
rect 15120 18816 15148 18856
rect 15378 18844 15384 18856
rect 15436 18844 15442 18896
rect 20438 18844 20444 18896
rect 20496 18884 20502 18896
rect 20625 18887 20683 18893
rect 20625 18884 20637 18887
rect 20496 18856 20637 18884
rect 20496 18844 20502 18856
rect 20625 18853 20637 18856
rect 20671 18853 20683 18887
rect 20625 18847 20683 18853
rect 20809 18887 20867 18893
rect 20809 18853 20821 18887
rect 20855 18884 20867 18887
rect 20990 18884 20996 18896
rect 20855 18856 20996 18884
rect 20855 18853 20867 18856
rect 20809 18847 20867 18853
rect 20990 18844 20996 18856
rect 21048 18844 21054 18896
rect 14599 18788 15148 18816
rect 14599 18785 14611 18788
rect 14553 18779 14611 18785
rect 15194 18776 15200 18828
rect 15252 18816 15258 18828
rect 15252 18788 17264 18816
rect 15252 18776 15258 18788
rect 7984 18720 8156 18748
rect 7984 18708 7990 18720
rect 9214 18708 9220 18760
rect 9272 18748 9278 18760
rect 9309 18751 9367 18757
rect 9309 18748 9321 18751
rect 9272 18720 9321 18748
rect 9272 18708 9278 18720
rect 9309 18717 9321 18720
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 11054 18708 11060 18760
rect 11112 18748 11118 18760
rect 11149 18751 11207 18757
rect 11149 18748 11161 18751
rect 11112 18720 11161 18748
rect 11112 18708 11118 18720
rect 11149 18717 11161 18720
rect 11195 18748 11207 18751
rect 11422 18748 11428 18760
rect 11195 18720 11428 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 11422 18708 11428 18720
rect 11480 18748 11486 18760
rect 12529 18751 12587 18757
rect 11480 18720 12296 18748
rect 11480 18708 11486 18720
rect 7834 18680 7840 18692
rect 7524 18652 7696 18680
rect 7795 18652 7840 18680
rect 7524 18640 7530 18652
rect 7834 18640 7840 18652
rect 7892 18640 7898 18692
rect 12268 18680 12296 18720
rect 12529 18717 12541 18751
rect 12575 18717 12587 18751
rect 12529 18711 12587 18717
rect 12544 18680 12572 18711
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 14090 18748 14096 18760
rect 13780 18720 14096 18748
rect 13780 18708 13786 18720
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 16666 18748 16672 18760
rect 16627 18720 16672 18748
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 16761 18751 16819 18757
rect 16761 18717 16773 18751
rect 16807 18717 16819 18751
rect 16761 18711 16819 18717
rect 14274 18680 14280 18692
rect 11624 18652 12112 18680
rect 12268 18652 12572 18680
rect 13924 18652 14280 18680
rect 8570 18612 8576 18624
rect 6012 18584 8576 18612
rect 8570 18572 8576 18584
rect 8628 18572 8634 18624
rect 8757 18615 8815 18621
rect 8757 18581 8769 18615
rect 8803 18612 8815 18615
rect 11624 18612 11652 18652
rect 11974 18612 11980 18624
rect 8803 18584 11652 18612
rect 11935 18584 11980 18612
rect 8803 18581 8815 18584
rect 8757 18575 8815 18581
rect 11974 18572 11980 18584
rect 12032 18572 12038 18624
rect 12084 18612 12112 18652
rect 13924 18612 13952 18652
rect 14274 18640 14280 18652
rect 14332 18640 14338 18692
rect 15930 18680 15936 18692
rect 15843 18652 15936 18680
rect 15930 18640 15936 18652
rect 15988 18680 15994 18692
rect 16776 18680 16804 18711
rect 17236 18689 17264 18788
rect 17310 18776 17316 18828
rect 17368 18816 17374 18828
rect 17405 18819 17463 18825
rect 17405 18816 17417 18819
rect 17368 18788 17417 18816
rect 17368 18776 17374 18788
rect 17405 18785 17417 18788
rect 17451 18785 17463 18819
rect 17405 18779 17463 18785
rect 17497 18819 17555 18825
rect 17497 18785 17509 18819
rect 17543 18816 17555 18819
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 17543 18788 17877 18816
rect 17543 18785 17555 18788
rect 17497 18779 17555 18785
rect 17865 18785 17877 18788
rect 17911 18785 17923 18819
rect 17865 18779 17923 18785
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18141 18819 18199 18825
rect 18141 18816 18153 18819
rect 18104 18788 18153 18816
rect 18104 18776 18110 18788
rect 18141 18785 18153 18788
rect 18187 18785 18199 18819
rect 18141 18779 18199 18785
rect 18601 18819 18659 18825
rect 18601 18785 18613 18819
rect 18647 18785 18659 18819
rect 18601 18779 18659 18785
rect 19061 18819 19119 18825
rect 19061 18785 19073 18819
rect 19107 18785 19119 18819
rect 20070 18816 20076 18828
rect 20031 18788 20076 18816
rect 19061 18779 19119 18785
rect 17954 18708 17960 18760
rect 18012 18748 18018 18760
rect 18616 18748 18644 18779
rect 19076 18748 19104 18779
rect 20070 18776 20076 18788
rect 20128 18776 20134 18828
rect 20254 18776 20260 18828
rect 20312 18816 20318 18828
rect 21177 18819 21235 18825
rect 21177 18816 21189 18819
rect 20312 18788 21189 18816
rect 20312 18776 20318 18788
rect 21177 18785 21189 18788
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 18012 18720 18644 18748
rect 18708 18720 19104 18748
rect 18012 18708 18018 18720
rect 15988 18652 16804 18680
rect 17221 18683 17279 18689
rect 15988 18640 15994 18652
rect 17221 18649 17233 18683
rect 17267 18649 17279 18683
rect 18708 18680 18736 18720
rect 17221 18643 17279 18649
rect 17328 18652 18736 18680
rect 18785 18683 18843 18689
rect 12084 18584 13952 18612
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 16209 18615 16267 18621
rect 16209 18612 16221 18615
rect 14056 18584 16221 18612
rect 14056 18572 14062 18584
rect 16209 18581 16221 18584
rect 16255 18581 16267 18615
rect 16209 18575 16267 18581
rect 16298 18572 16304 18624
rect 16356 18612 16362 18624
rect 17328 18612 17356 18652
rect 18785 18649 18797 18683
rect 18831 18680 18843 18683
rect 20622 18680 20628 18692
rect 18831 18652 20628 18680
rect 18831 18649 18843 18652
rect 18785 18643 18843 18649
rect 20622 18640 20628 18652
rect 20680 18640 20686 18692
rect 21358 18680 21364 18692
rect 21319 18652 21364 18680
rect 21358 18640 21364 18652
rect 21416 18640 21422 18692
rect 16356 18584 17356 18612
rect 18325 18615 18383 18621
rect 16356 18572 16362 18584
rect 18325 18581 18337 18615
rect 18371 18612 18383 18615
rect 19150 18612 19156 18624
rect 18371 18584 19156 18612
rect 18371 18581 18383 18584
rect 18325 18575 18383 18581
rect 19150 18572 19156 18584
rect 19208 18572 19214 18624
rect 19245 18615 19303 18621
rect 19245 18581 19257 18615
rect 19291 18612 19303 18615
rect 19518 18612 19524 18624
rect 19291 18584 19524 18612
rect 19291 18581 19303 18584
rect 19245 18575 19303 18581
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 1104 18522 21896 18544
rect 1104 18470 4447 18522
rect 4499 18470 4511 18522
rect 4563 18470 4575 18522
rect 4627 18470 4639 18522
rect 4691 18470 11378 18522
rect 11430 18470 11442 18522
rect 11494 18470 11506 18522
rect 11558 18470 11570 18522
rect 11622 18470 18308 18522
rect 18360 18470 18372 18522
rect 18424 18470 18436 18522
rect 18488 18470 18500 18522
rect 18552 18470 21896 18522
rect 1104 18448 21896 18470
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 7466 18408 7472 18420
rect 6687 18380 7472 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 7466 18368 7472 18380
rect 7524 18408 7530 18420
rect 7834 18408 7840 18420
rect 7524 18380 7840 18408
rect 7524 18368 7530 18380
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 8018 18368 8024 18420
rect 8076 18408 8082 18420
rect 13538 18408 13544 18420
rect 8076 18380 13544 18408
rect 8076 18368 8082 18380
rect 13538 18368 13544 18380
rect 13596 18368 13602 18420
rect 14829 18411 14887 18417
rect 14829 18377 14841 18411
rect 14875 18408 14887 18411
rect 16666 18408 16672 18420
rect 14875 18380 16672 18408
rect 14875 18377 14887 18380
rect 14829 18371 14887 18377
rect 16666 18368 16672 18380
rect 16724 18368 16730 18420
rect 17589 18411 17647 18417
rect 17589 18377 17601 18411
rect 17635 18408 17647 18411
rect 20254 18408 20260 18420
rect 17635 18380 20260 18408
rect 17635 18377 17647 18380
rect 17589 18371 17647 18377
rect 20254 18368 20260 18380
rect 20312 18368 20318 18420
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7558 18340 7564 18352
rect 7064 18312 7564 18340
rect 7064 18300 7070 18312
rect 7558 18300 7564 18312
rect 7616 18300 7622 18352
rect 9033 18343 9091 18349
rect 9033 18309 9045 18343
rect 9079 18340 9091 18343
rect 9674 18340 9680 18352
rect 9079 18312 9680 18340
rect 9079 18309 9091 18312
rect 9033 18303 9091 18309
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 10870 18340 10876 18352
rect 10831 18312 10876 18340
rect 10870 18300 10876 18312
rect 10928 18300 10934 18352
rect 12158 18300 12164 18352
rect 12216 18340 12222 18352
rect 15194 18340 15200 18352
rect 12216 18312 12480 18340
rect 12216 18300 12222 18312
rect 5353 18275 5411 18281
rect 5353 18241 5365 18275
rect 5399 18272 5411 18275
rect 6730 18272 6736 18284
rect 5399 18244 6736 18272
rect 5399 18241 5411 18244
rect 5353 18235 5411 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7374 18232 7380 18284
rect 7432 18272 7438 18284
rect 7432 18244 7788 18272
rect 7432 18232 7438 18244
rect 7653 18207 7711 18213
rect 7653 18173 7665 18207
rect 7699 18173 7711 18207
rect 7760 18204 7788 18244
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9953 18275 10011 18281
rect 9953 18272 9965 18275
rect 9364 18244 9965 18272
rect 9364 18232 9370 18244
rect 9953 18241 9965 18244
rect 9999 18241 10011 18275
rect 11882 18272 11888 18284
rect 9953 18235 10011 18241
rect 10060 18244 11888 18272
rect 10060 18204 10088 18244
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12066 18232 12072 18284
rect 12124 18272 12130 18284
rect 12452 18281 12480 18312
rect 13280 18312 15200 18340
rect 12345 18275 12403 18281
rect 12345 18272 12357 18275
rect 12124 18244 12357 18272
rect 12124 18232 12130 18244
rect 12345 18241 12357 18244
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 12437 18275 12495 18281
rect 12437 18241 12449 18275
rect 12483 18241 12495 18275
rect 12437 18235 12495 18241
rect 7760 18176 10088 18204
rect 7653 18167 7711 18173
rect 4985 18139 5043 18145
rect 4985 18105 4997 18139
rect 5031 18136 5043 18139
rect 5442 18136 5448 18148
rect 5031 18108 5448 18136
rect 5031 18105 5043 18108
rect 4985 18099 5043 18105
rect 5442 18096 5448 18108
rect 5500 18096 5506 18148
rect 6822 18136 6828 18148
rect 5644 18108 6828 18136
rect 5644 18080 5672 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 5626 18068 5632 18080
rect 5587 18040 5632 18068
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 6089 18071 6147 18077
rect 6089 18037 6101 18071
rect 6135 18068 6147 18071
rect 6362 18068 6368 18080
rect 6135 18040 6368 18068
rect 6135 18037 6147 18040
rect 6089 18031 6147 18037
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 7009 18071 7067 18077
rect 7009 18037 7021 18071
rect 7055 18068 7067 18071
rect 7098 18068 7104 18080
rect 7055 18040 7104 18068
rect 7055 18037 7067 18040
rect 7009 18031 7067 18037
rect 7098 18028 7104 18040
rect 7156 18028 7162 18080
rect 7377 18071 7435 18077
rect 7377 18037 7389 18071
rect 7423 18068 7435 18071
rect 7466 18068 7472 18080
rect 7423 18040 7472 18068
rect 7423 18037 7435 18040
rect 7377 18031 7435 18037
rect 7466 18028 7472 18040
rect 7524 18028 7530 18080
rect 7668 18068 7696 18167
rect 10134 18164 10140 18216
rect 10192 18204 10198 18216
rect 10689 18207 10747 18213
rect 10689 18204 10701 18207
rect 10192 18176 10701 18204
rect 10192 18164 10198 18176
rect 10689 18173 10701 18176
rect 10735 18173 10747 18207
rect 11146 18204 11152 18216
rect 11107 18176 11152 18204
rect 10689 18167 10747 18173
rect 11146 18164 11152 18176
rect 11204 18164 11210 18216
rect 13280 18204 13308 18312
rect 15194 18300 15200 18312
rect 15252 18300 15258 18352
rect 17773 18343 17831 18349
rect 17773 18340 17785 18343
rect 17052 18312 17785 18340
rect 13722 18272 13728 18284
rect 13683 18244 13728 18272
rect 13722 18232 13728 18244
rect 13780 18232 13786 18284
rect 14182 18272 14188 18284
rect 14143 18244 14188 18272
rect 14182 18232 14188 18244
rect 14240 18232 14246 18284
rect 14366 18272 14372 18284
rect 14327 18244 14372 18272
rect 14366 18232 14372 18244
rect 14424 18232 14430 18284
rect 11348 18176 13308 18204
rect 13541 18207 13599 18213
rect 7920 18139 7978 18145
rect 7920 18105 7932 18139
rect 7966 18136 7978 18139
rect 8846 18136 8852 18148
rect 7966 18108 8852 18136
rect 7966 18105 7978 18108
rect 7920 18099 7978 18105
rect 8846 18096 8852 18108
rect 8904 18096 8910 18148
rect 9214 18096 9220 18148
rect 9272 18136 9278 18148
rect 11238 18136 11244 18148
rect 9272 18108 11244 18136
rect 9272 18096 9278 18108
rect 11238 18096 11244 18108
rect 11296 18096 11302 18148
rect 8294 18068 8300 18080
rect 7668 18040 8300 18068
rect 8294 18028 8300 18040
rect 8352 18068 8358 18080
rect 9122 18068 9128 18080
rect 8352 18040 9128 18068
rect 8352 18028 8358 18040
rect 9122 18028 9128 18040
rect 9180 18028 9186 18080
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9490 18068 9496 18080
rect 9447 18040 9496 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 9766 18068 9772 18080
rect 9727 18040 9772 18068
rect 9766 18028 9772 18040
rect 9824 18028 9830 18080
rect 9858 18028 9864 18080
rect 9916 18068 9922 18080
rect 11348 18077 11376 18176
rect 13541 18173 13553 18207
rect 13587 18204 13599 18207
rect 15197 18207 15255 18213
rect 13587 18176 15148 18204
rect 13587 18173 13599 18176
rect 13541 18167 13599 18173
rect 13449 18139 13507 18145
rect 13449 18105 13461 18139
rect 13495 18136 13507 18139
rect 14734 18136 14740 18148
rect 13495 18108 14740 18136
rect 13495 18105 13507 18108
rect 13449 18099 13507 18105
rect 14734 18096 14740 18108
rect 14792 18096 14798 18148
rect 15120 18136 15148 18176
rect 15197 18173 15209 18207
rect 15243 18204 15255 18207
rect 15286 18204 15292 18216
rect 15243 18176 15292 18204
rect 15243 18173 15255 18176
rect 15197 18167 15255 18173
rect 15286 18164 15292 18176
rect 15344 18164 15350 18216
rect 15464 18207 15522 18213
rect 15464 18173 15476 18207
rect 15510 18204 15522 18207
rect 15930 18204 15936 18216
rect 15510 18176 15936 18204
rect 15510 18173 15522 18176
rect 15464 18167 15522 18173
rect 15930 18164 15936 18176
rect 15988 18164 15994 18216
rect 16022 18164 16028 18216
rect 16080 18204 16086 18216
rect 17052 18213 17080 18312
rect 17773 18309 17785 18312
rect 17819 18309 17831 18343
rect 17773 18303 17831 18309
rect 18892 18312 19840 18340
rect 17218 18232 17224 18284
rect 17276 18272 17282 18284
rect 17865 18275 17923 18281
rect 17865 18272 17877 18275
rect 17276 18244 17877 18272
rect 17276 18232 17282 18244
rect 17865 18241 17877 18244
rect 17911 18241 17923 18275
rect 17865 18235 17923 18241
rect 17037 18207 17095 18213
rect 17037 18204 17049 18207
rect 16080 18176 17049 18204
rect 16080 18164 16086 18176
rect 17037 18173 17049 18176
rect 17083 18173 17095 18207
rect 17402 18204 17408 18216
rect 17363 18176 17408 18204
rect 17037 18167 17095 18173
rect 17402 18164 17408 18176
rect 17460 18164 17466 18216
rect 17773 18207 17831 18213
rect 17773 18173 17785 18207
rect 17819 18204 17831 18207
rect 18892 18204 18920 18312
rect 19812 18281 19840 18312
rect 19613 18275 19671 18281
rect 19613 18272 19625 18275
rect 17819 18176 18920 18204
rect 18984 18244 19625 18272
rect 17819 18173 17831 18176
rect 17773 18167 17831 18173
rect 18984 18148 19012 18244
rect 19613 18241 19625 18244
rect 19659 18241 19671 18275
rect 19613 18235 19671 18241
rect 19797 18275 19855 18281
rect 19797 18241 19809 18275
rect 19843 18241 19855 18275
rect 19797 18235 19855 18241
rect 20622 18204 20628 18216
rect 20583 18176 20628 18204
rect 20622 18164 20628 18176
rect 20680 18164 20686 18216
rect 15746 18136 15752 18148
rect 15120 18108 15752 18136
rect 15746 18096 15752 18108
rect 15804 18096 15810 18148
rect 18132 18139 18190 18145
rect 18132 18105 18144 18139
rect 18178 18136 18190 18139
rect 18966 18136 18972 18148
rect 18178 18108 18972 18136
rect 18178 18105 18190 18108
rect 18132 18099 18190 18105
rect 18966 18096 18972 18108
rect 19024 18096 19030 18148
rect 19150 18096 19156 18148
rect 19208 18136 19214 18148
rect 21177 18139 21235 18145
rect 21177 18136 21189 18139
rect 19208 18108 21189 18136
rect 19208 18096 19214 18108
rect 21177 18105 21189 18108
rect 21223 18105 21235 18139
rect 21358 18136 21364 18148
rect 21319 18108 21364 18136
rect 21177 18099 21235 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 11333 18071 11391 18077
rect 9916 18040 9961 18068
rect 9916 18028 9922 18040
rect 11333 18037 11345 18071
rect 11379 18037 11391 18071
rect 11882 18068 11888 18080
rect 11843 18040 11888 18068
rect 11333 18031 11391 18037
rect 11882 18028 11888 18040
rect 11940 18028 11946 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12253 18071 12311 18077
rect 12253 18068 12265 18071
rect 12032 18040 12265 18068
rect 12032 18028 12038 18040
rect 12253 18037 12265 18040
rect 12299 18037 12311 18071
rect 12253 18031 12311 18037
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 12894 18068 12900 18080
rect 12492 18040 12900 18068
rect 12492 18028 12498 18040
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13078 18068 13084 18080
rect 13039 18040 13084 18068
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 14458 18028 14464 18080
rect 14516 18068 14522 18080
rect 16574 18068 16580 18080
rect 14516 18040 14561 18068
rect 16535 18040 16580 18068
rect 14516 18028 14522 18040
rect 16574 18028 16580 18040
rect 16632 18028 16638 18080
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 19245 18071 19303 18077
rect 19245 18068 19257 18071
rect 18932 18040 19257 18068
rect 18932 18028 18938 18040
rect 19245 18037 19257 18040
rect 19291 18037 19303 18071
rect 19886 18068 19892 18080
rect 19847 18040 19892 18068
rect 19245 18031 19303 18037
rect 19886 18028 19892 18040
rect 19944 18028 19950 18080
rect 20254 18068 20260 18080
rect 20215 18040 20260 18068
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20622 18028 20628 18080
rect 20680 18068 20686 18080
rect 20717 18071 20775 18077
rect 20717 18068 20729 18071
rect 20680 18040 20729 18068
rect 20680 18028 20686 18040
rect 20717 18037 20729 18040
rect 20763 18037 20775 18071
rect 20717 18031 20775 18037
rect 1104 17978 21896 18000
rect 1104 17926 7912 17978
rect 7964 17926 7976 17978
rect 8028 17926 8040 17978
rect 8092 17926 8104 17978
rect 8156 17926 14843 17978
rect 14895 17926 14907 17978
rect 14959 17926 14971 17978
rect 15023 17926 15035 17978
rect 15087 17926 21896 17978
rect 1104 17904 21896 17926
rect 4890 17824 4896 17876
rect 4948 17864 4954 17876
rect 5997 17867 6055 17873
rect 5997 17864 6009 17867
rect 4948 17836 6009 17864
rect 4948 17824 4954 17836
rect 5997 17833 6009 17836
rect 6043 17864 6055 17867
rect 6638 17864 6644 17876
rect 6043 17836 6644 17864
rect 6043 17833 6055 17836
rect 5997 17827 6055 17833
rect 6638 17824 6644 17836
rect 6696 17824 6702 17876
rect 6825 17867 6883 17873
rect 6825 17833 6837 17867
rect 6871 17864 6883 17867
rect 7006 17864 7012 17876
rect 6871 17836 7012 17864
rect 6871 17833 6883 17836
rect 6825 17827 6883 17833
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7248 17836 7849 17864
rect 7248 17824 7254 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 8757 17867 8815 17873
rect 8757 17833 8769 17867
rect 8803 17864 8815 17867
rect 9122 17864 9128 17876
rect 8803 17836 9128 17864
rect 8803 17833 8815 17836
rect 8757 17827 8815 17833
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 9306 17864 9312 17876
rect 9267 17836 9312 17864
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 12345 17867 12403 17873
rect 12345 17833 12357 17867
rect 12391 17864 12403 17867
rect 13078 17864 13084 17876
rect 12391 17836 13084 17864
rect 12391 17833 12403 17836
rect 12345 17827 12403 17833
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 13170 17824 13176 17876
rect 13228 17864 13234 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 13228 17836 13277 17864
rect 13228 17824 13234 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13265 17827 13323 17833
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 15013 17867 15071 17873
rect 15013 17864 15025 17867
rect 13771 17836 15025 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 15013 17833 15025 17836
rect 15059 17833 15071 17867
rect 17494 17864 17500 17876
rect 15013 17827 15071 17833
rect 15120 17836 17500 17864
rect 6086 17756 6092 17808
rect 6144 17796 6150 17808
rect 6144 17768 7972 17796
rect 6144 17756 6150 17768
rect 6638 17688 6644 17740
rect 6696 17728 6702 17740
rect 6696 17700 7880 17728
rect 6696 17688 6702 17700
rect 6457 17663 6515 17669
rect 6457 17629 6469 17663
rect 6503 17660 6515 17663
rect 7374 17660 7380 17672
rect 6503 17632 7380 17660
rect 6503 17629 6515 17632
rect 6457 17623 6515 17629
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 7558 17660 7564 17672
rect 7519 17632 7564 17660
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17629 7803 17663
rect 7745 17623 7803 17629
rect 7760 17592 7788 17623
rect 5828 17564 7788 17592
rect 7852 17592 7880 17700
rect 7944 17660 7972 17768
rect 8478 17756 8484 17808
rect 8536 17796 8542 17808
rect 10594 17796 10600 17808
rect 8536 17768 10600 17796
rect 8536 17756 8542 17768
rect 10594 17756 10600 17768
rect 10652 17756 10658 17808
rect 12434 17796 12440 17808
rect 11532 17768 12440 17796
rect 8573 17731 8631 17737
rect 8573 17697 8585 17731
rect 8619 17728 8631 17731
rect 8754 17728 8760 17740
rect 8619 17700 8760 17728
rect 8619 17697 8631 17700
rect 8573 17691 8631 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10422 17731 10480 17737
rect 10422 17728 10434 17731
rect 9732 17700 10434 17728
rect 9732 17688 9738 17700
rect 10422 17697 10434 17700
rect 10468 17697 10480 17731
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 10422 17691 10480 17697
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 11532 17737 11560 17768
rect 12434 17756 12440 17768
rect 12492 17756 12498 17808
rect 12526 17756 12532 17808
rect 12584 17796 12590 17808
rect 13357 17799 13415 17805
rect 13357 17796 13369 17799
rect 12584 17768 13369 17796
rect 12584 17756 12590 17768
rect 13357 17765 13369 17768
rect 13403 17765 13415 17799
rect 13357 17759 13415 17765
rect 13630 17756 13636 17808
rect 13688 17796 13694 17808
rect 15120 17796 15148 17836
rect 17494 17824 17500 17836
rect 17552 17824 17558 17876
rect 18966 17864 18972 17876
rect 18927 17836 18972 17864
rect 18966 17824 18972 17836
rect 19024 17824 19030 17876
rect 20165 17867 20223 17873
rect 20165 17833 20177 17867
rect 20211 17864 20223 17867
rect 20254 17864 20260 17876
rect 20211 17836 20260 17864
rect 20211 17833 20223 17836
rect 20165 17827 20223 17833
rect 20254 17824 20260 17836
rect 20312 17824 20318 17876
rect 13688 17768 15148 17796
rect 13688 17756 13694 17768
rect 15194 17756 15200 17808
rect 15252 17796 15258 17808
rect 15565 17799 15623 17805
rect 15565 17796 15577 17799
rect 15252 17768 15577 17796
rect 15252 17756 15258 17768
rect 15565 17765 15577 17768
rect 15611 17765 15623 17799
rect 16482 17796 16488 17808
rect 15565 17759 15623 17765
rect 15948 17768 16488 17796
rect 11517 17731 11575 17737
rect 11517 17697 11529 17731
rect 11563 17697 11575 17731
rect 14550 17728 14556 17740
rect 11517 17691 11575 17697
rect 11716 17700 14556 17728
rect 9582 17660 9588 17672
rect 7944 17632 9588 17660
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17660 10747 17663
rect 10962 17660 10968 17672
rect 10735 17632 10968 17660
rect 10735 17629 10747 17632
rect 10689 17623 10747 17629
rect 10962 17620 10968 17632
rect 11020 17620 11026 17672
rect 7852 17564 8800 17592
rect 5828 17536 5856 17564
rect 5721 17527 5779 17533
rect 5721 17493 5733 17527
rect 5767 17524 5779 17527
rect 5810 17524 5816 17536
rect 5767 17496 5816 17524
rect 5767 17493 5779 17496
rect 5721 17487 5779 17493
rect 5810 17484 5816 17496
rect 5868 17484 5874 17536
rect 7098 17524 7104 17536
rect 7059 17496 7104 17524
rect 7098 17484 7104 17496
rect 7156 17524 7162 17536
rect 7650 17524 7656 17536
rect 7156 17496 7656 17524
rect 7156 17484 7162 17496
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 8205 17527 8263 17533
rect 8205 17493 8217 17527
rect 8251 17524 8263 17527
rect 8662 17524 8668 17536
rect 8251 17496 8668 17524
rect 8251 17493 8263 17496
rect 8205 17487 8263 17493
rect 8662 17484 8668 17496
rect 8720 17484 8726 17536
rect 8772 17524 8800 17564
rect 11146 17552 11152 17604
rect 11204 17592 11210 17604
rect 11716 17601 11744 17700
rect 14550 17688 14556 17700
rect 14608 17688 14614 17740
rect 14921 17731 14979 17737
rect 14921 17697 14933 17731
rect 14967 17728 14979 17731
rect 15286 17728 15292 17740
rect 14967 17700 15292 17728
rect 14967 17697 14979 17700
rect 14921 17691 14979 17697
rect 15286 17688 15292 17700
rect 15344 17688 15350 17740
rect 12437 17663 12495 17669
rect 12437 17629 12449 17663
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 11701 17595 11759 17601
rect 11204 17564 11652 17592
rect 11204 17552 11210 17564
rect 10962 17524 10968 17536
rect 8772 17496 10968 17524
rect 10962 17484 10968 17496
rect 11020 17484 11026 17536
rect 11238 17524 11244 17536
rect 11199 17496 11244 17524
rect 11238 17484 11244 17496
rect 11296 17484 11302 17536
rect 11624 17524 11652 17564
rect 11701 17561 11713 17595
rect 11747 17561 11759 17595
rect 11974 17592 11980 17604
rect 11935 17564 11980 17592
rect 11701 17555 11759 17561
rect 11974 17552 11980 17564
rect 12032 17552 12038 17604
rect 12452 17592 12480 17623
rect 12526 17620 12532 17672
rect 12584 17660 12590 17672
rect 13173 17663 13231 17669
rect 12584 17632 12629 17660
rect 12584 17620 12590 17632
rect 13173 17629 13185 17663
rect 13219 17660 13231 17663
rect 13538 17660 13544 17672
rect 13219 17632 13544 17660
rect 13219 17629 13231 17632
rect 13173 17623 13231 17629
rect 13538 17620 13544 17632
rect 13596 17620 13602 17672
rect 14090 17620 14096 17672
rect 14148 17660 14154 17672
rect 15105 17663 15163 17669
rect 15105 17660 15117 17663
rect 14148 17632 15117 17660
rect 14148 17620 14154 17632
rect 15105 17629 15117 17632
rect 15151 17629 15163 17663
rect 15105 17623 15163 17629
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 15378 17660 15384 17672
rect 15252 17632 15384 17660
rect 15252 17620 15258 17632
rect 15378 17620 15384 17632
rect 15436 17620 15442 17672
rect 14553 17595 14611 17601
rect 14553 17592 14565 17595
rect 12452 17564 14565 17592
rect 14553 17561 14565 17564
rect 14599 17561 14611 17595
rect 14553 17555 14611 17561
rect 14642 17552 14648 17604
rect 14700 17592 14706 17604
rect 15010 17592 15016 17604
rect 14700 17564 15016 17592
rect 14700 17552 14706 17564
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 15948 17601 15976 17768
rect 16482 17756 16488 17768
rect 16540 17796 16546 17808
rect 17834 17799 17892 17805
rect 17834 17796 17846 17799
rect 16540 17768 17846 17796
rect 16540 17756 16546 17768
rect 17834 17765 17846 17768
rect 17880 17765 17892 17799
rect 17834 17759 17892 17765
rect 16574 17688 16580 17740
rect 16632 17728 16638 17740
rect 17034 17728 17040 17740
rect 17092 17737 17098 17740
rect 16632 17700 17040 17728
rect 16632 17688 16638 17700
rect 17034 17688 17040 17700
rect 17092 17691 17104 17737
rect 17092 17688 17098 17691
rect 17218 17688 17224 17740
rect 17276 17728 17282 17740
rect 17313 17731 17371 17737
rect 17313 17728 17325 17731
rect 17276 17700 17325 17728
rect 17276 17688 17282 17700
rect 17313 17697 17325 17700
rect 17359 17728 17371 17731
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 17359 17700 17601 17728
rect 17359 17697 17371 17700
rect 17313 17691 17371 17697
rect 17589 17697 17601 17700
rect 17635 17728 17647 17731
rect 18138 17728 18144 17740
rect 17635 17700 18144 17728
rect 17635 17697 17647 17700
rect 17589 17691 17647 17697
rect 18138 17688 18144 17700
rect 18196 17688 18202 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 21177 17731 21235 17737
rect 18932 17700 20392 17728
rect 18932 17688 18938 17700
rect 20254 17660 20260 17672
rect 20215 17632 20260 17660
rect 20254 17620 20260 17632
rect 20312 17620 20318 17672
rect 20364 17669 20392 17700
rect 21177 17697 21189 17731
rect 21223 17697 21235 17731
rect 21177 17691 21235 17697
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 15933 17595 15991 17601
rect 15933 17561 15945 17595
rect 15979 17561 15991 17595
rect 21192 17592 21220 17691
rect 21358 17592 21364 17604
rect 15933 17555 15991 17561
rect 18524 17564 21220 17592
rect 21319 17564 21364 17592
rect 12066 17524 12072 17536
rect 11624 17496 12072 17524
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 15470 17524 15476 17536
rect 12676 17496 15476 17524
rect 12676 17484 12682 17496
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 16206 17484 16212 17536
rect 16264 17524 16270 17536
rect 18524 17524 18552 17564
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 19794 17524 19800 17536
rect 16264 17496 18552 17524
rect 19755 17496 19800 17524
rect 16264 17484 16270 17496
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 1104 17434 21896 17456
rect 1104 17382 4447 17434
rect 4499 17382 4511 17434
rect 4563 17382 4575 17434
rect 4627 17382 4639 17434
rect 4691 17382 11378 17434
rect 11430 17382 11442 17434
rect 11494 17382 11506 17434
rect 11558 17382 11570 17434
rect 11622 17382 18308 17434
rect 18360 17382 18372 17434
rect 18424 17382 18436 17434
rect 18488 17382 18500 17434
rect 18552 17382 21896 17434
rect 1104 17360 21896 17382
rect 6086 17320 6092 17332
rect 6047 17292 6092 17320
rect 6086 17280 6092 17292
rect 6144 17280 6150 17332
rect 6638 17320 6644 17332
rect 6599 17292 6644 17320
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7558 17320 7564 17332
rect 6963 17292 7564 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7558 17280 7564 17292
rect 7616 17320 7622 17332
rect 8938 17320 8944 17332
rect 7616 17292 8944 17320
rect 7616 17280 7622 17292
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9217 17323 9275 17329
rect 9217 17289 9229 17323
rect 9263 17320 9275 17323
rect 9263 17292 9720 17320
rect 9263 17289 9275 17292
rect 9217 17283 9275 17289
rect 1578 17252 1584 17264
rect 1539 17224 1584 17252
rect 1578 17212 1584 17224
rect 1636 17212 1642 17264
rect 8662 17212 8668 17264
rect 8720 17252 8726 17264
rect 8720 17224 9628 17252
rect 8720 17212 8726 17224
rect 8294 17184 8300 17196
rect 8255 17156 8300 17184
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 9600 17193 9628 17224
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8772 17156 9137 17184
rect 6086 17116 6092 17128
rect 5736 17088 6092 17116
rect 1765 17051 1823 17057
rect 1765 17017 1777 17051
rect 1811 17048 1823 17051
rect 1811 17020 2268 17048
rect 1811 17017 1823 17020
rect 1765 17011 1823 17017
rect 2240 16992 2268 17020
rect 5736 16992 5764 17088
rect 6086 17076 6092 17088
rect 6144 17116 6150 17128
rect 8772 17116 8800 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9125 17147 9183 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17153 9551 17187
rect 9493 17147 9551 17153
rect 9585 17187 9643 17193
rect 9585 17153 9597 17187
rect 9631 17153 9643 17187
rect 9692 17184 9720 17292
rect 9858 17280 9864 17332
rect 9916 17320 9922 17332
rect 10045 17323 10103 17329
rect 10045 17320 10057 17323
rect 9916 17292 10057 17320
rect 9916 17280 9922 17292
rect 10045 17289 10057 17292
rect 10091 17289 10103 17323
rect 10045 17283 10103 17289
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 12250 17320 12256 17332
rect 10284 17292 12256 17320
rect 10284 17280 10290 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12437 17323 12495 17329
rect 12437 17289 12449 17323
rect 12483 17320 12495 17323
rect 13630 17320 13636 17332
rect 12483 17292 13636 17320
rect 12483 17289 12495 17292
rect 12437 17283 12495 17289
rect 13630 17280 13636 17292
rect 13688 17280 13694 17332
rect 14090 17320 14096 17332
rect 14051 17292 14096 17320
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14550 17320 14556 17332
rect 14507 17292 14556 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 14734 17320 14740 17332
rect 14695 17292 14740 17320
rect 14734 17280 14740 17292
rect 14792 17280 14798 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 16850 17320 16856 17332
rect 15528 17292 16856 17320
rect 15528 17280 15534 17292
rect 16850 17280 16856 17292
rect 16908 17280 16914 17332
rect 20254 17280 20260 17332
rect 20312 17320 20318 17332
rect 20533 17323 20591 17329
rect 20533 17320 20545 17323
rect 20312 17292 20545 17320
rect 20312 17280 20318 17292
rect 20533 17289 20545 17292
rect 20579 17289 20591 17323
rect 20533 17283 20591 17289
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 10321 17255 10379 17261
rect 10321 17252 10333 17255
rect 9824 17224 10333 17252
rect 9824 17212 9830 17224
rect 10321 17221 10333 17224
rect 10367 17221 10379 17255
rect 11146 17252 11152 17264
rect 10321 17215 10379 17221
rect 10520 17224 11152 17252
rect 10520 17184 10548 17224
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 11238 17212 11244 17264
rect 11296 17252 11302 17264
rect 12621 17255 12679 17261
rect 12621 17252 12633 17255
rect 11296 17224 12633 17252
rect 11296 17212 11302 17224
rect 12621 17221 12633 17224
rect 12667 17221 12679 17255
rect 12621 17215 12679 17221
rect 14182 17212 14188 17264
rect 14240 17252 14246 17264
rect 15841 17255 15899 17261
rect 15841 17252 15853 17255
rect 14240 17224 15853 17252
rect 14240 17212 14246 17224
rect 15841 17221 15853 17224
rect 15887 17221 15899 17255
rect 17126 17252 17132 17264
rect 15841 17215 15899 17221
rect 16316 17224 17132 17252
rect 10873 17187 10931 17193
rect 10873 17184 10885 17187
rect 9692 17156 10548 17184
rect 10612 17156 10885 17184
rect 9585 17147 9643 17153
rect 6144 17088 8800 17116
rect 8849 17119 8907 17125
rect 6144 17076 6150 17088
rect 8849 17085 8861 17119
rect 8895 17116 8907 17119
rect 9217 17119 9275 17125
rect 9217 17116 9229 17119
rect 8895 17088 9229 17116
rect 8895 17085 8907 17088
rect 8849 17079 8907 17085
rect 9217 17085 9229 17088
rect 9263 17085 9275 17119
rect 9508 17116 9536 17147
rect 9674 17116 9680 17128
rect 9508 17088 9680 17116
rect 9217 17079 9275 17085
rect 9674 17076 9680 17088
rect 9732 17116 9738 17128
rect 10612 17116 10640 17156
rect 10873 17153 10885 17156
rect 10919 17153 10931 17187
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 10873 17147 10931 17153
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 12158 17144 12164 17196
rect 12216 17184 12222 17196
rect 12710 17184 12716 17196
rect 12216 17156 12716 17184
rect 12216 17144 12222 17156
rect 12710 17144 12716 17156
rect 12768 17144 12774 17196
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 14792 17156 15301 17184
rect 14792 17144 14798 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15378 17144 15384 17196
rect 15436 17184 15442 17196
rect 16316 17184 16344 17224
rect 17126 17212 17132 17224
rect 17184 17252 17190 17264
rect 17184 17224 17816 17252
rect 17184 17212 17190 17224
rect 16482 17184 16488 17196
rect 15436 17156 16344 17184
rect 16443 17156 16488 17184
rect 15436 17144 15442 17156
rect 16482 17144 16488 17156
rect 16540 17144 16546 17196
rect 17034 17144 17040 17196
rect 17092 17184 17098 17196
rect 17681 17187 17739 17193
rect 17681 17184 17693 17187
rect 17092 17156 17693 17184
rect 17092 17144 17098 17156
rect 17681 17153 17693 17156
rect 17727 17153 17739 17187
rect 17681 17147 17739 17153
rect 9732 17088 10640 17116
rect 9732 17076 9738 17088
rect 10686 17076 10692 17128
rect 10744 17116 10750 17128
rect 10744 17088 10789 17116
rect 10744 17076 10750 17088
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 12253 17119 12311 17125
rect 12253 17116 12265 17119
rect 11020 17088 12265 17116
rect 11020 17076 11026 17088
rect 12253 17085 12265 17088
rect 12299 17085 12311 17119
rect 12253 17079 12311 17085
rect 12980 17119 13038 17125
rect 12980 17085 12992 17119
rect 13026 17116 13038 17119
rect 13538 17116 13544 17128
rect 13026 17088 13544 17116
rect 13026 17085 13038 17088
rect 12980 17079 13038 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 17402 17116 17408 17128
rect 14936 17088 17408 17116
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 8030 17051 8088 17057
rect 8030 17048 8042 17051
rect 7432 17020 8042 17048
rect 7432 17008 7438 17020
rect 8030 17017 8042 17020
rect 8076 17017 8088 17051
rect 8030 17011 8088 17017
rect 8938 17008 8944 17060
rect 8996 17048 9002 17060
rect 14936 17048 14964 17088
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 17589 17119 17647 17125
rect 17589 17085 17601 17119
rect 17635 17116 17647 17119
rect 17788 17116 17816 17224
rect 18138 17184 18144 17196
rect 18099 17156 18144 17184
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 20070 17184 20076 17196
rect 20031 17156 20076 17184
rect 19889 17147 19947 17153
rect 17635 17088 17816 17116
rect 18408 17119 18466 17125
rect 17635 17085 17647 17088
rect 17589 17079 17647 17085
rect 18408 17085 18420 17119
rect 18454 17116 18466 17119
rect 18874 17116 18880 17128
rect 18454 17088 18880 17116
rect 18454 17085 18466 17088
rect 18408 17079 18466 17085
rect 18874 17076 18880 17088
rect 18932 17076 18938 17128
rect 18966 17076 18972 17128
rect 19024 17116 19030 17128
rect 19904 17116 19932 17147
rect 20070 17144 20076 17156
rect 20128 17144 20134 17196
rect 19024 17088 19932 17116
rect 19024 17076 19030 17088
rect 21082 17076 21088 17128
rect 21140 17116 21146 17128
rect 21177 17119 21235 17125
rect 21177 17116 21189 17119
rect 21140 17088 21189 17116
rect 21140 17076 21146 17088
rect 21177 17085 21189 17088
rect 21223 17085 21235 17119
rect 21177 17079 21235 17085
rect 8996 17020 14964 17048
rect 8996 17008 9002 17020
rect 15010 17008 15016 17060
rect 15068 17048 15074 17060
rect 15197 17051 15255 17057
rect 15197 17048 15209 17051
rect 15068 17020 15209 17048
rect 15068 17008 15074 17020
rect 15197 17017 15209 17020
rect 15243 17017 15255 17051
rect 15562 17048 15568 17060
rect 15197 17011 15255 17017
rect 15304 17020 15568 17048
rect 2222 16980 2228 16992
rect 2183 16952 2228 16980
rect 2222 16940 2228 16952
rect 2280 16940 2286 16992
rect 5350 16980 5356 16992
rect 5311 16952 5356 16980
rect 5350 16940 5356 16952
rect 5408 16940 5414 16992
rect 5718 16980 5724 16992
rect 5679 16952 5724 16980
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 9030 16980 9036 16992
rect 8991 16952 9036 16980
rect 9030 16940 9036 16952
rect 9088 16940 9094 16992
rect 9125 16983 9183 16989
rect 9125 16949 9137 16983
rect 9171 16980 9183 16983
rect 9677 16983 9735 16989
rect 9677 16980 9689 16983
rect 9171 16952 9689 16980
rect 9171 16949 9183 16952
rect 9125 16943 9183 16949
rect 9677 16949 9689 16952
rect 9723 16949 9735 16983
rect 9677 16943 9735 16949
rect 9766 16940 9772 16992
rect 9824 16980 9830 16992
rect 10781 16983 10839 16989
rect 10781 16980 10793 16983
rect 9824 16952 10793 16980
rect 9824 16940 9830 16952
rect 10781 16949 10793 16952
rect 10827 16949 10839 16983
rect 10781 16943 10839 16949
rect 12621 16983 12679 16989
rect 12621 16949 12633 16983
rect 12667 16980 12679 16983
rect 13630 16980 13636 16992
rect 12667 16952 13636 16980
rect 12667 16949 12679 16952
rect 12621 16943 12679 16949
rect 13630 16940 13636 16952
rect 13688 16940 13694 16992
rect 15105 16983 15163 16989
rect 15105 16949 15117 16983
rect 15151 16980 15163 16983
rect 15304 16980 15332 17020
rect 15562 17008 15568 17020
rect 15620 17008 15626 17060
rect 16209 17051 16267 17057
rect 16209 17017 16221 17051
rect 16255 17048 16267 17051
rect 16255 17020 17172 17048
rect 16255 17017 16267 17020
rect 16209 17011 16267 17017
rect 15151 16952 15332 16980
rect 16301 16983 16359 16989
rect 15151 16949 15163 16952
rect 15105 16943 15163 16949
rect 16301 16949 16313 16983
rect 16347 16980 16359 16983
rect 16482 16980 16488 16992
rect 16347 16952 16488 16980
rect 16347 16949 16359 16952
rect 16301 16943 16359 16949
rect 16482 16940 16488 16952
rect 16540 16940 16546 16992
rect 17144 16989 17172 17020
rect 17218 17008 17224 17060
rect 17276 17048 17282 17060
rect 20070 17048 20076 17060
rect 17276 17020 20076 17048
rect 17276 17008 17282 17020
rect 20070 17008 20076 17020
rect 20128 17008 20134 17060
rect 17129 16983 17187 16989
rect 17129 16949 17141 16983
rect 17175 16949 17187 16983
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 17129 16943 17187 16949
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 19426 16940 19432 16992
rect 19484 16980 19490 16992
rect 19521 16983 19579 16989
rect 19521 16980 19533 16983
rect 19484 16952 19533 16980
rect 19484 16940 19490 16952
rect 19521 16949 19533 16952
rect 19567 16949 19579 16983
rect 20162 16980 20168 16992
rect 20123 16952 20168 16980
rect 19521 16943 19579 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 7912 16890
rect 7964 16838 7976 16890
rect 8028 16838 8040 16890
rect 8092 16838 8104 16890
rect 8156 16838 14843 16890
rect 14895 16838 14907 16890
rect 14959 16838 14971 16890
rect 15023 16838 15035 16890
rect 15087 16838 21896 16890
rect 1104 16816 21896 16838
rect 5718 16776 5724 16788
rect 5679 16748 5724 16776
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 6273 16779 6331 16785
rect 6273 16745 6285 16779
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8478 16776 8484 16788
rect 8343 16748 8484 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 6288 16708 6316 16739
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 8757 16779 8815 16785
rect 8757 16745 8769 16779
rect 8803 16776 8815 16779
rect 8938 16776 8944 16788
rect 8803 16748 8944 16776
rect 8803 16745 8815 16748
rect 8757 16739 8815 16745
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 9030 16736 9036 16788
rect 9088 16776 9094 16788
rect 9125 16779 9183 16785
rect 9125 16776 9137 16779
rect 9088 16748 9137 16776
rect 9088 16736 9094 16748
rect 9125 16745 9137 16748
rect 9171 16745 9183 16779
rect 9125 16739 9183 16745
rect 9677 16779 9735 16785
rect 9677 16745 9689 16779
rect 9723 16776 9735 16779
rect 9769 16779 9827 16785
rect 9769 16776 9781 16779
rect 9723 16748 9781 16776
rect 9723 16745 9735 16748
rect 9677 16739 9735 16745
rect 9769 16745 9781 16748
rect 9815 16745 9827 16779
rect 9769 16739 9827 16745
rect 10137 16779 10195 16785
rect 10137 16745 10149 16779
rect 10183 16776 10195 16779
rect 10686 16776 10692 16788
rect 10183 16748 10692 16776
rect 10183 16745 10195 16748
rect 10137 16739 10195 16745
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 13722 16776 13728 16788
rect 11072 16748 13728 16776
rect 10962 16708 10968 16720
rect 6288 16680 10968 16708
rect 10962 16668 10968 16680
rect 11020 16668 11026 16720
rect 5442 16640 5448 16652
rect 5403 16612 5448 16640
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 6089 16643 6147 16649
rect 6089 16609 6101 16643
rect 6135 16640 6147 16643
rect 7282 16640 7288 16652
rect 6135 16612 7288 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 7282 16600 7288 16612
rect 7340 16600 7346 16652
rect 7673 16643 7731 16649
rect 7673 16609 7685 16643
rect 7719 16640 7731 16643
rect 8570 16640 8576 16652
rect 7719 16612 8432 16640
rect 8531 16612 8576 16640
rect 7719 16609 7731 16612
rect 7673 16603 7731 16609
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16572 7987 16575
rect 8294 16572 8300 16584
rect 7975 16544 8300 16572
rect 7975 16541 7987 16544
rect 7929 16535 7987 16541
rect 8294 16532 8300 16544
rect 8352 16532 8358 16584
rect 8404 16572 8432 16612
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 9490 16640 9496 16652
rect 8680 16612 9352 16640
rect 9451 16612 9496 16640
rect 8680 16572 8708 16612
rect 8404 16544 8708 16572
rect 9324 16572 9352 16612
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9769 16643 9827 16649
rect 9769 16609 9781 16643
rect 9815 16640 9827 16643
rect 11072 16640 11100 16748
rect 13722 16736 13728 16748
rect 13780 16736 13786 16788
rect 13817 16779 13875 16785
rect 13817 16745 13829 16779
rect 13863 16776 13875 16779
rect 13906 16776 13912 16788
rect 13863 16748 13912 16776
rect 13863 16745 13875 16748
rect 13817 16739 13875 16745
rect 13906 16736 13912 16748
rect 13964 16736 13970 16788
rect 14274 16736 14280 16788
rect 14332 16776 14338 16788
rect 14461 16779 14519 16785
rect 14461 16776 14473 16779
rect 14332 16748 14473 16776
rect 14332 16736 14338 16748
rect 14461 16745 14473 16748
rect 14507 16776 14519 16779
rect 14921 16779 14979 16785
rect 14921 16776 14933 16779
rect 14507 16748 14933 16776
rect 14507 16745 14519 16748
rect 14461 16739 14519 16745
rect 14921 16745 14933 16748
rect 14967 16745 14979 16779
rect 15286 16776 15292 16788
rect 15247 16748 15292 16776
rect 14921 16739 14979 16745
rect 15286 16736 15292 16748
rect 15344 16736 15350 16788
rect 15562 16776 15568 16788
rect 15523 16748 15568 16776
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 16206 16776 16212 16788
rect 16167 16748 16212 16776
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 16482 16776 16488 16788
rect 16443 16748 16488 16776
rect 16482 16736 16488 16748
rect 16540 16736 16546 16788
rect 16850 16736 16856 16788
rect 16908 16776 16914 16788
rect 16945 16779 17003 16785
rect 16945 16776 16957 16779
rect 16908 16748 16957 16776
rect 16908 16736 16914 16748
rect 16945 16745 16957 16748
rect 16991 16745 17003 16779
rect 17494 16776 17500 16788
rect 17455 16748 17500 16776
rect 16945 16739 17003 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 17678 16736 17684 16788
rect 17736 16776 17742 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 17736 16748 18337 16776
rect 17736 16736 17742 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 18325 16739 18383 16745
rect 19797 16779 19855 16785
rect 19797 16745 19809 16779
rect 19843 16776 19855 16779
rect 19886 16776 19892 16788
rect 19843 16748 19892 16776
rect 19843 16745 19855 16748
rect 19797 16739 19855 16745
rect 19886 16736 19892 16748
rect 19944 16736 19950 16788
rect 11698 16668 11704 16720
rect 11756 16708 11762 16720
rect 11974 16708 11980 16720
rect 11756 16680 11980 16708
rect 11756 16668 11762 16680
rect 11974 16668 11980 16680
rect 12032 16668 12038 16720
rect 12526 16668 12532 16720
rect 12584 16708 12590 16720
rect 17957 16711 18015 16717
rect 17957 16708 17969 16711
rect 12584 16680 17969 16708
rect 12584 16668 12590 16680
rect 17957 16677 17969 16680
rect 18003 16708 18015 16711
rect 18785 16711 18843 16717
rect 18785 16708 18797 16711
rect 18003 16680 18797 16708
rect 18003 16677 18015 16680
rect 17957 16671 18015 16677
rect 18785 16677 18797 16680
rect 18831 16677 18843 16711
rect 18785 16671 18843 16677
rect 19518 16668 19524 16720
rect 19576 16708 19582 16720
rect 21177 16711 21235 16717
rect 21177 16708 21189 16711
rect 19576 16680 21189 16708
rect 19576 16668 19582 16680
rect 21177 16677 21189 16680
rect 21223 16677 21235 16711
rect 21177 16671 21235 16677
rect 9815 16612 11100 16640
rect 9815 16609 9827 16612
rect 9769 16603 9827 16609
rect 11238 16600 11244 16652
rect 11296 16640 11302 16652
rect 11618 16643 11676 16649
rect 11618 16640 11630 16643
rect 11296 16612 11630 16640
rect 11296 16600 11302 16612
rect 11618 16609 11630 16612
rect 11664 16609 11676 16643
rect 11618 16603 11676 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 12158 16640 12164 16652
rect 11931 16612 12164 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 12417 16643 12475 16649
rect 12417 16640 12429 16643
rect 12268 16612 12429 16640
rect 10226 16572 10232 16584
rect 9324 16544 10232 16572
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 12268 16572 12296 16612
rect 12417 16609 12429 16612
rect 12463 16609 12475 16643
rect 12417 16603 12475 16609
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16640 14059 16643
rect 14274 16640 14280 16652
rect 14047 16612 14280 16640
rect 14047 16609 14059 16612
rect 14001 16603 14059 16609
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 14550 16600 14556 16652
rect 14608 16640 14614 16652
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 14608 16612 14841 16640
rect 14608 16600 14614 16612
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 14918 16600 14924 16652
rect 14976 16640 14982 16652
rect 16025 16643 16083 16649
rect 16025 16640 16037 16643
rect 14976 16612 16037 16640
rect 14976 16600 14982 16612
rect 16025 16609 16037 16612
rect 16071 16609 16083 16643
rect 16025 16603 16083 16609
rect 16853 16643 16911 16649
rect 16853 16609 16865 16643
rect 16899 16609 16911 16643
rect 18690 16640 18696 16652
rect 18651 16612 18696 16640
rect 16853 16603 16911 16609
rect 11900 16544 12296 16572
rect 6546 16504 6552 16516
rect 6507 16476 6552 16504
rect 6546 16464 6552 16476
rect 6604 16464 6610 16516
rect 8312 16504 8340 16532
rect 8570 16504 8576 16516
rect 8312 16476 8576 16504
rect 8570 16464 8576 16476
rect 8628 16464 8634 16516
rect 8938 16464 8944 16516
rect 8996 16504 9002 16516
rect 9306 16504 9312 16516
rect 8996 16476 9312 16504
rect 8996 16464 9002 16476
rect 9306 16464 9312 16476
rect 9364 16464 9370 16516
rect 5994 16396 6000 16448
rect 6052 16436 6058 16448
rect 8294 16436 8300 16448
rect 6052 16408 8300 16436
rect 6052 16396 6058 16408
rect 8294 16396 8300 16408
rect 8352 16436 8358 16448
rect 9674 16436 9680 16448
rect 8352 16408 9680 16436
rect 8352 16396 8358 16408
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9766 16396 9772 16448
rect 9824 16436 9830 16448
rect 10505 16439 10563 16445
rect 10505 16436 10517 16439
rect 9824 16408 10517 16436
rect 9824 16396 9830 16408
rect 10505 16405 10517 16408
rect 10551 16436 10563 16439
rect 11900 16436 11928 16544
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 14461 16575 14519 16581
rect 14461 16572 14473 16575
rect 13412 16544 14473 16572
rect 13412 16532 13418 16544
rect 14461 16541 14473 16544
rect 14507 16541 14519 16575
rect 14734 16572 14740 16584
rect 14647 16544 14740 16572
rect 14461 16535 14519 16541
rect 14734 16532 14740 16544
rect 14792 16572 14798 16584
rect 15010 16572 15016 16584
rect 14792 16544 15016 16572
rect 14792 16532 14798 16544
rect 15010 16532 15016 16544
rect 15068 16532 15074 16584
rect 16206 16532 16212 16584
rect 16264 16572 16270 16584
rect 16868 16572 16896 16603
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 20622 16640 20628 16652
rect 20583 16612 20628 16640
rect 20622 16600 20628 16612
rect 20680 16600 20686 16652
rect 21358 16640 21364 16652
rect 21319 16612 21364 16640
rect 21358 16600 21364 16612
rect 21416 16600 21422 16652
rect 16264 16544 16896 16572
rect 16264 16532 16270 16544
rect 17034 16532 17040 16584
rect 17092 16572 17098 16584
rect 18969 16575 19027 16581
rect 17092 16544 17137 16572
rect 17092 16532 17098 16544
rect 18969 16541 18981 16575
rect 19015 16572 19027 16575
rect 19426 16572 19432 16584
rect 19015 16544 19432 16572
rect 19015 16541 19027 16544
rect 18969 16535 19027 16541
rect 19426 16532 19432 16544
rect 19484 16532 19490 16584
rect 13538 16504 13544 16516
rect 13451 16476 13544 16504
rect 13538 16464 13544 16476
rect 13596 16504 13602 16516
rect 14752 16504 14780 16532
rect 13596 16476 14780 16504
rect 13596 16464 13602 16476
rect 15470 16464 15476 16516
rect 15528 16504 15534 16516
rect 16298 16504 16304 16516
rect 15528 16476 16304 16504
rect 15528 16464 15534 16476
rect 16298 16464 16304 16476
rect 16356 16464 16362 16516
rect 10551 16408 11928 16436
rect 10551 16405 10563 16408
rect 10505 16399 10563 16405
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 12434 16436 12440 16448
rect 12124 16408 12440 16436
rect 12124 16396 12130 16408
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 19794 16436 19800 16448
rect 12860 16408 19800 16436
rect 12860 16396 12866 16408
rect 19794 16396 19800 16408
rect 19852 16396 19858 16448
rect 20254 16436 20260 16448
rect 20215 16408 20260 16436
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 20806 16436 20812 16448
rect 20767 16408 20812 16436
rect 20806 16396 20812 16408
rect 20864 16396 20870 16448
rect 1104 16346 21896 16368
rect 1104 16294 4447 16346
rect 4499 16294 4511 16346
rect 4563 16294 4575 16346
rect 4627 16294 4639 16346
rect 4691 16294 11378 16346
rect 11430 16294 11442 16346
rect 11494 16294 11506 16346
rect 11558 16294 11570 16346
rect 11622 16294 18308 16346
rect 18360 16294 18372 16346
rect 18424 16294 18436 16346
rect 18488 16294 18500 16346
rect 18552 16294 21896 16346
rect 1104 16272 21896 16294
rect 5994 16232 6000 16244
rect 5955 16204 6000 16232
rect 5994 16192 6000 16204
rect 6052 16192 6058 16244
rect 7006 16192 7012 16244
rect 7064 16232 7070 16244
rect 8665 16235 8723 16241
rect 8665 16232 8677 16235
rect 7064 16204 8677 16232
rect 7064 16192 7070 16204
rect 8665 16201 8677 16204
rect 8711 16201 8723 16235
rect 8665 16195 8723 16201
rect 10226 16192 10232 16244
rect 10284 16232 10290 16244
rect 12342 16232 12348 16244
rect 10284 16204 12348 16232
rect 10284 16192 10290 16204
rect 12342 16192 12348 16204
rect 12400 16232 12406 16244
rect 13081 16235 13139 16241
rect 13081 16232 13093 16235
rect 12400 16204 13093 16232
rect 12400 16192 12406 16204
rect 13081 16201 13093 16204
rect 13127 16201 13139 16235
rect 15470 16232 15476 16244
rect 13081 16195 13139 16201
rect 13556 16204 15476 16232
rect 11333 16167 11391 16173
rect 11333 16133 11345 16167
rect 11379 16164 11391 16167
rect 13556 16164 13584 16204
rect 15470 16192 15476 16204
rect 15528 16192 15534 16244
rect 15746 16232 15752 16244
rect 15707 16204 15752 16232
rect 15746 16192 15752 16204
rect 15804 16192 15810 16244
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 17126 16232 17132 16244
rect 17083 16204 17132 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 17126 16192 17132 16204
rect 17184 16192 17190 16244
rect 20162 16232 20168 16244
rect 17420 16204 20168 16232
rect 11379 16136 13584 16164
rect 11379 16133 11391 16136
rect 11333 16127 11391 16133
rect 15562 16124 15568 16176
rect 15620 16164 15626 16176
rect 17313 16167 17371 16173
rect 17313 16164 17325 16167
rect 15620 16136 17325 16164
rect 15620 16124 15626 16136
rect 17313 16133 17325 16136
rect 17359 16133 17371 16167
rect 17313 16127 17371 16133
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 8404 16068 9321 16096
rect 5350 16028 5356 16040
rect 5263 16000 5356 16028
rect 5350 15988 5356 16000
rect 5408 16028 5414 16040
rect 6454 16028 6460 16040
rect 5408 16000 6460 16028
rect 5408 15988 5414 16000
rect 6454 15988 6460 16000
rect 6512 15988 6518 16040
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 8214 16031 8272 16037
rect 8214 16028 8226 16031
rect 6604 16000 8226 16028
rect 6604 15988 6610 16000
rect 8214 15997 8226 16000
rect 8260 16028 8272 16031
rect 8404 16028 8432 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 10226 16096 10232 16108
rect 10187 16068 10232 16096
rect 9309 16059 9367 16065
rect 10226 16056 10232 16068
rect 10284 16056 10290 16108
rect 10318 16056 10324 16108
rect 10376 16096 10382 16108
rect 10376 16068 10421 16096
rect 10376 16056 10382 16068
rect 11238 16056 11244 16108
rect 11296 16096 11302 16108
rect 12342 16096 12348 16108
rect 11296 16068 12348 16096
rect 11296 16056 11302 16068
rect 12342 16056 12348 16068
rect 12400 16096 12406 16108
rect 12437 16099 12495 16105
rect 12437 16096 12449 16099
rect 12400 16068 12449 16096
rect 12400 16056 12406 16068
rect 12437 16065 12449 16068
rect 12483 16065 12495 16099
rect 14458 16096 14464 16108
rect 14419 16068 14464 16096
rect 12437 16059 12495 16065
rect 14458 16056 14464 16068
rect 14516 16056 14522 16108
rect 14734 16056 14740 16108
rect 14792 16096 14798 16108
rect 14829 16099 14887 16105
rect 14829 16096 14841 16099
rect 14792 16068 14841 16096
rect 14792 16056 14798 16068
rect 14829 16065 14841 16068
rect 14875 16065 14887 16099
rect 14829 16059 14887 16065
rect 15010 16056 15016 16108
rect 15068 16096 15074 16108
rect 16301 16099 16359 16105
rect 16301 16096 16313 16099
rect 15068 16068 16313 16096
rect 15068 16056 15074 16068
rect 16301 16065 16313 16068
rect 16347 16065 16359 16099
rect 16301 16059 16359 16065
rect 8260 16000 8432 16028
rect 8481 16031 8539 16037
rect 8260 15997 8272 16000
rect 8214 15991 8272 15997
rect 8481 15997 8493 16031
rect 8527 16028 8539 16031
rect 8570 16028 8576 16040
rect 8527 16000 8576 16028
rect 8527 15997 8539 16000
rect 8481 15991 8539 15997
rect 8570 15988 8576 16000
rect 8628 15988 8634 16040
rect 8665 16031 8723 16037
rect 8665 15997 8677 16031
rect 8711 16028 8723 16031
rect 9125 16031 9183 16037
rect 9125 16028 9137 16031
rect 8711 16000 9137 16028
rect 8711 15997 8723 16000
rect 8665 15991 8723 15997
rect 9125 15997 9137 16000
rect 9171 15997 9183 16031
rect 9125 15991 9183 15997
rect 9674 15988 9680 16040
rect 9732 16028 9738 16040
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 9732 16000 10425 16028
rect 9732 15988 9738 16000
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 11149 16031 11207 16037
rect 11149 15997 11161 16031
rect 11195 16028 11207 16031
rect 11882 16028 11888 16040
rect 11195 16000 11888 16028
rect 11195 15997 11207 16000
rect 11149 15991 11207 15997
rect 11882 15988 11888 16000
rect 11940 15988 11946 16040
rect 12158 15988 12164 16040
rect 12216 16028 12222 16040
rect 12216 16000 12480 16028
rect 12216 15988 12222 16000
rect 5718 15960 5724 15972
rect 5679 15932 5724 15960
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 8110 15960 8116 15972
rect 6748 15932 8116 15960
rect 4985 15895 5043 15901
rect 4985 15861 4997 15895
rect 5031 15892 5043 15895
rect 5534 15892 5540 15904
rect 5031 15864 5540 15892
rect 5031 15861 5043 15864
rect 4985 15855 5043 15861
rect 5534 15852 5540 15864
rect 5592 15852 5598 15904
rect 6362 15852 6368 15904
rect 6420 15892 6426 15904
rect 6748 15901 6776 15932
rect 8110 15920 8116 15932
rect 8168 15920 8174 15972
rect 8386 15920 8392 15972
rect 8444 15960 8450 15972
rect 9217 15963 9275 15969
rect 9217 15960 9229 15963
rect 8444 15932 9229 15960
rect 8444 15920 8450 15932
rect 9217 15929 9229 15932
rect 9263 15929 9275 15963
rect 12345 15963 12403 15969
rect 12345 15960 12357 15963
rect 9217 15923 9275 15929
rect 10796 15932 12357 15960
rect 6733 15895 6791 15901
rect 6733 15892 6745 15895
rect 6420 15864 6745 15892
rect 6420 15852 6426 15864
rect 6733 15861 6745 15864
rect 6779 15861 6791 15895
rect 6733 15855 6791 15861
rect 7101 15895 7159 15901
rect 7101 15861 7113 15895
rect 7147 15892 7159 15895
rect 8478 15892 8484 15904
rect 7147 15864 8484 15892
rect 7147 15861 7159 15864
rect 7101 15855 7159 15861
rect 8478 15852 8484 15864
rect 8536 15852 8542 15904
rect 8570 15852 8576 15904
rect 8628 15892 8634 15904
rect 10796 15901 10824 15932
rect 12345 15929 12357 15932
rect 12391 15929 12403 15963
rect 12452 15960 12480 16000
rect 12526 15988 12532 16040
rect 12584 16028 12590 16040
rect 12584 16000 14320 16028
rect 12584 15988 12590 16000
rect 13262 15960 13268 15972
rect 12452 15932 13268 15960
rect 12345 15923 12403 15929
rect 13262 15920 13268 15932
rect 13320 15920 13326 15972
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14194 15963 14252 15969
rect 14194 15960 14206 15963
rect 14148 15932 14206 15960
rect 14148 15920 14154 15932
rect 14194 15929 14206 15932
rect 14240 15929 14252 15963
rect 14292 15960 14320 16000
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16209 16031 16267 16037
rect 16209 16028 16221 16031
rect 15712 16000 16221 16028
rect 15712 15988 15718 16000
rect 16209 15997 16221 16000
rect 16255 16028 16267 16031
rect 17420 16028 17448 16204
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 19705 16167 19763 16173
rect 19705 16133 19717 16167
rect 19751 16164 19763 16167
rect 20346 16164 20352 16176
rect 19751 16136 20352 16164
rect 19751 16133 19763 16136
rect 19705 16127 19763 16133
rect 20346 16124 20352 16136
rect 20404 16164 20410 16176
rect 20404 16136 20668 16164
rect 20404 16124 20410 16136
rect 17862 16096 17868 16108
rect 17823 16068 17868 16096
rect 17862 16056 17868 16068
rect 17920 16096 17926 16108
rect 17920 16068 18460 16096
rect 17920 16056 17926 16068
rect 17678 16028 17684 16040
rect 16255 16000 17448 16028
rect 17639 16000 17684 16028
rect 16255 15997 16267 16000
rect 16209 15991 16267 15997
rect 17678 15988 17684 16000
rect 17736 15988 17742 16040
rect 18138 15988 18144 16040
rect 18196 16028 18202 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18196 16000 18337 16028
rect 18196 15988 18202 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18432 16028 18460 16068
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 20640 16105 20668 16136
rect 20533 16099 20591 16105
rect 20533 16096 20545 16099
rect 20220 16068 20545 16096
rect 20220 16056 20226 16068
rect 20533 16065 20545 16068
rect 20579 16065 20591 16099
rect 20533 16059 20591 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 20625 16059 20683 16065
rect 18581 16031 18639 16037
rect 18581 16028 18593 16031
rect 18432 16000 18593 16028
rect 18325 15991 18383 15997
rect 18581 15997 18593 16000
rect 18627 15997 18639 16031
rect 18581 15991 18639 15997
rect 19518 15988 19524 16040
rect 19576 16028 19582 16040
rect 21177 16031 21235 16037
rect 21177 16028 21189 16031
rect 19576 16000 21189 16028
rect 19576 15988 19582 16000
rect 21177 15997 21189 16000
rect 21223 15997 21235 16031
rect 21177 15991 21235 15997
rect 17954 15960 17960 15972
rect 14292 15932 17960 15960
rect 14194 15923 14252 15929
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 19334 15920 19340 15972
rect 19392 15960 19398 15972
rect 20441 15963 20499 15969
rect 20441 15960 20453 15963
rect 19392 15932 20453 15960
rect 19392 15920 19398 15932
rect 20441 15929 20453 15932
rect 20487 15929 20499 15963
rect 21358 15960 21364 15972
rect 21319 15932 21364 15960
rect 20441 15923 20499 15929
rect 21358 15920 21364 15932
rect 21416 15920 21422 15972
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8628 15864 8769 15892
rect 8628 15852 8634 15864
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 8757 15855 8815 15861
rect 10781 15895 10839 15901
rect 10781 15861 10793 15895
rect 10827 15861 10839 15895
rect 10781 15855 10839 15861
rect 11054 15852 11060 15904
rect 11112 15892 11118 15904
rect 11885 15895 11943 15901
rect 11885 15892 11897 15895
rect 11112 15864 11897 15892
rect 11112 15852 11118 15864
rect 11885 15861 11897 15864
rect 11931 15861 11943 15895
rect 11885 15855 11943 15861
rect 11974 15852 11980 15904
rect 12032 15892 12038 15904
rect 12253 15895 12311 15901
rect 12253 15892 12265 15895
rect 12032 15864 12265 15892
rect 12032 15852 12038 15864
rect 12253 15861 12265 15864
rect 12299 15861 12311 15895
rect 12253 15855 12311 15861
rect 13998 15852 14004 15904
rect 14056 15892 14062 15904
rect 15013 15895 15071 15901
rect 15013 15892 15025 15895
rect 14056 15864 15025 15892
rect 14056 15852 14062 15864
rect 15013 15861 15025 15864
rect 15059 15861 15071 15895
rect 15013 15855 15071 15861
rect 15105 15895 15163 15901
rect 15105 15861 15117 15895
rect 15151 15892 15163 15895
rect 15286 15892 15292 15904
rect 15151 15864 15292 15892
rect 15151 15861 15163 15864
rect 15105 15855 15163 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 15470 15892 15476 15904
rect 15431 15864 15476 15892
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16114 15892 16120 15904
rect 16075 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 16206 15852 16212 15904
rect 16264 15892 16270 15904
rect 17034 15892 17040 15904
rect 16264 15864 17040 15892
rect 16264 15852 16270 15864
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 17773 15895 17831 15901
rect 17773 15861 17785 15895
rect 17819 15892 17831 15895
rect 19610 15892 19616 15904
rect 17819 15864 19616 15892
rect 17819 15861 17831 15864
rect 17773 15855 17831 15861
rect 19610 15852 19616 15864
rect 19668 15852 19674 15904
rect 20073 15895 20131 15901
rect 20073 15861 20085 15895
rect 20119 15892 20131 15895
rect 20254 15892 20260 15904
rect 20119 15864 20260 15892
rect 20119 15861 20131 15864
rect 20073 15855 20131 15861
rect 20254 15852 20260 15864
rect 20312 15852 20318 15904
rect 1104 15802 21896 15824
rect 1104 15750 7912 15802
rect 7964 15750 7976 15802
rect 8028 15750 8040 15802
rect 8092 15750 8104 15802
rect 8156 15750 14843 15802
rect 14895 15750 14907 15802
rect 14959 15750 14971 15802
rect 15023 15750 15035 15802
rect 15087 15750 21896 15802
rect 1104 15728 21896 15750
rect 5718 15688 5724 15700
rect 5679 15660 5724 15688
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 6089 15691 6147 15697
rect 6089 15657 6101 15691
rect 6135 15688 6147 15691
rect 6638 15688 6644 15700
rect 6135 15660 6644 15688
rect 6135 15657 6147 15660
rect 6089 15651 6147 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 7101 15691 7159 15697
rect 7101 15657 7113 15691
rect 7147 15688 7159 15691
rect 8294 15688 8300 15700
rect 7147 15660 8300 15688
rect 7147 15657 7159 15660
rect 7101 15651 7159 15657
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8662 15648 8668 15700
rect 8720 15688 8726 15700
rect 9122 15688 9128 15700
rect 8720 15660 9128 15688
rect 8720 15648 8726 15660
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 11238 15648 11244 15700
rect 11296 15688 11302 15700
rect 11333 15691 11391 15697
rect 11333 15688 11345 15691
rect 11296 15660 11345 15688
rect 11296 15648 11302 15660
rect 11333 15657 11345 15660
rect 11379 15657 11391 15691
rect 11333 15651 11391 15657
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 12066 15688 12072 15700
rect 12023 15660 12072 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 12066 15648 12072 15660
rect 12124 15648 12130 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 12713 15691 12771 15697
rect 12713 15688 12725 15691
rect 12492 15660 12725 15688
rect 12492 15648 12498 15660
rect 12713 15657 12725 15660
rect 12759 15688 12771 15691
rect 12894 15688 12900 15700
rect 12759 15660 12900 15688
rect 12759 15657 12771 15660
rect 12713 15651 12771 15657
rect 12894 15648 12900 15660
rect 12952 15648 12958 15700
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 13998 15688 14004 15700
rect 13959 15660 14004 15688
rect 13998 15648 14004 15660
rect 14056 15648 14062 15700
rect 15286 15688 15292 15700
rect 15247 15660 15292 15688
rect 15286 15648 15292 15660
rect 15344 15648 15350 15700
rect 16117 15691 16175 15697
rect 16117 15657 16129 15691
rect 16163 15688 16175 15691
rect 16942 15688 16948 15700
rect 16163 15660 16804 15688
rect 16903 15660 16948 15688
rect 16163 15657 16175 15660
rect 16117 15651 16175 15657
rect 6733 15623 6791 15629
rect 6733 15589 6745 15623
rect 6779 15620 6791 15623
rect 9309 15623 9367 15629
rect 9309 15620 9321 15623
rect 6779 15592 9321 15620
rect 6779 15589 6791 15592
rect 6733 15583 6791 15589
rect 9309 15589 9321 15592
rect 9355 15589 9367 15623
rect 12802 15620 12808 15632
rect 9309 15583 9367 15589
rect 12406 15592 12808 15620
rect 8478 15552 8484 15564
rect 8536 15561 8542 15564
rect 8536 15555 8559 15561
rect 6564 15524 8484 15552
rect 6564 15493 6592 15524
rect 8478 15512 8484 15524
rect 8547 15552 8559 15555
rect 8662 15552 8668 15564
rect 8547 15524 8668 15552
rect 8547 15521 8559 15524
rect 8536 15515 8559 15521
rect 8536 15512 8542 15515
rect 8662 15512 8668 15524
rect 8720 15512 8726 15564
rect 10226 15561 10232 15564
rect 10220 15552 10232 15561
rect 10139 15524 10232 15552
rect 10220 15515 10232 15524
rect 10284 15552 10290 15564
rect 11793 15555 11851 15561
rect 10284 15524 11008 15552
rect 10226 15512 10232 15515
rect 10284 15512 10290 15524
rect 6549 15487 6607 15493
rect 6549 15453 6561 15487
rect 6595 15453 6607 15487
rect 6549 15447 6607 15453
rect 8757 15487 8815 15493
rect 8757 15453 8769 15487
rect 8803 15484 8815 15487
rect 9582 15484 9588 15496
rect 8803 15456 9588 15484
rect 8803 15453 8815 15456
rect 8757 15447 8815 15453
rect 9582 15444 9588 15456
rect 9640 15484 9646 15496
rect 9953 15487 10011 15493
rect 9953 15484 9965 15487
rect 9640 15456 9965 15484
rect 9640 15444 9646 15456
rect 9953 15453 9965 15456
rect 9999 15453 10011 15487
rect 9953 15447 10011 15453
rect 10980 15428 11008 15524
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12406 15552 12434 15592
rect 12802 15580 12808 15592
rect 12860 15580 12866 15632
rect 16776 15620 16804 15660
rect 16942 15648 16948 15660
rect 17000 15648 17006 15700
rect 17313 15691 17371 15697
rect 17313 15657 17325 15691
rect 17359 15688 17371 15691
rect 17862 15688 17868 15700
rect 17359 15660 17868 15688
rect 17359 15657 17371 15660
rect 17313 15651 17371 15657
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 18690 15648 18696 15700
rect 18748 15688 18754 15700
rect 18969 15691 19027 15697
rect 18969 15688 18981 15691
rect 18748 15660 18981 15688
rect 18748 15648 18754 15660
rect 18969 15657 18981 15660
rect 19015 15657 19027 15691
rect 18969 15651 19027 15657
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19668 15660 19809 15688
rect 19668 15648 19674 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 19797 15651 19855 15657
rect 16850 15620 16856 15632
rect 12995 15592 16436 15620
rect 16763 15592 16856 15620
rect 12618 15552 12624 15564
rect 11839 15524 12434 15552
rect 12579 15524 12624 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12897 15487 12955 15493
rect 12897 15453 12909 15487
rect 12943 15484 12955 15487
rect 12995 15484 13023 15592
rect 13262 15512 13268 15564
rect 13320 15552 13326 15564
rect 13633 15555 13691 15561
rect 13320 15524 13492 15552
rect 13320 15512 13326 15524
rect 12943 15456 13023 15484
rect 13357 15487 13415 15493
rect 12943 15453 12955 15456
rect 12897 15447 12955 15453
rect 13357 15453 13369 15487
rect 13403 15453 13415 15487
rect 13464 15484 13492 15524
rect 13633 15521 13645 15555
rect 13679 15552 13691 15555
rect 14090 15552 14096 15564
rect 13679 15524 14096 15552
rect 13679 15521 13691 15524
rect 13633 15515 13691 15521
rect 14090 15512 14096 15524
rect 14148 15512 14154 15564
rect 14921 15555 14979 15561
rect 14200 15524 14780 15552
rect 14200 15484 14228 15524
rect 13464 15456 14228 15484
rect 14645 15487 14703 15493
rect 13357 15447 13415 15453
rect 14645 15453 14657 15487
rect 14691 15453 14703 15487
rect 14645 15447 14703 15453
rect 5534 15376 5540 15428
rect 5592 15416 5598 15428
rect 5592 15388 7512 15416
rect 5592 15376 5598 15388
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 6638 15348 6644 15360
rect 6420 15320 6644 15348
rect 6420 15308 6426 15320
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 7374 15348 7380 15360
rect 7335 15320 7380 15348
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 7484 15348 7512 15388
rect 10962 15376 10968 15428
rect 11020 15416 11026 15428
rect 12912 15416 12940 15447
rect 11020 15388 12940 15416
rect 13372 15416 13400 15447
rect 13814 15416 13820 15428
rect 13372 15388 13820 15416
rect 11020 15376 11026 15388
rect 13814 15376 13820 15388
rect 13872 15416 13878 15428
rect 14660 15416 14688 15447
rect 13872 15388 14688 15416
rect 14752 15416 14780 15524
rect 14921 15521 14933 15555
rect 14967 15552 14979 15555
rect 15286 15552 15292 15564
rect 14967 15524 15292 15552
rect 14967 15521 14979 15524
rect 14921 15515 14979 15521
rect 15286 15512 15292 15524
rect 15344 15512 15350 15564
rect 16206 15552 16212 15564
rect 16167 15524 16212 15552
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 14829 15487 14887 15493
rect 14829 15453 14841 15487
rect 14875 15484 14887 15487
rect 15194 15484 15200 15496
rect 14875 15456 15200 15484
rect 14875 15453 14887 15456
rect 14829 15447 14887 15453
rect 15194 15444 15200 15456
rect 15252 15444 15258 15496
rect 16114 15484 16120 15496
rect 15304 15456 16120 15484
rect 15304 15416 15332 15456
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 16408 15493 16436 15592
rect 16850 15580 16856 15592
rect 16908 15620 16914 15632
rect 18448 15623 18506 15629
rect 16908 15592 17724 15620
rect 16908 15580 16914 15592
rect 16761 15555 16819 15561
rect 16761 15521 16773 15555
rect 16807 15521 16819 15555
rect 17696 15552 17724 15592
rect 18448 15589 18460 15623
rect 18494 15620 18506 15623
rect 19426 15620 19432 15632
rect 18494 15592 19432 15620
rect 18494 15589 18506 15592
rect 18448 15583 18506 15589
rect 19426 15580 19432 15592
rect 19484 15620 19490 15632
rect 19484 15592 20392 15620
rect 19484 15580 19490 15592
rect 20165 15555 20223 15561
rect 20165 15552 20177 15555
rect 17696 15524 20177 15552
rect 16761 15515 16819 15521
rect 20165 15521 20177 15524
rect 20211 15521 20223 15555
rect 20165 15515 20223 15521
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15484 16451 15487
rect 16574 15484 16580 15496
rect 16439 15456 16580 15484
rect 16439 15453 16451 15456
rect 16393 15447 16451 15453
rect 16574 15444 16580 15456
rect 16632 15444 16638 15496
rect 14752 15388 15332 15416
rect 13872 15376 13878 15388
rect 15930 15376 15936 15428
rect 15988 15416 15994 15428
rect 16776 15416 16804 15515
rect 18693 15487 18751 15493
rect 18693 15453 18705 15487
rect 18739 15484 18751 15487
rect 19426 15484 19432 15496
rect 18739 15456 19432 15484
rect 18739 15453 18751 15456
rect 18693 15447 18751 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 20364 15493 20392 15592
rect 20806 15580 20812 15632
rect 20864 15620 20870 15632
rect 21177 15623 21235 15629
rect 21177 15620 21189 15623
rect 20864 15592 21189 15620
rect 20864 15580 20870 15592
rect 21177 15589 21189 15592
rect 21223 15589 21235 15623
rect 21177 15583 21235 15589
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15453 20315 15487
rect 20257 15447 20315 15453
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 15988 15388 16804 15416
rect 15988 15376 15994 15388
rect 12066 15348 12072 15360
rect 7484 15320 12072 15348
rect 12066 15308 12072 15320
rect 12124 15308 12130 15360
rect 12250 15348 12256 15360
rect 12211 15320 12256 15348
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 14458 15308 14464 15360
rect 14516 15348 14522 15360
rect 15102 15348 15108 15360
rect 14516 15320 15108 15348
rect 14516 15308 14522 15320
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 15746 15348 15752 15360
rect 15707 15320 15752 15348
rect 15746 15308 15752 15320
rect 15804 15308 15810 15360
rect 16022 15308 16028 15360
rect 16080 15348 16086 15360
rect 20272 15348 20300 15447
rect 21266 15348 21272 15360
rect 16080 15320 20300 15348
rect 21227 15320 21272 15348
rect 16080 15308 16086 15320
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 4447 15258
rect 4499 15206 4511 15258
rect 4563 15206 4575 15258
rect 4627 15206 4639 15258
rect 4691 15206 11378 15258
rect 11430 15206 11442 15258
rect 11494 15206 11506 15258
rect 11558 15206 11570 15258
rect 11622 15206 18308 15258
rect 18360 15206 18372 15258
rect 18424 15206 18436 15258
rect 18488 15206 18500 15258
rect 18552 15206 21896 15258
rect 1104 15184 21896 15206
rect 7377 15147 7435 15153
rect 7377 15113 7389 15147
rect 7423 15144 7435 15147
rect 9674 15144 9680 15156
rect 7423 15116 9680 15144
rect 7423 15113 7435 15116
rect 7377 15107 7435 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 11054 15144 11060 15156
rect 10143 15116 11060 15144
rect 7834 15076 7840 15088
rect 7795 15048 7840 15076
rect 7834 15036 7840 15048
rect 7892 15036 7898 15088
rect 9309 15079 9367 15085
rect 9309 15045 9321 15079
rect 9355 15076 9367 15079
rect 9766 15076 9772 15088
rect 9355 15048 9628 15076
rect 9355 15045 9367 15048
rect 9309 15039 9367 15045
rect 8570 15008 8576 15020
rect 8531 14980 8576 15008
rect 8570 14968 8576 14980
rect 8628 14968 8634 15020
rect 8662 14968 8668 15020
rect 8720 15008 8726 15020
rect 8720 14980 8765 15008
rect 8720 14968 8726 14980
rect 7650 14940 7656 14952
rect 7611 14912 7656 14940
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 9125 14943 9183 14949
rect 9125 14909 9137 14943
rect 9171 14909 9183 14943
rect 9600 14940 9628 15048
rect 9692 15048 9772 15076
rect 9692 15017 9720 15048
rect 9766 15036 9772 15048
rect 9824 15036 9830 15088
rect 10143 15076 10171 15116
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15144 11391 15147
rect 11974 15144 11980 15156
rect 11379 15116 11980 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12526 15104 12532 15156
rect 12584 15144 12590 15156
rect 18141 15147 18199 15153
rect 18141 15144 18153 15147
rect 12584 15116 18153 15144
rect 12584 15104 12590 15116
rect 18141 15113 18153 15116
rect 18187 15113 18199 15147
rect 18141 15107 18199 15113
rect 18509 15147 18567 15153
rect 18509 15113 18521 15147
rect 18555 15144 18567 15147
rect 18555 15116 21220 15144
rect 18555 15113 18567 15116
rect 18509 15107 18567 15113
rect 9876 15048 10171 15076
rect 10321 15079 10379 15085
rect 9876 15017 9904 15048
rect 10321 15045 10333 15079
rect 10367 15076 10379 15079
rect 11882 15076 11888 15088
rect 10367 15048 11888 15076
rect 10367 15045 10379 15048
rect 10321 15039 10379 15045
rect 11882 15036 11888 15048
rect 11940 15036 11946 15088
rect 14734 15036 14740 15088
rect 14792 15076 14798 15088
rect 14921 15079 14979 15085
rect 14921 15076 14933 15079
rect 14792 15048 14933 15076
rect 14792 15036 14798 15048
rect 14921 15045 14933 15048
rect 14967 15045 14979 15079
rect 16574 15076 16580 15088
rect 16535 15048 16580 15076
rect 14921 15039 14979 15045
rect 9677 15011 9735 15017
rect 9677 14977 9689 15011
rect 9723 14977 9735 15011
rect 9677 14971 9735 14977
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 10781 15011 10839 15017
rect 10781 14977 10793 15011
rect 10827 15008 10839 15011
rect 10962 15008 10968 15020
rect 10827 14980 10968 15008
rect 10827 14977 10839 14980
rect 10781 14971 10839 14977
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 12342 14968 12348 15020
rect 12400 15008 12406 15020
rect 12437 15011 12495 15017
rect 12437 15008 12449 15011
rect 12400 14980 12449 15008
rect 12400 14968 12406 14980
rect 12437 14977 12449 14980
rect 12483 14977 12495 15011
rect 12437 14971 12495 14977
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 12676 14980 12909 15008
rect 12676 14968 12682 14980
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 14936 15008 14964 15039
rect 16574 15036 16580 15048
rect 16632 15036 16638 15088
rect 16666 15036 16672 15088
rect 16724 15076 16730 15088
rect 16724 15048 19656 15076
rect 16724 15036 16730 15048
rect 19628 15020 19656 15048
rect 14936 14980 15332 15008
rect 12897 14971 12955 14977
rect 10505 14943 10563 14949
rect 9600 14912 9812 14940
rect 9125 14903 9183 14909
rect 6641 14875 6699 14881
rect 6641 14841 6653 14875
rect 6687 14872 6699 14875
rect 7742 14872 7748 14884
rect 6687 14844 7748 14872
rect 6687 14841 6699 14844
rect 6641 14835 6699 14841
rect 7742 14832 7748 14844
rect 7800 14872 7806 14884
rect 9140 14872 9168 14903
rect 9784 14884 9812 14912
rect 10505 14909 10517 14943
rect 10551 14940 10563 14943
rect 10873 14943 10931 14949
rect 10873 14940 10885 14943
rect 10551 14912 10885 14940
rect 10551 14909 10563 14912
rect 10505 14903 10563 14909
rect 10873 14909 10885 14912
rect 10919 14940 10931 14943
rect 12250 14940 12256 14952
rect 10919 14912 12112 14940
rect 12211 14912 12256 14940
rect 10919 14909 10931 14912
rect 10873 14903 10931 14909
rect 9674 14872 9680 14884
rect 7800 14844 8524 14872
rect 9140 14844 9680 14872
rect 7800 14832 7806 14844
rect 7006 14804 7012 14816
rect 6967 14776 7012 14804
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 8113 14807 8171 14813
rect 8113 14773 8125 14807
rect 8159 14804 8171 14807
rect 8386 14804 8392 14816
rect 8159 14776 8392 14804
rect 8159 14773 8171 14776
rect 8113 14767 8171 14773
rect 8386 14764 8392 14776
rect 8444 14764 8450 14816
rect 8496 14813 8524 14844
rect 9674 14832 9680 14844
rect 9732 14832 9738 14884
rect 9766 14832 9772 14884
rect 9824 14832 9830 14884
rect 9950 14832 9956 14884
rect 10008 14872 10014 14884
rect 10008 14844 10053 14872
rect 10008 14832 10014 14844
rect 10226 14832 10232 14884
rect 10284 14872 10290 14884
rect 10284 14844 11928 14872
rect 10284 14832 10290 14844
rect 8481 14807 8539 14813
rect 8481 14773 8493 14807
rect 8527 14804 8539 14807
rect 10505 14807 10563 14813
rect 10505 14804 10517 14807
rect 8527 14776 10517 14804
rect 8527 14773 8539 14776
rect 8481 14767 8539 14773
rect 10505 14773 10517 14776
rect 10551 14773 10563 14807
rect 10505 14767 10563 14773
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11900 14813 11928 14844
rect 11885 14807 11943 14813
rect 11020 14776 11065 14804
rect 11020 14764 11026 14776
rect 11885 14773 11897 14807
rect 11931 14773 11943 14807
rect 12084 14804 12112 14912
rect 12250 14900 12256 14912
rect 12308 14900 12314 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 13630 14940 13636 14952
rect 13587 14912 13636 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 13630 14900 13636 14912
rect 13688 14900 13694 14952
rect 13814 14949 13820 14952
rect 13808 14940 13820 14949
rect 13775 14912 13820 14940
rect 13808 14903 13820 14912
rect 13814 14900 13820 14903
rect 13872 14900 13878 14952
rect 15102 14900 15108 14952
rect 15160 14940 15166 14952
rect 15197 14943 15255 14949
rect 15197 14940 15209 14943
rect 15160 14912 15209 14940
rect 15160 14900 15166 14912
rect 15197 14909 15209 14912
rect 15243 14909 15255 14943
rect 15304 14940 15332 14980
rect 16206 14968 16212 15020
rect 16264 15008 16270 15020
rect 18969 15011 19027 15017
rect 16264 14980 18460 15008
rect 16264 14968 16270 14980
rect 15453 14943 15511 14949
rect 15453 14940 15465 14943
rect 15304 14912 15465 14940
rect 15197 14903 15255 14909
rect 15453 14909 15465 14912
rect 15499 14909 15511 14943
rect 15453 14903 15511 14909
rect 15838 14900 15844 14952
rect 15896 14940 15902 14952
rect 17865 14943 17923 14949
rect 17865 14940 17877 14943
rect 15896 14912 17877 14940
rect 15896 14900 15902 14912
rect 17865 14909 17877 14912
rect 17911 14909 17923 14943
rect 17865 14903 17923 14909
rect 18141 14943 18199 14949
rect 18141 14909 18153 14943
rect 18187 14940 18199 14943
rect 18325 14943 18383 14949
rect 18325 14940 18337 14943
rect 18187 14912 18337 14940
rect 18187 14909 18199 14912
rect 18141 14903 18199 14909
rect 18325 14909 18337 14912
rect 18371 14909 18383 14943
rect 18432 14940 18460 14980
rect 18969 14977 18981 15011
rect 19015 15008 19027 15011
rect 19334 15008 19340 15020
rect 19015 14980 19340 15008
rect 19015 14977 19027 14980
rect 18969 14971 19027 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 19242 14940 19248 14952
rect 18432 14912 19248 14940
rect 18325 14903 18383 14909
rect 19242 14900 19248 14912
rect 19300 14900 19306 14952
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19484 14912 19656 14940
rect 19484 14900 19490 14912
rect 12158 14832 12164 14884
rect 12216 14872 12222 14884
rect 15562 14872 15568 14884
rect 12216 14844 15568 14872
rect 12216 14832 12222 14844
rect 15562 14832 15568 14844
rect 15620 14832 15626 14884
rect 16206 14832 16212 14884
rect 16264 14872 16270 14884
rect 17129 14875 17187 14881
rect 17129 14872 17141 14875
rect 16264 14844 17141 14872
rect 16264 14832 16270 14844
rect 17129 14841 17141 14844
rect 17175 14841 17187 14875
rect 19518 14872 19524 14884
rect 17129 14835 17187 14841
rect 18064 14844 19524 14872
rect 12250 14804 12256 14816
rect 12084 14776 12256 14804
rect 11885 14767 11943 14773
rect 12250 14764 12256 14776
rect 12308 14764 12314 14816
rect 12345 14807 12403 14813
rect 12345 14773 12357 14807
rect 12391 14804 12403 14807
rect 15746 14804 15752 14816
rect 12391 14776 15752 14804
rect 12391 14773 12403 14776
rect 12345 14767 12403 14773
rect 15746 14764 15752 14776
rect 15804 14764 15810 14816
rect 15838 14764 15844 14816
rect 15896 14804 15902 14816
rect 17954 14804 17960 14816
rect 15896 14776 17960 14804
rect 15896 14764 15902 14776
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 18064 14813 18092 14844
rect 19518 14832 19524 14844
rect 19576 14832 19582 14884
rect 19628 14872 19656 14912
rect 20346 14900 20352 14952
rect 20404 14949 20410 14952
rect 21192 14949 21220 15116
rect 20404 14940 20416 14949
rect 20625 14943 20683 14949
rect 20404 14912 20449 14940
rect 20404 14903 20416 14912
rect 20625 14909 20637 14943
rect 20671 14909 20683 14943
rect 20625 14903 20683 14909
rect 21177 14943 21235 14949
rect 21177 14909 21189 14943
rect 21223 14909 21235 14943
rect 21177 14903 21235 14909
rect 20404 14900 20410 14903
rect 20640 14872 20668 14903
rect 21358 14872 21364 14884
rect 19628 14844 20668 14872
rect 21319 14844 21364 14872
rect 21358 14832 21364 14844
rect 21416 14832 21422 14884
rect 18049 14807 18107 14813
rect 18049 14773 18061 14807
rect 18095 14773 18107 14807
rect 19242 14804 19248 14816
rect 19203 14776 19248 14804
rect 18049 14767 18107 14773
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 1104 14714 21896 14736
rect 1104 14662 7912 14714
rect 7964 14662 7976 14714
rect 8028 14662 8040 14714
rect 8092 14662 8104 14714
rect 8156 14662 14843 14714
rect 14895 14662 14907 14714
rect 14959 14662 14971 14714
rect 15023 14662 15035 14714
rect 15087 14662 21896 14714
rect 1104 14640 21896 14662
rect 5534 14560 5540 14612
rect 5592 14600 5598 14612
rect 5629 14603 5687 14609
rect 5629 14600 5641 14603
rect 5592 14572 5641 14600
rect 5592 14560 5598 14572
rect 5629 14569 5641 14572
rect 5675 14600 5687 14603
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5675 14572 6009 14600
rect 5675 14569 5687 14572
rect 5629 14563 5687 14569
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6454 14600 6460 14612
rect 6236 14572 6460 14600
rect 6236 14560 6242 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 7282 14560 7288 14612
rect 7340 14600 7346 14612
rect 7469 14603 7527 14609
rect 7469 14600 7481 14603
rect 7340 14572 7481 14600
rect 7340 14560 7346 14572
rect 7469 14569 7481 14572
rect 7515 14569 7527 14603
rect 7469 14563 7527 14569
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 7708 14572 7941 14600
rect 7708 14560 7714 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 8386 14600 8392 14612
rect 8347 14572 8392 14600
rect 7929 14563 7987 14569
rect 8386 14560 8392 14572
rect 8444 14560 8450 14612
rect 12897 14603 12955 14609
rect 12897 14600 12909 14603
rect 8496 14572 12909 14600
rect 2682 14492 2688 14544
rect 2740 14532 2746 14544
rect 8496 14532 8524 14572
rect 12897 14569 12909 14572
rect 12943 14569 12955 14603
rect 12897 14563 12955 14569
rect 13357 14603 13415 14609
rect 13357 14569 13369 14603
rect 13403 14600 13415 14603
rect 13538 14600 13544 14612
rect 13403 14572 13544 14600
rect 13403 14569 13415 14572
rect 13357 14563 13415 14569
rect 13538 14560 13544 14572
rect 13596 14560 13602 14612
rect 13906 14560 13912 14612
rect 13964 14600 13970 14612
rect 14185 14603 14243 14609
rect 14185 14600 14197 14603
rect 13964 14572 14197 14600
rect 13964 14560 13970 14572
rect 14185 14569 14197 14572
rect 14231 14569 14243 14603
rect 14185 14563 14243 14569
rect 14274 14560 14280 14612
rect 14332 14600 14338 14612
rect 14369 14603 14427 14609
rect 14369 14600 14381 14603
rect 14332 14572 14381 14600
rect 14332 14560 14338 14572
rect 14369 14569 14381 14572
rect 14415 14569 14427 14603
rect 14369 14563 14427 14569
rect 14921 14603 14979 14609
rect 14921 14569 14933 14603
rect 14967 14600 14979 14603
rect 16666 14600 16672 14612
rect 14967 14572 16672 14600
rect 14967 14569 14979 14572
rect 14921 14563 14979 14569
rect 16666 14560 16672 14572
rect 16724 14560 16730 14612
rect 17310 14560 17316 14612
rect 17368 14600 17374 14612
rect 18325 14603 18383 14609
rect 17368 14572 18276 14600
rect 17368 14560 17374 14572
rect 2740 14504 8524 14532
rect 2740 14492 2746 14504
rect 9214 14492 9220 14544
rect 9272 14532 9278 14544
rect 10962 14532 10968 14544
rect 9272 14504 10968 14532
rect 9272 14492 9278 14504
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11517 14535 11575 14541
rect 11517 14501 11529 14535
rect 11563 14532 11575 14535
rect 11698 14532 11704 14544
rect 11563 14504 11704 14532
rect 11563 14501 11575 14504
rect 11517 14495 11575 14501
rect 11698 14492 11704 14504
rect 11756 14492 11762 14544
rect 15378 14532 15384 14544
rect 11992 14504 15384 14532
rect 7650 14464 7656 14476
rect 7611 14436 7656 14464
rect 7650 14424 7656 14436
rect 7708 14424 7714 14476
rect 8294 14464 8300 14476
rect 8255 14436 8300 14464
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 9493 14467 9551 14473
rect 9493 14433 9505 14467
rect 9539 14464 9551 14467
rect 9582 14464 9588 14476
rect 9539 14436 9588 14464
rect 9539 14433 9551 14436
rect 9493 14427 9551 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 9760 14467 9818 14473
rect 9760 14433 9772 14467
rect 9806 14464 9818 14467
rect 11992 14464 12020 14504
rect 15378 14492 15384 14504
rect 15436 14492 15442 14544
rect 15565 14535 15623 14541
rect 15565 14501 15577 14535
rect 15611 14532 15623 14535
rect 18248 14532 18276 14572
rect 18325 14569 18337 14603
rect 18371 14600 18383 14603
rect 18371 14572 21220 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 15611 14504 15792 14532
rect 18248 14504 18644 14532
rect 15611 14501 15623 14504
rect 15565 14495 15623 14501
rect 12158 14464 12164 14476
rect 9806 14436 12020 14464
rect 12119 14436 12164 14464
rect 9806 14433 9818 14436
rect 9760 14427 9818 14433
rect 12158 14424 12164 14436
rect 12216 14424 12222 14476
rect 12989 14467 13047 14473
rect 12989 14464 13001 14467
rect 12406 14436 13001 14464
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 8481 14399 8539 14405
rect 8481 14396 8493 14399
rect 7432 14368 8493 14396
rect 7432 14356 7438 14368
rect 8481 14365 8493 14368
rect 8527 14365 8539 14399
rect 8481 14359 8539 14365
rect 11238 14356 11244 14408
rect 11296 14396 11302 14408
rect 11609 14399 11667 14405
rect 11609 14396 11621 14399
rect 11296 14368 11621 14396
rect 11296 14356 11302 14368
rect 11609 14365 11621 14368
rect 11655 14365 11667 14399
rect 11609 14359 11667 14365
rect 11701 14399 11759 14405
rect 11701 14365 11713 14399
rect 11747 14365 11759 14399
rect 11701 14359 11759 14365
rect 7193 14331 7251 14337
rect 7193 14297 7205 14331
rect 7239 14328 7251 14331
rect 8846 14328 8852 14340
rect 7239 14300 8852 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 8846 14288 8852 14300
rect 8904 14288 8910 14340
rect 11716 14328 11744 14359
rect 12066 14356 12072 14408
rect 12124 14396 12130 14408
rect 12406 14396 12434 14436
rect 12989 14433 13001 14436
rect 13035 14433 13047 14467
rect 12989 14427 13047 14433
rect 13817 14467 13875 14473
rect 13817 14433 13829 14467
rect 13863 14464 13875 14467
rect 14182 14464 14188 14476
rect 13863 14436 14188 14464
rect 13863 14433 13875 14436
rect 13817 14427 13875 14433
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14737 14467 14795 14473
rect 14737 14464 14749 14467
rect 14323 14436 14749 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 14737 14433 14749 14436
rect 14783 14433 14795 14467
rect 15764 14464 15792 14504
rect 16114 14464 16120 14476
rect 15764 14436 16120 14464
rect 14737 14427 14795 14433
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 16482 14424 16488 14476
rect 16540 14464 16546 14476
rect 17598 14467 17656 14473
rect 17598 14464 17610 14467
rect 16540 14436 17610 14464
rect 16540 14424 16546 14436
rect 17598 14433 17610 14436
rect 17644 14433 17656 14467
rect 18138 14464 18144 14476
rect 18099 14436 18144 14464
rect 17598 14427 17656 14433
rect 18138 14424 18144 14436
rect 18196 14424 18202 14476
rect 18616 14473 18644 14504
rect 20346 14492 20352 14544
rect 20404 14532 20410 14544
rect 21192 14541 21220 14572
rect 21177 14535 21235 14541
rect 20404 14504 20576 14532
rect 20404 14492 20410 14504
rect 18601 14467 18659 14473
rect 18601 14433 18613 14467
rect 18647 14433 18659 14467
rect 18601 14427 18659 14433
rect 19061 14467 19119 14473
rect 19061 14433 19073 14467
rect 19107 14433 19119 14467
rect 19061 14427 19119 14433
rect 12802 14396 12808 14408
rect 12124 14368 12434 14396
rect 12715 14368 12808 14396
rect 12124 14356 12130 14368
rect 12802 14356 12808 14368
rect 12860 14396 12866 14408
rect 14458 14396 14464 14408
rect 12860 14368 14464 14396
rect 12860 14356 12866 14368
rect 14458 14356 14464 14368
rect 14516 14356 14522 14408
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15841 14399 15899 14405
rect 15841 14365 15853 14399
rect 15887 14365 15899 14399
rect 17862 14396 17868 14408
rect 17823 14368 17868 14396
rect 15841 14359 15899 14365
rect 10428 14300 11744 14328
rect 12345 14331 12403 14337
rect 6825 14263 6883 14269
rect 6825 14229 6837 14263
rect 6871 14260 6883 14263
rect 7374 14260 7380 14272
rect 6871 14232 7380 14260
rect 6871 14229 6883 14232
rect 6825 14223 6883 14229
rect 7374 14220 7380 14232
rect 7432 14220 7438 14272
rect 7834 14220 7840 14272
rect 7892 14260 7898 14272
rect 8570 14260 8576 14272
rect 7892 14232 8576 14260
rect 7892 14220 7898 14232
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9217 14263 9275 14269
rect 9217 14229 9229 14263
rect 9263 14260 9275 14263
rect 9306 14260 9312 14272
rect 9263 14232 9312 14260
rect 9263 14229 9275 14232
rect 9217 14223 9275 14229
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9490 14220 9496 14272
rect 9548 14260 9554 14272
rect 10428 14260 10456 14300
rect 12345 14297 12357 14331
rect 12391 14328 12403 14331
rect 13906 14328 13912 14340
rect 12391 14300 13912 14328
rect 12391 14297 12403 14300
rect 12345 14291 12403 14297
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 14001 14331 14059 14337
rect 14001 14297 14013 14331
rect 14047 14328 14059 14331
rect 14642 14328 14648 14340
rect 14047 14300 14648 14328
rect 14047 14297 14059 14300
rect 14001 14291 14059 14297
rect 14642 14288 14648 14300
rect 14700 14288 14706 14340
rect 15194 14328 15200 14340
rect 15155 14300 15200 14328
rect 15194 14288 15200 14300
rect 15252 14288 15258 14340
rect 15378 14288 15384 14340
rect 15436 14328 15442 14340
rect 15856 14328 15884 14359
rect 17862 14356 17868 14368
rect 17920 14356 17926 14408
rect 17954 14356 17960 14408
rect 18012 14396 18018 14408
rect 19076 14396 19104 14427
rect 19334 14424 19340 14476
rect 19392 14464 19398 14476
rect 20438 14464 20444 14476
rect 19392 14436 20444 14464
rect 19392 14424 19398 14436
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 20548 14464 20576 14504
rect 21177 14501 21189 14535
rect 21223 14501 21235 14535
rect 21177 14495 21235 14501
rect 20548 14436 20668 14464
rect 20530 14396 20536 14408
rect 18012 14368 19104 14396
rect 20491 14368 20536 14396
rect 18012 14356 18018 14368
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 20640 14405 20668 14436
rect 20625 14399 20683 14405
rect 20625 14365 20637 14399
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 16485 14331 16543 14337
rect 16485 14328 16497 14331
rect 15436 14300 16497 14328
rect 15436 14288 15442 14300
rect 16485 14297 16497 14300
rect 16531 14297 16543 14331
rect 16485 14291 16543 14297
rect 19245 14331 19303 14337
rect 19245 14297 19257 14331
rect 19291 14328 19303 14331
rect 21174 14328 21180 14340
rect 19291 14300 21180 14328
rect 19291 14297 19303 14300
rect 19245 14291 19303 14297
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 21358 14328 21364 14340
rect 21319 14300 21364 14328
rect 21358 14288 21364 14300
rect 21416 14288 21422 14340
rect 9548 14232 10456 14260
rect 10873 14263 10931 14269
rect 9548 14220 9554 14232
rect 10873 14229 10885 14263
rect 10919 14260 10931 14263
rect 11054 14260 11060 14272
rect 10919 14232 11060 14260
rect 10919 14229 10931 14232
rect 10873 14223 10931 14229
rect 11054 14220 11060 14232
rect 11112 14220 11118 14272
rect 11146 14220 11152 14272
rect 11204 14260 11210 14272
rect 18782 14260 18788 14272
rect 11204 14232 11249 14260
rect 18743 14232 18788 14260
rect 11204 14220 11210 14232
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 19334 14220 19340 14272
rect 19392 14260 19398 14272
rect 19613 14263 19671 14269
rect 19613 14260 19625 14263
rect 19392 14232 19625 14260
rect 19392 14220 19398 14232
rect 19613 14229 19625 14232
rect 19659 14229 19671 14263
rect 19613 14223 19671 14229
rect 20073 14263 20131 14269
rect 20073 14229 20085 14263
rect 20119 14260 20131 14263
rect 20346 14260 20352 14272
rect 20119 14232 20352 14260
rect 20119 14229 20131 14232
rect 20073 14223 20131 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 1104 14170 21896 14192
rect 1104 14118 4447 14170
rect 4499 14118 4511 14170
rect 4563 14118 4575 14170
rect 4627 14118 4639 14170
rect 4691 14118 11378 14170
rect 11430 14118 11442 14170
rect 11494 14118 11506 14170
rect 11558 14118 11570 14170
rect 11622 14118 18308 14170
rect 18360 14118 18372 14170
rect 18424 14118 18436 14170
rect 18488 14118 18500 14170
rect 18552 14118 21896 14170
rect 1104 14096 21896 14118
rect 6086 14016 6092 14068
rect 6144 14056 6150 14068
rect 7101 14059 7159 14065
rect 7101 14056 7113 14059
rect 6144 14028 7113 14056
rect 6144 14016 6150 14028
rect 7101 14025 7113 14028
rect 7147 14025 7159 14059
rect 7101 14019 7159 14025
rect 7561 14059 7619 14065
rect 7561 14025 7573 14059
rect 7607 14056 7619 14059
rect 7742 14056 7748 14068
rect 7607 14028 7748 14056
rect 7607 14025 7619 14028
rect 7561 14019 7619 14025
rect 7742 14016 7748 14028
rect 7800 14016 7806 14068
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8389 14059 8447 14065
rect 8389 14056 8401 14059
rect 8352 14028 8401 14056
rect 8352 14016 8358 14028
rect 8389 14025 8401 14028
rect 8435 14056 8447 14059
rect 8754 14056 8760 14068
rect 8435 14028 8760 14056
rect 8435 14025 8447 14028
rect 8389 14019 8447 14025
rect 8754 14016 8760 14028
rect 8812 14016 8818 14068
rect 9309 14059 9367 14065
rect 9309 14025 9321 14059
rect 9355 14056 9367 14059
rect 10686 14056 10692 14068
rect 9355 14028 10692 14056
rect 9355 14025 9367 14028
rect 9309 14019 9367 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 12158 14056 12164 14068
rect 12119 14028 12164 14056
rect 12158 14016 12164 14028
rect 12216 14016 12222 14068
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14090 14056 14096 14068
rect 14051 14028 14096 14056
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 17862 14016 17868 14068
rect 17920 14056 17926 14068
rect 19886 14056 19892 14068
rect 17920 14028 18552 14056
rect 19847 14028 19892 14056
rect 17920 14016 17926 14028
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 7834 13988 7840 14000
rect 5224 13960 7840 13988
rect 5224 13948 5230 13960
rect 7834 13948 7840 13960
rect 7892 13948 7898 14000
rect 9490 13948 9496 14000
rect 9548 13988 9554 14000
rect 9585 13991 9643 13997
rect 9585 13988 9597 13991
rect 9548 13960 9597 13988
rect 9548 13948 9554 13960
rect 9585 13957 9597 13960
rect 9631 13957 9643 13991
rect 9585 13951 9643 13957
rect 11333 13991 11391 13997
rect 11333 13957 11345 13991
rect 11379 13988 11391 13991
rect 12434 13988 12440 14000
rect 11379 13960 12440 13988
rect 11379 13957 11391 13960
rect 11333 13951 11391 13957
rect 12434 13948 12440 13960
rect 12492 13948 12498 14000
rect 16022 13948 16028 14000
rect 16080 13988 16086 14000
rect 16482 13988 16488 14000
rect 16080 13960 16488 13988
rect 16080 13948 16086 13960
rect 16482 13948 16488 13960
rect 16540 13988 16546 14000
rect 17129 13991 17187 13997
rect 17129 13988 17141 13991
rect 16540 13960 17141 13988
rect 16540 13948 16546 13960
rect 17129 13957 17141 13960
rect 17175 13957 17187 13991
rect 17129 13951 17187 13957
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 5500 13892 6837 13920
rect 5500 13880 5506 13892
rect 6825 13889 6837 13892
rect 6871 13920 6883 13923
rect 9950 13920 9956 13932
rect 6871 13892 9956 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 14737 13923 14795 13929
rect 11624 13892 12480 13920
rect 11624 13864 11652 13892
rect 12452 13864 12480 13892
rect 14737 13889 14749 13923
rect 14783 13920 14795 13923
rect 15378 13920 15384 13932
rect 14783 13892 15384 13920
rect 14783 13889 14795 13892
rect 14737 13883 14795 13889
rect 7650 13812 7656 13864
rect 7708 13852 7714 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7708 13824 8217 13852
rect 7708 13812 7714 13824
rect 8205 13821 8217 13824
rect 8251 13821 8263 13855
rect 8846 13852 8852 13864
rect 8807 13824 8852 13852
rect 8205 13815 8263 13821
rect 8220 13716 8248 13815
rect 8846 13812 8852 13824
rect 8904 13812 8910 13864
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 10410 13852 10416 13864
rect 9171 13824 10416 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10612 13824 10977 13852
rect 10318 13744 10324 13796
rect 10376 13784 10382 13796
rect 10612 13784 10640 13824
rect 10965 13821 10977 13824
rect 11011 13852 11023 13855
rect 11606 13852 11612 13864
rect 11011 13824 11612 13852
rect 11011 13821 11023 13824
rect 10965 13815 11023 13821
rect 11606 13812 11612 13824
rect 11664 13812 11670 13864
rect 11882 13812 11888 13864
rect 11940 13852 11946 13864
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11940 13824 11989 13852
rect 11940 13812 11946 13824
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 12434 13852 12440 13864
rect 12347 13824 12440 13852
rect 11977 13815 12035 13821
rect 12434 13812 12440 13824
rect 12492 13812 12498 13864
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 14752 13852 14780 13883
rect 15378 13880 15384 13892
rect 15436 13880 15442 13932
rect 18524 13929 18552 14028
rect 19886 14016 19892 14028
rect 19944 14016 19950 14068
rect 19242 13948 19248 14000
rect 19300 13988 19306 14000
rect 19300 13960 20484 13988
rect 19300 13948 19306 13960
rect 16393 13923 16451 13929
rect 16393 13889 16405 13923
rect 16439 13889 16451 13923
rect 16393 13883 16451 13889
rect 18509 13923 18567 13929
rect 18509 13889 18521 13923
rect 18555 13920 18567 13923
rect 19426 13920 19432 13932
rect 18555 13892 19432 13920
rect 18555 13889 18567 13892
rect 18509 13883 18567 13889
rect 16298 13852 16304 13864
rect 14516 13824 14780 13852
rect 16259 13824 16304 13852
rect 14516 13812 14522 13824
rect 16298 13812 16304 13824
rect 16356 13812 16362 13864
rect 16408 13796 16436 13883
rect 19426 13880 19432 13892
rect 19484 13880 19490 13932
rect 19521 13923 19579 13929
rect 19521 13889 19533 13923
rect 19567 13920 19579 13923
rect 19610 13920 19616 13932
rect 19567 13892 19616 13920
rect 19567 13889 19579 13892
rect 19521 13883 19579 13889
rect 19610 13880 19616 13892
rect 19668 13880 19674 13932
rect 20346 13920 20352 13932
rect 20307 13892 20352 13920
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 20456 13929 20484 13960
rect 20441 13923 20499 13929
rect 20441 13889 20453 13923
rect 20487 13889 20499 13923
rect 20441 13883 20499 13889
rect 18782 13812 18788 13864
rect 18840 13852 18846 13864
rect 21177 13855 21235 13861
rect 21177 13852 21189 13855
rect 18840 13824 21189 13852
rect 18840 13812 18846 13824
rect 21177 13821 21189 13824
rect 21223 13821 21235 13855
rect 21358 13852 21364 13864
rect 21319 13824 21364 13852
rect 21177 13815 21235 13821
rect 21358 13812 21364 13824
rect 21416 13812 21422 13864
rect 10376 13756 10640 13784
rect 10376 13744 10382 13756
rect 10686 13744 10692 13796
rect 10744 13793 10750 13796
rect 10744 13784 10756 13793
rect 12704 13787 12762 13793
rect 10744 13756 10789 13784
rect 10744 13747 10756 13756
rect 12704 13753 12716 13787
rect 12750 13784 12762 13787
rect 12802 13784 12808 13796
rect 12750 13756 12808 13784
rect 12750 13753 12762 13756
rect 12704 13747 12762 13753
rect 10744 13744 10750 13747
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 14550 13784 14556 13796
rect 14463 13756 14556 13784
rect 14550 13744 14556 13756
rect 14608 13784 14614 13796
rect 15194 13784 15200 13796
rect 14608 13756 15200 13784
rect 14608 13744 14614 13756
rect 15194 13744 15200 13756
rect 15252 13744 15258 13796
rect 16206 13784 16212 13796
rect 16167 13756 16212 13784
rect 16206 13744 16212 13756
rect 16264 13744 16270 13796
rect 16390 13784 16396 13796
rect 16303 13756 16396 13784
rect 16390 13744 16396 13756
rect 16448 13784 16454 13796
rect 17862 13784 17868 13796
rect 16448 13756 17868 13784
rect 16448 13744 16454 13756
rect 17862 13744 17868 13756
rect 17920 13784 17926 13796
rect 18242 13787 18300 13793
rect 18242 13784 18254 13787
rect 17920 13756 18254 13784
rect 17920 13744 17926 13756
rect 18242 13753 18254 13756
rect 18288 13753 18300 13787
rect 20254 13784 20260 13796
rect 20215 13756 20260 13784
rect 18242 13747 18300 13753
rect 20254 13744 20260 13756
rect 20312 13744 20318 13796
rect 8665 13719 8723 13725
rect 8665 13716 8677 13719
rect 8220 13688 8677 13716
rect 8665 13685 8677 13688
rect 8711 13685 8723 13719
rect 8665 13679 8723 13685
rect 8938 13676 8944 13728
rect 8996 13716 9002 13728
rect 12526 13716 12532 13728
rect 8996 13688 12532 13716
rect 8996 13676 9002 13688
rect 12526 13676 12532 13688
rect 12584 13676 12590 13728
rect 13354 13676 13360 13728
rect 13412 13716 13418 13728
rect 14182 13716 14188 13728
rect 13412 13688 14188 13716
rect 13412 13676 13418 13688
rect 14182 13676 14188 13688
rect 14240 13716 14246 13728
rect 14461 13719 14519 13725
rect 14461 13716 14473 13719
rect 14240 13688 14473 13716
rect 14240 13676 14246 13688
rect 14461 13685 14473 13688
rect 14507 13685 14519 13719
rect 14461 13679 14519 13685
rect 14734 13676 14740 13728
rect 14792 13716 14798 13728
rect 15105 13719 15163 13725
rect 15105 13716 15117 13719
rect 14792 13688 15117 13716
rect 14792 13676 14798 13688
rect 15105 13685 15117 13688
rect 15151 13685 15163 13719
rect 15838 13716 15844 13728
rect 15799 13688 15844 13716
rect 15105 13679 15163 13685
rect 15838 13676 15844 13688
rect 15896 13676 15902 13728
rect 18874 13716 18880 13728
rect 18835 13688 18880 13716
rect 18874 13676 18880 13688
rect 18932 13676 18938 13728
rect 19242 13716 19248 13728
rect 19203 13688 19248 13716
rect 19242 13676 19248 13688
rect 19300 13676 19306 13728
rect 19337 13719 19395 13725
rect 19337 13685 19349 13719
rect 19383 13716 19395 13719
rect 19702 13716 19708 13728
rect 19383 13688 19708 13716
rect 19383 13685 19395 13688
rect 19337 13679 19395 13685
rect 19702 13676 19708 13688
rect 19760 13676 19766 13728
rect 1104 13626 21896 13648
rect 1104 13574 7912 13626
rect 7964 13574 7976 13626
rect 8028 13574 8040 13626
rect 8092 13574 8104 13626
rect 8156 13574 14843 13626
rect 14895 13574 14907 13626
rect 14959 13574 14971 13626
rect 15023 13574 15035 13626
rect 15087 13574 21896 13626
rect 1104 13552 21896 13574
rect 6730 13512 6736 13524
rect 6691 13484 6736 13512
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 8757 13515 8815 13521
rect 8757 13481 8769 13515
rect 8803 13512 8815 13515
rect 8803 13484 14228 13512
rect 8803 13481 8815 13484
rect 8757 13475 8815 13481
rect 7469 13447 7527 13453
rect 7469 13413 7481 13447
rect 7515 13444 7527 13447
rect 7742 13444 7748 13456
rect 7515 13416 7748 13444
rect 7515 13413 7527 13416
rect 7469 13407 7527 13413
rect 7742 13404 7748 13416
rect 7800 13404 7806 13456
rect 8938 13404 8944 13456
rect 8996 13444 9002 13456
rect 9125 13447 9183 13453
rect 9125 13444 9137 13447
rect 8996 13416 9137 13444
rect 8996 13404 9002 13416
rect 9125 13413 9137 13416
rect 9171 13413 9183 13447
rect 9125 13407 9183 13413
rect 9858 13404 9864 13456
rect 9916 13444 9922 13456
rect 10778 13444 10784 13456
rect 9916 13416 10784 13444
rect 9916 13404 9922 13416
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 11054 13404 11060 13456
rect 11112 13444 11118 13456
rect 11342 13447 11400 13453
rect 11342 13444 11354 13447
rect 11112 13416 11354 13444
rect 11112 13404 11118 13416
rect 11342 13413 11354 13416
rect 11388 13444 11400 13447
rect 11388 13416 12204 13444
rect 11388 13413 11400 13416
rect 11342 13407 11400 13413
rect 6730 13336 6736 13388
rect 6788 13376 6794 13388
rect 7098 13376 7104 13388
rect 6788 13348 7104 13376
rect 6788 13336 6794 13348
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 8294 13376 8300 13388
rect 8255 13348 8300 13376
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 8573 13379 8631 13385
rect 8573 13345 8585 13379
rect 8619 13376 8631 13379
rect 8956 13376 8984 13404
rect 8619 13348 8984 13376
rect 9493 13379 9551 13385
rect 8619 13345 8631 13348
rect 8573 13339 8631 13345
rect 9493 13345 9505 13379
rect 9539 13376 9551 13379
rect 10042 13376 10048 13388
rect 9539 13348 10048 13376
rect 9539 13345 9551 13348
rect 9493 13339 9551 13345
rect 10042 13336 10048 13348
rect 10100 13336 10106 13388
rect 11606 13376 11612 13388
rect 11567 13348 11612 13376
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 12176 13376 12204 13416
rect 12250 13404 12256 13456
rect 12308 13444 12314 13456
rect 14200 13444 14228 13484
rect 14274 13472 14280 13524
rect 14332 13512 14338 13524
rect 14553 13515 14611 13521
rect 14553 13512 14565 13515
rect 14332 13484 14565 13512
rect 14332 13472 14338 13484
rect 14553 13481 14565 13484
rect 14599 13481 14611 13515
rect 14553 13475 14611 13481
rect 15381 13515 15439 13521
rect 15381 13481 15393 13515
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 15749 13515 15807 13521
rect 15749 13481 15761 13515
rect 15795 13512 15807 13515
rect 15838 13512 15844 13524
rect 15795 13484 15844 13512
rect 15795 13481 15807 13484
rect 15749 13475 15807 13481
rect 12308 13416 12353 13444
rect 14200 13416 14780 13444
rect 12308 13404 12314 13416
rect 13633 13379 13691 13385
rect 12176 13348 12480 13376
rect 7837 13311 7895 13317
rect 7837 13277 7849 13311
rect 7883 13308 7895 13311
rect 10226 13308 10232 13320
rect 7883 13280 10232 13308
rect 7883 13277 7895 13280
rect 7837 13271 7895 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 11790 13268 11796 13320
rect 11848 13308 11854 13320
rect 12158 13308 12164 13320
rect 11848 13280 12164 13308
rect 11848 13268 11854 13280
rect 12158 13268 12164 13280
rect 12216 13308 12222 13320
rect 12452 13317 12480 13348
rect 13633 13345 13645 13379
rect 13679 13376 13691 13379
rect 14642 13376 14648 13388
rect 13679 13348 14648 13376
rect 13679 13345 13691 13348
rect 13633 13339 13691 13345
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12216 13280 12357 13308
rect 12216 13268 12222 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12437 13311 12495 13317
rect 12437 13277 12449 13311
rect 12483 13277 12495 13311
rect 12437 13271 12495 13277
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13044 13280 13737 13308
rect 13044 13268 13050 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 13909 13311 13967 13317
rect 13909 13277 13921 13311
rect 13955 13308 13967 13311
rect 14090 13308 14096 13320
rect 13955 13280 14096 13308
rect 13955 13277 13967 13280
rect 13909 13271 13967 13277
rect 14090 13268 14096 13280
rect 14148 13268 14154 13320
rect 14752 13308 14780 13416
rect 14921 13379 14979 13385
rect 14921 13345 14933 13379
rect 14967 13376 14979 13379
rect 15396 13376 15424 13475
rect 15838 13472 15844 13484
rect 15896 13472 15902 13524
rect 16390 13512 16396 13524
rect 16351 13484 16396 13512
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 16942 13472 16948 13524
rect 17000 13512 17006 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 17000 13484 18429 13512
rect 17000 13472 17006 13484
rect 18417 13481 18429 13484
rect 18463 13481 18475 13515
rect 18417 13475 18475 13481
rect 19242 13472 19248 13524
rect 19300 13512 19306 13524
rect 20073 13515 20131 13521
rect 20073 13512 20085 13515
rect 19300 13484 20085 13512
rect 19300 13472 19306 13484
rect 20073 13481 20085 13484
rect 20119 13481 20131 13515
rect 20073 13475 20131 13481
rect 17402 13444 17408 13456
rect 14967 13348 15424 13376
rect 15488 13416 17408 13444
rect 14967 13345 14979 13348
rect 14921 13339 14979 13345
rect 15488 13308 15516 13416
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 17586 13404 17592 13456
rect 17644 13444 17650 13456
rect 20162 13444 20168 13456
rect 17644 13416 20168 13444
rect 17644 13404 17650 13416
rect 20162 13404 20168 13416
rect 20220 13404 20226 13456
rect 21174 13444 21180 13456
rect 21135 13416 21180 13444
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13376 15899 13379
rect 17034 13376 17040 13388
rect 15887 13348 17040 13376
rect 15887 13345 15899 13348
rect 15841 13339 15899 13345
rect 17034 13336 17040 13348
rect 17092 13336 17098 13388
rect 17126 13336 17132 13388
rect 17184 13376 17190 13388
rect 17506 13379 17564 13385
rect 17506 13376 17518 13379
rect 17184 13348 17518 13376
rect 17184 13336 17190 13348
rect 17506 13345 17518 13348
rect 17552 13376 17564 13379
rect 19245 13379 19303 13385
rect 17552 13348 18092 13376
rect 17552 13345 17564 13348
rect 17506 13339 17564 13345
rect 16022 13308 16028 13320
rect 14752 13280 15516 13308
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 17770 13308 17776 13320
rect 17731 13280 17776 13308
rect 17770 13268 17776 13280
rect 17828 13268 17834 13320
rect 9674 13240 9680 13252
rect 9635 13212 9680 13240
rect 9674 13200 9680 13212
rect 9732 13200 9738 13252
rect 16574 13240 16580 13252
rect 11624 13212 16580 13240
rect 7101 13175 7159 13181
rect 7101 13141 7113 13175
rect 7147 13172 7159 13175
rect 7374 13172 7380 13184
rect 7147 13144 7380 13172
rect 7147 13141 7159 13144
rect 7101 13135 7159 13141
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 8386 13172 8392 13184
rect 8159 13144 8392 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 8386 13132 8392 13144
rect 8444 13132 8450 13184
rect 10229 13175 10287 13181
rect 10229 13141 10241 13175
rect 10275 13172 10287 13175
rect 10686 13172 10692 13184
rect 10275 13144 10692 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10686 13132 10692 13144
rect 10744 13132 10750 13184
rect 10870 13132 10876 13184
rect 10928 13172 10934 13184
rect 11624 13172 11652 13212
rect 16574 13200 16580 13212
rect 16632 13200 16638 13252
rect 17954 13240 17960 13252
rect 17788 13212 17960 13240
rect 11882 13172 11888 13184
rect 10928 13144 11652 13172
rect 11843 13144 11888 13172
rect 10928 13132 10934 13144
rect 11882 13132 11888 13144
rect 11940 13132 11946 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12897 13175 12955 13181
rect 12897 13172 12909 13175
rect 12032 13144 12909 13172
rect 12032 13132 12038 13144
rect 12897 13141 12909 13144
rect 12943 13141 12955 13175
rect 13262 13172 13268 13184
rect 13223 13144 13268 13172
rect 12897 13135 12955 13141
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 15105 13175 15163 13181
rect 15105 13141 15117 13175
rect 15151 13172 15163 13175
rect 17788 13172 17816 13212
rect 17954 13200 17960 13212
rect 18012 13200 18018 13252
rect 18064 13240 18092 13348
rect 19245 13345 19257 13379
rect 19291 13376 19303 13379
rect 20441 13379 20499 13385
rect 20441 13376 20453 13379
rect 19291 13348 20453 13376
rect 19291 13345 19303 13348
rect 19245 13339 19303 13345
rect 20441 13345 20453 13348
rect 20487 13345 20499 13379
rect 20441 13339 20499 13345
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13345 20591 13379
rect 20533 13339 20591 13345
rect 18138 13268 18144 13320
rect 18196 13308 18202 13320
rect 18509 13311 18567 13317
rect 18509 13308 18521 13311
rect 18196 13280 18521 13308
rect 18196 13268 18202 13280
rect 18509 13277 18521 13280
rect 18555 13277 18567 13311
rect 18509 13271 18567 13277
rect 18601 13311 18659 13317
rect 18601 13277 18613 13311
rect 18647 13277 18659 13311
rect 18601 13271 18659 13277
rect 19797 13311 19855 13317
rect 19797 13277 19809 13311
rect 19843 13308 19855 13311
rect 20070 13308 20076 13320
rect 19843 13280 20076 13308
rect 19843 13277 19855 13280
rect 19797 13271 19855 13277
rect 18616 13240 18644 13271
rect 20070 13268 20076 13280
rect 20128 13308 20134 13320
rect 20548 13308 20576 13339
rect 20128 13280 20576 13308
rect 20717 13311 20775 13317
rect 20128 13268 20134 13280
rect 20717 13277 20729 13311
rect 20763 13277 20775 13311
rect 20717 13271 20775 13277
rect 18064 13212 18644 13240
rect 20622 13200 20628 13252
rect 20680 13240 20686 13252
rect 20732 13240 20760 13271
rect 21358 13240 21364 13252
rect 20680 13212 20760 13240
rect 21319 13212 21364 13240
rect 20680 13200 20686 13212
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 18046 13172 18052 13184
rect 15151 13144 17816 13172
rect 18007 13144 18052 13172
rect 15151 13141 15163 13144
rect 15105 13135 15163 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 1104 13082 21896 13104
rect 1104 13030 4447 13082
rect 4499 13030 4511 13082
rect 4563 13030 4575 13082
rect 4627 13030 4639 13082
rect 4691 13030 11378 13082
rect 11430 13030 11442 13082
rect 11494 13030 11506 13082
rect 11558 13030 11570 13082
rect 11622 13030 18308 13082
rect 18360 13030 18372 13082
rect 18424 13030 18436 13082
rect 18488 13030 18500 13082
rect 18552 13030 21896 13082
rect 1104 13008 21896 13030
rect 7009 12971 7067 12977
rect 7009 12937 7021 12971
rect 7055 12968 7067 12971
rect 7742 12968 7748 12980
rect 7055 12940 7748 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 7837 12971 7895 12977
rect 7837 12937 7849 12971
rect 7883 12968 7895 12971
rect 10870 12968 10876 12980
rect 7883 12940 10876 12968
rect 7883 12937 7895 12940
rect 7837 12931 7895 12937
rect 10870 12928 10876 12940
rect 10928 12928 10934 12980
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11296 12940 11345 12968
rect 11296 12928 11302 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 11425 12971 11483 12977
rect 11425 12937 11437 12971
rect 11471 12968 11483 12971
rect 11974 12968 11980 12980
rect 11471 12940 11980 12968
rect 11471 12937 11483 12940
rect 11425 12931 11483 12937
rect 11974 12928 11980 12940
rect 12032 12968 12038 12980
rect 14277 12971 14335 12977
rect 14277 12968 14289 12971
rect 12032 12940 14289 12968
rect 12032 12928 12038 12940
rect 14277 12937 14289 12940
rect 14323 12937 14335 12971
rect 15197 12971 15255 12977
rect 14277 12931 14335 12937
rect 14384 12940 14688 12968
rect 5074 12860 5080 12912
rect 5132 12900 5138 12912
rect 6822 12900 6828 12912
rect 5132 12872 6828 12900
rect 5132 12860 5138 12872
rect 6822 12860 6828 12872
rect 6880 12900 6886 12912
rect 7285 12903 7343 12909
rect 7285 12900 7297 12903
rect 6880 12872 7297 12900
rect 6880 12860 6886 12872
rect 7285 12869 7297 12872
rect 7331 12900 7343 12903
rect 7650 12900 7656 12912
rect 7331 12872 7656 12900
rect 7331 12869 7343 12872
rect 7285 12863 7343 12869
rect 7650 12860 7656 12872
rect 7708 12860 7714 12912
rect 9858 12900 9864 12912
rect 9819 12872 9864 12900
rect 9858 12860 9864 12872
rect 9916 12860 9922 12912
rect 9950 12860 9956 12912
rect 10008 12900 10014 12912
rect 10137 12903 10195 12909
rect 10137 12900 10149 12903
rect 10008 12872 10149 12900
rect 10008 12860 10014 12872
rect 10137 12869 10149 12872
rect 10183 12869 10195 12903
rect 10137 12863 10195 12869
rect 10226 12860 10232 12912
rect 10284 12900 10290 12912
rect 12158 12900 12164 12912
rect 10284 12872 12164 12900
rect 10284 12860 10290 12872
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 14384 12900 14412 12940
rect 12406 12872 14412 12900
rect 10778 12832 10784 12844
rect 10739 12804 10784 12832
rect 10778 12792 10784 12804
rect 10836 12792 10842 12844
rect 10873 12835 10931 12841
rect 10873 12801 10885 12835
rect 10919 12832 10931 12835
rect 11882 12832 11888 12844
rect 10919 12804 11888 12832
rect 10919 12801 10931 12804
rect 10873 12795 10931 12801
rect 11882 12792 11888 12804
rect 11940 12792 11946 12844
rect 7282 12724 7288 12776
rect 7340 12764 7346 12776
rect 7653 12767 7711 12773
rect 7653 12764 7665 12767
rect 7340 12736 7665 12764
rect 7340 12724 7346 12736
rect 7653 12733 7665 12736
rect 7699 12733 7711 12767
rect 7653 12727 7711 12733
rect 9237 12767 9295 12773
rect 9237 12733 9249 12767
rect 9283 12764 9295 12767
rect 9398 12764 9404 12776
rect 9283 12736 9404 12764
rect 9283 12733 9295 12736
rect 9237 12727 9295 12733
rect 9398 12724 9404 12736
rect 9456 12724 9462 12776
rect 9493 12767 9551 12773
rect 9493 12733 9505 12767
rect 9539 12764 9551 12767
rect 9582 12764 9588 12776
rect 9539 12736 9588 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 8386 12656 8392 12708
rect 8444 12696 8450 12708
rect 9508 12696 9536 12727
rect 9582 12724 9588 12736
rect 9640 12724 9646 12776
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 12406 12764 12434 12872
rect 14458 12860 14464 12912
rect 14516 12900 14522 12912
rect 14660 12900 14688 12940
rect 15197 12937 15209 12971
rect 15243 12968 15255 12971
rect 15286 12968 15292 12980
rect 15243 12940 15292 12968
rect 15243 12937 15255 12940
rect 15197 12931 15255 12937
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 18874 12968 18880 12980
rect 15672 12940 18880 12968
rect 15672 12900 15700 12940
rect 18874 12928 18880 12940
rect 18932 12928 18938 12980
rect 19702 12928 19708 12980
rect 19760 12968 19766 12980
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 19760 12940 20453 12968
rect 19760 12928 19766 12940
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20441 12931 20499 12937
rect 14516 12872 14596 12900
rect 14660 12872 15700 12900
rect 18509 12903 18567 12909
rect 14516 12860 14522 12872
rect 13081 12835 13139 12841
rect 13081 12801 13093 12835
rect 13127 12832 13139 12835
rect 14090 12832 14096 12844
rect 13127 12804 13952 12832
rect 14051 12804 14096 12832
rect 13127 12801 13139 12804
rect 13081 12795 13139 12801
rect 10367 12736 12434 12764
rect 12805 12767 12863 12773
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 12805 12733 12817 12767
rect 12851 12764 12863 12767
rect 13262 12764 13268 12776
rect 12851 12736 13268 12764
rect 12851 12733 12863 12736
rect 12805 12727 12863 12733
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13924 12764 13952 12804
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14568 12841 14596 12872
rect 18509 12869 18521 12903
rect 18555 12869 18567 12903
rect 18509 12863 18567 12869
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12801 14611 12835
rect 14553 12795 14611 12801
rect 16206 12792 16212 12844
rect 16264 12832 16270 12844
rect 16301 12835 16359 12841
rect 16301 12832 16313 12835
rect 16264 12804 16313 12832
rect 16264 12792 16270 12804
rect 16301 12801 16313 12804
rect 16347 12801 16359 12835
rect 16301 12795 16359 12801
rect 17126 12792 17132 12844
rect 17184 12832 17190 12844
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17184 12804 17509 12832
rect 17184 12792 17190 12804
rect 17497 12801 17509 12804
rect 17543 12832 17555 12835
rect 18524 12832 18552 12863
rect 17543 12804 18552 12832
rect 17543 12801 17555 12804
rect 17497 12795 17555 12801
rect 20622 12792 20628 12844
rect 20680 12832 20686 12844
rect 20993 12835 21051 12841
rect 20993 12832 21005 12835
rect 20680 12804 21005 12832
rect 20680 12792 20686 12804
rect 20993 12801 21005 12804
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 14458 12764 14464 12776
rect 13924 12736 14464 12764
rect 14458 12724 14464 12736
rect 14516 12724 14522 12776
rect 14734 12724 14740 12776
rect 14792 12764 14798 12776
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14792 12736 14841 12764
rect 14792 12724 14798 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 15010 12724 15016 12776
rect 15068 12764 15074 12776
rect 16945 12767 17003 12773
rect 16945 12764 16957 12767
rect 15068 12736 16957 12764
rect 15068 12724 15074 12736
rect 16945 12733 16957 12736
rect 16991 12764 17003 12767
rect 17402 12764 17408 12776
rect 16991 12736 17408 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 17402 12724 17408 12736
rect 17460 12724 17466 12776
rect 17678 12764 17684 12776
rect 17639 12736 17684 12764
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 19610 12724 19616 12776
rect 19668 12773 19674 12776
rect 19668 12764 19680 12773
rect 19889 12767 19947 12773
rect 19668 12736 19713 12764
rect 19668 12727 19680 12736
rect 19889 12733 19901 12767
rect 19935 12733 19947 12767
rect 19889 12727 19947 12733
rect 19668 12724 19674 12727
rect 8444 12668 9536 12696
rect 8444 12656 8450 12668
rect 10410 12656 10416 12708
rect 10468 12696 10474 12708
rect 13817 12699 13875 12705
rect 10468 12668 12480 12696
rect 10468 12656 10474 12668
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7650 12628 7656 12640
rect 6972 12600 7656 12628
rect 6972 12588 6978 12600
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 8113 12631 8171 12637
rect 8113 12597 8125 12631
rect 8159 12628 8171 12631
rect 8478 12628 8484 12640
rect 8159 12600 8484 12628
rect 8159 12597 8171 12600
rect 8113 12591 8171 12597
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 9858 12588 9864 12640
rect 9916 12628 9922 12640
rect 10870 12628 10876 12640
rect 9916 12600 10876 12628
rect 9916 12588 9922 12600
rect 10870 12588 10876 12600
rect 10928 12628 10934 12640
rect 10965 12631 11023 12637
rect 10965 12628 10977 12631
rect 10928 12600 10977 12628
rect 10928 12588 10934 12600
rect 10965 12597 10977 12600
rect 11011 12597 11023 12631
rect 10965 12591 11023 12597
rect 11146 12588 11152 12640
rect 11204 12628 11210 12640
rect 11425 12631 11483 12637
rect 11425 12628 11437 12631
rect 11204 12600 11437 12628
rect 11204 12588 11210 12600
rect 11425 12597 11437 12600
rect 11471 12597 11483 12631
rect 11882 12628 11888 12640
rect 11843 12600 11888 12628
rect 11425 12591 11483 12597
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 12452 12637 12480 12668
rect 13817 12665 13829 12699
rect 13863 12696 13875 12699
rect 13863 12668 15792 12696
rect 13863 12665 13875 12668
rect 13817 12659 13875 12665
rect 12437 12631 12495 12637
rect 12437 12597 12449 12631
rect 12483 12597 12495 12631
rect 12437 12591 12495 12597
rect 12897 12631 12955 12637
rect 12897 12597 12909 12631
rect 12943 12628 12955 12631
rect 13449 12631 13507 12637
rect 13449 12628 13461 12631
rect 12943 12600 13461 12628
rect 12943 12597 12955 12600
rect 12897 12591 12955 12597
rect 13449 12597 13461 12600
rect 13495 12597 13507 12631
rect 13449 12591 13507 12597
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 15764 12637 15792 12668
rect 15838 12656 15844 12708
rect 15896 12696 15902 12708
rect 16209 12699 16267 12705
rect 16209 12696 16221 12699
rect 15896 12668 16221 12696
rect 15896 12656 15902 12668
rect 16209 12665 16221 12668
rect 16255 12665 16267 12699
rect 17420 12696 17448 12724
rect 17586 12696 17592 12708
rect 17420 12668 17592 12696
rect 16209 12659 16267 12665
rect 17586 12656 17592 12668
rect 17644 12656 17650 12708
rect 19426 12656 19432 12708
rect 19484 12696 19490 12708
rect 19904 12696 19932 12727
rect 20070 12696 20076 12708
rect 19484 12668 20076 12696
rect 19484 12656 19490 12668
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 14277 12631 14335 12637
rect 13964 12600 14009 12628
rect 13964 12588 13970 12600
rect 14277 12597 14289 12631
rect 14323 12628 14335 12631
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14323 12600 14749 12628
rect 14323 12597 14335 12600
rect 14277 12591 14335 12597
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 15749 12631 15807 12637
rect 15749 12597 15761 12631
rect 15795 12597 15807 12631
rect 16114 12628 16120 12640
rect 16075 12600 16120 12628
rect 15749 12591 15807 12597
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 16758 12588 16764 12640
rect 16816 12628 16822 12640
rect 17773 12631 17831 12637
rect 17773 12628 17785 12631
rect 16816 12600 17785 12628
rect 16816 12588 16822 12600
rect 17773 12597 17785 12600
rect 17819 12597 17831 12631
rect 17773 12591 17831 12597
rect 17954 12588 17960 12640
rect 18012 12628 18018 12640
rect 18141 12631 18199 12637
rect 18141 12628 18153 12631
rect 18012 12600 18153 12628
rect 18012 12588 18018 12600
rect 18141 12597 18153 12600
rect 18187 12597 18199 12631
rect 18141 12591 18199 12597
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 20809 12631 20867 12637
rect 20809 12628 20821 12631
rect 20772 12600 20821 12628
rect 20772 12588 20778 12600
rect 20809 12597 20821 12600
rect 20855 12597 20867 12631
rect 20809 12591 20867 12597
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 20956 12600 21001 12628
rect 20956 12588 20962 12600
rect 1104 12538 21896 12560
rect 1104 12486 7912 12538
rect 7964 12486 7976 12538
rect 8028 12486 8040 12538
rect 8092 12486 8104 12538
rect 8156 12486 14843 12538
rect 14895 12486 14907 12538
rect 14959 12486 14971 12538
rect 15023 12486 15035 12538
rect 15087 12486 21896 12538
rect 1104 12464 21896 12486
rect 6086 12384 6092 12436
rect 6144 12424 6150 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6144 12396 6929 12424
rect 6144 12384 6150 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 7837 12427 7895 12433
rect 7837 12393 7849 12427
rect 7883 12424 7895 12427
rect 10226 12424 10232 12436
rect 7883 12396 10232 12424
rect 7883 12393 7895 12396
rect 7837 12387 7895 12393
rect 6932 12356 6960 12387
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 11698 12424 11704 12436
rect 11659 12396 11704 12424
rect 11698 12384 11704 12396
rect 11756 12384 11762 12436
rect 11790 12384 11796 12436
rect 11848 12424 11854 12436
rect 13814 12424 13820 12436
rect 11848 12396 13820 12424
rect 11848 12384 11854 12396
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 14090 12384 14096 12436
rect 14148 12424 14154 12436
rect 14550 12424 14556 12436
rect 14148 12396 14556 12424
rect 14148 12384 14154 12396
rect 14550 12384 14556 12396
rect 14608 12384 14614 12436
rect 16298 12384 16304 12436
rect 16356 12424 16362 12436
rect 16485 12427 16543 12433
rect 16485 12424 16497 12427
rect 16356 12396 16497 12424
rect 16356 12384 16362 12396
rect 16485 12393 16497 12396
rect 16531 12393 16543 12427
rect 16485 12387 16543 12393
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 16945 12427 17003 12433
rect 16945 12424 16957 12427
rect 16908 12396 16957 12424
rect 16908 12384 16914 12396
rect 16945 12393 16957 12396
rect 16991 12393 17003 12427
rect 16945 12387 17003 12393
rect 17034 12384 17040 12436
rect 17092 12424 17098 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17092 12396 17509 12424
rect 17092 12384 17098 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 17865 12427 17923 12433
rect 17865 12393 17877 12427
rect 17911 12424 17923 12427
rect 18046 12424 18052 12436
rect 17911 12396 18052 12424
rect 17911 12393 17923 12396
rect 17865 12387 17923 12393
rect 18046 12384 18052 12396
rect 18104 12384 18110 12436
rect 18969 12427 19027 12433
rect 18969 12393 18981 12427
rect 19015 12424 19027 12427
rect 19150 12424 19156 12436
rect 19015 12396 19156 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19150 12384 19156 12396
rect 19208 12384 19214 12436
rect 19610 12384 19616 12436
rect 19668 12424 19674 12436
rect 19889 12427 19947 12433
rect 19889 12424 19901 12427
rect 19668 12396 19901 12424
rect 19668 12384 19674 12396
rect 19889 12393 19901 12396
rect 19935 12393 19947 12427
rect 19889 12387 19947 12393
rect 6932 12328 8688 12356
rect 7653 12291 7711 12297
rect 7653 12257 7665 12291
rect 7699 12288 7711 12291
rect 7742 12288 7748 12300
rect 7699 12260 7748 12288
rect 7699 12257 7711 12260
rect 7653 12251 7711 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 8110 12288 8116 12300
rect 8071 12260 8116 12288
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 8294 12248 8300 12300
rect 8352 12288 8358 12300
rect 8573 12291 8631 12297
rect 8573 12288 8585 12291
rect 8352 12260 8585 12288
rect 8352 12248 8358 12260
rect 8573 12257 8585 12260
rect 8619 12257 8631 12291
rect 8660 12288 8688 12328
rect 9398 12316 9404 12368
rect 9456 12356 9462 12368
rect 11333 12359 11391 12365
rect 9456 12328 11192 12356
rect 9456 12316 9462 12328
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 8660 12260 9597 12288
rect 8573 12251 8631 12257
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 9677 12291 9735 12297
rect 9677 12257 9689 12291
rect 9723 12288 9735 12291
rect 10318 12288 10324 12300
rect 9723 12260 10324 12288
rect 9723 12257 9735 12260
rect 9677 12251 9735 12257
rect 2222 12180 2228 12232
rect 2280 12220 2286 12232
rect 7098 12220 7104 12232
rect 2280 12192 7104 12220
rect 2280 12180 2286 12192
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7377 12223 7435 12229
rect 7377 12189 7389 12223
rect 7423 12220 7435 12223
rect 8128 12220 8156 12248
rect 7423 12192 8156 12220
rect 7423 12189 7435 12192
rect 7377 12183 7435 12189
rect 8478 12180 8484 12232
rect 8536 12220 8542 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8536 12192 9413 12220
rect 8536 12180 8542 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9600 12220 9628 12251
rect 10318 12248 10324 12260
rect 10376 12248 10382 12300
rect 10505 12291 10563 12297
rect 10505 12257 10517 12291
rect 10551 12288 10563 12291
rect 10870 12288 10876 12300
rect 10551 12260 10876 12288
rect 10551 12257 10563 12260
rect 10505 12251 10563 12257
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11164 12288 11192 12328
rect 11333 12325 11345 12359
rect 11379 12356 11391 12359
rect 11882 12356 11888 12368
rect 11379 12328 11888 12356
rect 11379 12325 11391 12328
rect 11333 12319 11391 12325
rect 11882 12316 11888 12328
rect 11940 12316 11946 12368
rect 13538 12356 13544 12368
rect 12406 12328 13544 12356
rect 12406 12288 12434 12328
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 18230 12356 18236 12368
rect 13780 12328 18236 12356
rect 13780 12316 13786 12328
rect 18230 12316 18236 12328
rect 18288 12316 18294 12368
rect 20070 12316 20076 12368
rect 20128 12356 20134 12368
rect 20128 12328 21312 12356
rect 20128 12316 20134 12328
rect 12526 12288 12532 12300
rect 11164 12260 12434 12288
rect 12487 12260 12532 12288
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 12796 12291 12854 12297
rect 12796 12257 12808 12291
rect 12842 12288 12854 12291
rect 13262 12288 13268 12300
rect 12842 12260 13268 12288
rect 12842 12257 12854 12260
rect 12796 12251 12854 12257
rect 13262 12248 13268 12260
rect 13320 12248 13326 12300
rect 13998 12248 14004 12300
rect 14056 12288 14062 12300
rect 15666 12291 15724 12297
rect 15666 12288 15678 12291
rect 14056 12260 15678 12288
rect 14056 12248 14062 12260
rect 15666 12257 15678 12260
rect 15712 12288 15724 12291
rect 15933 12291 15991 12297
rect 15712 12260 15884 12288
rect 15712 12257 15724 12260
rect 15666 12251 15724 12257
rect 10686 12220 10692 12232
rect 9600 12192 10692 12220
rect 9401 12183 9459 12189
rect 10686 12180 10692 12192
rect 10744 12180 10750 12232
rect 10778 12180 10784 12232
rect 10836 12220 10842 12232
rect 11057 12223 11115 12229
rect 11057 12220 11069 12223
rect 10836 12192 11069 12220
rect 10836 12180 10842 12192
rect 11057 12189 11069 12192
rect 11103 12189 11115 12223
rect 11057 12183 11115 12189
rect 11241 12223 11299 12229
rect 11241 12189 11253 12223
rect 11287 12220 11299 12223
rect 11698 12220 11704 12232
rect 11287 12192 11704 12220
rect 11287 12189 11299 12192
rect 11241 12183 11299 12189
rect 11698 12180 11704 12192
rect 11756 12180 11762 12232
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 12434 12220 12440 12232
rect 12299 12192 12440 12220
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 12434 12180 12440 12192
rect 12492 12180 12498 12232
rect 14734 12220 14740 12232
rect 13648 12192 14740 12220
rect 8754 12152 8760 12164
rect 8715 12124 8760 12152
rect 8754 12112 8760 12124
rect 8812 12112 8818 12164
rect 9030 12112 9036 12164
rect 9088 12152 9094 12164
rect 9214 12152 9220 12164
rect 9088 12124 9220 12152
rect 9088 12112 9094 12124
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 11974 12152 11980 12164
rect 9968 12124 11980 12152
rect 6270 12044 6276 12096
rect 6328 12084 6334 12096
rect 6914 12084 6920 12096
rect 6328 12056 6920 12084
rect 6328 12044 6334 12056
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 8297 12087 8355 12093
rect 8297 12053 8309 12087
rect 8343 12084 8355 12087
rect 9968 12084 9996 12124
rect 11974 12112 11980 12124
rect 12032 12112 12038 12164
rect 8343 12056 9996 12084
rect 10045 12087 10103 12093
rect 8343 12053 8355 12056
rect 8297 12047 8355 12053
rect 10045 12053 10057 12087
rect 10091 12084 10103 12087
rect 10502 12084 10508 12096
rect 10091 12056 10508 12084
rect 10091 12053 10103 12056
rect 10045 12047 10103 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 10689 12087 10747 12093
rect 10689 12053 10701 12087
rect 10735 12084 10747 12087
rect 13648 12084 13676 12192
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15856 12220 15884 12260
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16574 12288 16580 12300
rect 15979 12260 16580 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16574 12248 16580 12260
rect 16632 12248 16638 12300
rect 16853 12291 16911 12297
rect 16853 12257 16865 12291
rect 16899 12288 16911 12291
rect 17034 12288 17040 12300
rect 16899 12260 17040 12288
rect 16899 12257 16911 12260
rect 16853 12251 16911 12257
rect 17034 12248 17040 12260
rect 17092 12248 17098 12300
rect 17862 12248 17868 12300
rect 17920 12288 17926 12300
rect 18874 12288 18880 12300
rect 17920 12260 18092 12288
rect 18835 12260 18880 12288
rect 17920 12248 17926 12260
rect 16206 12220 16212 12232
rect 15856 12192 16212 12220
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 17126 12220 17132 12232
rect 17087 12192 17132 12220
rect 17126 12180 17132 12192
rect 17184 12180 17190 12232
rect 17954 12220 17960 12232
rect 17915 12192 17960 12220
rect 17954 12180 17960 12192
rect 18012 12180 18018 12232
rect 18064 12229 18092 12260
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 20622 12248 20628 12300
rect 20680 12288 20686 12300
rect 21284 12297 21312 12328
rect 21002 12291 21060 12297
rect 21002 12288 21014 12291
rect 20680 12260 21014 12288
rect 20680 12248 20686 12260
rect 21002 12257 21014 12260
rect 21048 12257 21060 12291
rect 21002 12251 21060 12257
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12257 21327 12291
rect 21269 12251 21327 12257
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12189 18107 12223
rect 18049 12183 18107 12189
rect 18966 12180 18972 12232
rect 19024 12220 19030 12232
rect 19061 12223 19119 12229
rect 19061 12220 19073 12223
rect 19024 12192 19073 12220
rect 19024 12180 19030 12192
rect 19061 12189 19073 12192
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 13722 12112 13728 12164
rect 13780 12152 13786 12164
rect 18782 12152 18788 12164
rect 13780 12124 14688 12152
rect 13780 12112 13786 12124
rect 10735 12056 13676 12084
rect 13909 12087 13967 12093
rect 10735 12053 10747 12056
rect 10689 12047 10747 12053
rect 13909 12053 13921 12087
rect 13955 12084 13967 12087
rect 13998 12084 14004 12096
rect 13955 12056 14004 12084
rect 13955 12053 13967 12056
rect 13909 12047 13967 12053
rect 13998 12044 14004 12056
rect 14056 12044 14062 12096
rect 14660 12084 14688 12124
rect 15948 12124 18788 12152
rect 15948 12084 15976 12124
rect 18782 12112 18788 12124
rect 18840 12112 18846 12164
rect 14660 12056 15976 12084
rect 16574 12044 16580 12096
rect 16632 12084 16638 12096
rect 18509 12087 18567 12093
rect 18509 12084 18521 12087
rect 16632 12056 18521 12084
rect 16632 12044 16638 12056
rect 18509 12053 18521 12056
rect 18555 12053 18567 12087
rect 18509 12047 18567 12053
rect 1104 11994 21896 12016
rect 1104 11942 4447 11994
rect 4499 11942 4511 11994
rect 4563 11942 4575 11994
rect 4627 11942 4639 11994
rect 4691 11942 11378 11994
rect 11430 11942 11442 11994
rect 11494 11942 11506 11994
rect 11558 11942 11570 11994
rect 11622 11942 18308 11994
rect 18360 11942 18372 11994
rect 18424 11942 18436 11994
rect 18488 11942 18500 11994
rect 18552 11942 21896 11994
rect 1104 11920 21896 11942
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9306 11880 9312 11892
rect 8812 11852 9312 11880
rect 8812 11840 8818 11852
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 10042 11880 10048 11892
rect 10003 11852 10048 11880
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10226 11840 10232 11892
rect 10284 11880 10290 11892
rect 11790 11880 11796 11892
rect 10284 11852 11796 11880
rect 10284 11840 10290 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12526 11880 12532 11892
rect 11900 11852 12532 11880
rect 9766 11812 9772 11824
rect 9679 11784 9772 11812
rect 9766 11772 9772 11784
rect 9824 11812 9830 11824
rect 9824 11784 10640 11812
rect 9824 11772 9830 11784
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 10502 11744 10508 11756
rect 10463 11716 10508 11744
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10612 11753 10640 11784
rect 11900 11753 11928 11852
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 13262 11880 13268 11892
rect 13223 11852 13268 11880
rect 13262 11840 13268 11852
rect 13320 11840 13326 11892
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14458 11840 14464 11892
rect 14516 11880 14522 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 14516 11852 16129 11880
rect 14516 11840 14522 11852
rect 16117 11849 16129 11852
rect 16163 11880 16175 11883
rect 16482 11880 16488 11892
rect 16163 11852 16488 11880
rect 16163 11849 16175 11852
rect 16117 11843 16175 11849
rect 16482 11840 16488 11852
rect 16540 11840 16546 11892
rect 17310 11880 17316 11892
rect 17271 11852 17316 11880
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 19886 11880 19892 11892
rect 18340 11852 19892 11880
rect 13814 11772 13820 11824
rect 13872 11812 13878 11824
rect 13872 11784 14320 11812
rect 13872 11772 13878 11784
rect 10597 11747 10655 11753
rect 10597 11713 10609 11747
rect 10643 11713 10655 11747
rect 10597 11707 10655 11713
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 13320 11716 14105 11744
rect 13320 11704 13326 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 14292 11688 14320 11784
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 18340 11812 18368 11852
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 19981 11883 20039 11889
rect 19981 11849 19993 11883
rect 20027 11880 20039 11883
rect 20622 11880 20628 11892
rect 20027 11852 20628 11880
rect 20027 11849 20039 11852
rect 19981 11843 20039 11849
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 16356 11784 18368 11812
rect 16356 11772 16362 11784
rect 14550 11704 14556 11756
rect 14608 11744 14614 11756
rect 14608 11716 14872 11744
rect 14608 11704 14614 11716
rect 8478 11636 8484 11688
rect 8536 11676 8542 11688
rect 8645 11679 8703 11685
rect 8645 11676 8657 11679
rect 8536 11648 8657 11676
rect 8536 11636 8542 11648
rect 8645 11645 8657 11648
rect 8691 11645 8703 11679
rect 8645 11639 8703 11645
rect 9214 11636 9220 11688
rect 9272 11676 9278 11688
rect 10226 11676 10232 11688
rect 9272 11648 10232 11676
rect 9272 11636 9278 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 10962 11676 10968 11688
rect 10336 11648 10968 11676
rect 7374 11568 7380 11620
rect 7432 11608 7438 11620
rect 10336 11608 10364 11648
rect 10962 11636 10968 11648
rect 11020 11636 11026 11688
rect 11974 11636 11980 11688
rect 12032 11676 12038 11688
rect 12032 11648 14136 11676
rect 12032 11636 12038 11648
rect 14108 11620 14136 11648
rect 14274 11636 14280 11688
rect 14332 11636 14338 11688
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 14737 11679 14795 11685
rect 14737 11676 14749 11679
rect 14424 11648 14749 11676
rect 14424 11636 14430 11648
rect 14737 11645 14749 11648
rect 14783 11645 14795 11679
rect 14844 11676 14872 11716
rect 15746 11704 15752 11756
rect 15804 11744 15810 11756
rect 15804 11716 17264 11744
rect 15804 11704 15810 11716
rect 14993 11679 15051 11685
rect 14993 11676 15005 11679
rect 14844 11648 15005 11676
rect 14737 11639 14795 11645
rect 14993 11645 15005 11648
rect 15039 11645 15051 11679
rect 14993 11639 15051 11645
rect 15470 11636 15476 11688
rect 15528 11676 15534 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 15528 11648 17141 11676
rect 15528 11636 15534 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 17236 11676 17264 11716
rect 19352 11716 19840 11744
rect 19352 11688 19380 11716
rect 18598 11676 18604 11688
rect 17236 11648 18604 11676
rect 17129 11639 17187 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 18966 11636 18972 11688
rect 19024 11685 19030 11688
rect 19024 11676 19036 11685
rect 19245 11679 19303 11685
rect 19024 11648 19069 11676
rect 19024 11639 19036 11648
rect 19245 11645 19257 11679
rect 19291 11676 19303 11679
rect 19334 11676 19340 11688
rect 19291 11648 19340 11676
rect 19291 11645 19303 11648
rect 19245 11639 19303 11645
rect 19024 11636 19030 11639
rect 19334 11636 19340 11648
rect 19392 11636 19398 11688
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11645 19763 11679
rect 19812 11676 19840 11716
rect 21361 11679 21419 11685
rect 21361 11676 21373 11679
rect 19812 11648 21373 11676
rect 19705 11639 19763 11645
rect 21361 11645 21373 11648
rect 21407 11645 21419 11679
rect 21361 11639 21419 11645
rect 7432 11580 10364 11608
rect 10413 11611 10471 11617
rect 7432 11568 7438 11580
rect 10413 11577 10425 11611
rect 10459 11608 10471 11611
rect 11057 11611 11115 11617
rect 11057 11608 11069 11611
rect 10459 11580 11069 11608
rect 10459 11577 10471 11580
rect 10413 11571 10471 11577
rect 11057 11577 11069 11580
rect 11103 11577 11115 11611
rect 11057 11571 11115 11577
rect 12152 11611 12210 11617
rect 12152 11577 12164 11611
rect 12198 11608 12210 11611
rect 13078 11608 13084 11620
rect 12198 11580 13084 11608
rect 12198 11577 12210 11580
rect 12152 11571 12210 11577
rect 13078 11568 13084 11580
rect 13136 11608 13142 11620
rect 13814 11608 13820 11620
rect 13136 11580 13820 11608
rect 13136 11568 13142 11580
rect 13814 11568 13820 11580
rect 13872 11568 13878 11620
rect 14090 11568 14096 11620
rect 14148 11568 14154 11620
rect 14642 11568 14648 11620
rect 14700 11608 14706 11620
rect 16393 11611 16451 11617
rect 16393 11608 16405 11611
rect 14700 11580 16405 11608
rect 14700 11568 14706 11580
rect 16393 11577 16405 11580
rect 16439 11577 16451 11611
rect 19720 11608 19748 11639
rect 21174 11617 21180 11620
rect 16393 11571 16451 11577
rect 16684 11580 19748 11608
rect 21116 11611 21180 11617
rect 8113 11543 8171 11549
rect 8113 11509 8125 11543
rect 8159 11540 8171 11543
rect 8202 11540 8208 11552
rect 8159 11512 8208 11540
rect 8159 11509 8171 11512
rect 8113 11503 8171 11509
rect 8202 11500 8208 11512
rect 8260 11500 8266 11552
rect 8846 11500 8852 11552
rect 8904 11540 8910 11552
rect 13630 11540 13636 11552
rect 8904 11512 13636 11540
rect 8904 11500 8910 11512
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13780 11512 13921 11540
rect 13780 11500 13786 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 13909 11503 13967 11509
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 14550 11540 14556 11552
rect 14047 11512 14556 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 15746 11540 15752 11552
rect 14792 11512 15752 11540
rect 14792 11500 14798 11512
rect 15746 11500 15752 11512
rect 15804 11500 15810 11552
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16684 11540 16712 11580
rect 21116 11577 21128 11611
rect 21162 11577 21180 11611
rect 21116 11571 21180 11577
rect 21174 11568 21180 11571
rect 21232 11568 21238 11620
rect 17862 11540 17868 11552
rect 15896 11512 16712 11540
rect 17823 11512 17868 11540
rect 15896 11500 15902 11512
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 19150 11540 19156 11552
rect 18196 11512 19156 11540
rect 18196 11500 18202 11512
rect 19150 11500 19156 11512
rect 19208 11500 19214 11552
rect 19518 11540 19524 11552
rect 19479 11512 19524 11540
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 1104 11450 21896 11472
rect 1104 11398 7912 11450
rect 7964 11398 7976 11450
rect 8028 11398 8040 11450
rect 8092 11398 8104 11450
rect 8156 11398 14843 11450
rect 14895 11398 14907 11450
rect 14959 11398 14971 11450
rect 15023 11398 15035 11450
rect 15087 11398 21896 11450
rect 1104 11376 21896 11398
rect 7101 11339 7159 11345
rect 7101 11305 7113 11339
rect 7147 11336 7159 11339
rect 7374 11336 7380 11348
rect 7147 11308 7380 11336
rect 7147 11305 7159 11308
rect 7101 11299 7159 11305
rect 7374 11296 7380 11308
rect 7432 11296 7438 11348
rect 8202 11336 8208 11348
rect 8115 11308 8208 11336
rect 8128 11209 8156 11308
rect 8202 11296 8208 11308
rect 8260 11336 8266 11348
rect 11606 11336 11612 11348
rect 8260 11308 11612 11336
rect 8260 11296 8266 11308
rect 11606 11296 11612 11308
rect 11664 11296 11670 11348
rect 11701 11339 11759 11345
rect 11701 11305 11713 11339
rect 11747 11336 11759 11339
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 11747 11308 12449 11336
rect 11747 11305 11759 11308
rect 11701 11299 11759 11305
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 13722 11336 13728 11348
rect 13683 11308 13728 11336
rect 12437 11299 12495 11305
rect 13722 11296 13728 11308
rect 13780 11296 13786 11348
rect 14274 11296 14280 11348
rect 14332 11336 14338 11348
rect 16114 11336 16120 11348
rect 14332 11308 16120 11336
rect 14332 11296 14338 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16482 11296 16488 11348
rect 16540 11336 16546 11348
rect 16540 11308 16712 11336
rect 16540 11296 16546 11308
rect 8481 11271 8539 11277
rect 8481 11237 8493 11271
rect 8527 11268 8539 11271
rect 9398 11268 9404 11280
rect 8527 11240 9404 11268
rect 8527 11237 8539 11240
rect 8481 11231 8539 11237
rect 9398 11228 9404 11240
rect 9456 11228 9462 11280
rect 9576 11271 9634 11277
rect 9576 11237 9588 11271
rect 9622 11268 9634 11271
rect 9766 11268 9772 11280
rect 9622 11240 9772 11268
rect 9622 11237 9634 11240
rect 9576 11231 9634 11237
rect 9766 11228 9772 11240
rect 9824 11228 9830 11280
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 13357 11271 13415 11277
rect 13357 11268 13369 11271
rect 12308 11240 13369 11268
rect 12308 11228 12314 11240
rect 13357 11237 13369 11240
rect 13403 11237 13415 11271
rect 16684 11268 16712 11308
rect 17034 11296 17040 11348
rect 17092 11336 17098 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 17092 11308 18521 11336
rect 17092 11296 17098 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 18509 11299 18567 11305
rect 18598 11296 18604 11348
rect 18656 11336 18662 11348
rect 20806 11336 20812 11348
rect 18656 11308 20812 11336
rect 18656 11296 18662 11308
rect 20806 11296 20812 11308
rect 20864 11296 20870 11348
rect 21174 11336 21180 11348
rect 21135 11308 21180 11336
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 16822 11271 16880 11277
rect 16822 11268 16834 11271
rect 16684 11240 16834 11268
rect 13357 11231 13415 11237
rect 16822 11237 16834 11240
rect 16868 11237 16880 11271
rect 20042 11271 20100 11277
rect 20042 11268 20054 11271
rect 16822 11231 16880 11237
rect 18524 11240 20054 11268
rect 8113 11203 8171 11209
rect 8113 11169 8125 11203
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 10778 11200 10784 11212
rect 8619 11172 10784 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 7837 11135 7895 11141
rect 7837 11101 7849 11135
rect 7883 11132 7895 11135
rect 8588 11132 8616 11163
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11020 11172 11253 11200
rect 11020 11160 11026 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 12066 11200 12072 11212
rect 11379 11172 12072 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 12342 11200 12348 11212
rect 12303 11172 12348 11200
rect 12342 11160 12348 11172
rect 12400 11160 12406 11212
rect 13630 11160 13636 11212
rect 13688 11200 13694 11212
rect 14553 11203 14611 11209
rect 14553 11200 14565 11203
rect 13688 11172 14565 11200
rect 13688 11160 13694 11172
rect 14553 11169 14565 11172
rect 14599 11169 14611 11203
rect 16298 11200 16304 11212
rect 16259 11172 16304 11200
rect 14553 11163 14611 11169
rect 16298 11160 16304 11172
rect 16356 11160 16362 11212
rect 17862 11160 17868 11212
rect 17920 11200 17926 11212
rect 18524 11200 18552 11240
rect 20042 11237 20054 11240
rect 20088 11237 20100 11271
rect 20042 11231 20100 11237
rect 17920 11172 18552 11200
rect 17920 11160 17926 11172
rect 18782 11160 18788 11212
rect 18840 11200 18846 11212
rect 18877 11203 18935 11209
rect 18877 11200 18889 11203
rect 18840 11172 18889 11200
rect 18840 11160 18846 11172
rect 18877 11169 18889 11172
rect 18923 11169 18935 11203
rect 18877 11163 18935 11169
rect 18969 11203 19027 11209
rect 18969 11169 18981 11203
rect 19015 11200 19027 11203
rect 19702 11200 19708 11212
rect 19015 11172 19708 11200
rect 19015 11169 19027 11172
rect 18969 11163 19027 11169
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 9030 11132 9036 11144
rect 7883 11104 8616 11132
rect 8680 11104 9036 11132
rect 7883 11101 7895 11104
rect 7837 11095 7895 11101
rect 7469 11067 7527 11073
rect 7469 11033 7481 11067
rect 7515 11064 7527 11067
rect 8297 11067 8355 11073
rect 7515 11036 8248 11064
rect 7515 11033 7527 11036
rect 7469 11027 7527 11033
rect 4798 10956 4804 11008
rect 4856 10996 4862 11008
rect 5626 10996 5632 11008
rect 4856 10968 5632 10996
rect 4856 10956 4862 10968
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 8220 10996 8248 11036
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 8481 11067 8539 11073
rect 8481 11064 8493 11067
rect 8343 11036 8493 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 8481 11033 8493 11036
rect 8527 11033 8539 11067
rect 8680 11064 8708 11104
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 11057 11135 11115 11141
rect 11057 11132 11069 11135
rect 9309 11095 9367 11101
rect 10704 11104 11069 11132
rect 8481 11027 8539 11033
rect 8588 11036 8708 11064
rect 8757 11067 8815 11073
rect 8386 10996 8392 11008
rect 8220 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10996 8450 11008
rect 8588 10996 8616 11036
rect 8757 11033 8769 11067
rect 8803 11064 8815 11067
rect 9214 11064 9220 11076
rect 8803 11036 9220 11064
rect 8803 11033 8815 11036
rect 8757 11027 8815 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 8444 10968 8616 10996
rect 9324 10996 9352 11095
rect 10318 11024 10324 11076
rect 10376 11064 10382 11076
rect 10594 11064 10600 11076
rect 10376 11036 10600 11064
rect 10376 11024 10382 11036
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 10704 11008 10732 11104
rect 11057 11101 11069 11104
rect 11103 11101 11115 11135
rect 11057 11095 11115 11101
rect 12621 11135 12679 11141
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 13078 11132 13084 11144
rect 13039 11104 13084 11132
rect 12621 11095 12679 11101
rect 10870 11024 10876 11076
rect 10928 11064 10934 11076
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 10928 11036 11989 11064
rect 10928 11024 10934 11036
rect 11977 11033 11989 11036
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 9950 10996 9956 11008
rect 9324 10968 9956 10996
rect 8444 10956 8450 10968
rect 9950 10956 9956 10968
rect 10008 10956 10014 11008
rect 10686 10996 10692 11008
rect 10647 10968 10692 10996
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12636 10996 12664 11095
rect 13078 11092 13084 11104
rect 13136 11092 13142 11144
rect 13262 11132 13268 11144
rect 13223 11104 13268 11132
rect 13262 11092 13268 11104
rect 13320 11092 13326 11144
rect 16485 11135 16543 11141
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16531 11104 16589 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 19058 11132 19064 11144
rect 19019 11104 19064 11132
rect 16577 11095 16635 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19797 11135 19855 11141
rect 19797 11132 19809 11135
rect 19392 11104 19809 11132
rect 19392 11092 19398 11104
rect 19797 11101 19809 11104
rect 19843 11101 19855 11135
rect 19797 11095 19855 11101
rect 11756 10968 12664 10996
rect 11756 10956 11762 10968
rect 14366 10956 14372 11008
rect 14424 10996 14430 11008
rect 16485 10999 16543 11005
rect 16485 10996 16497 10999
rect 14424 10968 16497 10996
rect 14424 10956 14430 10968
rect 16485 10965 16497 10968
rect 16531 10965 16543 10999
rect 17954 10996 17960 11008
rect 17915 10968 17960 10996
rect 16485 10959 16543 10965
rect 17954 10956 17960 10968
rect 18012 10956 18018 11008
rect 1104 10906 21896 10928
rect 1104 10854 4447 10906
rect 4499 10854 4511 10906
rect 4563 10854 4575 10906
rect 4627 10854 4639 10906
rect 4691 10854 11378 10906
rect 11430 10854 11442 10906
rect 11494 10854 11506 10906
rect 11558 10854 11570 10906
rect 11622 10854 18308 10906
rect 18360 10854 18372 10906
rect 18424 10854 18436 10906
rect 18488 10854 18500 10906
rect 18552 10854 21896 10906
rect 1104 10832 21896 10854
rect 1762 10752 1768 10804
rect 1820 10792 1826 10804
rect 7374 10792 7380 10804
rect 1820 10764 7380 10792
rect 1820 10752 1826 10764
rect 7374 10752 7380 10764
rect 7432 10752 7438 10804
rect 8665 10795 8723 10801
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 12250 10792 12256 10804
rect 8711 10764 12256 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 12250 10752 12256 10764
rect 12308 10752 12314 10804
rect 13173 10795 13231 10801
rect 13173 10761 13185 10795
rect 13219 10792 13231 10795
rect 13262 10792 13268 10804
rect 13219 10764 13268 10792
rect 13219 10761 13231 10764
rect 13173 10755 13231 10761
rect 13262 10752 13268 10764
rect 13320 10752 13326 10804
rect 13906 10752 13912 10804
rect 13964 10792 13970 10804
rect 14737 10795 14795 10801
rect 14737 10792 14749 10795
rect 13964 10764 14749 10792
rect 13964 10752 13970 10764
rect 14737 10761 14749 10764
rect 14783 10761 14795 10795
rect 17862 10792 17868 10804
rect 14737 10755 14795 10761
rect 16040 10764 17868 10792
rect 10870 10684 10876 10736
rect 10928 10724 10934 10736
rect 15838 10724 15844 10736
rect 10928 10696 15844 10724
rect 10928 10684 10934 10696
rect 15838 10684 15844 10696
rect 15896 10684 15902 10736
rect 12069 10659 12127 10665
rect 12069 10625 12081 10659
rect 12115 10656 12127 10659
rect 12342 10656 12348 10668
rect 12115 10628 12348 10656
rect 12115 10625 12127 10628
rect 12069 10619 12127 10625
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 12618 10656 12624 10668
rect 12531 10628 12624 10656
rect 12618 10616 12624 10628
rect 12676 10656 12682 10668
rect 13541 10659 13599 10665
rect 13541 10656 13553 10659
rect 12676 10628 13553 10656
rect 12676 10616 12682 10628
rect 13541 10625 13553 10628
rect 13587 10625 13599 10659
rect 13998 10656 14004 10668
rect 13541 10619 13599 10625
rect 13648 10628 14004 10656
rect 8481 10591 8539 10597
rect 8481 10557 8493 10591
rect 8527 10588 8539 10591
rect 8570 10588 8576 10600
rect 8527 10560 8576 10588
rect 8527 10557 8539 10560
rect 8481 10551 8539 10557
rect 8570 10548 8576 10560
rect 8628 10548 8634 10600
rect 8846 10548 8852 10600
rect 8904 10588 8910 10600
rect 8941 10591 8999 10597
rect 8941 10588 8953 10591
rect 8904 10560 8953 10588
rect 8904 10548 8910 10560
rect 8941 10557 8953 10560
rect 8987 10557 8999 10591
rect 8941 10551 8999 10557
rect 9401 10591 9459 10597
rect 9401 10557 9413 10591
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 9861 10591 9919 10597
rect 9861 10557 9873 10591
rect 9907 10588 9919 10591
rect 9950 10588 9956 10600
rect 9907 10560 9956 10588
rect 9907 10557 9919 10560
rect 9861 10551 9919 10557
rect 8205 10523 8263 10529
rect 8205 10489 8217 10523
rect 8251 10520 8263 10523
rect 9416 10520 9444 10551
rect 9950 10548 9956 10560
rect 10008 10548 10014 10600
rect 10128 10591 10186 10597
rect 10128 10557 10140 10591
rect 10174 10588 10186 10591
rect 10686 10588 10692 10600
rect 10174 10560 10692 10588
rect 10174 10557 10186 10560
rect 10128 10551 10186 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 13648 10588 13676 10628
rect 13998 10616 14004 10628
rect 14056 10656 14062 10668
rect 16040 10665 16068 10764
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 18877 10795 18935 10801
rect 18877 10761 18889 10795
rect 18923 10792 18935 10795
rect 18966 10792 18972 10804
rect 18923 10764 18972 10792
rect 18923 10761 18935 10764
rect 18877 10755 18935 10761
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 20533 10795 20591 10801
rect 20533 10761 20545 10795
rect 20579 10792 20591 10795
rect 20898 10792 20904 10804
rect 20579 10764 20904 10792
rect 20579 10761 20591 10764
rect 20533 10755 20591 10761
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 16577 10727 16635 10733
rect 16577 10693 16589 10727
rect 16623 10724 16635 10727
rect 18782 10724 18788 10736
rect 16623 10696 18788 10724
rect 16623 10693 16635 10696
rect 16577 10687 16635 10693
rect 18782 10684 18788 10696
rect 18840 10684 18846 10736
rect 15289 10659 15347 10665
rect 15289 10656 15301 10659
rect 14056 10628 15301 10656
rect 14056 10616 14062 10628
rect 15289 10625 15301 10628
rect 15335 10625 15347 10659
rect 15289 10619 15347 10625
rect 16025 10659 16083 10665
rect 16025 10625 16037 10659
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 17034 10656 17040 10668
rect 16163 10628 17040 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 17034 10616 17040 10628
rect 17092 10616 17098 10668
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10625 17279 10659
rect 17402 10656 17408 10668
rect 17363 10628 17408 10656
rect 17221 10619 17279 10625
rect 11112 10560 13676 10588
rect 13725 10591 13783 10597
rect 11112 10548 11118 10560
rect 13725 10557 13737 10591
rect 13771 10588 13783 10591
rect 13814 10588 13820 10600
rect 13771 10560 13820 10588
rect 13771 10557 13783 10560
rect 13725 10551 13783 10557
rect 13814 10548 13820 10560
rect 13872 10548 13878 10600
rect 14642 10548 14648 10600
rect 14700 10588 14706 10600
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 14700 10560 15209 10588
rect 14700 10548 14706 10560
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10588 16267 10591
rect 16574 10588 16580 10600
rect 16255 10560 16580 10588
rect 16255 10557 16267 10560
rect 16209 10551 16267 10557
rect 16574 10548 16580 10560
rect 16632 10548 16638 10600
rect 17236 10588 17264 10619
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 18874 10656 18880 10668
rect 18647 10628 18880 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 21174 10656 21180 10668
rect 21135 10628 21180 10656
rect 21174 10616 21180 10628
rect 21232 10616 21238 10668
rect 17310 10588 17316 10600
rect 17236 10560 17316 10588
rect 17310 10548 17316 10560
rect 17368 10548 17374 10600
rect 20257 10591 20315 10597
rect 20257 10588 20269 10591
rect 19352 10560 20269 10588
rect 19352 10532 19380 10560
rect 20257 10557 20269 10560
rect 20303 10557 20315 10591
rect 20257 10551 20315 10557
rect 15286 10520 15292 10532
rect 8251 10492 15292 10520
rect 8251 10489 8263 10492
rect 8205 10483 8263 10489
rect 15286 10480 15292 10492
rect 15344 10480 15350 10532
rect 19334 10480 19340 10532
rect 19392 10480 19398 10532
rect 20012 10523 20070 10529
rect 20012 10489 20024 10523
rect 20058 10520 20070 10523
rect 20346 10520 20352 10532
rect 20058 10492 20352 10520
rect 20058 10489 20070 10492
rect 20012 10483 20070 10489
rect 20346 10480 20352 10492
rect 20404 10480 20410 10532
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 4304 10424 7757 10452
rect 4304 10412 4310 10424
rect 7745 10421 7757 10424
rect 7791 10452 7803 10455
rect 8846 10452 8852 10464
rect 7791 10424 8852 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9122 10452 9128 10464
rect 9083 10424 9128 10452
rect 9122 10412 9128 10424
rect 9180 10412 9186 10464
rect 9582 10452 9588 10464
rect 9543 10424 9588 10452
rect 9582 10412 9588 10424
rect 9640 10412 9646 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 11054 10452 11060 10464
rect 9916 10424 11060 10452
rect 9916 10412 9922 10424
rect 11054 10412 11060 10424
rect 11112 10412 11118 10464
rect 11241 10455 11299 10461
rect 11241 10421 11253 10455
rect 11287 10452 11299 10455
rect 11698 10452 11704 10464
rect 11287 10424 11704 10452
rect 11287 10421 11299 10424
rect 11241 10415 11299 10421
rect 11698 10412 11704 10424
rect 11756 10412 11762 10464
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 12710 10452 12716 10464
rect 12492 10424 12716 10452
rect 12492 10412 12498 10424
rect 12710 10412 12716 10424
rect 12768 10412 12774 10464
rect 12802 10412 12808 10464
rect 12860 10452 12866 10464
rect 13817 10455 13875 10461
rect 12860 10424 12905 10452
rect 12860 10412 12866 10424
rect 13817 10421 13829 10455
rect 13863 10452 13875 10455
rect 13998 10452 14004 10464
rect 13863 10424 14004 10452
rect 13863 10421 13875 10424
rect 13817 10415 13875 10421
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 14182 10452 14188 10464
rect 14143 10424 14188 10452
rect 14182 10412 14188 10424
rect 14240 10412 14246 10464
rect 14734 10412 14740 10464
rect 14792 10452 14798 10464
rect 15105 10455 15163 10461
rect 15105 10452 15117 10455
rect 14792 10424 15117 10452
rect 14792 10412 14798 10424
rect 15105 10421 15117 10424
rect 15151 10421 15163 10455
rect 15105 10415 15163 10421
rect 16666 10412 16672 10464
rect 16724 10452 16730 10464
rect 17497 10455 17555 10461
rect 17497 10452 17509 10455
rect 16724 10424 17509 10452
rect 16724 10412 16730 10424
rect 17497 10421 17509 10424
rect 17543 10421 17555 10455
rect 17497 10415 17555 10421
rect 17865 10455 17923 10461
rect 17865 10421 17877 10455
rect 17911 10452 17923 10455
rect 18230 10452 18236 10464
rect 17911 10424 18236 10452
rect 17911 10421 17923 10424
rect 17865 10415 17923 10421
rect 18230 10412 18236 10424
rect 18288 10412 18294 10464
rect 20898 10452 20904 10464
rect 20859 10424 20904 10452
rect 20898 10412 20904 10424
rect 20956 10412 20962 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21082 10452 21088 10464
rect 21039 10424 21088 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 1104 10362 21896 10384
rect 1104 10310 7912 10362
rect 7964 10310 7976 10362
rect 8028 10310 8040 10362
rect 8092 10310 8104 10362
rect 8156 10310 14843 10362
rect 14895 10310 14907 10362
rect 14959 10310 14971 10362
rect 15023 10310 15035 10362
rect 15087 10310 21896 10362
rect 1104 10288 21896 10310
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 8846 10248 8852 10260
rect 8444 10220 8852 10248
rect 8444 10208 8450 10220
rect 8846 10208 8852 10220
rect 8904 10208 8910 10260
rect 9217 10251 9275 10257
rect 9217 10217 9229 10251
rect 9263 10248 9275 10251
rect 10045 10251 10103 10257
rect 10045 10248 10057 10251
rect 9263 10220 10057 10248
rect 9263 10217 9275 10220
rect 9217 10211 9275 10217
rect 10045 10217 10057 10220
rect 10091 10217 10103 10251
rect 10045 10211 10103 10217
rect 10137 10251 10195 10257
rect 10137 10217 10149 10251
rect 10183 10248 10195 10251
rect 10410 10248 10416 10260
rect 10183 10220 10416 10248
rect 10183 10217 10195 10220
rect 10137 10211 10195 10217
rect 10410 10208 10416 10220
rect 10468 10208 10474 10260
rect 10505 10251 10563 10257
rect 10505 10217 10517 10251
rect 10551 10217 10563 10251
rect 10505 10211 10563 10217
rect 10689 10251 10747 10257
rect 10689 10217 10701 10251
rect 10735 10248 10747 10251
rect 12161 10251 12219 10257
rect 10735 10220 12020 10248
rect 10735 10217 10747 10220
rect 10689 10211 10747 10217
rect 9122 10140 9128 10192
rect 9180 10180 9186 10192
rect 10520 10180 10548 10211
rect 11992 10180 12020 10220
rect 12161 10217 12173 10251
rect 12207 10248 12219 10251
rect 13817 10251 13875 10257
rect 12207 10220 12434 10248
rect 12207 10217 12219 10220
rect 12161 10211 12219 10217
rect 12253 10183 12311 10189
rect 12253 10180 12265 10183
rect 9180 10152 10272 10180
rect 10520 10152 11928 10180
rect 11992 10152 12265 10180
rect 9180 10140 9186 10152
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8803 10084 9321 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 9309 10081 9321 10084
rect 9355 10112 9367 10115
rect 10244 10112 10272 10152
rect 10870 10112 10876 10124
rect 9355 10084 9996 10112
rect 10244 10084 10876 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 8297 9911 8355 9917
rect 8297 9908 8309 9911
rect 4856 9880 8309 9908
rect 4856 9868 4862 9880
rect 8297 9877 8309 9880
rect 8343 9908 8355 9911
rect 9217 9911 9275 9917
rect 9217 9908 9229 9911
rect 8343 9880 9229 9908
rect 8343 9877 8355 9880
rect 8297 9871 8355 9877
rect 9217 9877 9229 9880
rect 9263 9877 9275 9911
rect 9490 9908 9496 9920
rect 9451 9880 9496 9908
rect 9217 9871 9275 9877
rect 9490 9868 9496 9880
rect 9548 9868 9554 9920
rect 9968 9908 9996 10084
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 11054 10121 11060 10124
rect 11048 10075 11060 10121
rect 11112 10112 11118 10124
rect 11790 10112 11796 10124
rect 11112 10084 11796 10112
rect 11054 10072 11060 10075
rect 11112 10072 11118 10084
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 11900 10112 11928 10152
rect 12253 10149 12265 10152
rect 12299 10149 12311 10183
rect 12406 10180 12434 10220
rect 13817 10217 13829 10251
rect 13863 10248 13875 10251
rect 13906 10248 13912 10260
rect 13863 10220 13912 10248
rect 13863 10217 13875 10220
rect 13817 10211 13875 10217
rect 13906 10208 13912 10220
rect 13964 10208 13970 10260
rect 14182 10208 14188 10260
rect 14240 10248 14246 10260
rect 14921 10251 14979 10257
rect 14921 10248 14933 10251
rect 14240 10220 14933 10248
rect 14240 10208 14246 10220
rect 14921 10217 14933 10220
rect 14967 10217 14979 10251
rect 15930 10248 15936 10260
rect 15891 10220 15936 10248
rect 14921 10211 14979 10217
rect 15930 10208 15936 10220
rect 15988 10208 15994 10260
rect 16117 10251 16175 10257
rect 16117 10217 16129 10251
rect 16163 10248 16175 10251
rect 18230 10248 18236 10260
rect 16163 10220 17908 10248
rect 18191 10220 18236 10248
rect 16163 10217 16175 10220
rect 16117 10211 16175 10217
rect 12618 10180 12624 10192
rect 12406 10152 12624 10180
rect 12253 10143 12311 10149
rect 12618 10140 12624 10152
rect 12676 10189 12682 10192
rect 12676 10183 12740 10189
rect 12676 10149 12694 10183
rect 12728 10180 12740 10183
rect 12728 10152 12769 10180
rect 12728 10149 12740 10152
rect 12676 10143 12740 10149
rect 12676 10140 12682 10143
rect 12986 10112 12992 10124
rect 11900 10084 12992 10112
rect 12986 10072 12992 10084
rect 13044 10072 13050 10124
rect 13924 10112 13952 10208
rect 14366 10140 14372 10192
rect 14424 10180 14430 10192
rect 17681 10183 17739 10189
rect 17681 10180 17693 10183
rect 14424 10152 15700 10180
rect 14424 10140 14430 10152
rect 13924 10084 15148 10112
rect 10042 10004 10048 10056
rect 10100 10044 10106 10056
rect 10686 10044 10692 10056
rect 10100 10016 10692 10044
rect 10100 10004 10106 10016
rect 10686 10004 10692 10016
rect 10744 10044 10750 10056
rect 10781 10047 10839 10053
rect 10781 10044 10793 10047
rect 10744 10016 10793 10044
rect 10744 10004 10750 10016
rect 10781 10013 10793 10016
rect 10827 10013 10839 10047
rect 10781 10007 10839 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10044 12311 10047
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 12299 10016 12449 10044
rect 12299 10013 12311 10016
rect 12253 10007 12311 10013
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 13538 10004 13544 10056
rect 13596 10044 13602 10056
rect 15010 10044 15016 10056
rect 13596 10016 14872 10044
rect 14971 10016 15016 10044
rect 13596 10004 13602 10016
rect 14550 9976 14556 9988
rect 13740 9948 13952 9976
rect 14511 9948 14556 9976
rect 13740 9908 13768 9948
rect 9968 9880 13768 9908
rect 13924 9908 13952 9948
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 14844 9976 14872 10016
rect 15010 10004 15016 10016
rect 15068 10004 15074 10056
rect 15120 10053 15148 10084
rect 15105 10047 15163 10053
rect 15105 10013 15117 10047
rect 15151 10013 15163 10047
rect 15672 10044 15700 10152
rect 15764 10152 17693 10180
rect 15764 10121 15792 10152
rect 17681 10149 17693 10152
rect 17727 10149 17739 10183
rect 17880 10180 17908 10220
rect 18230 10208 18236 10220
rect 18288 10208 18294 10260
rect 18690 10208 18696 10260
rect 18748 10248 18754 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 18748 10220 18889 10248
rect 18748 10208 18754 10220
rect 18877 10217 18889 10220
rect 18923 10217 18935 10251
rect 18877 10211 18935 10217
rect 19702 10208 19708 10260
rect 19760 10248 19766 10260
rect 19797 10251 19855 10257
rect 19797 10248 19809 10251
rect 19760 10220 19809 10248
rect 19760 10208 19766 10220
rect 19797 10217 19809 10220
rect 19843 10217 19855 10251
rect 20990 10248 20996 10260
rect 20951 10220 20996 10248
rect 19797 10211 19855 10217
rect 20990 10208 20996 10220
rect 21048 10208 21054 10260
rect 20162 10180 20168 10192
rect 17880 10152 20168 10180
rect 17681 10143 17739 10149
rect 20162 10140 20168 10152
rect 20220 10140 20226 10192
rect 15749 10115 15807 10121
rect 15749 10081 15761 10115
rect 15795 10081 15807 10115
rect 15749 10075 15807 10081
rect 16476 10115 16534 10121
rect 16476 10081 16488 10115
rect 16522 10112 16534 10115
rect 17954 10112 17960 10124
rect 16522 10084 17960 10112
rect 16522 10081 16534 10084
rect 16476 10075 16534 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 19061 10115 19119 10121
rect 19061 10112 19073 10115
rect 18840 10084 19073 10112
rect 18840 10072 18846 10084
rect 19061 10081 19073 10084
rect 19107 10081 19119 10115
rect 20806 10112 20812 10124
rect 20767 10084 20812 10112
rect 19061 10075 19119 10081
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 16022 10044 16028 10056
rect 15672 10016 16028 10044
rect 15105 10007 15163 10013
rect 16022 10004 16028 10016
rect 16080 10044 16086 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 16080 10016 16221 10044
rect 16080 10004 16086 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18325 10047 18383 10053
rect 18325 10044 18337 10047
rect 18196 10016 18337 10044
rect 18196 10004 18202 10016
rect 18325 10013 18337 10016
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18509 10047 18567 10053
rect 18509 10013 18521 10047
rect 18555 10044 18567 10047
rect 18598 10044 18604 10056
rect 18555 10016 18604 10044
rect 18555 10013 18567 10016
rect 18509 10007 18567 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 20254 10044 20260 10056
rect 20215 10016 20260 10044
rect 20254 10004 20260 10016
rect 20312 10004 20318 10056
rect 20346 10004 20352 10056
rect 20404 10044 20410 10056
rect 20404 10016 20449 10044
rect 20404 10004 20410 10016
rect 16117 9979 16175 9985
rect 16117 9976 16129 9979
rect 14844 9948 16129 9976
rect 16117 9945 16129 9948
rect 16163 9945 16175 9979
rect 17954 9976 17960 9988
rect 16117 9939 16175 9945
rect 17328 9948 17960 9976
rect 17328 9908 17356 9948
rect 17954 9936 17960 9948
rect 18012 9936 18018 9988
rect 13924 9880 17356 9908
rect 17402 9868 17408 9920
rect 17460 9908 17466 9920
rect 17589 9911 17647 9917
rect 17589 9908 17601 9911
rect 17460 9880 17601 9908
rect 17460 9868 17466 9880
rect 17589 9877 17601 9880
rect 17635 9877 17647 9911
rect 17589 9871 17647 9877
rect 17681 9911 17739 9917
rect 17681 9877 17693 9911
rect 17727 9908 17739 9911
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17727 9880 17877 9908
rect 17727 9877 17739 9880
rect 17681 9871 17739 9877
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 21266 9908 21272 9920
rect 21227 9880 21272 9908
rect 17865 9871 17923 9877
rect 21266 9868 21272 9880
rect 21324 9868 21330 9920
rect 1104 9818 21896 9840
rect 1104 9766 4447 9818
rect 4499 9766 4511 9818
rect 4563 9766 4575 9818
rect 4627 9766 4639 9818
rect 4691 9766 11378 9818
rect 11430 9766 11442 9818
rect 11494 9766 11506 9818
rect 11558 9766 11570 9818
rect 11622 9766 18308 9818
rect 18360 9766 18372 9818
rect 18424 9766 18436 9818
rect 18488 9766 18500 9818
rect 18552 9766 21896 9818
rect 1104 9744 21896 9766
rect 7374 9664 7380 9716
rect 7432 9704 7438 9716
rect 8021 9707 8079 9713
rect 8021 9704 8033 9707
rect 7432 9676 8033 9704
rect 7432 9664 7438 9676
rect 8021 9673 8033 9676
rect 8067 9673 8079 9707
rect 8021 9667 8079 9673
rect 9490 9664 9496 9716
rect 9548 9704 9554 9716
rect 13538 9704 13544 9716
rect 9548 9676 13544 9704
rect 9548 9664 9554 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 14642 9704 14648 9716
rect 13648 9676 14648 9704
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 9677 9639 9735 9645
rect 9677 9636 9689 9639
rect 9640 9608 9689 9636
rect 9640 9596 9646 9608
rect 9677 9605 9689 9608
rect 9723 9605 9735 9639
rect 9677 9599 9735 9605
rect 10137 9639 10195 9645
rect 10137 9605 10149 9639
rect 10183 9605 10195 9639
rect 11885 9639 11943 9645
rect 11885 9636 11897 9639
rect 10137 9599 10195 9605
rect 10888 9608 11897 9636
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10152 9568 10180 9599
rect 10100 9540 10180 9568
rect 10100 9528 10106 9540
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10505 9571 10563 9577
rect 10505 9568 10517 9571
rect 10376 9540 10517 9568
rect 10376 9528 10382 9540
rect 10505 9537 10517 9540
rect 10551 9537 10563 9571
rect 10505 9531 10563 9537
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9490 9500 9496 9512
rect 9263 9472 9496 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 9674 9460 9680 9512
rect 9732 9500 9738 9512
rect 9858 9500 9864 9512
rect 9732 9472 9864 9500
rect 9732 9460 9738 9472
rect 9858 9460 9864 9472
rect 9916 9460 9922 9512
rect 9953 9503 10011 9509
rect 9953 9469 9965 9503
rect 9999 9500 10011 9503
rect 10888 9500 10916 9608
rect 11885 9605 11897 9608
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 13262 9596 13268 9648
rect 13320 9636 13326 9648
rect 13648 9636 13676 9676
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 16022 9664 16028 9716
rect 16080 9704 16086 9716
rect 18509 9707 18567 9713
rect 16080 9676 17080 9704
rect 16080 9664 16086 9676
rect 13320 9608 13676 9636
rect 13725 9639 13783 9645
rect 13320 9596 13326 9608
rect 13725 9605 13737 9639
rect 13771 9636 13783 9639
rect 15010 9636 15016 9648
rect 13771 9608 15016 9636
rect 13771 9605 13783 9608
rect 13725 9599 13783 9605
rect 15010 9596 15016 9608
rect 15068 9596 15074 9648
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12618 9528 12624 9580
rect 12676 9568 12682 9580
rect 13081 9571 13139 9577
rect 13081 9568 13093 9571
rect 12676 9540 13093 9568
rect 12676 9528 12682 9540
rect 13081 9537 13093 9540
rect 13127 9537 13139 9571
rect 13081 9531 13139 9537
rect 13909 9571 13967 9577
rect 13909 9537 13921 9571
rect 13955 9568 13967 9571
rect 14550 9568 14556 9580
rect 13955 9540 14556 9568
rect 13955 9537 13967 9540
rect 13909 9531 13967 9537
rect 14550 9528 14556 9540
rect 14608 9528 14614 9580
rect 15378 9528 15384 9580
rect 15436 9568 15442 9580
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15436 9540 15577 9568
rect 15436 9528 15442 9540
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 16577 9571 16635 9577
rect 16577 9537 16589 9571
rect 16623 9568 16635 9571
rect 16666 9568 16672 9580
rect 16623 9540 16672 9568
rect 16623 9537 16635 9540
rect 16577 9531 16635 9537
rect 16666 9528 16672 9540
rect 16724 9528 16730 9580
rect 17052 9568 17080 9676
rect 18509 9673 18521 9707
rect 18555 9704 18567 9707
rect 18598 9704 18604 9716
rect 18555 9676 18604 9704
rect 18555 9673 18567 9676
rect 18509 9667 18567 9673
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 20165 9707 20223 9713
rect 20165 9673 20177 9707
rect 20211 9704 20223 9707
rect 20346 9704 20352 9716
rect 20211 9676 20352 9704
rect 20211 9673 20223 9676
rect 20165 9667 20223 9673
rect 20346 9664 20352 9676
rect 20404 9664 20410 9716
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 17052 9540 17141 9568
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 18616 9568 18644 9664
rect 20990 9568 20996 9580
rect 18616 9540 18920 9568
rect 20951 9540 20996 9568
rect 17129 9531 17187 9537
rect 9999 9472 10916 9500
rect 11793 9503 11851 9509
rect 9999 9469 10011 9472
rect 9953 9463 10011 9469
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12253 9503 12311 9509
rect 12253 9500 12265 9503
rect 11839 9472 12265 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12253 9469 12265 9472
rect 12299 9469 12311 9503
rect 17034 9500 17040 9512
rect 12253 9463 12311 9469
rect 12360 9472 17040 9500
rect 9398 9392 9404 9444
rect 9456 9432 9462 9444
rect 12360 9432 12388 9472
rect 17034 9460 17040 9472
rect 17092 9460 17098 9512
rect 17144 9500 17172 9531
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 17144 9472 18797 9500
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 18892 9500 18920 9540
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 19041 9503 19099 9509
rect 19041 9500 19053 9503
rect 18892 9472 19053 9500
rect 18785 9463 18843 9469
rect 19041 9469 19053 9472
rect 19087 9469 19099 9503
rect 19041 9463 19099 9469
rect 9456 9404 12388 9432
rect 9456 9392 9462 9404
rect 12434 9392 12440 9444
rect 12492 9432 12498 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 12492 9404 13921 9432
rect 12492 9392 12498 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14369 9435 14427 9441
rect 14369 9401 14381 9435
rect 14415 9432 14427 9435
rect 14415 9404 15056 9432
rect 14415 9401 14427 9404
rect 14369 9395 14427 9401
rect 8386 9364 8392 9376
rect 8347 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8662 9324 8668 9376
rect 8720 9364 8726 9376
rect 8849 9367 8907 9373
rect 8849 9364 8861 9367
rect 8720 9336 8861 9364
rect 8720 9324 8726 9336
rect 8849 9333 8861 9336
rect 8895 9364 8907 9367
rect 9030 9364 9036 9376
rect 8895 9336 9036 9364
rect 8895 9333 8907 9336
rect 8849 9327 8907 9333
rect 9030 9324 9036 9336
rect 9088 9364 9094 9376
rect 10689 9367 10747 9373
rect 10689 9364 10701 9367
rect 9088 9336 10701 9364
rect 9088 9324 9094 9336
rect 10689 9333 10701 9336
rect 10735 9333 10747 9367
rect 10689 9327 10747 9333
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11149 9367 11207 9373
rect 10836 9336 10881 9364
rect 10836 9324 10842 9336
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11793 9367 11851 9373
rect 11793 9364 11805 9367
rect 11195 9336 11805 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11793 9333 11805 9336
rect 11839 9333 11851 9367
rect 11793 9327 11851 9333
rect 12066 9324 12072 9376
rect 12124 9364 12130 9376
rect 12345 9367 12403 9373
rect 12345 9364 12357 9367
rect 12124 9336 12357 9364
rect 12124 9324 12130 9336
rect 12345 9333 12357 9336
rect 12391 9333 12403 9367
rect 12345 9327 12403 9333
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 13262 9364 13268 9376
rect 12584 9336 13268 9364
rect 12584 9324 12590 9336
rect 13262 9324 13268 9336
rect 13320 9324 13326 9376
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13998 9364 14004 9376
rect 13412 9336 13457 9364
rect 13959 9336 14004 9364
rect 13412 9324 13418 9336
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 14274 9324 14280 9376
rect 14332 9364 14338 9376
rect 15028 9373 15056 9404
rect 15102 9392 15108 9444
rect 15160 9432 15166 9444
rect 17402 9441 17408 9444
rect 15473 9435 15531 9441
rect 15473 9432 15485 9435
rect 15160 9404 15485 9432
rect 15160 9392 15166 9404
rect 15473 9401 15485 9404
rect 15519 9401 15531 9435
rect 17396 9432 17408 9441
rect 17363 9404 17408 9432
rect 15473 9395 15531 9401
rect 17396 9395 17408 9404
rect 17402 9392 17408 9395
rect 17460 9392 17466 9444
rect 18800 9432 18828 9463
rect 20162 9460 20168 9512
rect 20220 9500 20226 9512
rect 20901 9503 20959 9509
rect 20901 9500 20913 9503
rect 20220 9472 20913 9500
rect 20220 9460 20226 9472
rect 20901 9469 20913 9472
rect 20947 9469 20959 9503
rect 20901 9463 20959 9469
rect 19334 9432 19340 9444
rect 18800 9404 19340 9432
rect 19334 9392 19340 9404
rect 19392 9392 19398 9444
rect 14461 9367 14519 9373
rect 14461 9364 14473 9367
rect 14332 9336 14473 9364
rect 14332 9324 14338 9336
rect 14461 9333 14473 9336
rect 14507 9333 14519 9367
rect 14461 9327 14519 9333
rect 15013 9367 15071 9373
rect 15013 9333 15025 9367
rect 15059 9333 15071 9367
rect 15013 9327 15071 9333
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15381 9367 15439 9373
rect 15381 9364 15393 9367
rect 15344 9336 15393 9364
rect 15344 9324 15350 9336
rect 15381 9333 15393 9336
rect 15427 9364 15439 9367
rect 15654 9364 15660 9376
rect 15427 9336 15660 9364
rect 15427 9333 15439 9336
rect 15381 9327 15439 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 16114 9364 16120 9376
rect 16075 9336 16120 9364
rect 16114 9324 16120 9336
rect 16172 9324 16178 9376
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16942 9364 16948 9376
rect 16632 9336 16948 9364
rect 16632 9324 16638 9336
rect 16942 9324 16948 9336
rect 17000 9324 17006 9376
rect 19150 9324 19156 9376
rect 19208 9364 19214 9376
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 19208 9336 20453 9364
rect 19208 9324 19214 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 20806 9364 20812 9376
rect 20767 9336 20812 9364
rect 20441 9327 20499 9333
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 1104 9274 21896 9296
rect 1104 9222 7912 9274
rect 7964 9222 7976 9274
rect 8028 9222 8040 9274
rect 8092 9222 8104 9274
rect 8156 9222 14843 9274
rect 14895 9222 14907 9274
rect 14959 9222 14971 9274
rect 15023 9222 15035 9274
rect 15087 9222 21896 9274
rect 1104 9200 21896 9222
rect 9490 9120 9496 9172
rect 9548 9160 9554 9172
rect 10870 9160 10876 9172
rect 9548 9132 10876 9160
rect 9548 9120 9554 9132
rect 10870 9120 10876 9132
rect 10928 9120 10934 9172
rect 11054 9160 11060 9172
rect 11015 9132 11060 9160
rect 11054 9120 11060 9132
rect 11112 9120 11118 9172
rect 11146 9120 11152 9172
rect 11204 9160 11210 9172
rect 11790 9160 11796 9172
rect 11204 9132 11796 9160
rect 11204 9120 11210 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 12066 9160 12072 9172
rect 12027 9132 12072 9160
rect 12066 9120 12072 9132
rect 12124 9120 12130 9172
rect 13633 9163 13691 9169
rect 13633 9129 13645 9163
rect 13679 9160 13691 9163
rect 13998 9160 14004 9172
rect 13679 9132 14004 9160
rect 13679 9129 13691 9132
rect 13633 9123 13691 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 15933 9163 15991 9169
rect 15933 9160 15945 9163
rect 14608 9132 15945 9160
rect 14608 9120 14614 9132
rect 15933 9129 15945 9132
rect 15979 9160 15991 9163
rect 16117 9163 16175 9169
rect 16117 9160 16129 9163
rect 15979 9132 16129 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16117 9129 16129 9132
rect 16163 9129 16175 9163
rect 16117 9123 16175 9129
rect 16209 9163 16267 9169
rect 16209 9129 16221 9163
rect 16255 9129 16267 9163
rect 16209 9123 16267 9129
rect 6362 9052 6368 9104
rect 6420 9092 6426 9104
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 6420 9064 8309 9092
rect 6420 9052 6426 9064
rect 8297 9061 8309 9064
rect 8343 9092 8355 9095
rect 9398 9092 9404 9104
rect 8343 9064 9404 9092
rect 8343 9061 8355 9064
rect 8297 9055 8355 9061
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 10686 9092 10692 9104
rect 9508 9064 10692 9092
rect 6270 8984 6276 9036
rect 6328 9024 6334 9036
rect 7190 9024 7196 9036
rect 6328 8996 7196 9024
rect 6328 8984 6334 8996
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 8757 9027 8815 9033
rect 8757 8993 8769 9027
rect 8803 9024 8815 9027
rect 9122 9024 9128 9036
rect 8803 8996 9128 9024
rect 8803 8993 8815 8996
rect 8757 8987 8815 8993
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 7466 8916 7472 8968
rect 7524 8956 7530 8968
rect 7650 8956 7656 8968
rect 7524 8928 7656 8956
rect 7524 8916 7530 8928
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9508 8956 9536 9064
rect 10686 9052 10692 9064
rect 10744 9052 10750 9104
rect 10778 9052 10784 9104
rect 10836 9092 10842 9104
rect 12345 9095 12403 9101
rect 12345 9092 12357 9095
rect 10836 9064 12357 9092
rect 10836 9052 10842 9064
rect 12345 9061 12357 9064
rect 12391 9061 12403 9095
rect 12345 9055 12403 9061
rect 13541 9095 13599 9101
rect 13541 9061 13553 9095
rect 13587 9092 13599 9095
rect 16224 9092 16252 9123
rect 16298 9120 16304 9172
rect 16356 9160 16362 9172
rect 16669 9163 16727 9169
rect 16669 9160 16681 9163
rect 16356 9132 16681 9160
rect 16356 9120 16362 9132
rect 16669 9129 16681 9132
rect 16715 9129 16727 9163
rect 17494 9160 17500 9172
rect 17455 9132 17500 9160
rect 16669 9123 16727 9129
rect 17494 9120 17500 9132
rect 17552 9120 17558 9172
rect 17957 9163 18015 9169
rect 17957 9129 17969 9163
rect 18003 9129 18015 9163
rect 17957 9123 18015 9129
rect 13587 9064 16252 9092
rect 13587 9061 13599 9064
rect 13541 9055 13599 9061
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17589 9095 17647 9101
rect 17589 9092 17601 9095
rect 17092 9064 17601 9092
rect 17092 9052 17098 9064
rect 17589 9061 17601 9064
rect 17635 9061 17647 9095
rect 17972 9092 18000 9123
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18233 9163 18291 9169
rect 18233 9160 18245 9163
rect 18196 9132 18245 9160
rect 18196 9120 18202 9132
rect 18233 9129 18245 9132
rect 18279 9129 18291 9163
rect 18233 9123 18291 9129
rect 20806 9120 20812 9172
rect 20864 9160 20870 9172
rect 20993 9163 21051 9169
rect 20993 9160 21005 9163
rect 20864 9132 21005 9160
rect 20864 9120 20870 9132
rect 20993 9129 21005 9132
rect 21039 9129 21051 9163
rect 20993 9123 21051 9129
rect 18601 9095 18659 9101
rect 18601 9092 18613 9095
rect 17972 9064 18613 9092
rect 17589 9055 17647 9061
rect 18601 9061 18613 9064
rect 18647 9061 18659 9095
rect 18601 9055 18659 9061
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9933 9027 9991 9033
rect 9933 9024 9945 9027
rect 9640 8996 9945 9024
rect 9640 8984 9646 8996
rect 9933 8993 9945 8996
rect 9979 9024 9991 9027
rect 10318 9024 10324 9036
rect 9979 8996 10324 9024
rect 9979 8993 9991 8996
rect 9933 8987 9991 8993
rect 10318 8984 10324 8996
rect 10376 9024 10382 9036
rect 11698 9024 11704 9036
rect 10376 8996 11468 9024
rect 11659 8996 11704 9024
rect 10376 8984 10382 8996
rect 11440 8965 11468 8996
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 14366 8984 14372 9036
rect 14424 9024 14430 9036
rect 14826 9033 14832 9036
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14424 8996 14565 9024
rect 14424 8984 14430 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14820 9024 14832 9033
rect 14739 8996 14832 9024
rect 14553 8987 14611 8993
rect 14820 8987 14832 8996
rect 14884 9024 14890 9036
rect 15378 9024 15384 9036
rect 14884 8996 15384 9024
rect 14826 8984 14832 8987
rect 14884 8984 14890 8996
rect 15378 8984 15384 8996
rect 15436 8984 15442 9036
rect 15562 8984 15568 9036
rect 15620 9024 15626 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 15620 8996 16589 9024
rect 15620 8984 15626 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 17402 8984 17408 9036
rect 17460 9024 17466 9036
rect 17460 8996 18828 9024
rect 17460 8984 17466 8996
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 9456 8928 9689 8956
rect 9456 8916 9462 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 11425 8959 11483 8965
rect 11425 8925 11437 8959
rect 11471 8925 11483 8959
rect 11425 8919 11483 8925
rect 11609 8959 11667 8965
rect 11609 8925 11621 8959
rect 11655 8956 11667 8959
rect 12066 8956 12072 8968
rect 11655 8928 12072 8956
rect 11655 8925 11667 8928
rect 11609 8919 11667 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 13722 8956 13728 8968
rect 12406 8928 13308 8956
rect 13683 8928 13728 8956
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8573 8891 8631 8897
rect 8573 8888 8585 8891
rect 8168 8860 8585 8888
rect 8168 8848 8174 8860
rect 8573 8857 8585 8860
rect 8619 8857 8631 8891
rect 12406 8888 12434 8928
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 8573 8851 8631 8857
rect 10612 8860 12434 8888
rect 12636 8860 13185 8888
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7708 8792 7849 8820
rect 7708 8780 7714 8792
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8720 8792 9137 8820
rect 8720 8780 8726 8792
rect 9125 8789 9137 8792
rect 9171 8820 9183 8823
rect 10612 8820 10640 8860
rect 9171 8792 10640 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 12636 8820 12664 8860
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13280 8888 13308 8928
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 13998 8916 14004 8968
rect 14056 8956 14062 8968
rect 14458 8956 14464 8968
rect 14056 8928 14464 8956
rect 14056 8916 14062 8928
rect 14458 8916 14464 8928
rect 14516 8916 14522 8968
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8925 16819 8959
rect 16761 8919 16819 8925
rect 17313 8959 17371 8965
rect 17313 8925 17325 8959
rect 17359 8956 17371 8959
rect 18046 8956 18052 8968
rect 17359 8928 18052 8956
rect 17359 8925 17371 8928
rect 17313 8919 17371 8925
rect 14366 8888 14372 8900
rect 13280 8860 14372 8888
rect 13173 8851 13231 8857
rect 14366 8848 14372 8860
rect 14424 8848 14430 8900
rect 16117 8891 16175 8897
rect 16117 8857 16129 8891
rect 16163 8888 16175 8891
rect 16776 8888 16804 8919
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18690 8956 18696 8968
rect 18651 8928 18696 8956
rect 18690 8916 18696 8928
rect 18748 8916 18754 8968
rect 18800 8965 18828 8996
rect 20162 8984 20168 9036
rect 20220 9024 20226 9036
rect 20349 9027 20407 9033
rect 20349 9024 20361 9027
rect 20220 8996 20361 9024
rect 20220 8984 20226 8996
rect 20349 8993 20361 8996
rect 20395 8993 20407 9027
rect 20349 8987 20407 8993
rect 18785 8959 18843 8965
rect 18785 8925 18797 8959
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 19058 8916 19064 8968
rect 19116 8956 19122 8968
rect 20441 8959 20499 8965
rect 20441 8956 20453 8959
rect 19116 8928 20453 8956
rect 19116 8916 19122 8928
rect 20441 8925 20453 8928
rect 20487 8925 20499 8959
rect 20441 8919 20499 8925
rect 20625 8959 20683 8965
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 20990 8956 20996 8968
rect 20671 8928 20996 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 20990 8916 20996 8928
rect 21048 8916 21054 8968
rect 16163 8860 16804 8888
rect 16163 8857 16175 8860
rect 16117 8851 16175 8857
rect 12802 8820 12808 8832
rect 10744 8792 12664 8820
rect 12763 8792 12808 8820
rect 10744 8780 10750 8792
rect 12802 8780 12808 8792
rect 12860 8780 12866 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 18782 8820 18788 8832
rect 14516 8792 18788 8820
rect 14516 8780 14522 8792
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 19518 8780 19524 8832
rect 19576 8820 19582 8832
rect 19613 8823 19671 8829
rect 19613 8820 19625 8823
rect 19576 8792 19625 8820
rect 19576 8780 19582 8792
rect 19613 8789 19625 8792
rect 19659 8789 19671 8823
rect 19978 8820 19984 8832
rect 19939 8792 19984 8820
rect 19613 8783 19671 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 1104 8730 21896 8752
rect 1104 8678 4447 8730
rect 4499 8678 4511 8730
rect 4563 8678 4575 8730
rect 4627 8678 4639 8730
rect 4691 8678 11378 8730
rect 11430 8678 11442 8730
rect 11494 8678 11506 8730
rect 11558 8678 11570 8730
rect 11622 8678 18308 8730
rect 18360 8678 18372 8730
rect 18424 8678 18436 8730
rect 18488 8678 18500 8730
rect 18552 8678 21896 8730
rect 1104 8656 21896 8678
rect 7190 8616 7196 8628
rect 7151 8588 7196 8616
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 8389 8619 8447 8625
rect 8389 8585 8401 8619
rect 8435 8616 8447 8619
rect 9398 8616 9404 8628
rect 8435 8588 9404 8616
rect 8435 8585 8447 8588
rect 8389 8579 8447 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9582 8616 9588 8628
rect 9543 8588 9588 8616
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9674 8576 9680 8628
rect 9732 8616 9738 8628
rect 9732 8588 11100 8616
rect 9732 8576 9738 8588
rect 8849 8551 8907 8557
rect 8849 8517 8861 8551
rect 8895 8517 8907 8551
rect 8849 8511 8907 8517
rect 9309 8551 9367 8557
rect 9309 8517 9321 8551
rect 9355 8548 9367 8551
rect 9950 8548 9956 8560
rect 9355 8520 9956 8548
rect 9355 8517 9367 8520
rect 9309 8511 9367 8517
rect 8864 8480 8892 8511
rect 9950 8508 9956 8520
rect 10008 8508 10014 8560
rect 10962 8508 10968 8560
rect 11020 8508 11026 8560
rect 11072 8548 11100 8588
rect 11146 8576 11152 8628
rect 11204 8616 11210 8628
rect 13446 8616 13452 8628
rect 11204 8588 13452 8616
rect 11204 8576 11210 8588
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 13722 8616 13728 8628
rect 13587 8588 13728 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 13814 8576 13820 8628
rect 13872 8616 13878 8628
rect 14274 8616 14280 8628
rect 13872 8588 13917 8616
rect 14235 8588 14280 8616
rect 13872 8576 13878 8588
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 17954 8616 17960 8628
rect 14424 8588 17960 8616
rect 14424 8576 14430 8588
rect 17954 8576 17960 8588
rect 18012 8576 18018 8628
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 18690 8616 18696 8628
rect 18371 8588 18696 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 18690 8576 18696 8588
rect 18748 8576 18754 8628
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 19613 8619 19671 8625
rect 19613 8616 19625 8619
rect 19300 8588 19625 8616
rect 19300 8576 19306 8588
rect 19613 8585 19625 8588
rect 19659 8616 19671 8619
rect 19797 8619 19855 8625
rect 19797 8616 19809 8619
rect 19659 8588 19809 8616
rect 19659 8585 19671 8588
rect 19613 8579 19671 8585
rect 19797 8585 19809 8588
rect 19843 8585 19855 8619
rect 19797 8579 19855 8585
rect 11072 8520 12204 8548
rect 8864 8452 9996 8480
rect 7742 8372 7748 8424
rect 7800 8412 7806 8424
rect 8110 8412 8116 8424
rect 7800 8384 8116 8412
rect 7800 8372 7806 8384
rect 8110 8372 8116 8384
rect 8168 8412 8174 8424
rect 8205 8415 8263 8421
rect 8205 8412 8217 8415
rect 8168 8384 8217 8412
rect 8168 8372 8174 8384
rect 8205 8381 8217 8384
rect 8251 8381 8263 8415
rect 8662 8412 8668 8424
rect 8623 8384 8668 8412
rect 8205 8375 8263 8381
rect 8662 8372 8668 8384
rect 8720 8372 8726 8424
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9968 8412 9996 8452
rect 10980 8421 11008 8508
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11241 8483 11299 8489
rect 11241 8480 11253 8483
rect 11112 8452 11253 8480
rect 11112 8440 11118 8452
rect 11241 8449 11253 8452
rect 11287 8449 11299 8483
rect 12176 8480 12204 8520
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 18785 8551 18843 8557
rect 18785 8548 18797 8551
rect 18196 8520 18797 8548
rect 18196 8508 18202 8520
rect 18785 8517 18797 8520
rect 18831 8517 18843 8551
rect 19978 8548 19984 8560
rect 18785 8511 18843 8517
rect 19260 8520 19984 8548
rect 13633 8483 13691 8489
rect 12176 8452 12296 8480
rect 11241 8443 11299 8449
rect 10965 8415 11023 8421
rect 9968 8384 10916 8412
rect 10888 8356 10916 8384
rect 10965 8381 10977 8415
rect 11011 8412 11023 8415
rect 12161 8415 12219 8421
rect 12161 8412 12173 8415
rect 11011 8384 12173 8412
rect 11011 8381 11023 8384
rect 10965 8375 11023 8381
rect 12161 8381 12173 8384
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 7561 8347 7619 8353
rect 7561 8313 7573 8347
rect 7607 8344 7619 8347
rect 8478 8344 8484 8356
rect 7607 8316 8484 8344
rect 7607 8313 7619 8316
rect 7561 8307 7619 8313
rect 8478 8304 8484 8316
rect 8536 8344 8542 8356
rect 8754 8344 8760 8356
rect 8536 8316 8760 8344
rect 8536 8304 8542 8316
rect 8754 8304 8760 8316
rect 8812 8344 8818 8356
rect 10134 8344 10140 8356
rect 8812 8316 10140 8344
rect 8812 8304 8818 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10778 8353 10784 8356
rect 10720 8347 10784 8353
rect 10720 8313 10732 8347
rect 10766 8313 10784 8347
rect 10720 8307 10784 8313
rect 10778 8304 10784 8307
rect 10836 8304 10842 8356
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11330 8344 11336 8356
rect 10928 8316 11336 8344
rect 10928 8304 10934 8316
rect 11330 8304 11336 8316
rect 11388 8304 11394 8356
rect 12268 8344 12296 8452
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 13679 8452 14596 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 12434 8421 12440 8424
rect 12428 8375 12440 8421
rect 12492 8412 12498 8424
rect 14001 8415 14059 8421
rect 12492 8384 12528 8412
rect 12434 8372 12440 8375
rect 12492 8372 12498 8384
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14458 8412 14464 8424
rect 14047 8384 14464 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 14568 8412 14596 8452
rect 14642 8440 14648 8492
rect 14700 8480 14706 8492
rect 14826 8480 14832 8492
rect 14700 8452 14832 8480
rect 14700 8440 14706 8452
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 15562 8480 15568 8492
rect 15519 8452 15568 8480
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 16393 8483 16451 8489
rect 16393 8480 16405 8483
rect 15804 8452 16405 8480
rect 15804 8440 15810 8452
rect 16393 8449 16405 8452
rect 16439 8449 16451 8483
rect 17773 8483 17831 8489
rect 16393 8443 16451 8449
rect 16776 8452 17264 8480
rect 16776 8412 16804 8452
rect 14568 8384 16804 8412
rect 16850 8372 16856 8424
rect 16908 8412 16914 8424
rect 17129 8415 17187 8421
rect 17129 8412 17141 8415
rect 16908 8384 17141 8412
rect 16908 8372 16914 8384
rect 17129 8381 17141 8384
rect 17175 8381 17187 8415
rect 17236 8412 17264 8452
rect 17773 8449 17785 8483
rect 17819 8480 17831 8483
rect 18046 8480 18052 8492
rect 17819 8452 18052 8480
rect 17819 8449 17831 8452
rect 17773 8443 17831 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 19260 8489 19288 8520
rect 19978 8508 19984 8520
rect 20036 8508 20042 8560
rect 19245 8483 19303 8489
rect 19245 8449 19257 8483
rect 19291 8449 19303 8483
rect 19245 8443 19303 8449
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8480 19487 8483
rect 19613 8483 19671 8489
rect 19613 8480 19625 8483
rect 19475 8452 19625 8480
rect 19475 8449 19487 8452
rect 19429 8443 19487 8449
rect 19613 8449 19625 8452
rect 19659 8449 19671 8483
rect 19613 8443 19671 8449
rect 17957 8415 18015 8421
rect 17957 8412 17969 8415
rect 17236 8384 17969 8412
rect 17129 8375 17187 8381
rect 17957 8381 17969 8384
rect 18003 8412 18015 8415
rect 18782 8412 18788 8424
rect 18003 8384 18788 8412
rect 18003 8381 18015 8384
rect 17957 8375 18015 8381
rect 18782 8372 18788 8384
rect 18840 8372 18846 8424
rect 19150 8412 19156 8424
rect 19111 8384 19156 8412
rect 19150 8372 19156 8384
rect 19208 8372 19214 8424
rect 19334 8372 19340 8424
rect 19392 8412 19398 8424
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 19392 8384 21189 8412
rect 19392 8372 19398 8384
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 21177 8375 21235 8381
rect 12268 8316 12848 8344
rect 7190 8236 7196 8288
rect 7248 8276 7254 8288
rect 7466 8276 7472 8288
rect 7248 8248 7472 8276
rect 7248 8236 7254 8248
rect 7466 8236 7472 8248
rect 7524 8276 7530 8288
rect 7837 8279 7895 8285
rect 7837 8276 7849 8279
rect 7524 8248 7849 8276
rect 7524 8236 7530 8248
rect 7837 8245 7849 8248
rect 7883 8245 7895 8279
rect 7837 8239 7895 8245
rect 10962 8236 10968 8288
rect 11020 8276 11026 8288
rect 11701 8279 11759 8285
rect 11701 8276 11713 8279
rect 11020 8248 11713 8276
rect 11020 8236 11026 8248
rect 11701 8245 11713 8248
rect 11747 8276 11759 8279
rect 11790 8276 11796 8288
rect 11747 8248 11796 8276
rect 11747 8245 11759 8248
rect 11701 8239 11759 8245
rect 11790 8236 11796 8248
rect 11848 8236 11854 8288
rect 12820 8276 12848 8316
rect 12894 8304 12900 8356
rect 12952 8344 12958 8356
rect 14645 8347 14703 8353
rect 14645 8344 14657 8347
rect 12952 8316 14657 8344
rect 12952 8304 12958 8316
rect 14645 8313 14657 8316
rect 14691 8313 14703 8347
rect 14645 8307 14703 8313
rect 14737 8347 14795 8353
rect 14737 8313 14749 8347
rect 14783 8344 14795 8347
rect 14826 8344 14832 8356
rect 14783 8316 14832 8344
rect 14783 8313 14795 8316
rect 14737 8307 14795 8313
rect 14826 8304 14832 8316
rect 14884 8304 14890 8356
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 16209 8347 16267 8353
rect 16209 8344 16221 8347
rect 16080 8316 16221 8344
rect 16080 8304 16086 8316
rect 16209 8313 16221 8316
rect 16255 8313 16267 8347
rect 16209 8307 16267 8313
rect 16301 8347 16359 8353
rect 16301 8313 16313 8347
rect 16347 8344 16359 8347
rect 17586 8344 17592 8356
rect 16347 8316 17592 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 17586 8304 17592 8316
rect 17644 8304 17650 8356
rect 20622 8344 20628 8356
rect 17696 8316 20628 8344
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 12820 8248 13645 8276
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 14550 8236 14556 8288
rect 14608 8276 14614 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 14608 8248 15853 8276
rect 14608 8236 14614 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 17313 8279 17371 8285
rect 17313 8245 17325 8279
rect 17359 8276 17371 8279
rect 17696 8276 17724 8316
rect 20622 8304 20628 8316
rect 20680 8304 20686 8356
rect 20990 8353 20996 8356
rect 20932 8347 20996 8353
rect 20932 8313 20944 8347
rect 20978 8313 20996 8347
rect 20932 8307 20996 8313
rect 20990 8304 20996 8307
rect 21048 8304 21054 8356
rect 17359 8248 17724 8276
rect 17865 8279 17923 8285
rect 17359 8245 17371 8248
rect 17313 8239 17371 8245
rect 17865 8245 17877 8279
rect 17911 8276 17923 8279
rect 18046 8276 18052 8288
rect 17911 8248 18052 8276
rect 17911 8245 17923 8248
rect 17865 8239 17923 8245
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 19242 8276 19248 8288
rect 19024 8248 19248 8276
rect 19024 8236 19030 8248
rect 19242 8236 19248 8248
rect 19300 8236 19306 8288
rect 1104 8186 21896 8208
rect 1104 8134 7912 8186
rect 7964 8134 7976 8186
rect 8028 8134 8040 8186
rect 8092 8134 8104 8186
rect 8156 8134 14843 8186
rect 14895 8134 14907 8186
rect 14959 8134 14971 8186
rect 15023 8134 15035 8186
rect 15087 8134 21896 8186
rect 1104 8112 21896 8134
rect 7006 8072 7012 8084
rect 6967 8044 7012 8072
rect 7006 8032 7012 8044
rect 7064 8032 7070 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 9180 8044 9321 8072
rect 9180 8032 9186 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 9916 8044 10149 8072
rect 9916 8032 9922 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10689 8075 10747 8081
rect 10689 8072 10701 8075
rect 10284 8044 10701 8072
rect 10284 8032 10290 8044
rect 10689 8041 10701 8044
rect 10735 8072 10747 8075
rect 10962 8072 10968 8084
rect 10735 8044 10968 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10962 8032 10968 8044
rect 11020 8032 11026 8084
rect 11057 8075 11115 8081
rect 11057 8041 11069 8075
rect 11103 8072 11115 8075
rect 11698 8072 11704 8084
rect 11103 8044 11704 8072
rect 11103 8041 11115 8044
rect 11057 8035 11115 8041
rect 11698 8032 11704 8044
rect 11756 8032 11762 8084
rect 12066 8072 12072 8084
rect 12027 8044 12072 8072
rect 12066 8032 12072 8044
rect 12124 8032 12130 8084
rect 12342 8032 12348 8084
rect 12400 8072 12406 8084
rect 12400 8044 14596 8072
rect 12400 8032 12406 8044
rect 7837 8007 7895 8013
rect 7837 7973 7849 8007
rect 7883 8004 7895 8007
rect 11790 8004 11796 8016
rect 7883 7976 11796 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 8588 7945 8616 7976
rect 11790 7964 11796 7976
rect 11848 7964 11854 8016
rect 12796 8007 12854 8013
rect 12796 7973 12808 8007
rect 12842 8004 12854 8007
rect 13722 8004 13728 8016
rect 12842 7976 13728 8004
rect 12842 7973 12854 7976
rect 12796 7967 12854 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 14458 8004 14464 8016
rect 14419 7976 14464 8004
rect 14458 7964 14464 7976
rect 14516 7964 14522 8016
rect 14568 8004 14596 8044
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 14921 8075 14979 8081
rect 14921 8072 14933 8075
rect 14700 8044 14933 8072
rect 14700 8032 14706 8044
rect 14921 8041 14933 8044
rect 14967 8041 14979 8075
rect 17678 8072 17684 8084
rect 17639 8044 17684 8072
rect 14921 8035 14979 8041
rect 17678 8032 17684 8044
rect 17736 8032 17742 8084
rect 18782 8072 18788 8084
rect 18743 8044 18788 8072
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 20990 8032 20996 8084
rect 21048 8072 21054 8084
rect 21177 8075 21235 8081
rect 21177 8072 21189 8075
rect 21048 8044 21189 8072
rect 21048 8032 21054 8044
rect 21177 8041 21189 8044
rect 21223 8041 21235 8075
rect 21177 8035 21235 8041
rect 17862 8004 17868 8016
rect 14568 7976 17868 8004
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 8113 7939 8171 7945
rect 8113 7936 8125 7939
rect 7515 7908 8125 7936
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 8113 7905 8125 7908
rect 8159 7905 8171 7939
rect 8113 7899 8171 7905
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7905 8631 7939
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 8573 7899 8631 7905
rect 8128 7800 8156 7899
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 10778 7936 10784 7948
rect 10520 7908 10784 7936
rect 8846 7828 8852 7880
rect 8904 7868 8910 7880
rect 9030 7868 9036 7880
rect 8904 7840 9036 7868
rect 8904 7828 8910 7840
rect 9030 7828 9036 7840
rect 9088 7828 9094 7880
rect 9766 7868 9772 7880
rect 9727 7840 9772 7868
rect 9766 7828 9772 7840
rect 9824 7828 9830 7880
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7868 10011 7871
rect 10042 7868 10048 7880
rect 9999 7840 10048 7868
rect 9999 7837 10011 7840
rect 9953 7831 10011 7837
rect 10042 7828 10048 7840
rect 10100 7828 10106 7880
rect 10520 7877 10548 7908
rect 10778 7896 10784 7908
rect 10836 7936 10842 7948
rect 10836 7908 11192 7936
rect 10836 7896 10842 7908
rect 11164 7880 11192 7908
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 11701 7939 11759 7945
rect 11701 7936 11713 7939
rect 11388 7908 11713 7936
rect 11388 7896 11394 7908
rect 11701 7905 11713 7908
rect 11747 7905 11759 7939
rect 11701 7899 11759 7905
rect 15746 7896 15752 7948
rect 15804 7936 15810 7948
rect 16034 7939 16092 7945
rect 16034 7936 16046 7939
rect 15804 7908 16046 7936
rect 15804 7896 15810 7908
rect 16034 7905 16046 7908
rect 16080 7905 16092 7939
rect 17770 7936 17776 7948
rect 17731 7908 17776 7936
rect 16034 7899 16092 7905
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 18046 7896 18052 7948
rect 18104 7936 18110 7948
rect 18693 7939 18751 7945
rect 18693 7936 18705 7939
rect 18104 7908 18705 7936
rect 18104 7896 18110 7908
rect 18693 7905 18705 7908
rect 18739 7905 18751 7939
rect 18693 7899 18751 7905
rect 19334 7896 19340 7948
rect 19392 7936 19398 7948
rect 19797 7939 19855 7945
rect 19797 7936 19809 7939
rect 19392 7908 19809 7936
rect 19392 7896 19398 7908
rect 19797 7905 19809 7908
rect 19843 7905 19855 7939
rect 19797 7899 19855 7905
rect 20064 7939 20122 7945
rect 20064 7905 20076 7939
rect 20110 7936 20122 7939
rect 20530 7936 20536 7948
rect 20110 7908 20536 7936
rect 20110 7905 20122 7908
rect 20064 7899 20122 7905
rect 20530 7896 20536 7908
rect 20588 7896 20594 7948
rect 10505 7871 10563 7877
rect 10505 7837 10517 7871
rect 10551 7837 10563 7871
rect 10505 7831 10563 7837
rect 10597 7871 10655 7877
rect 10597 7837 10609 7871
rect 10643 7837 10655 7871
rect 10597 7831 10655 7837
rect 9858 7800 9864 7812
rect 8128 7772 9864 7800
rect 9858 7760 9864 7772
rect 9916 7760 9922 7812
rect 10137 7803 10195 7809
rect 10137 7769 10149 7803
rect 10183 7800 10195 7803
rect 10612 7800 10640 7831
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 11425 7871 11483 7877
rect 11425 7868 11437 7871
rect 11204 7840 11437 7868
rect 11204 7828 11210 7840
rect 11425 7837 11437 7840
rect 11471 7837 11483 7871
rect 11425 7831 11483 7837
rect 11609 7871 11667 7877
rect 11609 7837 11621 7871
rect 11655 7868 11667 7871
rect 11790 7868 11796 7880
rect 11655 7840 11796 7868
rect 11655 7837 11667 7840
rect 11609 7831 11667 7837
rect 11790 7828 11796 7840
rect 11848 7828 11854 7880
rect 12526 7868 12532 7880
rect 12487 7840 12532 7868
rect 12526 7828 12532 7840
rect 12584 7828 12590 7880
rect 16298 7868 16304 7880
rect 16259 7840 16304 7868
rect 16298 7828 16304 7840
rect 16356 7828 16362 7880
rect 16390 7828 16396 7880
rect 16448 7868 16454 7880
rect 16853 7871 16911 7877
rect 16853 7868 16865 7871
rect 16448 7840 16865 7868
rect 16448 7828 16454 7840
rect 16853 7837 16865 7840
rect 16899 7837 16911 7871
rect 16853 7831 16911 7837
rect 17310 7828 17316 7880
rect 17368 7868 17374 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17368 7840 17509 7868
rect 17368 7828 17374 7840
rect 17497 7837 17509 7840
rect 17543 7868 17555 7871
rect 18509 7871 18567 7877
rect 18509 7868 18521 7871
rect 17543 7840 18521 7868
rect 17543 7837 17555 7840
rect 17497 7831 17555 7837
rect 18509 7837 18521 7840
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 12066 7800 12072 7812
rect 10183 7772 12072 7800
rect 10183 7769 10195 7772
rect 10137 7763 10195 7769
rect 12066 7760 12072 7772
rect 12124 7760 12130 7812
rect 13740 7772 14118 7800
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8757 7735 8815 7741
rect 8757 7701 8769 7735
rect 8803 7732 8815 7735
rect 13740 7732 13768 7772
rect 13906 7732 13912 7744
rect 8803 7704 13768 7732
rect 13867 7704 13912 7732
rect 8803 7701 8815 7704
rect 8757 7695 8815 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14090 7732 14118 7772
rect 16316 7772 19840 7800
rect 16316 7732 16344 7772
rect 14090 7704 16344 7732
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18966 7732 18972 7744
rect 18187 7704 18972 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 19150 7732 19156 7744
rect 19111 7704 19156 7732
rect 19150 7692 19156 7704
rect 19208 7692 19214 7744
rect 19812 7732 19840 7772
rect 20990 7732 20996 7744
rect 19812 7704 20996 7732
rect 20990 7692 20996 7704
rect 21048 7692 21054 7744
rect 1104 7642 21896 7664
rect 1104 7590 4447 7642
rect 4499 7590 4511 7642
rect 4563 7590 4575 7642
rect 4627 7590 4639 7642
rect 4691 7590 11378 7642
rect 11430 7590 11442 7642
rect 11494 7590 11506 7642
rect 11558 7590 11570 7642
rect 11622 7590 18308 7642
rect 18360 7590 18372 7642
rect 18424 7590 18436 7642
rect 18488 7590 18500 7642
rect 18552 7590 21896 7642
rect 1104 7568 21896 7590
rect 7377 7531 7435 7537
rect 7377 7497 7389 7531
rect 7423 7528 7435 7531
rect 7650 7528 7656 7540
rect 7423 7500 7656 7528
rect 7423 7497 7435 7500
rect 7377 7491 7435 7497
rect 7650 7488 7656 7500
rect 7708 7528 7714 7540
rect 9493 7531 9551 7537
rect 7708 7500 9168 7528
rect 7708 7488 7714 7500
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 7009 7463 7067 7469
rect 7009 7460 7021 7463
rect 6880 7432 7021 7460
rect 6880 7420 6886 7432
rect 7009 7429 7021 7432
rect 7055 7460 7067 7463
rect 8110 7460 8116 7472
rect 7055 7432 8116 7460
rect 7055 7429 7067 7432
rect 7009 7423 7067 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 9140 7392 9168 7500
rect 9493 7497 9505 7531
rect 9539 7528 9551 7531
rect 10042 7528 10048 7540
rect 9539 7500 10048 7528
rect 9539 7497 9551 7500
rect 9493 7491 9551 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 11146 7528 11152 7540
rect 11107 7500 11152 7528
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 11440 7500 11836 7528
rect 11440 7472 11468 7500
rect 11422 7420 11428 7472
rect 11480 7420 11486 7472
rect 11514 7420 11520 7472
rect 11572 7460 11578 7472
rect 11808 7460 11836 7500
rect 12250 7488 12256 7540
rect 12308 7528 12314 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 12308 7500 12357 7528
rect 12308 7488 12314 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12437 7531 12495 7537
rect 12437 7497 12449 7531
rect 12483 7528 12495 7531
rect 15105 7531 15163 7537
rect 12483 7500 14596 7528
rect 12483 7497 12495 7500
rect 12437 7491 12495 7497
rect 14458 7460 14464 7472
rect 11572 7432 11744 7460
rect 11808 7432 14464 7460
rect 11572 7420 11578 7432
rect 9140 7364 9904 7392
rect 9876 7336 9904 7364
rect 11054 7352 11060 7404
rect 11112 7352 11118 7404
rect 11716 7392 11744 7432
rect 14458 7420 14464 7432
rect 14516 7420 14522 7472
rect 14568 7460 14596 7500
rect 15105 7497 15117 7531
rect 15151 7528 15163 7531
rect 15746 7528 15752 7540
rect 15151 7500 15752 7528
rect 15151 7497 15163 7500
rect 15105 7491 15163 7497
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 16356 7500 16528 7528
rect 16356 7488 16362 7500
rect 15470 7460 15476 7472
rect 14568 7432 15476 7460
rect 15470 7420 15476 7432
rect 15528 7420 15534 7472
rect 13173 7395 13231 7401
rect 13173 7392 13185 7395
rect 11716 7364 13185 7392
rect 13173 7361 13185 7364
rect 13219 7361 13231 7395
rect 13173 7355 13231 7361
rect 13906 7352 13912 7404
rect 13964 7392 13970 7404
rect 16500 7401 16528 7500
rect 16592 7500 17141 7528
rect 14185 7395 14243 7401
rect 14185 7392 14197 7395
rect 13964 7364 14197 7392
rect 13964 7352 13970 7364
rect 14185 7361 14197 7364
rect 14231 7361 14243 7395
rect 14185 7355 14243 7361
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 7742 7284 7748 7336
rect 7800 7324 7806 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7800 7296 7849 7324
rect 7800 7284 7806 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 8113 7327 8171 7333
rect 8113 7293 8125 7327
rect 8159 7324 8171 7327
rect 9769 7327 9827 7333
rect 9769 7324 9781 7327
rect 8159 7296 9781 7324
rect 8159 7293 8171 7296
rect 8113 7287 8171 7293
rect 9769 7293 9781 7296
rect 9815 7293 9827 7327
rect 9769 7287 9827 7293
rect 7558 7148 7564 7200
rect 7616 7188 7622 7200
rect 7653 7191 7711 7197
rect 7653 7188 7665 7191
rect 7616 7160 7665 7188
rect 7616 7148 7622 7160
rect 7653 7157 7665 7160
rect 7699 7188 7711 7191
rect 8128 7188 8156 7287
rect 8380 7259 8438 7265
rect 8380 7225 8392 7259
rect 8426 7256 8438 7259
rect 9030 7256 9036 7268
rect 8426 7228 9036 7256
rect 8426 7225 8438 7228
rect 8380 7219 8438 7225
rect 9030 7216 9036 7228
rect 9088 7216 9094 7268
rect 9784 7256 9812 7287
rect 9858 7284 9864 7336
rect 9916 7284 9922 7336
rect 10042 7333 10048 7336
rect 10036 7324 10048 7333
rect 10003 7296 10048 7324
rect 10036 7287 10048 7296
rect 10042 7284 10048 7287
rect 10100 7284 10106 7336
rect 10410 7284 10416 7336
rect 10468 7324 10474 7336
rect 11072 7324 11100 7352
rect 10468 7296 11100 7324
rect 11977 7327 12035 7333
rect 10468 7284 10474 7296
rect 11977 7293 11989 7327
rect 12023 7324 12035 7327
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 12023 7296 12173 7324
rect 12023 7293 12035 7296
rect 11977 7287 12035 7293
rect 12161 7293 12173 7296
rect 12207 7324 12219 7327
rect 12437 7327 12495 7333
rect 12437 7324 12449 7327
rect 12207 7296 12449 7324
rect 12207 7293 12219 7296
rect 12161 7287 12219 7293
rect 12437 7293 12449 7296
rect 12483 7293 12495 7327
rect 12437 7287 12495 7293
rect 12526 7284 12532 7336
rect 12584 7324 12590 7336
rect 12802 7324 12808 7336
rect 12584 7296 12808 7324
rect 12584 7284 12590 7296
rect 12802 7284 12808 7296
rect 12860 7284 12866 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14001 7327 14059 7333
rect 14001 7324 14013 7327
rect 13872 7296 14013 7324
rect 13872 7284 13878 7296
rect 14001 7293 14013 7296
rect 14047 7293 14059 7327
rect 14001 7287 14059 7293
rect 14829 7327 14887 7333
rect 14829 7293 14841 7327
rect 14875 7293 14887 7327
rect 16206 7324 16212 7336
rect 16264 7333 16270 7336
rect 16264 7327 16287 7333
rect 16139 7296 16212 7324
rect 14829 7287 14887 7293
rect 10962 7256 10968 7268
rect 9784 7228 10968 7256
rect 10962 7216 10968 7228
rect 11020 7216 11026 7268
rect 12986 7256 12992 7268
rect 11440 7228 12664 7256
rect 12947 7228 12992 7256
rect 7699 7160 8156 7188
rect 7699 7157 7711 7160
rect 7653 7151 7711 7157
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 11440 7188 11468 7228
rect 12636 7197 12664 7228
rect 12986 7216 12992 7228
rect 13044 7216 13050 7268
rect 13354 7216 13360 7268
rect 13412 7256 13418 7268
rect 14093 7259 14151 7265
rect 14093 7256 14105 7259
rect 13412 7228 14105 7256
rect 13412 7216 13418 7228
rect 14093 7225 14105 7228
rect 14139 7225 14151 7259
rect 14844 7256 14872 7287
rect 16206 7284 16212 7296
rect 16275 7324 16287 7327
rect 16592 7324 16620 7500
rect 17129 7497 17141 7500
rect 17175 7528 17187 7531
rect 17175 7500 18552 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 18524 7460 18552 7500
rect 18524 7432 19380 7460
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 19352 7401 19380 7432
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 19024 7364 19257 7392
rect 19024 7352 19030 7364
rect 19245 7361 19257 7364
rect 19291 7361 19303 7395
rect 19245 7355 19303 7361
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7361 19395 7395
rect 19337 7355 19395 7361
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20441 7395 20499 7401
rect 20441 7392 20453 7395
rect 20128 7364 20453 7392
rect 20128 7352 20134 7364
rect 20441 7361 20453 7364
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 16275 7296 16620 7324
rect 18509 7327 18567 7333
rect 16275 7293 16287 7296
rect 16264 7287 16287 7293
rect 18509 7293 18521 7327
rect 18555 7324 18567 7327
rect 18874 7324 18880 7336
rect 18555 7296 18880 7324
rect 18555 7293 18567 7296
rect 18509 7287 18567 7293
rect 16264 7284 16270 7287
rect 18874 7284 18880 7296
rect 18932 7284 18938 7336
rect 19150 7324 19156 7336
rect 19111 7296 19156 7324
rect 19150 7284 19156 7296
rect 19208 7284 19214 7336
rect 17126 7256 17132 7268
rect 14844 7228 17132 7256
rect 14093 7219 14151 7225
rect 17126 7216 17132 7228
rect 17184 7216 17190 7268
rect 17310 7216 17316 7268
rect 17368 7256 17374 7268
rect 18242 7259 18300 7265
rect 18242 7256 18254 7259
rect 17368 7228 18254 7256
rect 17368 7216 17374 7228
rect 18242 7225 18254 7228
rect 18288 7225 18300 7259
rect 18242 7219 18300 7225
rect 8260 7160 11468 7188
rect 11885 7191 11943 7197
rect 8260 7148 8266 7160
rect 11885 7157 11897 7191
rect 11931 7188 11943 7191
rect 11977 7191 12035 7197
rect 11977 7188 11989 7191
rect 11931 7160 11989 7188
rect 11931 7157 11943 7160
rect 11885 7151 11943 7157
rect 11977 7157 11989 7160
rect 12023 7157 12035 7191
rect 11977 7151 12035 7157
rect 12621 7191 12679 7197
rect 12621 7157 12633 7191
rect 12667 7157 12679 7191
rect 13078 7188 13084 7200
rect 13039 7160 13084 7188
rect 12621 7151 12679 7157
rect 13078 7148 13084 7160
rect 13136 7148 13142 7200
rect 13630 7188 13636 7200
rect 13591 7160 13636 7188
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 14182 7148 14188 7200
rect 14240 7188 14246 7200
rect 14645 7191 14703 7197
rect 14645 7188 14657 7191
rect 14240 7160 14657 7188
rect 14240 7148 14246 7160
rect 14645 7157 14657 7160
rect 14691 7157 14703 7191
rect 14645 7151 14703 7157
rect 17586 7148 17592 7200
rect 17644 7188 17650 7200
rect 18785 7191 18843 7197
rect 18785 7188 18797 7191
rect 17644 7160 18797 7188
rect 17644 7148 17650 7160
rect 18785 7157 18797 7160
rect 18831 7157 18843 7191
rect 19886 7188 19892 7200
rect 19847 7160 19892 7188
rect 18785 7151 18843 7157
rect 19886 7148 19892 7160
rect 19944 7148 19950 7200
rect 20254 7188 20260 7200
rect 20215 7160 20260 7188
rect 20254 7148 20260 7160
rect 20312 7148 20318 7200
rect 20346 7148 20352 7200
rect 20404 7188 20410 7200
rect 20898 7188 20904 7200
rect 20404 7160 20449 7188
rect 20859 7160 20904 7188
rect 20404 7148 20410 7160
rect 20898 7148 20904 7160
rect 20956 7148 20962 7200
rect 1104 7098 21896 7120
rect 1104 7046 7912 7098
rect 7964 7046 7976 7098
rect 8028 7046 8040 7098
rect 8092 7046 8104 7098
rect 8156 7046 14843 7098
rect 14895 7046 14907 7098
rect 14959 7046 14971 7098
rect 15023 7046 15035 7098
rect 15087 7046 21896 7098
rect 1104 7024 21896 7046
rect 9674 6944 9680 6996
rect 9732 6984 9738 6996
rect 10045 6987 10103 6993
rect 10045 6984 10057 6987
rect 9732 6956 10057 6984
rect 9732 6944 9738 6956
rect 10045 6953 10057 6956
rect 10091 6953 10103 6987
rect 10045 6947 10103 6953
rect 10318 6944 10324 6996
rect 10376 6984 10382 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10376 6956 10885 6984
rect 10376 6944 10382 6956
rect 10873 6953 10885 6956
rect 10919 6984 10931 6987
rect 11330 6984 11336 6996
rect 10919 6956 11336 6984
rect 10919 6953 10931 6956
rect 10873 6947 10931 6953
rect 11330 6944 11336 6956
rect 11388 6944 11394 6996
rect 11514 6984 11520 6996
rect 11475 6956 11520 6984
rect 11514 6944 11520 6956
rect 11572 6984 11578 6996
rect 11790 6984 11796 6996
rect 11572 6956 11796 6984
rect 11572 6944 11578 6956
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12400 6956 13492 6984
rect 12400 6944 12406 6956
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 11425 6919 11483 6925
rect 8352 6888 11008 6916
rect 8352 6876 8358 6888
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6808 6610 6860
rect 7009 6851 7067 6857
rect 7009 6817 7021 6851
rect 7055 6848 7067 6851
rect 7650 6848 7656 6860
rect 7055 6820 7656 6848
rect 7055 6817 7067 6820
rect 7009 6811 7067 6817
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 8110 6848 8116 6860
rect 8071 6820 8116 6848
rect 8110 6808 8116 6820
rect 8168 6808 8174 6860
rect 10980 6857 11008 6888
rect 11425 6885 11437 6919
rect 11471 6916 11483 6919
rect 12434 6916 12440 6928
rect 11471 6888 12440 6916
rect 11471 6885 11483 6888
rect 11425 6879 11483 6885
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 13170 6916 13176 6928
rect 12544 6888 13176 6916
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 8803 6820 9689 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 9677 6811 9735 6817
rect 10965 6851 11023 6857
rect 10965 6817 10977 6851
rect 11011 6848 11023 6851
rect 12544 6848 12572 6888
rect 13170 6876 13176 6888
rect 13228 6876 13234 6928
rect 13464 6916 13492 6956
rect 13538 6944 13544 6996
rect 13596 6984 13602 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13596 6956 13645 6984
rect 13596 6944 13602 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 16390 6984 16396 6996
rect 16351 6956 16396 6984
rect 13633 6947 13691 6953
rect 16390 6944 16396 6956
rect 16448 6944 16454 6996
rect 16482 6944 16488 6996
rect 16540 6984 16546 6996
rect 18877 6987 18935 6993
rect 16540 6956 18276 6984
rect 16540 6944 16546 6956
rect 14921 6919 14979 6925
rect 14921 6916 14933 6919
rect 13464 6888 14933 6916
rect 14921 6885 14933 6888
rect 14967 6916 14979 6919
rect 16114 6916 16120 6928
rect 14967 6888 16120 6916
rect 14967 6885 14979 6888
rect 14921 6879 14979 6885
rect 16114 6876 16120 6888
rect 16172 6916 16178 6928
rect 17405 6919 17463 6925
rect 17405 6916 17417 6919
rect 16172 6888 17417 6916
rect 16172 6876 16178 6888
rect 17405 6885 17417 6888
rect 17451 6885 17463 6919
rect 17405 6879 17463 6885
rect 18248 6916 18276 6956
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 20898 6984 20904 6996
rect 18923 6956 20904 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 20898 6944 20904 6956
rect 20956 6944 20962 6996
rect 19058 6916 19064 6928
rect 18248 6888 19064 6916
rect 11011 6820 12572 6848
rect 11011 6817 11023 6820
rect 10965 6811 11023 6817
rect 12618 6808 12624 6860
rect 12676 6857 12682 6860
rect 12676 6848 12688 6857
rect 12676 6820 12721 6848
rect 12676 6811 12688 6820
rect 12676 6808 12682 6811
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 12897 6851 12955 6857
rect 12897 6848 12909 6851
rect 12860 6820 12909 6848
rect 12860 6808 12866 6820
rect 12897 6817 12909 6820
rect 12943 6817 12955 6851
rect 12897 6811 12955 6817
rect 13814 6808 13820 6860
rect 13872 6848 13878 6860
rect 14734 6848 14740 6860
rect 13872 6820 14740 6848
rect 13872 6808 13878 6820
rect 14734 6808 14740 6820
rect 14792 6808 14798 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15565 6851 15623 6857
rect 15565 6848 15577 6851
rect 15252 6820 15577 6848
rect 15252 6808 15258 6820
rect 15565 6817 15577 6820
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 17494 6848 17500 6860
rect 16264 6820 16620 6848
rect 17455 6820 17500 6848
rect 16264 6808 16270 6820
rect 7377 6783 7435 6789
rect 7377 6749 7389 6783
rect 7423 6780 7435 6783
rect 8128 6780 8156 6808
rect 7423 6752 8156 6780
rect 7423 6749 7435 6752
rect 7377 6743 7435 6749
rect 9030 6740 9036 6792
rect 9088 6780 9094 6792
rect 9401 6783 9459 6789
rect 9401 6780 9413 6783
rect 9088 6752 9413 6780
rect 9088 6740 9094 6752
rect 9401 6749 9413 6752
rect 9447 6749 9459 6783
rect 9582 6780 9588 6792
rect 9543 6752 9588 6780
rect 9401 6743 9459 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10502 6780 10508 6792
rect 10376 6752 10508 6780
rect 10376 6740 10382 6752
rect 10502 6740 10508 6752
rect 10560 6740 10566 6792
rect 10870 6740 10876 6792
rect 10928 6780 10934 6792
rect 11057 6783 11115 6789
rect 11057 6780 11069 6783
rect 10928 6752 11069 6780
rect 10928 6740 10934 6752
rect 11057 6749 11069 6752
rect 11103 6749 11115 6783
rect 13725 6783 13783 6789
rect 13725 6780 13737 6783
rect 11057 6743 11115 6749
rect 12912 6752 13737 6780
rect 12912 6724 12940 6752
rect 13725 6749 13737 6752
rect 13771 6749 13783 6783
rect 13906 6780 13912 6792
rect 13867 6752 13912 6780
rect 13725 6743 13783 6749
rect 13906 6740 13912 6752
rect 13964 6740 13970 6792
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 16592 6789 16620 6820
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 18248 6857 18276 6888
rect 19058 6876 19064 6888
rect 19116 6876 19122 6928
rect 20070 6925 20076 6928
rect 20064 6916 20076 6925
rect 19352 6888 20076 6916
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6817 18291 6851
rect 19352 6848 19380 6888
rect 20064 6879 20076 6888
rect 20070 6876 20076 6879
rect 20128 6876 20134 6928
rect 18233 6811 18291 6817
rect 18616 6820 19380 6848
rect 15013 6783 15071 6789
rect 15013 6780 15025 6783
rect 14148 6752 15025 6780
rect 14148 6740 14154 6752
rect 15013 6749 15025 6752
rect 15059 6749 15071 6783
rect 15013 6743 15071 6749
rect 15105 6783 15163 6789
rect 15105 6749 15117 6783
rect 15151 6749 15163 6783
rect 15105 6743 15163 6749
rect 16485 6783 16543 6789
rect 16485 6749 16497 6783
rect 16531 6749 16543 6783
rect 16485 6743 16543 6749
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6749 16635 6783
rect 16577 6743 16635 6749
rect 8754 6672 8760 6724
rect 8812 6712 8818 6724
rect 10686 6712 10692 6724
rect 8812 6684 10692 6712
rect 8812 6672 8818 6684
rect 10686 6672 10692 6684
rect 10744 6672 10750 6724
rect 10778 6672 10784 6724
rect 10836 6712 10842 6724
rect 11425 6715 11483 6721
rect 11425 6712 11437 6715
rect 10836 6684 11437 6712
rect 10836 6672 10842 6684
rect 11425 6681 11437 6684
rect 11471 6681 11483 6715
rect 11425 6675 11483 6681
rect 12894 6672 12900 6724
rect 12952 6672 12958 6724
rect 13354 6712 13360 6724
rect 13096 6684 13360 6712
rect 6270 6644 6276 6656
rect 6231 6616 6276 6644
rect 6270 6604 6276 6616
rect 6328 6604 6334 6656
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 9398 6644 9404 6656
rect 8343 6616 9404 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 10502 6644 10508 6656
rect 10463 6616 10508 6644
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 11146 6604 11152 6656
rect 11204 6644 11210 6656
rect 13096 6644 13124 6684
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 13924 6712 13952 6740
rect 15120 6712 15148 6743
rect 16022 6712 16028 6724
rect 13924 6684 15148 6712
rect 15983 6684 16028 6712
rect 16022 6672 16028 6684
rect 16080 6672 16086 6724
rect 16500 6712 16528 6743
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 18616 6789 18644 6820
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17368 6752 17601 6780
rect 17368 6740 17374 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6749 18659 6783
rect 18782 6780 18788 6792
rect 18743 6752 18788 6780
rect 18601 6743 18659 6749
rect 18782 6740 18788 6752
rect 18840 6740 18846 6792
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 18932 6752 19809 6780
rect 18932 6740 18938 6752
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 17037 6715 17095 6721
rect 17037 6712 17049 6715
rect 16500 6684 17049 6712
rect 17037 6681 17049 6684
rect 17083 6681 17095 6715
rect 17037 6675 17095 6681
rect 13262 6644 13268 6656
rect 11204 6616 13124 6644
rect 13223 6616 13268 6644
rect 11204 6604 11210 6616
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 13446 6604 13452 6656
rect 13504 6644 13510 6656
rect 14553 6647 14611 6653
rect 14553 6644 14565 6647
rect 13504 6616 14565 6644
rect 13504 6604 13510 6616
rect 14553 6613 14565 6616
rect 14599 6613 14611 6647
rect 14553 6607 14611 6613
rect 15749 6647 15807 6653
rect 15749 6613 15761 6647
rect 15795 6644 15807 6647
rect 17770 6644 17776 6656
rect 15795 6616 17776 6644
rect 15795 6613 15807 6616
rect 15749 6607 15807 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 17954 6604 17960 6656
rect 18012 6644 18018 6656
rect 18049 6647 18107 6653
rect 18049 6644 18061 6647
rect 18012 6616 18061 6644
rect 18012 6604 18018 6616
rect 18049 6613 18061 6616
rect 18095 6613 18107 6647
rect 18049 6607 18107 6613
rect 19245 6647 19303 6653
rect 19245 6613 19257 6647
rect 19291 6644 19303 6647
rect 19978 6644 19984 6656
rect 19291 6616 19984 6644
rect 19291 6613 19303 6616
rect 19245 6607 19303 6613
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 21177 6647 21235 6653
rect 21177 6644 21189 6647
rect 20588 6616 21189 6644
rect 20588 6604 20594 6616
rect 21177 6613 21189 6616
rect 21223 6613 21235 6647
rect 21177 6607 21235 6613
rect 1104 6554 21896 6576
rect 1104 6502 4447 6554
rect 4499 6502 4511 6554
rect 4563 6502 4575 6554
rect 4627 6502 4639 6554
rect 4691 6502 11378 6554
rect 11430 6502 11442 6554
rect 11494 6502 11506 6554
rect 11558 6502 11570 6554
rect 11622 6502 18308 6554
rect 18360 6502 18372 6554
rect 18424 6502 18436 6554
rect 18488 6502 18500 6554
rect 18552 6502 21896 6554
rect 1104 6480 21896 6502
rect 9125 6443 9183 6449
rect 9125 6440 9137 6443
rect 7668 6412 9137 6440
rect 6914 6332 6920 6384
rect 6972 6372 6978 6384
rect 7282 6372 7288 6384
rect 6972 6344 7288 6372
rect 6972 6332 6978 6344
rect 7282 6332 7288 6344
rect 7340 6372 7346 6384
rect 7668 6372 7696 6412
rect 9125 6409 9137 6412
rect 9171 6409 9183 6443
rect 9125 6403 9183 6409
rect 9309 6443 9367 6449
rect 9309 6409 9321 6443
rect 9355 6440 9367 6443
rect 9582 6440 9588 6452
rect 9355 6412 9588 6440
rect 9355 6409 9367 6412
rect 9309 6403 9367 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 13354 6440 13360 6452
rect 12268 6412 13360 6440
rect 7340 6344 7696 6372
rect 7340 6332 7346 6344
rect 8846 6332 8852 6384
rect 8904 6372 8910 6384
rect 12268 6372 12296 6412
rect 13354 6400 13360 6412
rect 13412 6400 13418 6452
rect 13556 6412 14596 6440
rect 8904 6344 12296 6372
rect 12805 6375 12863 6381
rect 8904 6332 8910 6344
rect 12805 6341 12817 6375
rect 12851 6372 12863 6375
rect 12986 6372 12992 6384
rect 12851 6344 12992 6372
rect 12851 6341 12863 6344
rect 12805 6335 12863 6341
rect 12986 6332 12992 6344
rect 13044 6332 13050 6384
rect 13170 6332 13176 6384
rect 13228 6372 13234 6384
rect 13556 6372 13584 6412
rect 13228 6344 13584 6372
rect 13228 6332 13234 6344
rect 7558 6264 7564 6316
rect 7616 6304 7622 6316
rect 7653 6307 7711 6313
rect 7653 6304 7665 6307
rect 7616 6276 7665 6304
rect 7616 6264 7622 6276
rect 7653 6273 7665 6276
rect 7699 6273 7711 6307
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 7653 6267 7711 6273
rect 8772 6276 9873 6304
rect 2222 6196 2228 6248
rect 2280 6236 2286 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 2280 6208 6929 6236
rect 2280 6196 2286 6208
rect 6917 6205 6929 6208
rect 6963 6236 6975 6239
rect 7374 6236 7380 6248
rect 6963 6208 7380 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8772 6236 8800 6276
rect 9861 6273 9873 6276
rect 9907 6304 9919 6307
rect 10870 6304 10876 6316
rect 9907 6276 10876 6304
rect 9907 6273 9919 6276
rect 9861 6267 9919 6273
rect 10870 6264 10876 6276
rect 10928 6264 10934 6316
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12161 6307 12219 6313
rect 12161 6304 12173 6307
rect 12023 6276 12173 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 12161 6273 12173 6276
rect 12207 6273 12219 6307
rect 12161 6267 12219 6273
rect 12345 6307 12403 6313
rect 12345 6273 12357 6307
rect 12391 6304 12403 6307
rect 13446 6304 13452 6316
rect 12391 6276 13452 6304
rect 12391 6273 12403 6276
rect 12345 6267 12403 6273
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 8312 6208 8800 6236
rect 5810 6128 5816 6180
rect 5868 6168 5874 6180
rect 5868 6140 7696 6168
rect 5868 6128 5874 6140
rect 6086 6100 6092 6112
rect 6047 6072 6092 6100
rect 6086 6060 6092 6072
rect 6144 6060 6150 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6641 6103 6699 6109
rect 6641 6100 6653 6103
rect 6328 6072 6653 6100
rect 6328 6060 6334 6072
rect 6641 6069 6653 6072
rect 6687 6100 6699 6103
rect 6914 6100 6920 6112
rect 6687 6072 6920 6100
rect 6687 6069 6699 6072
rect 6641 6063 6699 6069
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 7668 6100 7696 6140
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 7920 6171 7978 6177
rect 7920 6168 7932 6171
rect 7800 6140 7932 6168
rect 7800 6128 7806 6140
rect 7920 6137 7932 6140
rect 7966 6168 7978 6171
rect 8312 6168 8340 6208
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 13722 6236 13728 6248
rect 9456 6208 13728 6236
rect 9456 6196 9462 6208
rect 13722 6196 13728 6208
rect 13780 6196 13786 6248
rect 14366 6196 14372 6248
rect 14424 6236 14430 6248
rect 14461 6239 14519 6245
rect 14461 6236 14473 6239
rect 14424 6208 14473 6236
rect 14424 6196 14430 6208
rect 14461 6205 14473 6208
rect 14507 6205 14519 6239
rect 14568 6236 14596 6412
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 19702 6440 19708 6452
rect 14884 6412 19708 6440
rect 14884 6400 14890 6412
rect 19702 6400 19708 6412
rect 19760 6400 19766 6452
rect 20070 6400 20076 6452
rect 20128 6400 20134 6452
rect 20254 6400 20260 6452
rect 20312 6440 20318 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 20312 6412 20637 6440
rect 20312 6400 20318 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 20088 6372 20116 6400
rect 20349 6375 20407 6381
rect 20349 6372 20361 6375
rect 20088 6344 20361 6372
rect 20349 6341 20361 6344
rect 20395 6341 20407 6375
rect 20349 6335 20407 6341
rect 15286 6304 15292 6316
rect 15247 6276 15292 6304
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 15930 6264 15936 6316
rect 15988 6304 15994 6316
rect 16298 6304 16304 6316
rect 15988 6276 16304 6304
rect 15988 6264 15994 6276
rect 16298 6264 16304 6276
rect 16356 6304 16362 6316
rect 16356 6276 16896 6304
rect 16356 6264 16362 6276
rect 15565 6239 15623 6245
rect 15565 6236 15577 6239
rect 14568 6208 15577 6236
rect 14461 6199 14519 6205
rect 15565 6205 15577 6208
rect 15611 6205 15623 6239
rect 15565 6199 15623 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16868 6236 16896 6276
rect 20070 6264 20076 6316
rect 20128 6304 20134 6316
rect 21177 6307 21235 6313
rect 21177 6304 21189 6307
rect 20128 6276 21189 6304
rect 20128 6264 20134 6276
rect 21177 6273 21189 6276
rect 21223 6273 21235 6307
rect 21177 6267 21235 6273
rect 17313 6239 17371 6245
rect 17313 6236 17325 6239
rect 16868 6208 17325 6236
rect 16209 6199 16267 6205
rect 17313 6205 17325 6208
rect 17359 6205 17371 6239
rect 17313 6199 17371 6205
rect 7966 6140 8340 6168
rect 7966 6137 7978 6140
rect 7920 6131 7978 6137
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 9769 6171 9827 6177
rect 9769 6168 9781 6171
rect 9640 6140 9781 6168
rect 9640 6128 9646 6140
rect 9769 6137 9781 6140
rect 9815 6137 9827 6171
rect 9769 6131 9827 6137
rect 9858 6128 9864 6180
rect 9916 6168 9922 6180
rect 10686 6168 10692 6180
rect 9916 6140 10692 6168
rect 9916 6128 9922 6140
rect 10686 6128 10692 6140
rect 10744 6128 10750 6180
rect 11793 6171 11851 6177
rect 11793 6137 11805 6171
rect 11839 6168 11851 6171
rect 12342 6168 12348 6180
rect 11839 6140 12348 6168
rect 11839 6137 11851 6140
rect 11793 6131 11851 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12437 6171 12495 6177
rect 12437 6137 12449 6171
rect 12483 6168 12495 6171
rect 12483 6140 13584 6168
rect 12483 6137 12495 6140
rect 12437 6131 12495 6137
rect 8846 6100 8852 6112
rect 7668 6072 8852 6100
rect 8846 6060 8852 6072
rect 8904 6060 8910 6112
rect 9030 6100 9036 6112
rect 8991 6072 9036 6100
rect 9030 6060 9036 6072
rect 9088 6060 9094 6112
rect 9125 6103 9183 6109
rect 9125 6069 9137 6103
rect 9171 6100 9183 6103
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9171 6072 9689 6100
rect 9171 6069 9183 6072
rect 9125 6063 9183 6069
rect 9677 6069 9689 6072
rect 9723 6069 9735 6103
rect 9677 6063 9735 6069
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 10321 6103 10379 6109
rect 10321 6100 10333 6103
rect 10100 6072 10333 6100
rect 10100 6060 10106 6072
rect 10321 6069 10333 6072
rect 10367 6069 10379 6103
rect 10778 6100 10784 6112
rect 10739 6072 10784 6100
rect 10321 6063 10379 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 11977 6103 12035 6109
rect 11977 6069 11989 6103
rect 12023 6100 12035 6103
rect 12618 6100 12624 6112
rect 12023 6072 12624 6100
rect 12023 6069 12035 6072
rect 11977 6063 12035 6069
rect 12618 6060 12624 6072
rect 12676 6100 12682 6112
rect 13081 6103 13139 6109
rect 13081 6100 13093 6103
rect 12676 6072 13093 6100
rect 12676 6060 12682 6072
rect 13081 6069 13093 6072
rect 13127 6100 13139 6103
rect 13170 6100 13176 6112
rect 13127 6072 13176 6100
rect 13127 6069 13139 6072
rect 13081 6063 13139 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13556 6100 13584 6140
rect 13906 6128 13912 6180
rect 13964 6168 13970 6180
rect 14194 6171 14252 6177
rect 14194 6168 14206 6171
rect 13964 6140 14206 6168
rect 13964 6128 13970 6140
rect 14194 6137 14206 6140
rect 14240 6137 14252 6171
rect 14194 6131 14252 6137
rect 14550 6128 14556 6180
rect 14608 6168 14614 6180
rect 16224 6168 16252 6199
rect 18874 6196 18880 6248
rect 18932 6236 18938 6248
rect 18969 6239 19027 6245
rect 18969 6236 18981 6239
rect 18932 6208 18981 6236
rect 18932 6196 18938 6208
rect 18969 6205 18981 6208
rect 19015 6205 19027 6239
rect 19236 6239 19294 6245
rect 19236 6236 19248 6239
rect 18969 6199 19027 6205
rect 19168 6208 19248 6236
rect 14608 6140 16252 6168
rect 14608 6128 14614 6140
rect 17402 6128 17408 6180
rect 17460 6168 17466 6180
rect 17558 6171 17616 6177
rect 17558 6168 17570 6171
rect 17460 6140 17570 6168
rect 17460 6128 17466 6140
rect 17558 6137 17570 6140
rect 17604 6137 17616 6171
rect 18782 6168 18788 6180
rect 17558 6131 17616 6137
rect 18616 6140 18788 6168
rect 14737 6103 14795 6109
rect 14737 6100 14749 6103
rect 13556 6072 14749 6100
rect 14737 6069 14749 6072
rect 14783 6069 14795 6103
rect 15470 6100 15476 6112
rect 15431 6072 15476 6100
rect 14737 6063 14795 6069
rect 15470 6060 15476 6072
rect 15528 6060 15534 6112
rect 15933 6103 15991 6109
rect 15933 6069 15945 6103
rect 15979 6100 15991 6103
rect 16206 6100 16212 6112
rect 15979 6072 16212 6100
rect 15979 6069 15991 6072
rect 15933 6063 15991 6069
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 16390 6100 16396 6112
rect 16351 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 17037 6103 17095 6109
rect 17037 6069 17049 6103
rect 17083 6100 17095 6103
rect 18616 6100 18644 6140
rect 18782 6128 18788 6140
rect 18840 6128 18846 6180
rect 17083 6072 18644 6100
rect 18693 6103 18751 6109
rect 17083 6069 17095 6072
rect 17037 6063 17095 6069
rect 18693 6069 18705 6103
rect 18739 6100 18751 6103
rect 19168 6100 19196 6208
rect 19236 6205 19248 6208
rect 19282 6236 19294 6239
rect 20088 6236 20116 6264
rect 20990 6236 20996 6248
rect 19282 6208 20116 6236
rect 20951 6208 20996 6236
rect 19282 6205 19294 6208
rect 19236 6199 19294 6205
rect 20990 6196 20996 6208
rect 21048 6196 21054 6248
rect 21082 6100 21088 6112
rect 18739 6072 19196 6100
rect 21043 6072 21088 6100
rect 18739 6069 18751 6072
rect 18693 6063 18751 6069
rect 21082 6060 21088 6072
rect 21140 6060 21146 6112
rect 1104 6010 21896 6032
rect 1104 5958 7912 6010
rect 7964 5958 7976 6010
rect 8028 5958 8040 6010
rect 8092 5958 8104 6010
rect 8156 5958 14843 6010
rect 14895 5958 14907 6010
rect 14959 5958 14971 6010
rect 15023 5958 15035 6010
rect 15087 5958 21896 6010
rect 1104 5936 21896 5958
rect 1765 5899 1823 5905
rect 1765 5865 1777 5899
rect 1811 5865 1823 5899
rect 5810 5896 5816 5908
rect 5771 5868 5816 5896
rect 1765 5859 1823 5865
rect 1780 5828 1808 5859
rect 5810 5856 5816 5868
rect 5868 5856 5874 5908
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6319 5868 7696 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 6794 5831 6852 5837
rect 6794 5828 6806 5831
rect 1780 5800 6806 5828
rect 6794 5797 6806 5800
rect 6840 5797 6852 5831
rect 7668 5828 7696 5868
rect 7742 5856 7748 5908
rect 7800 5896 7806 5908
rect 7929 5899 7987 5905
rect 7929 5896 7941 5899
rect 7800 5868 7941 5896
rect 7800 5856 7806 5868
rect 7929 5865 7941 5868
rect 7975 5865 7987 5899
rect 8754 5896 8760 5908
rect 8715 5868 8760 5896
rect 7929 5859 7987 5865
rect 8754 5856 8760 5868
rect 8812 5856 8818 5908
rect 9585 5899 9643 5905
rect 9585 5865 9597 5899
rect 9631 5896 9643 5899
rect 9766 5896 9772 5908
rect 9631 5868 9772 5896
rect 9631 5865 9643 5868
rect 9585 5859 9643 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 9953 5899 10011 5905
rect 9953 5865 9965 5899
rect 9999 5896 10011 5899
rect 10502 5896 10508 5908
rect 9999 5868 10508 5896
rect 9999 5865 10011 5868
rect 9953 5859 10011 5865
rect 10502 5856 10508 5868
rect 10560 5856 10566 5908
rect 10686 5856 10692 5908
rect 10744 5896 10750 5908
rect 10744 5868 12434 5896
rect 10744 5856 10750 5868
rect 8386 5828 8392 5840
rect 7668 5800 8392 5828
rect 6794 5791 6852 5797
rect 8386 5788 8392 5800
rect 8444 5788 8450 5840
rect 10042 5788 10048 5840
rect 10100 5828 10106 5840
rect 10100 5800 10145 5828
rect 10100 5788 10106 5800
rect 11790 5788 11796 5840
rect 11848 5837 11854 5840
rect 11848 5828 11860 5837
rect 12406 5828 12434 5868
rect 12618 5856 12624 5908
rect 12676 5896 12682 5908
rect 12802 5896 12808 5908
rect 12676 5868 12808 5896
rect 12676 5856 12682 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 12986 5896 12992 5908
rect 12943 5868 12992 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 12986 5856 12992 5868
rect 13044 5856 13050 5908
rect 13078 5856 13084 5908
rect 13136 5896 13142 5908
rect 13173 5899 13231 5905
rect 13173 5896 13185 5899
rect 13136 5868 13185 5896
rect 13136 5856 13142 5868
rect 13173 5865 13185 5868
rect 13219 5865 13231 5899
rect 13173 5859 13231 5865
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13630 5896 13636 5908
rect 13587 5868 13636 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13722 5856 13728 5908
rect 13780 5896 13786 5908
rect 15933 5899 15991 5905
rect 13780 5868 15884 5896
rect 13780 5856 13786 5868
rect 15470 5828 15476 5840
rect 11848 5800 11893 5828
rect 12406 5800 15476 5828
rect 11848 5791 11860 5800
rect 11848 5788 11854 5791
rect 15470 5788 15476 5800
rect 15528 5788 15534 5840
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5760 1642 5772
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1636 5732 2053 5760
rect 1636 5720 1642 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 2041 5723 2099 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 7558 5760 7564 5772
rect 6595 5732 7564 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7742 5720 7748 5772
rect 7800 5760 7806 5772
rect 8202 5760 8208 5772
rect 7800 5732 8208 5760
rect 7800 5720 7806 5732
rect 8202 5720 8208 5732
rect 8260 5720 8266 5772
rect 8297 5763 8355 5769
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8573 5763 8631 5769
rect 8573 5760 8585 5763
rect 8343 5732 8585 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 8573 5729 8585 5732
rect 8619 5760 8631 5763
rect 12069 5763 12127 5769
rect 8619 5732 10824 5760
rect 8619 5729 8631 5732
rect 8573 5723 8631 5729
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 10137 5695 10195 5701
rect 10137 5692 10149 5695
rect 9088 5664 10149 5692
rect 9088 5652 9094 5664
rect 10137 5661 10149 5664
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10686 5652 10692 5704
rect 10744 5652 10750 5704
rect 10704 5624 10732 5652
rect 7484 5596 10732 5624
rect 7484 5568 7512 5596
rect 6086 5516 6092 5568
rect 6144 5556 6150 5568
rect 7466 5556 7472 5568
rect 6144 5528 7472 5556
rect 6144 5516 6150 5528
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 9309 5559 9367 5565
rect 9309 5525 9321 5559
rect 9355 5556 9367 5559
rect 10134 5556 10140 5568
rect 9355 5528 10140 5556
rect 9355 5525 9367 5528
rect 9309 5519 9367 5525
rect 10134 5516 10140 5528
rect 10192 5516 10198 5568
rect 10686 5556 10692 5568
rect 10647 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10796 5556 10824 5732
rect 12069 5729 12081 5763
rect 12115 5760 12127 5763
rect 12618 5760 12624 5772
rect 12115 5732 12624 5760
rect 12115 5729 12127 5732
rect 12069 5723 12127 5729
rect 12618 5720 12624 5732
rect 12676 5720 12682 5772
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5729 12771 5763
rect 12713 5723 12771 5729
rect 12526 5692 12532 5704
rect 12084 5664 12532 5692
rect 12084 5636 12112 5664
rect 12526 5652 12532 5664
rect 12584 5652 12590 5704
rect 12066 5584 12072 5636
rect 12124 5584 12130 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12728 5624 12756 5723
rect 13262 5720 13268 5772
rect 13320 5760 13326 5772
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 13320 5732 13645 5760
rect 13320 5720 13326 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5760 14611 5763
rect 14734 5760 14740 5772
rect 14599 5732 14740 5760
rect 14599 5729 14611 5732
rect 14553 5723 14611 5729
rect 14734 5720 14740 5732
rect 14792 5720 14798 5772
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15562 5760 15568 5772
rect 15252 5732 15424 5760
rect 15523 5732 15568 5760
rect 15252 5720 15258 5732
rect 13170 5652 13176 5704
rect 13228 5692 13234 5704
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13228 5664 13737 5692
rect 13228 5652 13234 5664
rect 13725 5661 13737 5664
rect 13771 5661 13783 5695
rect 15286 5692 15292 5704
rect 15247 5664 15292 5692
rect 13725 5655 13783 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15396 5692 15424 5732
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 15856 5760 15884 5868
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 15979 5868 16681 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 17310 5896 17316 5908
rect 17271 5868 17316 5896
rect 16669 5859 16727 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17862 5856 17868 5908
rect 17920 5896 17926 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 17920 5868 20177 5896
rect 17920 5856 17926 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 20165 5859 20223 5865
rect 20346 5856 20352 5908
rect 20404 5896 20410 5908
rect 20533 5899 20591 5905
rect 20533 5896 20545 5899
rect 20404 5868 20545 5896
rect 20404 5856 20410 5868
rect 20533 5865 20545 5868
rect 20579 5865 20591 5899
rect 20533 5859 20591 5865
rect 16206 5788 16212 5840
rect 16264 5828 16270 5840
rect 16577 5831 16635 5837
rect 16577 5828 16589 5831
rect 16264 5800 16589 5828
rect 16264 5788 16270 5800
rect 16577 5797 16589 5800
rect 16623 5797 16635 5831
rect 16577 5791 16635 5797
rect 18448 5831 18506 5837
rect 18448 5797 18460 5831
rect 18494 5828 18506 5831
rect 19794 5828 19800 5840
rect 18494 5800 19800 5828
rect 18494 5797 18506 5800
rect 18448 5791 18506 5797
rect 19794 5788 19800 5800
rect 19852 5788 19858 5840
rect 20070 5788 20076 5840
rect 20128 5788 20134 5840
rect 20622 5788 20628 5840
rect 20680 5828 20686 5840
rect 21177 5831 21235 5837
rect 21177 5828 21189 5831
rect 20680 5800 21189 5828
rect 20680 5788 20686 5800
rect 21177 5797 21189 5800
rect 21223 5797 21235 5831
rect 21177 5791 21235 5797
rect 19153 5763 19211 5769
rect 19153 5760 19165 5763
rect 15856 5732 19165 5760
rect 19153 5729 19165 5732
rect 19199 5760 19211 5763
rect 20088 5760 20116 5788
rect 19199 5732 19334 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 15473 5695 15531 5701
rect 15473 5692 15485 5695
rect 15396 5664 15485 5692
rect 15473 5661 15485 5664
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 16482 5652 16488 5704
rect 16540 5692 16546 5704
rect 16761 5695 16819 5701
rect 16761 5692 16773 5695
rect 16540 5664 16773 5692
rect 16540 5652 16546 5664
rect 16761 5661 16773 5664
rect 16807 5661 16819 5695
rect 16761 5655 16819 5661
rect 18693 5695 18751 5701
rect 18693 5661 18705 5695
rect 18739 5692 18751 5695
rect 18874 5692 18880 5704
rect 18739 5664 18880 5692
rect 18739 5661 18751 5664
rect 18693 5655 18751 5661
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 14182 5624 14188 5636
rect 12492 5596 12537 5624
rect 12728 5596 14188 5624
rect 12492 5584 12498 5596
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 14568 5596 14872 5624
rect 14568 5556 14596 5596
rect 14734 5556 14740 5568
rect 10796 5528 14596 5556
rect 14695 5528 14740 5556
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 14844 5556 14872 5596
rect 16114 5584 16120 5636
rect 16172 5624 16178 5636
rect 16209 5627 16267 5633
rect 16209 5624 16221 5627
rect 16172 5596 16221 5624
rect 16172 5584 16178 5596
rect 16209 5593 16221 5596
rect 16255 5593 16267 5627
rect 19306 5624 19334 5732
rect 19996 5732 20116 5760
rect 19996 5701 20024 5732
rect 19981 5695 20039 5701
rect 19981 5661 19993 5695
rect 20027 5661 20039 5695
rect 19981 5655 20039 5661
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5661 20131 5695
rect 20073 5655 20131 5661
rect 20088 5624 20116 5655
rect 20990 5624 20996 5636
rect 19306 5596 20116 5624
rect 20951 5596 20996 5624
rect 16209 5587 16267 5593
rect 20990 5584 20996 5596
rect 21048 5584 21054 5636
rect 18690 5556 18696 5568
rect 14844 5528 18696 5556
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 18966 5556 18972 5568
rect 18927 5528 18972 5556
rect 18966 5516 18972 5528
rect 19024 5516 19030 5568
rect 1104 5466 21896 5488
rect 1104 5414 4447 5466
rect 4499 5414 4511 5466
rect 4563 5414 4575 5466
rect 4627 5414 4639 5466
rect 4691 5414 11378 5466
rect 11430 5414 11442 5466
rect 11494 5414 11506 5466
rect 11558 5414 11570 5466
rect 11622 5414 18308 5466
rect 18360 5414 18372 5466
rect 18424 5414 18436 5466
rect 18488 5414 18500 5466
rect 18552 5414 21896 5466
rect 1104 5392 21896 5414
rect 5718 5312 5724 5364
rect 5776 5352 5782 5364
rect 6641 5355 6699 5361
rect 6641 5352 6653 5355
rect 5776 5324 6653 5352
rect 5776 5312 5782 5324
rect 6641 5321 6653 5324
rect 6687 5352 6699 5355
rect 9214 5352 9220 5364
rect 6687 5324 9220 5352
rect 6687 5321 6699 5324
rect 6641 5315 6699 5321
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 10318 5352 10324 5364
rect 10279 5324 10324 5352
rect 10318 5312 10324 5324
rect 10376 5312 10382 5364
rect 10413 5355 10471 5361
rect 10413 5321 10425 5355
rect 10459 5352 10471 5355
rect 18598 5352 18604 5364
rect 10459 5324 18604 5352
rect 10459 5321 10471 5324
rect 10413 5315 10471 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 5997 5287 6055 5293
rect 5997 5284 6009 5287
rect 5868 5256 6009 5284
rect 5868 5244 5874 5256
rect 5997 5253 6009 5256
rect 6043 5253 6055 5287
rect 5997 5247 6055 5253
rect 7377 5287 7435 5293
rect 7377 5253 7389 5287
rect 7423 5284 7435 5287
rect 7558 5284 7564 5296
rect 7423 5256 7564 5284
rect 7423 5253 7435 5256
rect 7377 5247 7435 5253
rect 7558 5244 7564 5256
rect 7616 5244 7622 5296
rect 7745 5287 7803 5293
rect 7745 5253 7757 5287
rect 7791 5284 7803 5287
rect 8294 5284 8300 5296
rect 7791 5256 8300 5284
rect 7791 5253 7803 5256
rect 7745 5247 7803 5253
rect 8294 5244 8300 5256
rect 8352 5284 8358 5296
rect 9030 5284 9036 5296
rect 8352 5256 9036 5284
rect 8352 5244 8358 5256
rect 9030 5244 9036 5256
rect 9088 5284 9094 5296
rect 9306 5284 9312 5296
rect 9088 5256 9312 5284
rect 9088 5244 9094 5256
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 9861 5287 9919 5293
rect 9861 5253 9873 5287
rect 9907 5253 9919 5287
rect 9861 5247 9919 5253
rect 10505 5287 10563 5293
rect 10505 5253 10517 5287
rect 10551 5284 10563 5287
rect 12802 5284 12808 5296
rect 10551 5256 12808 5284
rect 10551 5253 10563 5256
rect 10505 5247 10563 5253
rect 8481 5219 8539 5225
rect 8481 5185 8493 5219
rect 8527 5216 8539 5219
rect 9876 5216 9904 5247
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 16117 5287 16175 5293
rect 16117 5253 16129 5287
rect 16163 5253 16175 5287
rect 16117 5247 16175 5253
rect 8527 5188 9720 5216
rect 9876 5188 10640 5216
rect 8527 5185 8539 5188
rect 8481 5179 8539 5185
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 8757 5151 8815 5157
rect 8757 5148 8769 5151
rect 8628 5120 8769 5148
rect 8628 5108 8634 5120
rect 8757 5117 8769 5120
rect 8803 5117 8815 5151
rect 8757 5111 8815 5117
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5148 9275 5151
rect 9306 5148 9312 5160
rect 9263 5120 9312 5148
rect 9263 5117 9275 5120
rect 9217 5111 9275 5117
rect 7009 5083 7067 5089
rect 7009 5049 7021 5083
rect 7055 5080 7067 5083
rect 7282 5080 7288 5092
rect 7055 5052 7288 5080
rect 7055 5049 7067 5052
rect 7009 5043 7067 5049
rect 7282 5040 7288 5052
rect 7340 5040 7346 5092
rect 8113 5083 8171 5089
rect 8113 5049 8125 5083
rect 8159 5080 8171 5083
rect 9232 5080 9260 5111
rect 9306 5108 9312 5120
rect 9364 5108 9370 5160
rect 9692 5157 9720 5188
rect 9677 5151 9735 5157
rect 9677 5117 9689 5151
rect 9723 5148 9735 5151
rect 9953 5151 10011 5157
rect 9953 5148 9965 5151
rect 9723 5120 9965 5148
rect 9723 5117 9735 5120
rect 9677 5111 9735 5117
rect 9953 5117 9965 5120
rect 9999 5117 10011 5151
rect 10134 5148 10140 5160
rect 10047 5120 10140 5148
rect 9953 5111 10011 5117
rect 10134 5108 10140 5120
rect 10192 5148 10198 5160
rect 10505 5151 10563 5157
rect 10505 5148 10517 5151
rect 10192 5120 10517 5148
rect 10192 5108 10198 5120
rect 10505 5117 10517 5120
rect 10551 5117 10563 5151
rect 10612 5148 10640 5188
rect 10686 5176 10692 5228
rect 10744 5216 10750 5228
rect 10781 5219 10839 5225
rect 10781 5216 10793 5219
rect 10744 5188 10793 5216
rect 10744 5176 10750 5188
rect 10781 5185 10793 5188
rect 10827 5216 10839 5219
rect 12526 5216 12532 5228
rect 10827 5188 12532 5216
rect 10827 5185 10839 5188
rect 10781 5179 10839 5185
rect 12526 5176 12532 5188
rect 12584 5176 12590 5228
rect 16132 5216 16160 5247
rect 17126 5244 17132 5296
rect 17184 5284 17190 5296
rect 19613 5287 19671 5293
rect 19613 5284 19625 5287
rect 17184 5256 19625 5284
rect 17184 5244 17190 5256
rect 19613 5253 19625 5256
rect 19659 5253 19671 5287
rect 19613 5247 19671 5253
rect 19794 5244 19800 5296
rect 19852 5284 19858 5296
rect 19852 5256 21220 5284
rect 19852 5244 19858 5256
rect 21192 5228 21220 5256
rect 16482 5216 16488 5228
rect 16132 5188 16488 5216
rect 16482 5176 16488 5188
rect 16540 5216 16546 5228
rect 17681 5219 17739 5225
rect 17681 5216 17693 5219
rect 16540 5188 17693 5216
rect 16540 5176 16546 5188
rect 17681 5185 17693 5188
rect 17727 5185 17739 5219
rect 17681 5179 17739 5185
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19944 5188 20085 5216
rect 19944 5176 19950 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20530 5216 20536 5228
rect 20303 5188 20536 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20530 5176 20536 5188
rect 20588 5176 20594 5228
rect 21174 5216 21180 5228
rect 21087 5188 21180 5216
rect 21174 5176 21180 5188
rect 21232 5176 21238 5228
rect 10873 5151 10931 5157
rect 10873 5148 10885 5151
rect 10612 5120 10885 5148
rect 10505 5111 10563 5117
rect 10873 5117 10885 5120
rect 10919 5148 10931 5151
rect 11698 5148 11704 5160
rect 10919 5120 11704 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11698 5108 11704 5120
rect 11756 5108 11762 5160
rect 11882 5108 11888 5160
rect 11940 5148 11946 5160
rect 12345 5151 12403 5157
rect 12345 5148 12357 5151
rect 11940 5120 12357 5148
rect 11940 5108 11946 5120
rect 12345 5117 12357 5120
rect 12391 5117 12403 5151
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 12345 5111 12403 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 14366 5108 14372 5160
rect 14424 5148 14430 5160
rect 14642 5148 14648 5160
rect 14424 5120 14648 5148
rect 14424 5108 14430 5120
rect 14642 5108 14648 5120
rect 14700 5148 14706 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14700 5120 14749 5148
rect 14700 5108 14706 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 15004 5151 15062 5157
rect 15004 5117 15016 5151
rect 15050 5148 15062 5151
rect 15286 5148 15292 5160
rect 15050 5120 15292 5148
rect 15050 5117 15062 5120
rect 15004 5111 15062 5117
rect 11146 5080 11152 5092
rect 8159 5052 9260 5080
rect 9416 5052 11152 5080
rect 8159 5049 8171 5052
rect 8113 5043 8171 5049
rect 8570 4972 8576 5024
rect 8628 5012 8634 5024
rect 9416 5021 9444 5052
rect 11146 5040 11152 5052
rect 11204 5040 11210 5092
rect 11422 5040 11428 5092
rect 11480 5080 11486 5092
rect 13348 5083 13406 5089
rect 11480 5052 12388 5080
rect 11480 5040 11486 5052
rect 8941 5015 8999 5021
rect 8941 5012 8953 5015
rect 8628 4984 8953 5012
rect 8628 4972 8634 4984
rect 8941 4981 8953 4984
rect 8987 4981 8999 5015
rect 8941 4975 8999 4981
rect 9401 5015 9459 5021
rect 9401 4981 9413 5015
rect 9447 4981 9459 5015
rect 9401 4975 9459 4981
rect 9953 5015 10011 5021
rect 9953 4981 9965 5015
rect 9999 5012 10011 5015
rect 10413 5015 10471 5021
rect 10413 5012 10425 5015
rect 9999 4984 10425 5012
rect 9999 4981 10011 4984
rect 9953 4975 10011 4981
rect 10413 4981 10425 4984
rect 10459 4981 10471 5015
rect 10962 5012 10968 5024
rect 10923 4984 10968 5012
rect 10413 4975 10471 4981
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11238 4972 11244 5024
rect 11296 5012 11302 5024
rect 11333 5015 11391 5021
rect 11333 5012 11345 5015
rect 11296 4984 11345 5012
rect 11296 4972 11302 4984
rect 11333 4981 11345 4984
rect 11379 4981 11391 5015
rect 11333 4975 11391 4981
rect 11698 4972 11704 5024
rect 11756 5012 11762 5024
rect 11885 5015 11943 5021
rect 11885 5012 11897 5015
rect 11756 4984 11897 5012
rect 11756 4972 11762 4984
rect 11885 4981 11897 4984
rect 11931 4981 11943 5015
rect 11885 4975 11943 4981
rect 12066 4972 12072 5024
rect 12124 5012 12130 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 12124 4984 12265 5012
rect 12124 4972 12130 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12360 5012 12388 5052
rect 13348 5049 13360 5083
rect 13394 5080 13406 5083
rect 13446 5080 13452 5092
rect 13394 5052 13452 5080
rect 13394 5049 13406 5052
rect 13348 5043 13406 5049
rect 13446 5040 13452 5052
rect 13504 5040 13510 5092
rect 12618 5012 12624 5024
rect 12360 4984 12624 5012
rect 12253 4975 12311 4981
rect 12618 4972 12624 4984
rect 12676 5012 12682 5024
rect 13078 5012 13084 5024
rect 12676 4984 13084 5012
rect 12676 4972 12682 4984
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 14461 5015 14519 5021
rect 14461 4981 14473 5015
rect 14507 5012 14519 5015
rect 15028 5012 15056 5111
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 19978 5148 19984 5160
rect 19939 5120 19984 5148
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 16577 5083 16635 5089
rect 16577 5049 16589 5083
rect 16623 5080 16635 5083
rect 17497 5083 17555 5089
rect 17497 5080 17509 5083
rect 16623 5052 17509 5080
rect 16623 5049 16635 5052
rect 16577 5043 16635 5049
rect 17497 5049 17509 5052
rect 17543 5049 17555 5083
rect 17497 5043 17555 5049
rect 17586 5040 17592 5092
rect 17644 5080 17650 5092
rect 18233 5083 18291 5089
rect 17644 5052 17689 5080
rect 17644 5040 17650 5052
rect 18233 5049 18245 5083
rect 18279 5080 18291 5083
rect 19242 5080 19248 5092
rect 18279 5052 19248 5080
rect 18279 5049 18291 5052
rect 18233 5043 18291 5049
rect 19242 5040 19248 5052
rect 19300 5040 19306 5092
rect 19337 5083 19395 5089
rect 19337 5049 19349 5083
rect 19383 5080 19395 5083
rect 20993 5083 21051 5089
rect 20993 5080 21005 5083
rect 19383 5052 21005 5080
rect 19383 5049 19395 5052
rect 19337 5043 19395 5049
rect 20993 5049 21005 5052
rect 21039 5049 21051 5083
rect 20993 5043 21051 5049
rect 17126 5012 17132 5024
rect 14507 4984 15056 5012
rect 17087 4984 17132 5012
rect 14507 4981 14519 4984
rect 14461 4975 14519 4981
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 18693 5015 18751 5021
rect 18693 4981 18705 5015
rect 18739 5012 18751 5015
rect 19058 5012 19064 5024
rect 18739 4984 19064 5012
rect 18739 4981 18751 4984
rect 18693 4975 18751 4981
rect 19058 4972 19064 4984
rect 19116 4972 19122 5024
rect 20622 5012 20628 5024
rect 20583 4984 20628 5012
rect 20622 4972 20628 4984
rect 20680 4972 20686 5024
rect 21082 4972 21088 5024
rect 21140 5012 21146 5024
rect 21140 4984 21185 5012
rect 21140 4972 21146 4984
rect 1104 4922 21896 4944
rect 1104 4870 7912 4922
rect 7964 4870 7976 4922
rect 8028 4870 8040 4922
rect 8092 4870 8104 4922
rect 8156 4870 14843 4922
rect 14895 4870 14907 4922
rect 14959 4870 14971 4922
rect 15023 4870 15035 4922
rect 15087 4870 21896 4922
rect 1104 4848 21896 4870
rect 6178 4808 6184 4820
rect 6139 4780 6184 4808
rect 6178 4768 6184 4780
rect 6236 4768 6242 4820
rect 6549 4811 6607 4817
rect 6549 4777 6561 4811
rect 6595 4808 6607 4811
rect 6914 4808 6920 4820
rect 6595 4780 6920 4808
rect 6595 4777 6607 4780
rect 6549 4771 6607 4777
rect 6914 4768 6920 4780
rect 6972 4768 6978 4820
rect 7285 4811 7343 4817
rect 7285 4777 7297 4811
rect 7331 4808 7343 4811
rect 8294 4808 8300 4820
rect 7331 4780 8300 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 8294 4768 8300 4780
rect 8352 4768 8358 4820
rect 8570 4768 8576 4820
rect 8628 4768 8634 4820
rect 9306 4768 9312 4820
rect 9364 4808 9370 4820
rect 17313 4811 17371 4817
rect 9364 4780 17264 4808
rect 9364 4768 9370 4780
rect 6825 4743 6883 4749
rect 6825 4709 6837 4743
rect 6871 4740 6883 4743
rect 7558 4740 7564 4752
rect 6871 4712 7564 4740
rect 6871 4709 6883 4712
rect 6825 4703 6883 4709
rect 7558 4700 7564 4712
rect 7616 4740 7622 4752
rect 8386 4740 8392 4752
rect 7616 4712 8392 4740
rect 7616 4700 7622 4712
rect 8386 4700 8392 4712
rect 8444 4700 8450 4752
rect 8588 4740 8616 4768
rect 11241 4743 11299 4749
rect 8588 4712 11192 4740
rect 8757 4675 8815 4681
rect 8757 4641 8769 4675
rect 8803 4672 8815 4675
rect 9306 4672 9312 4684
rect 8803 4644 9312 4672
rect 8803 4641 8815 4644
rect 8757 4635 8815 4641
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9858 4672 9864 4684
rect 9646 4644 9864 4672
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 9646 4604 9674 4644
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 10036 4675 10094 4681
rect 10036 4641 10048 4675
rect 10082 4672 10094 4675
rect 10594 4672 10600 4684
rect 10082 4644 10600 4672
rect 10082 4641 10094 4644
rect 10036 4635 10094 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11164 4672 11192 4712
rect 11241 4709 11253 4743
rect 11287 4740 11299 4743
rect 11670 4743 11728 4749
rect 11670 4740 11682 4743
rect 11287 4712 11682 4740
rect 11287 4709 11299 4712
rect 11241 4703 11299 4709
rect 11670 4709 11682 4712
rect 11716 4709 11728 4743
rect 14366 4740 14372 4752
rect 11670 4703 11728 4709
rect 11900 4712 14372 4740
rect 11900 4672 11928 4712
rect 14366 4700 14372 4712
rect 14424 4740 14430 4752
rect 14642 4740 14648 4752
rect 14424 4712 14648 4740
rect 14424 4700 14430 4712
rect 14642 4700 14648 4712
rect 14700 4700 14706 4752
rect 14734 4700 14740 4752
rect 14792 4740 14798 4752
rect 15013 4743 15071 4749
rect 15013 4740 15025 4743
rect 14792 4712 15025 4740
rect 14792 4700 14798 4712
rect 15013 4709 15025 4712
rect 15059 4709 15071 4743
rect 15013 4703 15071 4709
rect 16200 4743 16258 4749
rect 16200 4709 16212 4743
rect 16246 4740 16258 4743
rect 16482 4740 16488 4752
rect 16246 4712 16488 4740
rect 16246 4709 16258 4712
rect 16200 4703 16258 4709
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 17236 4740 17264 4780
rect 17313 4777 17325 4811
rect 17359 4808 17371 4811
rect 17402 4808 17408 4820
rect 17359 4780 17408 4808
rect 17359 4777 17371 4780
rect 17313 4771 17371 4777
rect 17402 4768 17408 4780
rect 17460 4768 17466 4820
rect 18138 4808 18144 4820
rect 17512 4780 18144 4808
rect 17512 4740 17540 4780
rect 18138 4768 18144 4780
rect 18196 4768 18202 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 19705 4811 19763 4817
rect 19705 4808 19717 4811
rect 18932 4780 19717 4808
rect 18932 4768 18938 4780
rect 19705 4777 19717 4780
rect 19751 4777 19763 4811
rect 21174 4808 21180 4820
rect 21135 4780 21180 4808
rect 19705 4771 19763 4777
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 17770 4740 17776 4752
rect 17236 4712 17540 4740
rect 17731 4712 17776 4740
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 18693 4743 18751 4749
rect 18693 4709 18705 4743
rect 18739 4740 18751 4743
rect 22094 4740 22100 4752
rect 18739 4712 22100 4740
rect 18739 4709 18751 4712
rect 18693 4703 18751 4709
rect 22094 4700 22100 4712
rect 22152 4700 22158 4752
rect 11164 4644 11928 4672
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 12492 4644 13369 4672
rect 12492 4632 12498 4644
rect 13357 4641 13369 4644
rect 13403 4641 13415 4675
rect 13906 4672 13912 4684
rect 13867 4644 13912 4672
rect 13357 4635 13415 4641
rect 13906 4632 13912 4644
rect 13964 4632 13970 4684
rect 15565 4675 15623 4681
rect 15565 4641 15577 4675
rect 15611 4641 15623 4675
rect 18506 4672 18512 4684
rect 18467 4644 18512 4672
rect 15565 4635 15623 4641
rect 6972 4576 9674 4604
rect 9769 4607 9827 4613
rect 6972 4564 6978 4576
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 11422 4604 11428 4616
rect 9769 4567 9827 4573
rect 10796 4576 11428 4604
rect 8846 4496 8852 4548
rect 8904 4536 8910 4548
rect 9398 4536 9404 4548
rect 8904 4508 9404 4536
rect 8904 4496 8910 4508
rect 9398 4496 9404 4508
rect 9456 4496 9462 4548
rect 7650 4468 7656 4480
rect 7611 4440 7656 4468
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8294 4468 8300 4480
rect 8067 4440 8300 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8389 4471 8447 4477
rect 8389 4437 8401 4471
rect 8435 4468 8447 4471
rect 8938 4468 8944 4480
rect 8435 4440 8944 4468
rect 8435 4437 8447 4440
rect 8389 4431 8447 4437
rect 8938 4428 8944 4440
rect 8996 4428 9002 4480
rect 9493 4471 9551 4477
rect 9493 4437 9505 4471
rect 9539 4468 9551 4471
rect 9674 4468 9680 4480
rect 9539 4440 9680 4468
rect 9539 4437 9551 4440
rect 9493 4431 9551 4437
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9784 4468 9812 4567
rect 10796 4468 10824 4576
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 15580 4604 15608 4635
rect 18506 4632 18512 4644
rect 18564 4632 18570 4684
rect 18782 4632 18788 4684
rect 18840 4672 18846 4684
rect 20070 4681 20076 4684
rect 19061 4675 19119 4681
rect 19061 4672 19073 4675
rect 18840 4644 19073 4672
rect 18840 4632 18846 4644
rect 19061 4641 19073 4644
rect 19107 4641 19119 4675
rect 19061 4635 19119 4641
rect 19705 4675 19763 4681
rect 19705 4641 19717 4675
rect 19751 4672 19763 4675
rect 19797 4675 19855 4681
rect 19797 4672 19809 4675
rect 19751 4644 19809 4672
rect 19751 4641 19763 4644
rect 19705 4635 19763 4641
rect 19797 4641 19809 4644
rect 19843 4641 19855 4675
rect 19797 4635 19855 4641
rect 20064 4635 20076 4681
rect 20128 4672 20134 4684
rect 20128 4644 20164 4672
rect 20070 4632 20076 4635
rect 20128 4632 20134 4644
rect 15930 4604 15936 4616
rect 12728 4576 15608 4604
rect 15891 4576 15936 4604
rect 11146 4536 11152 4548
rect 11059 4508 11152 4536
rect 11146 4496 11152 4508
rect 11204 4536 11210 4548
rect 11241 4539 11299 4545
rect 11241 4536 11253 4539
rect 11204 4508 11253 4536
rect 11204 4496 11210 4508
rect 11241 4505 11253 4508
rect 11287 4505 11299 4539
rect 11241 4499 11299 4505
rect 9784 4440 10824 4468
rect 10962 4428 10968 4480
rect 11020 4468 11026 4480
rect 12728 4468 12756 4576
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 18138 4564 18144 4616
rect 18196 4604 18202 4616
rect 18874 4604 18880 4616
rect 18196 4576 18880 4604
rect 18196 4564 18202 4576
rect 18874 4564 18880 4576
rect 18932 4564 18938 4616
rect 19150 4604 19156 4616
rect 19076 4576 19156 4604
rect 13170 4536 13176 4548
rect 13131 4508 13176 4536
rect 13170 4496 13176 4508
rect 13228 4496 13234 4548
rect 13722 4536 13728 4548
rect 13683 4508 13728 4536
rect 13722 4496 13728 4508
rect 13780 4496 13786 4548
rect 14734 4496 14740 4548
rect 14792 4536 14798 4548
rect 14829 4539 14887 4545
rect 14829 4536 14841 4539
rect 14792 4508 14841 4536
rect 14792 4496 14798 4508
rect 14829 4505 14841 4508
rect 14875 4505 14887 4539
rect 15378 4536 15384 4548
rect 15339 4508 15384 4536
rect 14829 4499 14887 4505
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 17034 4496 17040 4548
rect 17092 4536 17098 4548
rect 17589 4539 17647 4545
rect 17589 4536 17601 4539
rect 17092 4508 17601 4536
rect 17092 4496 17098 4508
rect 17589 4505 17601 4508
rect 17635 4505 17647 4539
rect 17589 4499 17647 4505
rect 11020 4440 12756 4468
rect 12805 4471 12863 4477
rect 11020 4428 11026 4440
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 13446 4468 13452 4480
rect 12851 4440 13452 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 13446 4428 13452 4440
rect 13504 4428 13510 4480
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 19076 4468 19104 4576
rect 19150 4564 19156 4576
rect 19208 4564 19214 4616
rect 14599 4440 19104 4468
rect 19153 4471 19211 4477
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 19153 4437 19165 4471
rect 19199 4468 19211 4471
rect 21542 4468 21548 4480
rect 19199 4440 21548 4468
rect 19199 4437 19211 4440
rect 19153 4431 19211 4437
rect 21542 4428 21548 4440
rect 21600 4428 21606 4480
rect 1104 4378 21896 4400
rect 1104 4326 4447 4378
rect 4499 4326 4511 4378
rect 4563 4326 4575 4378
rect 4627 4326 4639 4378
rect 4691 4326 11378 4378
rect 11430 4326 11442 4378
rect 11494 4326 11506 4378
rect 11558 4326 11570 4378
rect 11622 4326 18308 4378
rect 18360 4326 18372 4378
rect 18424 4326 18436 4378
rect 18488 4326 18500 4378
rect 18552 4326 21896 4378
rect 1104 4304 21896 4326
rect 5718 4264 5724 4276
rect 5679 4236 5724 4264
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9548 4236 9593 4264
rect 9548 4224 9554 4236
rect 10594 4224 10600 4276
rect 10652 4264 10658 4276
rect 18690 4264 18696 4276
rect 10652 4236 18696 4264
rect 10652 4224 10658 4236
rect 18690 4224 18696 4236
rect 18748 4224 18754 4276
rect 20717 4267 20775 4273
rect 20717 4233 20729 4267
rect 20763 4264 20775 4267
rect 21082 4264 21088 4276
rect 20763 4236 21088 4264
rect 20763 4233 20775 4236
rect 20717 4227 20775 4233
rect 21082 4224 21088 4236
rect 21140 4224 21146 4276
rect 8294 4156 8300 4208
rect 8352 4196 8358 4208
rect 9674 4196 9680 4208
rect 8352 4168 9680 4196
rect 8352 4156 8358 4168
rect 9674 4156 9680 4168
rect 9732 4156 9738 4208
rect 10042 4156 10048 4208
rect 10100 4196 10106 4208
rect 10502 4196 10508 4208
rect 10100 4168 10508 4196
rect 10100 4156 10106 4168
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 11146 4196 11152 4208
rect 10796 4168 11152 4196
rect 6546 4128 6552 4140
rect 6507 4100 6552 4128
rect 6546 4088 6552 4100
rect 6604 4088 6610 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4128 7711 4131
rect 10318 4128 10324 4140
rect 7699 4100 10324 4128
rect 7699 4097 7711 4100
rect 7653 4091 7711 4097
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 10796 4137 10824 4168
rect 11146 4156 11152 4168
rect 11204 4156 11210 4208
rect 12897 4199 12955 4205
rect 12897 4196 12909 4199
rect 11256 4168 12909 4196
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 11256 4128 11284 4168
rect 12897 4165 12909 4168
rect 12943 4165 12955 4199
rect 17402 4196 17408 4208
rect 12897 4159 12955 4165
rect 16408 4168 17408 4196
rect 12342 4128 12348 4140
rect 10781 4091 10839 4097
rect 10888 4100 11284 4128
rect 12303 4100 12348 4128
rect 6917 4063 6975 4069
rect 6917 4029 6929 4063
rect 6963 4060 6975 4063
rect 8018 4060 8024 4072
rect 6963 4032 8024 4060
rect 6963 4029 6975 4032
rect 6917 4023 6975 4029
rect 8018 4020 8024 4032
rect 8076 4020 8082 4072
rect 8294 4060 8300 4072
rect 8255 4032 8300 4060
rect 8294 4020 8300 4032
rect 8352 4020 8358 4072
rect 8757 4063 8815 4069
rect 8757 4029 8769 4063
rect 8803 4029 8815 4063
rect 8757 4023 8815 4029
rect 9217 4063 9275 4069
rect 9217 4029 9229 4063
rect 9263 4060 9275 4063
rect 9493 4063 9551 4069
rect 9493 4060 9505 4063
rect 9263 4032 9505 4060
rect 9263 4029 9275 4032
rect 9217 4023 9275 4029
rect 9493 4029 9505 4032
rect 9539 4029 9551 4063
rect 9493 4023 9551 4029
rect 9701 4063 9759 4069
rect 9701 4029 9713 4063
rect 9747 4060 9759 4063
rect 9950 4060 9956 4072
rect 9747 4032 9956 4060
rect 9747 4029 9759 4032
rect 9701 4023 9759 4029
rect 4154 3952 4160 4004
rect 4212 3992 4218 4004
rect 7193 3995 7251 4001
rect 7193 3992 7205 3995
rect 4212 3964 7205 3992
rect 4212 3952 4218 3964
rect 7193 3961 7205 3964
rect 7239 3992 7251 3995
rect 8772 3992 8800 4023
rect 9950 4020 9956 4032
rect 10008 4020 10014 4072
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10888 4060 10916 4100
rect 12342 4088 12348 4100
rect 12400 4088 12406 4140
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 13446 4128 13452 4140
rect 13407 4100 13452 4128
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 14550 4128 14556 4140
rect 14511 4100 14556 4128
rect 14550 4088 14556 4100
rect 14608 4088 14614 4140
rect 16206 4128 16212 4140
rect 16167 4100 16212 4128
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 16408 4137 16436 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 17494 4156 17500 4208
rect 17552 4196 17558 4208
rect 18138 4196 18144 4208
rect 17552 4168 18144 4196
rect 17552 4156 17558 4168
rect 18138 4156 18144 4168
rect 18196 4196 18202 4208
rect 19705 4199 19763 4205
rect 18196 4168 18368 4196
rect 18196 4156 18202 4168
rect 16393 4131 16451 4137
rect 16393 4097 16405 4131
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 16482 4088 16488 4140
rect 16540 4128 16546 4140
rect 18340 4137 18368 4168
rect 19705 4165 19717 4199
rect 19751 4165 19763 4199
rect 19705 4159 19763 4165
rect 17681 4131 17739 4137
rect 17681 4128 17693 4131
rect 16540 4100 17693 4128
rect 16540 4088 16546 4100
rect 17681 4097 17693 4100
rect 17727 4097 17739 4131
rect 17681 4091 17739 4097
rect 18325 4131 18383 4137
rect 18325 4097 18337 4131
rect 18371 4097 18383 4131
rect 19720 4128 19748 4159
rect 20070 4128 20076 4140
rect 19720 4100 20076 4128
rect 18325 4091 18383 4097
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 10192 4032 10237 4060
rect 10336 4032 10916 4060
rect 10965 4063 11023 4069
rect 10192 4020 10198 4032
rect 10336 3992 10364 4032
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11698 4060 11704 4072
rect 11011 4032 11704 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11698 4020 11704 4032
rect 11756 4020 11762 4072
rect 11793 4063 11851 4069
rect 11793 4029 11805 4063
rect 11839 4060 11851 4063
rect 13265 4063 13323 4069
rect 13265 4060 13277 4063
rect 11839 4032 13277 4060
rect 11839 4029 11851 4032
rect 11793 4023 11851 4029
rect 13265 4029 13277 4032
rect 13311 4029 13323 4063
rect 13265 4023 13323 4029
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14075 4063 14133 4069
rect 14075 4060 14087 4063
rect 13872 4032 14087 4060
rect 13872 4020 13878 4032
rect 14075 4029 14087 4032
rect 14121 4029 14133 4063
rect 14075 4023 14133 4029
rect 14274 4020 14280 4072
rect 14332 4060 14338 4072
rect 15013 4063 15071 4069
rect 15013 4060 15025 4063
rect 14332 4032 15025 4060
rect 14332 4020 14338 4032
rect 15013 4029 15025 4032
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 16117 4063 16175 4069
rect 16117 4029 16129 4063
rect 16163 4060 16175 4063
rect 17126 4060 17132 4072
rect 16163 4032 17132 4060
rect 16163 4029 16175 4032
rect 16117 4023 16175 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 21266 4060 21272 4072
rect 17276 4032 18276 4060
rect 21227 4032 21272 4060
rect 17276 4020 17282 4032
rect 7239 3964 8340 3992
rect 8772 3964 10364 3992
rect 10873 3995 10931 4001
rect 7239 3961 7251 3964
rect 7193 3955 7251 3961
rect 8312 3936 8340 3964
rect 10873 3961 10885 3995
rect 10919 3992 10931 3995
rect 10919 3964 11928 3992
rect 10919 3961 10931 3964
rect 10873 3955 10931 3961
rect 6089 3927 6147 3933
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 7282 3924 7288 3936
rect 6135 3896 7288 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8202 3924 8208 3936
rect 8067 3896 8208 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8294 3884 8300 3936
rect 8352 3884 8358 3936
rect 8478 3924 8484 3936
rect 8439 3896 8484 3924
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 8938 3924 8944 3936
rect 8899 3896 8944 3924
rect 8938 3884 8944 3896
rect 8996 3884 9002 3936
rect 9401 3927 9459 3933
rect 9401 3893 9413 3927
rect 9447 3924 9459 3927
rect 9766 3924 9772 3936
rect 9447 3896 9772 3924
rect 9447 3893 9459 3896
rect 9401 3887 9459 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3924 9919 3927
rect 10134 3924 10140 3936
rect 9907 3896 10140 3924
rect 9907 3893 9919 3896
rect 9861 3887 9919 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10321 3927 10379 3933
rect 10321 3893 10333 3927
rect 10367 3924 10379 3927
rect 10778 3924 10784 3936
rect 10367 3896 10784 3924
rect 10367 3893 10379 3896
rect 10321 3887 10379 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 11900 3933 11928 3964
rect 11974 3952 11980 4004
rect 12032 3992 12038 4004
rect 13357 3995 13415 4001
rect 13357 3992 13369 3995
rect 12032 3964 13369 3992
rect 12032 3952 12038 3964
rect 13357 3961 13369 3964
rect 13403 3961 13415 3995
rect 14642 3992 14648 4004
rect 14603 3964 14648 3992
rect 13357 3955 13415 3961
rect 14642 3952 14648 3964
rect 14700 3952 14706 4004
rect 15194 3992 15200 4004
rect 15155 3964 15200 3992
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 17313 3995 17371 4001
rect 17313 3992 17325 3995
rect 15344 3964 17325 3992
rect 15344 3952 15350 3964
rect 17313 3961 17325 3964
rect 17359 3961 17371 3995
rect 17313 3955 17371 3961
rect 17586 3952 17592 4004
rect 17644 3992 17650 4004
rect 17865 3995 17923 4001
rect 17865 3992 17877 3995
rect 17644 3964 17877 3992
rect 17644 3952 17650 3964
rect 17865 3961 17877 3964
rect 17911 3961 17923 3995
rect 17865 3955 17923 3961
rect 11333 3927 11391 3933
rect 11333 3893 11345 3927
rect 11379 3924 11391 3927
rect 11793 3927 11851 3933
rect 11793 3924 11805 3927
rect 11379 3896 11805 3924
rect 11379 3893 11391 3896
rect 11333 3887 11391 3893
rect 11793 3893 11805 3896
rect 11839 3893 11851 3927
rect 11793 3887 11851 3893
rect 11885 3927 11943 3933
rect 11885 3893 11897 3927
rect 11931 3893 11943 3927
rect 11885 3887 11943 3893
rect 12066 3884 12072 3936
rect 12124 3924 12130 3936
rect 12250 3924 12256 3936
rect 12124 3896 12256 3924
rect 12124 3884 12130 3896
rect 12250 3884 12256 3896
rect 12308 3884 12314 3936
rect 13998 3884 14004 3936
rect 14056 3924 14062 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 14056 3896 14565 3924
rect 14056 3884 14062 3896
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 15746 3924 15752 3936
rect 15707 3896 15752 3924
rect 14553 3887 14611 3893
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 17221 3927 17279 3933
rect 17221 3924 17233 3927
rect 16080 3896 17233 3924
rect 16080 3884 16086 3896
rect 17221 3893 17233 3896
rect 17267 3893 17279 3927
rect 18248 3924 18276 4032
rect 21266 4020 21272 4032
rect 21324 4020 21330 4072
rect 18592 3995 18650 4001
rect 18592 3961 18604 3995
rect 18638 3992 18650 3995
rect 18874 3992 18880 4004
rect 18638 3964 18880 3992
rect 18638 3961 18650 3964
rect 18592 3955 18650 3961
rect 18874 3952 18880 3964
rect 18932 3952 18938 4004
rect 21085 3995 21143 4001
rect 21085 3992 21097 3995
rect 20272 3964 21097 3992
rect 20272 3933 20300 3964
rect 21085 3961 21097 3964
rect 21131 3961 21143 3995
rect 21085 3955 21143 3961
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 18248 3896 20269 3924
rect 17221 3887 17279 3893
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20257 3887 20315 3893
rect 20346 3884 20352 3936
rect 20404 3924 20410 3936
rect 20404 3896 20449 3924
rect 20404 3884 20410 3896
rect 1104 3834 21896 3856
rect 1104 3782 7912 3834
rect 7964 3782 7976 3834
rect 8028 3782 8040 3834
rect 8092 3782 8104 3834
rect 8156 3782 14843 3834
rect 14895 3782 14907 3834
rect 14959 3782 14971 3834
rect 15023 3782 15035 3834
rect 15087 3782 21896 3834
rect 1104 3760 21896 3782
rect 5353 3723 5411 3729
rect 5353 3689 5365 3723
rect 5399 3720 5411 3723
rect 7006 3720 7012 3732
rect 5399 3692 7012 3720
rect 5399 3689 5411 3692
rect 5353 3683 5411 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7282 3680 7288 3732
rect 7340 3720 7346 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 7340 3692 7941 3720
rect 7340 3680 7346 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 9677 3723 9735 3729
rect 9677 3720 9689 3723
rect 7929 3683 7987 3689
rect 8266 3692 9689 3720
rect 6641 3655 6699 3661
rect 6641 3621 6653 3655
rect 6687 3652 6699 3655
rect 7190 3652 7196 3664
rect 6687 3624 7196 3652
rect 6687 3621 6699 3624
rect 6641 3615 6699 3621
rect 7190 3612 7196 3624
rect 7248 3652 7254 3664
rect 8266 3652 8294 3692
rect 9677 3689 9689 3692
rect 9723 3689 9735 3723
rect 9677 3683 9735 3689
rect 10413 3723 10471 3729
rect 10413 3689 10425 3723
rect 10459 3720 10471 3723
rect 10962 3720 10968 3732
rect 10459 3692 10968 3720
rect 10459 3689 10471 3692
rect 10413 3683 10471 3689
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 11238 3680 11244 3732
rect 11296 3720 11302 3732
rect 11517 3723 11575 3729
rect 11517 3720 11529 3723
rect 11296 3692 11529 3720
rect 11296 3680 11302 3692
rect 11517 3689 11529 3692
rect 11563 3689 11575 3723
rect 11517 3683 11575 3689
rect 11698 3680 11704 3732
rect 11756 3720 11762 3732
rect 12161 3723 12219 3729
rect 12161 3720 12173 3723
rect 11756 3692 12173 3720
rect 11756 3680 11762 3692
rect 12161 3689 12173 3692
rect 12207 3689 12219 3723
rect 13998 3720 14004 3732
rect 13959 3692 14004 3720
rect 12161 3683 12219 3689
rect 13998 3680 14004 3692
rect 14056 3680 14062 3732
rect 15746 3720 15752 3732
rect 14090 3692 15752 3720
rect 14090 3652 14118 3692
rect 15746 3680 15752 3692
rect 15804 3680 15810 3732
rect 15838 3680 15844 3732
rect 15896 3720 15902 3732
rect 16574 3720 16580 3732
rect 15896 3692 16580 3720
rect 15896 3680 15902 3692
rect 16574 3680 16580 3692
rect 16632 3680 16638 3732
rect 16669 3723 16727 3729
rect 16669 3689 16681 3723
rect 16715 3720 16727 3723
rect 18598 3720 18604 3732
rect 16715 3692 18604 3720
rect 16715 3689 16727 3692
rect 16669 3683 16727 3689
rect 18598 3680 18604 3692
rect 18656 3680 18662 3732
rect 18874 3720 18880 3732
rect 18835 3692 18880 3720
rect 18874 3680 18880 3692
rect 18932 3680 18938 3732
rect 19150 3680 19156 3732
rect 19208 3720 19214 3732
rect 20622 3720 20628 3732
rect 19208 3692 20628 3720
rect 19208 3680 19214 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 7248 3624 8294 3652
rect 8588 3624 14118 3652
rect 7248 3612 7254 3624
rect 4985 3587 5043 3593
rect 4985 3553 4997 3587
rect 5031 3584 5043 3587
rect 7742 3584 7748 3596
rect 5031 3556 7748 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 7742 3544 7748 3556
rect 7800 3544 7806 3596
rect 7926 3544 7932 3596
rect 7984 3584 7990 3596
rect 8588 3593 8616 3624
rect 14642 3612 14648 3664
rect 14700 3652 14706 3664
rect 14798 3655 14856 3661
rect 14798 3652 14810 3655
rect 14700 3624 14810 3652
rect 14700 3612 14706 3624
rect 14798 3621 14810 3624
rect 14844 3621 14856 3655
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 14798 3615 14856 3621
rect 15580 3624 19993 3652
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7984 3556 8125 3584
rect 7984 3544 7990 3556
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8113 3547 8171 3553
rect 8573 3587 8631 3593
rect 8573 3553 8585 3587
rect 8619 3553 8631 3587
rect 8846 3584 8852 3596
rect 8807 3556 8852 3584
rect 8573 3547 8631 3553
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 9030 3544 9036 3596
rect 9088 3584 9094 3596
rect 9309 3587 9367 3593
rect 9309 3584 9321 3587
rect 9088 3556 9321 3584
rect 9088 3544 9094 3556
rect 9309 3553 9321 3556
rect 9355 3553 9367 3587
rect 9309 3547 9367 3553
rect 9677 3587 9735 3593
rect 9677 3553 9689 3587
rect 9723 3584 9735 3587
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 9723 3556 9781 3584
rect 9723 3553 9735 3556
rect 9677 3547 9735 3553
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 10229 3587 10287 3593
rect 10229 3553 10241 3587
rect 10275 3584 10287 3587
rect 10502 3584 10508 3596
rect 10275 3556 10508 3584
rect 10275 3553 10287 3556
rect 10229 3547 10287 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 10686 3584 10692 3596
rect 10647 3556 10692 3584
rect 10686 3544 10692 3556
rect 10744 3544 10750 3596
rect 12434 3584 12440 3596
rect 10796 3556 12440 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5629 3519 5687 3525
rect 5629 3516 5641 3519
rect 5316 3488 5641 3516
rect 5316 3476 5322 3488
rect 5629 3485 5641 3488
rect 5675 3485 5687 3519
rect 5629 3479 5687 3485
rect 7834 3476 7840 3528
rect 7892 3516 7898 3528
rect 10042 3516 10048 3528
rect 7892 3488 10048 3516
rect 7892 3476 7898 3488
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 10796 3516 10824 3556
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 12802 3584 12808 3596
rect 12763 3556 12808 3584
rect 12802 3544 12808 3556
rect 12860 3544 12866 3596
rect 13633 3587 13691 3593
rect 13633 3584 13645 3587
rect 13004 3556 13645 3584
rect 10652 3488 10824 3516
rect 10652 3476 10658 3488
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 11241 3519 11299 3525
rect 11241 3516 11253 3519
rect 11204 3488 11253 3516
rect 11204 3476 11210 3488
rect 11241 3485 11253 3488
rect 11287 3485 11299 3519
rect 11241 3479 11299 3485
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3516 11483 3519
rect 11606 3516 11612 3528
rect 11471 3488 11612 3516
rect 11471 3485 11483 3488
rect 11425 3479 11483 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 12342 3476 12348 3528
rect 12400 3516 12406 3528
rect 13004 3516 13032 3556
rect 13633 3553 13645 3556
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 14366 3544 14372 3596
rect 14424 3584 14430 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14424 3556 14565 3584
rect 14424 3544 14430 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 12400 3488 13032 3516
rect 12400 3476 12406 3488
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13357 3519 13415 3525
rect 13357 3516 13369 3519
rect 13320 3488 13369 3516
rect 13320 3476 13326 3488
rect 13357 3485 13369 3488
rect 13403 3485 13415 3519
rect 13357 3479 13415 3485
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 14090 3516 14096 3528
rect 13587 3488 14096 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 1765 3451 1823 3457
rect 1765 3448 1777 3451
rect 1360 3420 1777 3448
rect 1360 3408 1366 3420
rect 1765 3417 1777 3420
rect 1811 3417 1823 3451
rect 1765 3411 1823 3417
rect 6546 3408 6552 3460
rect 6604 3448 6610 3460
rect 8110 3448 8116 3460
rect 6604 3420 8116 3448
rect 6604 3408 6610 3420
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8297 3451 8355 3457
rect 8297 3417 8309 3451
rect 8343 3448 8355 3451
rect 8343 3420 9352 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 5868 3352 6193 3380
rect 5868 3340 5874 3352
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6181 3343 6239 3349
rect 7009 3383 7067 3389
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7098 3380 7104 3392
rect 7055 3352 7104 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7098 3340 7104 3352
rect 7156 3340 7162 3392
rect 7282 3380 7288 3392
rect 7243 3352 7288 3380
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7616 3352 7757 3380
rect 7616 3340 7622 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7926 3380 7932 3392
rect 7887 3352 7932 3380
rect 7745 3343 7803 3349
rect 7926 3340 7932 3352
rect 7984 3340 7990 3392
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8386 3380 8392 3392
rect 8076 3352 8392 3380
rect 8076 3340 8082 3352
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8757 3383 8815 3389
rect 8757 3349 8769 3383
rect 8803 3380 8815 3383
rect 8849 3383 8907 3389
rect 8849 3380 8861 3383
rect 8803 3352 8861 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 8849 3349 8861 3352
rect 8895 3349 8907 3383
rect 9324 3380 9352 3420
rect 9398 3408 9404 3460
rect 9456 3448 9462 3460
rect 9493 3451 9551 3457
rect 9493 3448 9505 3451
rect 9456 3420 9505 3448
rect 9456 3408 9462 3420
rect 9493 3417 9505 3420
rect 9539 3417 9551 3451
rect 9493 3411 9551 3417
rect 9953 3451 10011 3457
rect 9953 3417 9965 3451
rect 9999 3448 10011 3451
rect 12618 3448 12624 3460
rect 9999 3420 12480 3448
rect 12579 3420 12624 3448
rect 9999 3417 10011 3420
rect 9953 3411 10011 3417
rect 10042 3380 10048 3392
rect 9324 3352 10048 3380
rect 8849 3343 8907 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 10873 3383 10931 3389
rect 10873 3349 10885 3383
rect 10919 3380 10931 3383
rect 11790 3380 11796 3392
rect 10919 3352 11796 3380
rect 10919 3349 10931 3352
rect 10873 3343 10931 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 11885 3383 11943 3389
rect 11885 3349 11897 3383
rect 11931 3380 11943 3383
rect 11974 3380 11980 3392
rect 11931 3352 11980 3380
rect 11931 3349 11943 3352
rect 11885 3343 11943 3349
rect 11974 3340 11980 3352
rect 12032 3340 12038 3392
rect 12452 3380 12480 3420
rect 12618 3408 12624 3420
rect 12676 3408 12682 3460
rect 15580 3380 15608 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 19981 3615 20039 3621
rect 20438 3612 20444 3664
rect 20496 3652 20502 3664
rect 20533 3655 20591 3661
rect 20533 3652 20545 3655
rect 20496 3624 20545 3652
rect 20496 3612 20502 3624
rect 20533 3621 20545 3624
rect 20579 3621 20591 3655
rect 20898 3652 20904 3664
rect 20533 3615 20591 3621
rect 20640 3624 20904 3652
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 17586 3584 17592 3596
rect 16448 3556 17592 3584
rect 16448 3544 16454 3556
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17764 3587 17822 3593
rect 17764 3553 17776 3587
rect 17810 3584 17822 3587
rect 18138 3584 18144 3596
rect 17810 3556 18144 3584
rect 17810 3553 17822 3556
rect 17764 3547 17822 3553
rect 18138 3544 18144 3556
rect 18196 3544 18202 3596
rect 18690 3544 18696 3596
rect 18748 3584 18754 3596
rect 20640 3584 20668 3624
rect 20898 3612 20904 3624
rect 20956 3652 20962 3664
rect 21269 3655 21327 3661
rect 21269 3652 21281 3655
rect 20956 3624 21281 3652
rect 20956 3612 20962 3624
rect 21269 3621 21281 3624
rect 21315 3621 21327 3655
rect 21269 3615 21327 3621
rect 18748 3556 20668 3584
rect 18748 3544 18754 3556
rect 20714 3544 20720 3596
rect 20772 3584 20778 3596
rect 20772 3556 20817 3584
rect 20772 3544 20778 3556
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 16761 3519 16819 3525
rect 16761 3516 16773 3519
rect 16632 3488 16773 3516
rect 16632 3476 16638 3488
rect 16761 3485 16773 3488
rect 16807 3485 16819 3519
rect 16942 3516 16948 3528
rect 16903 3488 16948 3516
rect 16761 3479 16819 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 17126 3476 17132 3528
rect 17184 3516 17190 3528
rect 17494 3516 17500 3528
rect 17184 3488 17500 3516
rect 17184 3476 17190 3488
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 20732 3516 20760 3544
rect 18524 3488 20760 3516
rect 15930 3380 15936 3392
rect 12452 3352 15608 3380
rect 15891 3352 15936 3380
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16298 3380 16304 3392
rect 16259 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 17310 3340 17316 3392
rect 17368 3380 17374 3392
rect 18524 3380 18552 3488
rect 19334 3408 19340 3460
rect 19392 3448 19398 3460
rect 19797 3451 19855 3457
rect 19797 3448 19809 3451
rect 19392 3420 19809 3448
rect 19392 3408 19398 3420
rect 19797 3417 19809 3420
rect 19843 3417 19855 3451
rect 19797 3411 19855 3417
rect 19150 3380 19156 3392
rect 17368 3352 18552 3380
rect 19111 3352 19156 3380
rect 17368 3340 17374 3352
rect 19150 3340 19156 3352
rect 19208 3340 19214 3392
rect 19242 3340 19248 3392
rect 19300 3380 19306 3392
rect 20806 3380 20812 3392
rect 19300 3352 20812 3380
rect 19300 3340 19306 3352
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 21174 3380 21180 3392
rect 21135 3352 21180 3380
rect 21174 3340 21180 3352
rect 21232 3340 21238 3392
rect 1104 3290 21896 3312
rect 1104 3238 4447 3290
rect 4499 3238 4511 3290
rect 4563 3238 4575 3290
rect 4627 3238 4639 3290
rect 4691 3238 11378 3290
rect 11430 3238 11442 3290
rect 11494 3238 11506 3290
rect 11558 3238 11570 3290
rect 11622 3238 18308 3290
rect 18360 3238 18372 3290
rect 18424 3238 18436 3290
rect 18488 3238 18500 3290
rect 18552 3238 21896 3290
rect 1104 3216 21896 3238
rect 4893 3179 4951 3185
rect 4893 3145 4905 3179
rect 4939 3176 4951 3179
rect 9306 3176 9312 3188
rect 4939 3148 9312 3176
rect 4939 3145 4951 3148
rect 4893 3139 4951 3145
rect 9306 3136 9312 3148
rect 9364 3136 9370 3188
rect 9766 3136 9772 3188
rect 9824 3176 9830 3188
rect 10597 3179 10655 3185
rect 10597 3176 10609 3179
rect 9824 3148 10609 3176
rect 9824 3136 9830 3148
rect 10597 3145 10609 3148
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10873 3179 10931 3185
rect 10873 3145 10885 3179
rect 10919 3176 10931 3179
rect 12802 3176 12808 3188
rect 10919 3148 12808 3176
rect 10919 3145 10931 3148
rect 10873 3139 10931 3145
rect 12802 3136 12808 3148
rect 12860 3136 12866 3188
rect 13262 3176 13268 3188
rect 13223 3148 13268 3176
rect 13262 3136 13268 3148
rect 13320 3136 13326 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14240 3148 14596 3176
rect 14240 3136 14246 3148
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 4430 3108 4436 3120
rect 1627 3080 2774 3108
rect 4391 3080 4436 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 2746 3040 2774 3080
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 6089 3111 6147 3117
rect 6089 3077 6101 3111
rect 6135 3108 6147 3111
rect 10502 3108 10508 3120
rect 6135 3080 10508 3108
rect 6135 3077 6147 3080
rect 6089 3071 6147 3077
rect 10502 3068 10508 3080
rect 10560 3068 10566 3120
rect 6914 3040 6920 3052
rect 2746 3012 6920 3040
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7834 3040 7840 3052
rect 7156 3012 7512 3040
rect 7795 3012 7840 3040
rect 7156 3000 7162 3012
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1302 2972 1308 2984
rect 900 2944 1308 2972
rect 900 2932 906 2944
rect 1302 2932 1308 2944
rect 1360 2972 1366 2984
rect 1397 2975 1455 2981
rect 1397 2972 1409 2975
rect 1360 2944 1409 2972
rect 1360 2932 1366 2944
rect 1397 2941 1409 2944
rect 1443 2941 1455 2975
rect 1397 2935 1455 2941
rect 1486 2932 1492 2984
rect 1544 2972 1550 2984
rect 1857 2975 1915 2981
rect 1857 2972 1869 2975
rect 1544 2944 1869 2972
rect 1544 2932 1550 2944
rect 1857 2941 1869 2944
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 1872 2904 1900 2935
rect 1946 2932 1952 2984
rect 2004 2972 2010 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2004 2944 2789 2972
rect 2004 2932 2010 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 4706 2972 4712 2984
rect 4619 2944 4712 2972
rect 2777 2935 2835 2941
rect 4706 2932 4712 2944
rect 4764 2972 4770 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 4764 2944 5549 2972
rect 4764 2932 4770 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 7006 2972 7012 2984
rect 6919 2944 7012 2972
rect 5537 2935 5595 2941
rect 7006 2932 7012 2944
rect 7064 2972 7070 2984
rect 7282 2972 7288 2984
rect 7064 2944 7288 2972
rect 7064 2932 7070 2944
rect 7282 2932 7288 2944
rect 7340 2932 7346 2984
rect 7484 2981 7512 3012
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 8110 3000 8116 3052
rect 8168 3040 8174 3052
rect 8168 3012 8892 3040
rect 8168 3000 8174 3012
rect 7469 2975 7527 2981
rect 7469 2941 7481 2975
rect 7515 2941 7527 2975
rect 7926 2972 7932 2984
rect 7887 2944 7932 2972
rect 7469 2935 7527 2941
rect 2317 2907 2375 2913
rect 2317 2904 2329 2907
rect 1872 2876 2329 2904
rect 2317 2873 2329 2876
rect 2363 2873 2375 2907
rect 2317 2867 2375 2873
rect 2498 2864 2504 2916
rect 2556 2904 2562 2916
rect 3053 2907 3111 2913
rect 3053 2904 3065 2907
rect 2556 2876 3065 2904
rect 2556 2864 2562 2876
rect 3053 2873 3065 2876
rect 3099 2873 3111 2907
rect 7484 2904 7512 2935
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 8018 2932 8024 2984
rect 8076 2972 8082 2984
rect 8389 2975 8447 2981
rect 8389 2972 8401 2975
rect 8076 2944 8401 2972
rect 8076 2932 8082 2944
rect 8389 2941 8401 2944
rect 8435 2941 8447 2975
rect 8389 2935 8447 2941
rect 8478 2932 8484 2984
rect 8536 2972 8542 2984
rect 8754 2972 8760 2984
rect 8536 2944 8760 2972
rect 8536 2932 8542 2944
rect 8754 2932 8760 2944
rect 8812 2932 8818 2984
rect 8864 2981 8892 3012
rect 8938 3000 8944 3052
rect 8996 3040 9002 3052
rect 8996 3012 9812 3040
rect 8996 3000 9002 3012
rect 8849 2975 8907 2981
rect 8849 2941 8861 2975
rect 8895 2941 8907 2975
rect 9306 2972 9312 2984
rect 9267 2944 9312 2972
rect 8849 2935 8907 2941
rect 9306 2932 9312 2944
rect 9364 2932 9370 2984
rect 9784 2981 9812 3012
rect 10134 3000 10140 3052
rect 10192 3040 10198 3052
rect 11885 3043 11943 3049
rect 10192 3012 11192 3040
rect 10192 3000 10198 3012
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2941 9827 2975
rect 9769 2935 9827 2941
rect 10042 2932 10048 2984
rect 10100 2972 10106 2984
rect 11164 2981 11192 3012
rect 11885 3009 11897 3043
rect 11931 3040 11943 3043
rect 13280 3040 13308 3136
rect 14568 3108 14596 3148
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 14921 3179 14979 3185
rect 14921 3176 14933 3179
rect 14700 3148 14933 3176
rect 14700 3136 14706 3148
rect 14921 3145 14933 3148
rect 14967 3145 14979 3179
rect 14921 3139 14979 3145
rect 15212 3148 18092 3176
rect 15212 3108 15240 3148
rect 14568 3080 15240 3108
rect 16577 3111 16635 3117
rect 16577 3077 16589 3111
rect 16623 3108 16635 3111
rect 16761 3111 16819 3117
rect 16761 3108 16773 3111
rect 16623 3080 16773 3108
rect 16623 3077 16635 3080
rect 16577 3071 16635 3077
rect 16761 3077 16773 3080
rect 16807 3108 16819 3111
rect 16942 3108 16948 3120
rect 16807 3080 16948 3108
rect 16807 3077 16819 3080
rect 16761 3071 16819 3077
rect 16942 3068 16948 3080
rect 17000 3068 17006 3120
rect 18064 3108 18092 3148
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 18509 3179 18567 3185
rect 18509 3176 18521 3179
rect 18196 3148 18521 3176
rect 18196 3136 18202 3148
rect 18509 3145 18521 3148
rect 18555 3145 18567 3179
rect 21174 3176 21180 3188
rect 18509 3139 18567 3145
rect 18708 3148 21180 3176
rect 18708 3108 18736 3148
rect 21174 3136 21180 3148
rect 21232 3136 21238 3188
rect 21358 3108 21364 3120
rect 18064 3080 18736 3108
rect 18800 3080 21364 3108
rect 15013 3043 15071 3049
rect 11931 3012 12020 3040
rect 13280 3012 13676 3040
rect 11931 3009 11943 3012
rect 11885 3003 11943 3009
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 10100 2944 10241 2972
rect 10100 2932 10106 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 10229 2935 10287 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10689 2975 10747 2981
rect 10689 2972 10701 2975
rect 10643 2944 10701 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 10689 2941 10701 2944
rect 10735 2941 10747 2975
rect 10689 2935 10747 2941
rect 11149 2975 11207 2981
rect 11149 2941 11161 2975
rect 11195 2941 11207 2975
rect 11149 2935 11207 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 11992 2972 12020 3012
rect 13078 2972 13084 2984
rect 11756 2944 11928 2972
rect 11992 2944 13084 2972
rect 11756 2932 11762 2944
rect 9214 2904 9220 2916
rect 7484 2876 9220 2904
rect 3053 2867 3111 2873
rect 9214 2864 9220 2876
rect 9272 2864 9278 2916
rect 11900 2904 11928 2944
rect 13078 2932 13084 2944
rect 13136 2972 13142 2984
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 13136 2944 13553 2972
rect 13136 2932 13142 2944
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13648 2972 13676 3012
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15102 3040 15108 3052
rect 15059 3012 15108 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 16666 3000 16672 3052
rect 16724 3040 16730 3052
rect 16724 3012 17264 3040
rect 16724 3000 16730 3012
rect 13797 2975 13855 2981
rect 13797 2972 13809 2975
rect 13648 2944 13809 2972
rect 13541 2935 13599 2941
rect 13797 2941 13809 2944
rect 13843 2941 13855 2975
rect 13797 2935 13855 2941
rect 14366 2932 14372 2984
rect 14424 2972 14430 2984
rect 15197 2975 15255 2981
rect 15197 2972 15209 2975
rect 14424 2944 15209 2972
rect 14424 2932 14430 2944
rect 15197 2941 15209 2944
rect 15243 2941 15255 2975
rect 15197 2935 15255 2941
rect 15464 2975 15522 2981
rect 15464 2941 15476 2975
rect 15510 2972 15522 2975
rect 15930 2972 15936 2984
rect 15510 2944 15936 2972
rect 15510 2941 15522 2944
rect 15464 2935 15522 2941
rect 12130 2907 12188 2913
rect 12130 2904 12142 2907
rect 9968 2876 11836 2904
rect 11900 2876 12142 2904
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 3142 2796 3148 2848
rect 3200 2836 3206 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 3200 2808 3433 2836
rect 3200 2796 3206 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 3602 2796 3608 2848
rect 3660 2836 3666 2848
rect 3973 2839 4031 2845
rect 3973 2836 3985 2839
rect 3660 2808 3985 2836
rect 3660 2796 3666 2808
rect 3973 2805 3985 2808
rect 4019 2836 4031 2839
rect 4154 2836 4160 2848
rect 4019 2808 4160 2836
rect 4019 2805 4031 2808
rect 3973 2799 4031 2805
rect 4154 2796 4160 2808
rect 4212 2796 4218 2848
rect 5166 2836 5172 2848
rect 5127 2808 5172 2836
rect 5166 2796 5172 2808
rect 5224 2796 5230 2848
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 6549 2839 6607 2845
rect 6549 2836 6561 2839
rect 6512 2808 6561 2836
rect 6512 2796 6518 2808
rect 6549 2805 6561 2808
rect 6595 2805 6607 2839
rect 6549 2799 6607 2805
rect 7193 2839 7251 2845
rect 7193 2805 7205 2839
rect 7239 2836 7251 2839
rect 7466 2836 7472 2848
rect 7239 2808 7472 2836
rect 7239 2805 7251 2808
rect 7193 2799 7251 2805
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 7653 2839 7711 2845
rect 7653 2805 7665 2839
rect 7699 2836 7711 2839
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 7699 2808 7849 2836
rect 7699 2805 7711 2808
rect 7653 2799 7711 2805
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 7837 2799 7895 2805
rect 8113 2839 8171 2845
rect 8113 2805 8125 2839
rect 8159 2836 8171 2839
rect 8478 2836 8484 2848
rect 8159 2808 8484 2836
rect 8159 2805 8171 2808
rect 8113 2799 8171 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 9030 2836 9036 2848
rect 8628 2808 8673 2836
rect 8991 2808 9036 2836
rect 8628 2796 8634 2808
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9493 2839 9551 2845
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9582 2836 9588 2848
rect 9539 2808 9588 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9968 2845 9996 2876
rect 9953 2839 10011 2845
rect 9953 2805 9965 2839
rect 9999 2805 10011 2839
rect 9953 2799 10011 2805
rect 10413 2839 10471 2845
rect 10413 2805 10425 2839
rect 10459 2836 10471 2839
rect 10686 2836 10692 2848
rect 10459 2808 10692 2836
rect 10459 2805 10471 2808
rect 10413 2799 10471 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 11333 2839 11391 2845
rect 11333 2805 11345 2839
rect 11379 2836 11391 2839
rect 11698 2836 11704 2848
rect 11379 2808 11704 2836
rect 11379 2805 11391 2808
rect 11333 2799 11391 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 11808 2836 11836 2876
rect 12130 2873 12142 2876
rect 12176 2873 12188 2907
rect 12130 2867 12188 2873
rect 12250 2864 12256 2916
rect 12308 2904 12314 2916
rect 13906 2904 13912 2916
rect 12308 2876 13912 2904
rect 12308 2864 12314 2876
rect 13906 2864 13912 2876
rect 13964 2864 13970 2916
rect 15212 2904 15240 2935
rect 15930 2932 15936 2944
rect 15988 2932 15994 2984
rect 17126 2972 17132 2984
rect 16592 2944 17132 2972
rect 16592 2904 16620 2944
rect 17126 2932 17132 2944
rect 17184 2932 17190 2984
rect 17236 2972 17264 3012
rect 18506 3000 18512 3052
rect 18564 3040 18570 3052
rect 18800 3040 18828 3080
rect 18564 3012 18828 3040
rect 18564 3000 18570 3012
rect 18874 3000 18880 3052
rect 18932 3040 18938 3052
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 18932 3012 19349 3040
rect 18932 3000 18938 3012
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 19337 3003 19395 3009
rect 19613 3043 19671 3049
rect 19613 3009 19625 3043
rect 19659 3040 19671 3043
rect 20533 3043 20591 3049
rect 20533 3040 20545 3043
rect 19659 3012 20545 3040
rect 19659 3009 19671 3012
rect 19613 3003 19671 3009
rect 20533 3009 20545 3012
rect 20579 3009 20591 3043
rect 20533 3003 20591 3009
rect 20806 3000 20812 3052
rect 20864 3040 20870 3052
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 20864 3012 21097 3040
rect 20864 3000 20870 3012
rect 21085 3009 21097 3012
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 17236 2944 18828 2972
rect 15212 2876 16620 2904
rect 16761 2907 16819 2913
rect 16761 2873 16773 2907
rect 16807 2904 16819 2907
rect 17374 2907 17432 2913
rect 17374 2904 17386 2907
rect 16807 2876 17386 2904
rect 16807 2873 16819 2876
rect 16761 2867 16819 2873
rect 17374 2873 17386 2876
rect 17420 2873 17432 2907
rect 18800 2904 18828 2944
rect 19058 2932 19064 2984
rect 19116 2972 19122 2984
rect 19153 2975 19211 2981
rect 19153 2972 19165 2975
rect 19116 2944 19165 2972
rect 19116 2932 19122 2944
rect 19153 2941 19165 2944
rect 19199 2941 19211 2975
rect 19153 2935 19211 2941
rect 19242 2932 19248 2984
rect 19300 2972 19306 2984
rect 19300 2944 19345 2972
rect 19300 2932 19306 2944
rect 20622 2932 20628 2984
rect 20680 2972 20686 2984
rect 21284 2981 21312 3080
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 20717 2975 20775 2981
rect 20717 2972 20729 2975
rect 20680 2944 20729 2972
rect 20680 2932 20686 2944
rect 20717 2941 20729 2944
rect 20763 2941 20775 2975
rect 20717 2935 20775 2941
rect 21269 2975 21327 2981
rect 21269 2941 21281 2975
rect 21315 2941 21327 2975
rect 21269 2935 21327 2941
rect 19613 2907 19671 2913
rect 19613 2904 19625 2907
rect 18800 2876 19625 2904
rect 17374 2867 17432 2873
rect 19613 2873 19625 2876
rect 19659 2873 19671 2907
rect 19794 2904 19800 2916
rect 19755 2876 19800 2904
rect 19613 2867 19671 2873
rect 19794 2864 19800 2876
rect 19852 2864 19858 2916
rect 19981 2907 20039 2913
rect 19981 2873 19993 2907
rect 20027 2873 20039 2907
rect 19981 2867 20039 2873
rect 15013 2839 15071 2845
rect 15013 2836 15025 2839
rect 11808 2808 15025 2836
rect 15013 2805 15025 2808
rect 15059 2805 15071 2839
rect 18782 2836 18788 2848
rect 18743 2808 18788 2836
rect 15013 2799 15071 2805
rect 18782 2796 18788 2808
rect 18840 2796 18846 2848
rect 19702 2796 19708 2848
rect 19760 2836 19766 2848
rect 19996 2836 20024 2867
rect 19760 2808 20024 2836
rect 19760 2796 19766 2808
rect 1104 2746 21896 2768
rect 1104 2694 7912 2746
rect 7964 2694 7976 2746
rect 8028 2694 8040 2746
rect 8092 2694 8104 2746
rect 8156 2694 14843 2746
rect 14895 2694 14907 2746
rect 14959 2694 14971 2746
rect 15023 2694 15035 2746
rect 15087 2694 21896 2746
rect 1104 2672 21896 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 4062 2632 4068 2644
rect 1627 2604 4068 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 4062 2592 4068 2604
rect 4120 2592 4126 2644
rect 4246 2632 4252 2644
rect 4207 2604 4252 2632
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4798 2632 4804 2644
rect 4759 2604 4804 2632
rect 4798 2592 4804 2604
rect 4856 2592 4862 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 8662 2632 8668 2644
rect 6963 2604 8668 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 8662 2592 8668 2604
rect 8720 2592 8726 2644
rect 9950 2592 9956 2644
rect 10008 2632 10014 2644
rect 10689 2635 10747 2641
rect 10689 2632 10701 2635
rect 10008 2604 10701 2632
rect 10008 2592 10014 2604
rect 10689 2601 10701 2604
rect 10735 2601 10747 2635
rect 11146 2632 11152 2644
rect 11107 2604 11152 2632
rect 10689 2595 10747 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 11885 2635 11943 2641
rect 11885 2601 11897 2635
rect 11931 2632 11943 2635
rect 11931 2604 12940 2632
rect 11931 2601 11943 2604
rect 11885 2595 11943 2601
rect 2222 2564 2228 2576
rect 2183 2536 2228 2564
rect 2222 2524 2228 2536
rect 2280 2524 2286 2576
rect 4154 2564 4160 2576
rect 4115 2536 4160 2564
rect 4154 2524 4160 2536
rect 4212 2524 4218 2576
rect 5537 2567 5595 2573
rect 5537 2533 5549 2567
rect 5583 2564 5595 2567
rect 6362 2564 6368 2576
rect 5583 2536 6368 2564
rect 5583 2533 5595 2536
rect 5537 2527 5595 2533
rect 6362 2524 6368 2536
rect 6420 2524 6426 2576
rect 7374 2524 7380 2576
rect 7432 2564 7438 2576
rect 7561 2567 7619 2573
rect 7561 2564 7573 2567
rect 7432 2536 7573 2564
rect 7432 2524 7438 2536
rect 7561 2533 7573 2536
rect 7607 2533 7619 2567
rect 7561 2527 7619 2533
rect 8389 2567 8447 2573
rect 8389 2533 8401 2567
rect 8435 2564 8447 2567
rect 9122 2564 9128 2576
rect 8435 2536 9128 2564
rect 8435 2533 8447 2536
rect 8389 2527 8447 2533
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 10134 2564 10140 2576
rect 9324 2536 10140 2564
rect 290 2456 296 2508
rect 348 2496 354 2508
rect 1394 2496 1400 2508
rect 348 2468 1400 2496
rect 348 2456 354 2468
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2041 2499 2099 2505
rect 2041 2496 2053 2499
rect 2004 2468 2053 2496
rect 2004 2456 2010 2468
rect 2041 2465 2053 2468
rect 2087 2465 2099 2499
rect 2498 2496 2504 2508
rect 2459 2468 2504 2496
rect 2041 2459 2099 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 3050 2456 3056 2508
rect 3108 2496 3114 2508
rect 3145 2499 3203 2505
rect 3145 2496 3157 2499
rect 3108 2468 3157 2496
rect 3108 2456 3114 2468
rect 3145 2465 3157 2468
rect 3191 2465 3203 2499
rect 4709 2499 4767 2505
rect 4709 2496 4721 2499
rect 3145 2459 3203 2465
rect 4172 2468 4721 2496
rect 4172 2440 4200 2468
rect 4709 2465 4721 2468
rect 4755 2496 4767 2499
rect 5166 2496 5172 2508
rect 4755 2468 5172 2496
rect 4755 2465 4767 2468
rect 4709 2459 4767 2465
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 5258 2456 5264 2508
rect 5316 2496 5322 2508
rect 5353 2499 5411 2505
rect 5353 2496 5365 2499
rect 5316 2468 5365 2496
rect 5316 2456 5322 2468
rect 5353 2465 5365 2468
rect 5399 2465 5411 2499
rect 5353 2459 5411 2465
rect 5810 2456 5816 2508
rect 5868 2496 5874 2508
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5868 2468 6009 2496
rect 5868 2456 5874 2468
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 6454 2456 6460 2508
rect 6512 2496 6518 2508
rect 6825 2499 6883 2505
rect 6825 2496 6837 2499
rect 6512 2468 6837 2496
rect 6512 2456 6518 2468
rect 6825 2465 6837 2468
rect 6871 2465 6883 2499
rect 6825 2459 6883 2465
rect 7650 2456 7656 2508
rect 7708 2496 7714 2508
rect 7745 2499 7803 2505
rect 7745 2496 7757 2499
rect 7708 2468 7757 2496
rect 7708 2456 7714 2468
rect 7745 2465 7757 2468
rect 7791 2465 7803 2499
rect 8202 2496 8208 2508
rect 8163 2468 8208 2496
rect 7745 2459 7803 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2496 8723 2499
rect 8938 2496 8944 2508
rect 8711 2468 8944 2496
rect 8711 2465 8723 2468
rect 8665 2459 8723 2465
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 9324 2428 9352 2536
rect 10134 2524 10140 2536
rect 10192 2524 10198 2576
rect 10229 2567 10287 2573
rect 10229 2533 10241 2567
rect 10275 2564 10287 2567
rect 10410 2564 10416 2576
rect 10275 2536 10416 2564
rect 10275 2533 10287 2536
rect 10229 2527 10287 2533
rect 10410 2524 10416 2536
rect 10468 2524 10474 2576
rect 11698 2524 11704 2576
rect 11756 2564 11762 2576
rect 12912 2573 12940 2604
rect 14550 2592 14556 2644
rect 14608 2632 14614 2644
rect 14737 2635 14795 2641
rect 14737 2632 14749 2635
rect 14608 2604 14749 2632
rect 14608 2592 14614 2604
rect 14737 2601 14749 2604
rect 14783 2601 14795 2635
rect 14737 2595 14795 2601
rect 15838 2592 15844 2644
rect 15896 2632 15902 2644
rect 16025 2635 16083 2641
rect 16025 2632 16037 2635
rect 15896 2604 16037 2632
rect 15896 2592 15902 2604
rect 16025 2601 16037 2604
rect 16071 2601 16083 2635
rect 16025 2595 16083 2601
rect 16485 2635 16543 2641
rect 16485 2601 16497 2635
rect 16531 2632 16543 2635
rect 16574 2632 16580 2644
rect 16531 2604 16580 2632
rect 16531 2601 16543 2604
rect 16485 2595 16543 2601
rect 16574 2592 16580 2604
rect 16632 2592 16638 2644
rect 17313 2635 17371 2641
rect 17313 2601 17325 2635
rect 17359 2632 17371 2635
rect 18506 2632 18512 2644
rect 17359 2604 18512 2632
rect 17359 2601 17371 2604
rect 17313 2595 17371 2601
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 18598 2592 18604 2644
rect 18656 2632 18662 2644
rect 20073 2635 20131 2641
rect 20073 2632 20085 2635
rect 18656 2604 20085 2632
rect 18656 2592 18662 2604
rect 20073 2601 20085 2604
rect 20119 2601 20131 2635
rect 20073 2595 20131 2601
rect 12253 2567 12311 2573
rect 12253 2564 12265 2567
rect 11756 2536 12265 2564
rect 11756 2524 11762 2536
rect 12253 2533 12265 2536
rect 12299 2533 12311 2567
rect 12253 2527 12311 2533
rect 12897 2567 12955 2573
rect 12897 2533 12909 2567
rect 12943 2533 12955 2567
rect 15289 2567 15347 2573
rect 12897 2527 12955 2533
rect 13372 2536 14136 2564
rect 9490 2496 9496 2508
rect 9451 2468 9496 2496
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 10045 2499 10103 2505
rect 10045 2496 10057 2499
rect 9824 2468 10057 2496
rect 9824 2456 9830 2468
rect 10045 2465 10057 2468
rect 10091 2496 10103 2499
rect 10318 2496 10324 2508
rect 10091 2468 10324 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 10594 2496 10600 2508
rect 10555 2468 10600 2496
rect 10594 2456 10600 2468
rect 10652 2456 10658 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 10928 2468 11253 2496
rect 10928 2456 10934 2468
rect 11241 2465 11253 2468
rect 11287 2496 11299 2499
rect 13372 2496 13400 2536
rect 11287 2468 13400 2496
rect 13449 2499 13507 2505
rect 11287 2465 11299 2468
rect 11241 2459 11299 2465
rect 13449 2465 13461 2499
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 14001 2499 14059 2505
rect 14001 2465 14013 2499
rect 14047 2465 14059 2499
rect 14108 2496 14136 2536
rect 15289 2533 15301 2567
rect 15335 2564 15347 2567
rect 17586 2564 17592 2576
rect 15335 2536 17592 2564
rect 15335 2533 15347 2536
rect 15289 2527 15347 2533
rect 17586 2524 17592 2536
rect 17644 2524 17650 2576
rect 18138 2564 18144 2576
rect 17696 2536 18144 2564
rect 14108 2468 16068 2496
rect 14001 2459 14059 2465
rect 5828 2400 9352 2428
rect 9677 2431 9735 2437
rect 2682 2292 2688 2304
rect 2643 2264 2688 2292
rect 2682 2252 2688 2264
rect 2740 2252 2746 2304
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 5828 2292 5856 2400
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 9723 2400 12204 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 11885 2363 11943 2369
rect 11885 2360 11897 2363
rect 8536 2332 11897 2360
rect 8536 2320 8542 2332
rect 11885 2329 11897 2332
rect 11931 2329 11943 2363
rect 12066 2360 12072 2372
rect 12027 2332 12072 2360
rect 11885 2323 11943 2329
rect 12066 2320 12072 2332
rect 12124 2320 12130 2372
rect 12176 2360 12204 2400
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 13464 2428 13492 2459
rect 12308 2400 13492 2428
rect 12308 2388 12314 2400
rect 12710 2360 12716 2372
rect 12176 2332 12716 2360
rect 12710 2320 12716 2332
rect 12768 2320 12774 2372
rect 14016 2360 14044 2459
rect 15930 2428 15936 2440
rect 15891 2400 15936 2428
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 16040 2428 16068 2468
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16172 2468 16217 2496
rect 16172 2456 16178 2468
rect 17696 2437 17724 2536
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18785 2567 18843 2573
rect 18785 2533 18797 2567
rect 18831 2564 18843 2567
rect 18966 2564 18972 2576
rect 18831 2536 18972 2564
rect 18831 2533 18843 2536
rect 18785 2527 18843 2533
rect 18966 2524 18972 2536
rect 19024 2524 19030 2576
rect 19058 2524 19064 2576
rect 19116 2564 19122 2576
rect 20533 2567 20591 2573
rect 20533 2564 20545 2567
rect 19116 2536 20545 2564
rect 19116 2524 19122 2536
rect 20533 2533 20545 2536
rect 20579 2533 20591 2567
rect 20533 2527 20591 2533
rect 20717 2567 20775 2573
rect 20717 2533 20729 2567
rect 20763 2564 20775 2567
rect 22005 2567 22063 2573
rect 22005 2564 22017 2567
rect 20763 2536 22017 2564
rect 20763 2533 20775 2536
rect 20717 2527 20775 2533
rect 22005 2533 22017 2536
rect 22051 2533 22063 2567
rect 22005 2527 22063 2533
rect 17954 2496 17960 2508
rect 17915 2468 17960 2496
rect 17954 2456 17960 2468
rect 18012 2456 18018 2508
rect 19429 2499 19487 2505
rect 19429 2465 19441 2499
rect 19475 2496 19487 2499
rect 19518 2496 19524 2508
rect 19475 2468 19524 2496
rect 19475 2465 19487 2468
rect 19429 2459 19487 2465
rect 19518 2456 19524 2468
rect 19576 2456 19582 2508
rect 16761 2431 16819 2437
rect 16761 2428 16773 2431
rect 16040 2400 16773 2428
rect 16761 2397 16773 2400
rect 16807 2397 16819 2431
rect 16761 2391 16819 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17862 2428 17868 2440
rect 17823 2400 17868 2428
rect 17681 2391 17739 2397
rect 17862 2388 17868 2400
rect 17920 2428 17926 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 17920 2400 19257 2428
rect 17920 2388 17926 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 12912 2332 14044 2360
rect 15473 2363 15531 2369
rect 3283 2264 5856 2292
rect 5905 2295 5963 2301
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 5905 2261 5917 2295
rect 5951 2292 5963 2295
rect 8294 2292 8300 2304
rect 5951 2264 8300 2292
rect 5951 2261 5963 2264
rect 5905 2255 5963 2261
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8846 2292 8852 2304
rect 8807 2264 8852 2292
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 10778 2252 10784 2304
rect 10836 2292 10842 2304
rect 12912 2292 12940 2332
rect 15473 2329 15485 2363
rect 15519 2360 15531 2363
rect 15519 2332 17724 2360
rect 15519 2329 15531 2332
rect 15473 2323 15531 2329
rect 10836 2264 12940 2292
rect 10836 2252 10842 2264
rect 12986 2252 12992 2304
rect 13044 2292 13050 2304
rect 13538 2292 13544 2304
rect 13044 2264 13089 2292
rect 13499 2264 13544 2292
rect 13044 2252 13050 2264
rect 13538 2252 13544 2264
rect 13596 2252 13602 2304
rect 14090 2292 14096 2304
rect 14051 2264 14096 2292
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 17696 2292 17724 2332
rect 17770 2320 17776 2372
rect 17828 2360 17834 2372
rect 18601 2363 18659 2369
rect 18601 2360 18613 2363
rect 17828 2332 18613 2360
rect 17828 2320 17834 2332
rect 18601 2329 18613 2332
rect 18647 2329 18659 2363
rect 18601 2323 18659 2329
rect 19150 2320 19156 2372
rect 19208 2360 19214 2372
rect 19208 2332 19380 2360
rect 19208 2320 19214 2332
rect 18138 2292 18144 2304
rect 17696 2264 18144 2292
rect 18138 2252 18144 2264
rect 18196 2252 18202 2304
rect 18325 2295 18383 2301
rect 18325 2261 18337 2295
rect 18371 2292 18383 2295
rect 19242 2292 19248 2304
rect 18371 2264 19248 2292
rect 18371 2261 18383 2264
rect 18325 2255 18383 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 19352 2292 19380 2332
rect 19426 2320 19432 2372
rect 19484 2360 19490 2372
rect 20732 2360 20760 2527
rect 21269 2499 21327 2505
rect 21269 2496 21281 2499
rect 19484 2332 20760 2360
rect 20824 2468 21281 2496
rect 19484 2320 19490 2332
rect 20824 2292 20852 2468
rect 21269 2465 21281 2468
rect 21315 2496 21327 2499
rect 22097 2499 22155 2505
rect 22097 2496 22109 2499
rect 21315 2468 22109 2496
rect 21315 2465 21327 2468
rect 21269 2459 21327 2465
rect 22097 2465 22109 2468
rect 22143 2465 22155 2499
rect 22097 2459 22155 2465
rect 21082 2360 21088 2372
rect 21043 2332 21088 2360
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 19352 2264 20852 2292
rect 1104 2202 21896 2224
rect 1104 2150 4447 2202
rect 4499 2150 4511 2202
rect 4563 2150 4575 2202
rect 4627 2150 4639 2202
rect 4691 2150 11378 2202
rect 11430 2150 11442 2202
rect 11494 2150 11506 2202
rect 11558 2150 11570 2202
rect 11622 2150 18308 2202
rect 18360 2150 18372 2202
rect 18424 2150 18436 2202
rect 18488 2150 18500 2202
rect 18552 2150 21896 2202
rect 1104 2128 21896 2150
rect 9030 2048 9036 2100
rect 9088 2088 9094 2100
rect 12250 2088 12256 2100
rect 9088 2060 12256 2088
rect 9088 2048 9094 2060
rect 12250 2048 12256 2060
rect 12308 2048 12314 2100
rect 14090 2048 14096 2100
rect 14148 2088 14154 2100
rect 19886 2088 19892 2100
rect 14148 2060 19892 2088
rect 14148 2048 14154 2060
rect 19886 2048 19892 2060
rect 19944 2048 19950 2100
rect 2038 1980 2044 2032
rect 2096 2020 2102 2032
rect 17954 2020 17960 2032
rect 2096 1992 17960 2020
rect 2096 1980 2102 1992
rect 17954 1980 17960 1992
rect 18012 1980 18018 2032
rect 8662 1912 8668 1964
rect 8720 1952 8726 1964
rect 9490 1952 9496 1964
rect 8720 1924 9496 1952
rect 8720 1912 8726 1924
rect 9490 1912 9496 1924
rect 9548 1912 9554 1964
rect 9858 1912 9864 1964
rect 9916 1952 9922 1964
rect 11422 1952 11428 1964
rect 9916 1924 11428 1952
rect 9916 1912 9922 1924
rect 11422 1912 11428 1924
rect 11480 1912 11486 1964
rect 16758 1912 16764 1964
rect 16816 1952 16822 1964
rect 21082 1952 21088 1964
rect 16816 1924 21088 1952
rect 16816 1912 16822 1924
rect 21082 1912 21088 1924
rect 21140 1912 21146 1964
rect 2682 1844 2688 1896
rect 2740 1884 2746 1896
rect 16114 1884 16120 1896
rect 2740 1856 16120 1884
rect 2740 1844 2746 1856
rect 16114 1844 16120 1856
rect 16172 1844 16178 1896
rect 13538 1776 13544 1828
rect 13596 1816 13602 1828
rect 20438 1816 20444 1828
rect 13596 1788 20444 1816
rect 13596 1776 13602 1788
rect 20438 1776 20444 1788
rect 20496 1776 20502 1828
rect 6178 1708 6184 1760
rect 6236 1748 6242 1760
rect 17862 1748 17868 1760
rect 6236 1720 17868 1748
rect 6236 1708 6242 1720
rect 17862 1708 17868 1720
rect 17920 1708 17926 1760
rect 8846 1640 8852 1692
rect 8904 1680 8910 1692
rect 16850 1680 16856 1692
rect 8904 1652 16856 1680
rect 8904 1640 8910 1652
rect 16850 1640 16856 1652
rect 16908 1640 16914 1692
rect 8938 1572 8944 1624
rect 8996 1612 9002 1624
rect 18046 1612 18052 1624
rect 8996 1584 18052 1612
rect 8996 1572 9002 1584
rect 18046 1572 18052 1584
rect 18104 1572 18110 1624
rect 12986 1504 12992 1556
rect 13044 1544 13050 1556
rect 22646 1544 22652 1556
rect 13044 1516 22652 1544
rect 13044 1504 13050 1516
rect 22646 1504 22652 1516
rect 22704 1504 22710 1556
rect 21910 1436 21916 1488
rect 21968 1476 21974 1488
rect 22097 1479 22155 1485
rect 22097 1476 22109 1479
rect 21968 1448 22109 1476
rect 21968 1436 21974 1448
rect 22097 1445 22109 1448
rect 22143 1445 22155 1479
rect 22097 1439 22155 1445
rect 22002 1408 22008 1420
rect 21963 1380 22008 1408
rect 22002 1368 22008 1380
rect 22060 1368 22066 1420
<< via1 >>
rect 4447 20646 4499 20698
rect 4511 20646 4563 20698
rect 4575 20646 4627 20698
rect 4639 20646 4691 20698
rect 11378 20646 11430 20698
rect 11442 20646 11494 20698
rect 11506 20646 11558 20698
rect 11570 20646 11622 20698
rect 18308 20646 18360 20698
rect 18372 20646 18424 20698
rect 18436 20646 18488 20698
rect 18500 20646 18552 20698
rect 848 20544 900 20596
rect 5080 20544 5132 20596
rect 8944 20544 8996 20596
rect 6000 20476 6052 20528
rect 7104 20476 7156 20528
rect 7564 20476 7616 20528
rect 8208 20476 8260 20528
rect 11428 20476 11480 20528
rect 12072 20519 12124 20528
rect 12072 20485 12081 20519
rect 12081 20485 12115 20519
rect 12115 20485 12124 20519
rect 12072 20476 12124 20485
rect 12256 20544 12308 20596
rect 12624 20519 12676 20528
rect 12624 20485 12633 20519
rect 12633 20485 12667 20519
rect 12667 20485 12676 20519
rect 12624 20476 12676 20485
rect 13176 20519 13228 20528
rect 13176 20485 13185 20519
rect 13185 20485 13219 20519
rect 13219 20485 13228 20519
rect 13176 20476 13228 20485
rect 13728 20519 13780 20528
rect 13728 20485 13737 20519
rect 13737 20485 13771 20519
rect 13771 20485 13780 20519
rect 13728 20476 13780 20485
rect 14464 20544 14516 20596
rect 18144 20544 18196 20596
rect 16396 20476 16448 20528
rect 17684 20476 17736 20528
rect 17960 20476 18012 20528
rect 18604 20476 18656 20528
rect 18972 20519 19024 20528
rect 18972 20485 18981 20519
rect 18981 20485 19015 20519
rect 19015 20485 19024 20519
rect 18972 20476 19024 20485
rect 19524 20519 19576 20528
rect 19524 20485 19533 20519
rect 19533 20485 19567 20519
rect 19567 20485 19576 20519
rect 19524 20476 19576 20485
rect 5172 20408 5224 20460
rect 6920 20408 6972 20460
rect 3056 20340 3108 20392
rect 3608 20340 3660 20392
rect 5264 20340 5316 20392
rect 5816 20340 5868 20392
rect 6460 20340 6512 20392
rect 10048 20408 10100 20460
rect 7564 20340 7616 20392
rect 1952 20272 2004 20324
rect 4896 20315 4948 20324
rect 4896 20281 4905 20315
rect 4905 20281 4939 20315
rect 4939 20281 4948 20315
rect 4896 20272 4948 20281
rect 7288 20272 7340 20324
rect 7472 20272 7524 20324
rect 8116 20340 8168 20392
rect 2688 20247 2740 20256
rect 2688 20213 2697 20247
rect 2697 20213 2731 20247
rect 2731 20213 2740 20247
rect 2688 20204 2740 20213
rect 4160 20204 4212 20256
rect 5908 20247 5960 20256
rect 5908 20213 5917 20247
rect 5917 20213 5951 20247
rect 5951 20213 5960 20247
rect 5908 20204 5960 20213
rect 7380 20204 7432 20256
rect 8392 20272 8444 20324
rect 8760 20340 8812 20392
rect 18788 20408 18840 20460
rect 10324 20340 10376 20392
rect 10784 20340 10836 20392
rect 10876 20340 10928 20392
rect 20444 20408 20496 20460
rect 8668 20204 8720 20256
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 9496 20247 9548 20256
rect 9496 20213 9505 20247
rect 9505 20213 9539 20247
rect 9539 20213 9548 20247
rect 9496 20204 9548 20213
rect 9864 20272 9916 20324
rect 10416 20272 10468 20324
rect 10508 20315 10560 20324
rect 10508 20281 10517 20315
rect 10517 20281 10551 20315
rect 10551 20281 10560 20315
rect 10508 20272 10560 20281
rect 11060 20272 11112 20324
rect 11704 20272 11756 20324
rect 12808 20315 12860 20324
rect 12808 20281 12817 20315
rect 12817 20281 12851 20315
rect 12851 20281 12860 20315
rect 12808 20272 12860 20281
rect 13728 20272 13780 20324
rect 13912 20315 13964 20324
rect 13912 20281 13921 20315
rect 13921 20281 13955 20315
rect 13955 20281 13964 20315
rect 13912 20272 13964 20281
rect 16120 20315 16172 20324
rect 9956 20204 10008 20256
rect 11152 20247 11204 20256
rect 11152 20213 11161 20247
rect 11161 20213 11195 20247
rect 11195 20213 11204 20247
rect 11152 20204 11204 20213
rect 16120 20281 16129 20315
rect 16129 20281 16163 20315
rect 16163 20281 16172 20315
rect 16120 20272 16172 20281
rect 16672 20315 16724 20324
rect 16672 20281 16681 20315
rect 16681 20281 16715 20315
rect 16715 20281 16724 20315
rect 16672 20272 16724 20281
rect 20168 20340 20220 20392
rect 17684 20315 17736 20324
rect 17684 20281 17693 20315
rect 17693 20281 17727 20315
rect 17727 20281 17736 20315
rect 17684 20272 17736 20281
rect 17960 20272 18012 20324
rect 18788 20315 18840 20324
rect 18788 20281 18797 20315
rect 18797 20281 18831 20315
rect 18831 20281 18840 20315
rect 18788 20272 18840 20281
rect 19432 20272 19484 20324
rect 20628 20315 20680 20324
rect 20628 20281 20637 20315
rect 20637 20281 20671 20315
rect 20671 20281 20680 20315
rect 20628 20272 20680 20281
rect 20812 20315 20864 20324
rect 20812 20281 20821 20315
rect 20821 20281 20855 20315
rect 20855 20281 20864 20315
rect 20812 20272 20864 20281
rect 21180 20315 21232 20324
rect 21180 20281 21189 20315
rect 21189 20281 21223 20315
rect 21223 20281 21232 20315
rect 21180 20272 21232 20281
rect 21456 20272 21508 20324
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 21088 20204 21140 20256
rect 7912 20102 7964 20154
rect 7976 20102 8028 20154
rect 8040 20102 8092 20154
rect 8104 20102 8156 20154
rect 14843 20102 14895 20154
rect 14907 20102 14959 20154
rect 14971 20102 15023 20154
rect 15035 20102 15087 20154
rect 2320 20043 2372 20052
rect 2320 20009 2329 20043
rect 2329 20009 2363 20043
rect 2363 20009 2372 20043
rect 2320 20000 2372 20009
rect 3056 20000 3108 20052
rect 3608 20000 3660 20052
rect 4160 20000 4212 20052
rect 1400 19932 1452 19984
rect 1952 19932 2004 19984
rect 7104 20000 7156 20052
rect 8208 20000 8260 20052
rect 8944 20000 8996 20052
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 2504 19864 2556 19916
rect 4804 19864 4856 19916
rect 6092 19907 6144 19916
rect 6092 19873 6101 19907
rect 6101 19873 6135 19907
rect 6135 19873 6144 19907
rect 6092 19864 6144 19873
rect 6552 19907 6604 19916
rect 6552 19873 6561 19907
rect 6561 19873 6595 19907
rect 6595 19873 6604 19907
rect 6552 19864 6604 19873
rect 7012 19907 7064 19916
rect 7012 19873 7021 19907
rect 7021 19873 7055 19907
rect 7055 19873 7064 19907
rect 7012 19864 7064 19873
rect 7656 19907 7708 19916
rect 7656 19873 7665 19907
rect 7665 19873 7699 19907
rect 7699 19873 7708 19907
rect 7656 19864 7708 19873
rect 8116 19907 8168 19916
rect 8116 19873 8125 19907
rect 8125 19873 8159 19907
rect 8159 19873 8168 19907
rect 8116 19864 8168 19873
rect 9772 19932 9824 19984
rect 10048 19932 10100 19984
rect 11428 20000 11480 20052
rect 8392 19864 8444 19916
rect 8576 19907 8628 19916
rect 8576 19873 8585 19907
rect 8585 19873 8619 19907
rect 8619 19873 8628 19907
rect 8576 19864 8628 19873
rect 9312 19864 9364 19916
rect 9588 19864 9640 19916
rect 10324 19864 10376 19916
rect 11060 19864 11112 19916
rect 2044 19796 2096 19848
rect 6644 19796 6696 19848
rect 6828 19796 6880 19848
rect 9864 19796 9916 19848
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 2780 19771 2832 19780
rect 2780 19737 2789 19771
rect 2789 19737 2823 19771
rect 2823 19737 2832 19771
rect 7196 19771 7248 19780
rect 2780 19728 2832 19737
rect 7196 19737 7205 19771
rect 7205 19737 7239 19771
rect 7239 19737 7248 19771
rect 7196 19728 7248 19737
rect 8116 19728 8168 19780
rect 10140 19728 10192 19780
rect 10232 19728 10284 19780
rect 12072 19932 12124 19984
rect 12900 19864 12952 19916
rect 13268 19796 13320 19848
rect 13728 20000 13780 20052
rect 13820 19864 13872 19916
rect 14464 20000 14516 20052
rect 14740 20000 14792 20052
rect 14280 19932 14332 19984
rect 15200 20000 15252 20052
rect 18788 20000 18840 20052
rect 21548 20000 21600 20052
rect 15384 19932 15436 19984
rect 15936 19932 15988 19984
rect 16396 19975 16448 19984
rect 16396 19941 16405 19975
rect 16405 19941 16439 19975
rect 16439 19941 16448 19975
rect 16396 19932 16448 19941
rect 16580 19932 16632 19984
rect 17040 19932 17092 19984
rect 19340 19932 19392 19984
rect 19892 19932 19944 19984
rect 14464 19864 14516 19916
rect 15200 19864 15252 19916
rect 16948 19907 17000 19916
rect 16948 19873 16957 19907
rect 16957 19873 16991 19907
rect 16991 19873 17000 19907
rect 16948 19864 17000 19873
rect 17500 19907 17552 19916
rect 17500 19873 17509 19907
rect 17509 19873 17543 19907
rect 17543 19873 17552 19907
rect 17500 19864 17552 19873
rect 18512 19907 18564 19916
rect 18512 19873 18521 19907
rect 18521 19873 18555 19907
rect 18555 19873 18564 19907
rect 18512 19864 18564 19873
rect 18604 19864 18656 19916
rect 19616 19864 19668 19916
rect 20536 19907 20588 19916
rect 20536 19873 20545 19907
rect 20545 19873 20579 19907
rect 20579 19873 20588 19907
rect 20536 19864 20588 19873
rect 19340 19796 19392 19848
rect 16672 19728 16724 19780
rect 21364 19771 21416 19780
rect 21364 19737 21373 19771
rect 21373 19737 21407 19771
rect 21407 19737 21416 19771
rect 21364 19728 21416 19737
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 6644 19660 6696 19712
rect 6828 19660 6880 19712
rect 7104 19660 7156 19712
rect 10324 19660 10376 19712
rect 11244 19660 11296 19712
rect 12348 19703 12400 19712
rect 12348 19669 12357 19703
rect 12357 19669 12391 19703
rect 12391 19669 12400 19703
rect 12348 19660 12400 19669
rect 14372 19660 14424 19712
rect 14556 19660 14608 19712
rect 22100 19660 22152 19712
rect 4447 19558 4499 19610
rect 4511 19558 4563 19610
rect 4575 19558 4627 19610
rect 4639 19558 4691 19610
rect 11378 19558 11430 19610
rect 11442 19558 11494 19610
rect 11506 19558 11558 19610
rect 11570 19558 11622 19610
rect 18308 19558 18360 19610
rect 18372 19558 18424 19610
rect 18436 19558 18488 19610
rect 18500 19558 18552 19610
rect 1952 19499 2004 19508
rect 1952 19465 1961 19499
rect 1961 19465 1995 19499
rect 1995 19465 2004 19499
rect 1952 19456 2004 19465
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 4804 19456 4856 19508
rect 6460 19456 6512 19508
rect 6644 19456 6696 19508
rect 12900 19456 12952 19508
rect 13268 19499 13320 19508
rect 13268 19465 13277 19499
rect 13277 19465 13311 19499
rect 13311 19465 13320 19499
rect 13268 19456 13320 19465
rect 296 19252 348 19304
rect 1676 19252 1728 19304
rect 5264 19252 5316 19304
rect 7288 19320 7340 19372
rect 7564 19320 7616 19372
rect 7104 19252 7156 19304
rect 7380 19252 7432 19304
rect 8852 19252 8904 19304
rect 9036 19295 9088 19304
rect 9036 19261 9045 19295
rect 9045 19261 9079 19295
rect 9079 19261 9088 19295
rect 9036 19252 9088 19261
rect 6552 19184 6604 19236
rect 9220 19252 9272 19304
rect 9680 19252 9732 19304
rect 10968 19320 11020 19372
rect 14740 19456 14792 19508
rect 17224 19456 17276 19508
rect 20628 19456 20680 19508
rect 16120 19388 16172 19440
rect 10600 19252 10652 19304
rect 6184 19116 6236 19168
rect 6276 19116 6328 19168
rect 7380 19159 7432 19168
rect 7380 19125 7389 19159
rect 7389 19125 7423 19159
rect 7423 19125 7432 19159
rect 7380 19116 7432 19125
rect 7748 19116 7800 19168
rect 8300 19159 8352 19168
rect 8300 19125 8309 19159
rect 8309 19125 8343 19159
rect 8343 19125 8352 19159
rect 8300 19116 8352 19125
rect 8760 19159 8812 19168
rect 8760 19125 8769 19159
rect 8769 19125 8803 19159
rect 8803 19125 8812 19159
rect 8760 19116 8812 19125
rect 9312 19116 9364 19168
rect 10048 19116 10100 19168
rect 10692 19184 10744 19236
rect 14280 19252 14332 19304
rect 18604 19320 18656 19372
rect 12164 19227 12216 19236
rect 12164 19193 12198 19227
rect 12198 19193 12216 19227
rect 12164 19184 12216 19193
rect 12348 19184 12400 19236
rect 12440 19184 12492 19236
rect 17040 19252 17092 19304
rect 17592 19252 17644 19304
rect 18420 19295 18472 19304
rect 18420 19261 18429 19295
rect 18429 19261 18463 19295
rect 18463 19261 18472 19295
rect 18420 19252 18472 19261
rect 19064 19252 19116 19304
rect 19432 19388 19484 19440
rect 19248 19252 19300 19304
rect 21088 19252 21140 19304
rect 11428 19116 11480 19168
rect 12716 19116 12768 19168
rect 14188 19116 14240 19168
rect 16580 19116 16632 19168
rect 17960 19116 18012 19168
rect 19708 19184 19760 19236
rect 19984 19227 20036 19236
rect 19984 19193 19993 19227
rect 19993 19193 20027 19227
rect 20027 19193 20036 19227
rect 19984 19184 20036 19193
rect 21364 19227 21416 19236
rect 21364 19193 21373 19227
rect 21373 19193 21407 19227
rect 21407 19193 21416 19227
rect 21364 19184 21416 19193
rect 19340 19116 19392 19168
rect 21088 19116 21140 19168
rect 7912 19014 7964 19066
rect 7976 19014 8028 19066
rect 8040 19014 8092 19066
rect 8104 19014 8156 19066
rect 14843 19014 14895 19066
rect 14907 19014 14959 19066
rect 14971 19014 15023 19066
rect 15035 19014 15087 19066
rect 5816 18912 5868 18964
rect 7012 18912 7064 18964
rect 6184 18844 6236 18896
rect 7472 18912 7524 18964
rect 10692 18955 10744 18964
rect 6092 18776 6144 18828
rect 6276 18708 6328 18760
rect 5264 18640 5316 18692
rect 5540 18572 5592 18624
rect 7472 18640 7524 18692
rect 7932 18708 7984 18760
rect 8484 18776 8536 18828
rect 9312 18844 9364 18896
rect 10692 18921 10701 18955
rect 10701 18921 10735 18955
rect 10735 18921 10744 18955
rect 10692 18912 10744 18921
rect 11244 18955 11296 18964
rect 11244 18921 11253 18955
rect 11253 18921 11287 18955
rect 11287 18921 11296 18955
rect 11244 18912 11296 18921
rect 12256 18912 12308 18964
rect 12808 18912 12860 18964
rect 13544 18912 13596 18964
rect 14188 18912 14240 18964
rect 16580 18955 16632 18964
rect 14004 18844 14056 18896
rect 16580 18921 16589 18955
rect 16589 18921 16623 18955
rect 16623 18921 16632 18955
rect 16580 18912 16632 18921
rect 16672 18912 16724 18964
rect 17684 18955 17736 18964
rect 17684 18921 17693 18955
rect 17693 18921 17727 18955
rect 17727 18921 17736 18955
rect 17684 18912 17736 18921
rect 19248 18912 19300 18964
rect 22652 18912 22704 18964
rect 11244 18776 11296 18828
rect 11336 18819 11388 18828
rect 11336 18785 11345 18819
rect 11345 18785 11379 18819
rect 11379 18785 11388 18819
rect 11336 18776 11388 18785
rect 12072 18776 12124 18828
rect 13452 18776 13504 18828
rect 15384 18844 15436 18896
rect 20444 18844 20496 18896
rect 20996 18844 21048 18896
rect 15200 18776 15252 18828
rect 9220 18708 9272 18760
rect 11060 18708 11112 18760
rect 11428 18708 11480 18760
rect 7840 18683 7892 18692
rect 7840 18649 7849 18683
rect 7849 18649 7883 18683
rect 7883 18649 7892 18683
rect 7840 18640 7892 18649
rect 13728 18708 13780 18760
rect 14096 18708 14148 18760
rect 16672 18751 16724 18760
rect 16672 18717 16681 18751
rect 16681 18717 16715 18751
rect 16715 18717 16724 18751
rect 16672 18708 16724 18717
rect 8576 18572 8628 18624
rect 11980 18615 12032 18624
rect 11980 18581 11989 18615
rect 11989 18581 12023 18615
rect 12023 18581 12032 18615
rect 11980 18572 12032 18581
rect 14280 18640 14332 18692
rect 15936 18683 15988 18692
rect 15936 18649 15945 18683
rect 15945 18649 15979 18683
rect 15979 18649 15988 18683
rect 17316 18776 17368 18828
rect 18052 18776 18104 18828
rect 20076 18819 20128 18828
rect 17960 18708 18012 18760
rect 20076 18785 20085 18819
rect 20085 18785 20119 18819
rect 20119 18785 20128 18819
rect 20076 18776 20128 18785
rect 20260 18776 20312 18828
rect 15936 18640 15988 18649
rect 14004 18572 14056 18624
rect 16304 18572 16356 18624
rect 20628 18640 20680 18692
rect 21364 18683 21416 18692
rect 21364 18649 21373 18683
rect 21373 18649 21407 18683
rect 21407 18649 21416 18683
rect 21364 18640 21416 18649
rect 19156 18572 19208 18624
rect 19524 18572 19576 18624
rect 4447 18470 4499 18522
rect 4511 18470 4563 18522
rect 4575 18470 4627 18522
rect 4639 18470 4691 18522
rect 11378 18470 11430 18522
rect 11442 18470 11494 18522
rect 11506 18470 11558 18522
rect 11570 18470 11622 18522
rect 18308 18470 18360 18522
rect 18372 18470 18424 18522
rect 18436 18470 18488 18522
rect 18500 18470 18552 18522
rect 7472 18368 7524 18420
rect 7840 18368 7892 18420
rect 8024 18368 8076 18420
rect 13544 18368 13596 18420
rect 16672 18368 16724 18420
rect 20260 18368 20312 18420
rect 7012 18300 7064 18352
rect 7564 18300 7616 18352
rect 9680 18300 9732 18352
rect 10876 18343 10928 18352
rect 10876 18309 10885 18343
rect 10885 18309 10919 18343
rect 10919 18309 10928 18343
rect 10876 18300 10928 18309
rect 12164 18300 12216 18352
rect 6736 18232 6788 18284
rect 7380 18232 7432 18284
rect 9312 18232 9364 18284
rect 11888 18232 11940 18284
rect 12072 18232 12124 18284
rect 5448 18096 5500 18148
rect 6828 18096 6880 18148
rect 5632 18071 5684 18080
rect 5632 18037 5641 18071
rect 5641 18037 5675 18071
rect 5675 18037 5684 18071
rect 5632 18028 5684 18037
rect 6368 18028 6420 18080
rect 7104 18028 7156 18080
rect 7472 18028 7524 18080
rect 10140 18164 10192 18216
rect 11152 18207 11204 18216
rect 11152 18173 11161 18207
rect 11161 18173 11195 18207
rect 11195 18173 11204 18207
rect 11152 18164 11204 18173
rect 15200 18300 15252 18352
rect 13728 18275 13780 18284
rect 13728 18241 13737 18275
rect 13737 18241 13771 18275
rect 13771 18241 13780 18275
rect 13728 18232 13780 18241
rect 14188 18275 14240 18284
rect 14188 18241 14197 18275
rect 14197 18241 14231 18275
rect 14231 18241 14240 18275
rect 14188 18232 14240 18241
rect 14372 18275 14424 18284
rect 14372 18241 14381 18275
rect 14381 18241 14415 18275
rect 14415 18241 14424 18275
rect 14372 18232 14424 18241
rect 8852 18096 8904 18148
rect 9220 18096 9272 18148
rect 11244 18096 11296 18148
rect 8300 18028 8352 18080
rect 9128 18028 9180 18080
rect 9496 18028 9548 18080
rect 9772 18071 9824 18080
rect 9772 18037 9781 18071
rect 9781 18037 9815 18071
rect 9815 18037 9824 18071
rect 9772 18028 9824 18037
rect 9864 18071 9916 18080
rect 9864 18037 9873 18071
rect 9873 18037 9907 18071
rect 9907 18037 9916 18071
rect 14740 18096 14792 18148
rect 15292 18164 15344 18216
rect 15936 18164 15988 18216
rect 16028 18164 16080 18216
rect 17224 18232 17276 18284
rect 17408 18207 17460 18216
rect 17408 18173 17417 18207
rect 17417 18173 17451 18207
rect 17451 18173 17460 18207
rect 17408 18164 17460 18173
rect 20628 18207 20680 18216
rect 20628 18173 20637 18207
rect 20637 18173 20671 18207
rect 20671 18173 20680 18207
rect 20628 18164 20680 18173
rect 15752 18096 15804 18148
rect 18972 18096 19024 18148
rect 19156 18096 19208 18148
rect 21364 18139 21416 18148
rect 21364 18105 21373 18139
rect 21373 18105 21407 18139
rect 21407 18105 21416 18139
rect 21364 18096 21416 18105
rect 9864 18028 9916 18037
rect 11888 18071 11940 18080
rect 11888 18037 11897 18071
rect 11897 18037 11931 18071
rect 11931 18037 11940 18071
rect 11888 18028 11940 18037
rect 11980 18028 12032 18080
rect 12440 18028 12492 18080
rect 12900 18028 12952 18080
rect 13084 18071 13136 18080
rect 13084 18037 13093 18071
rect 13093 18037 13127 18071
rect 13127 18037 13136 18071
rect 13084 18028 13136 18037
rect 14464 18071 14516 18080
rect 14464 18037 14473 18071
rect 14473 18037 14507 18071
rect 14507 18037 14516 18071
rect 16580 18071 16632 18080
rect 14464 18028 14516 18037
rect 16580 18037 16589 18071
rect 16589 18037 16623 18071
rect 16623 18037 16632 18071
rect 16580 18028 16632 18037
rect 18880 18028 18932 18080
rect 19892 18071 19944 18080
rect 19892 18037 19901 18071
rect 19901 18037 19935 18071
rect 19935 18037 19944 18071
rect 19892 18028 19944 18037
rect 20260 18071 20312 18080
rect 20260 18037 20269 18071
rect 20269 18037 20303 18071
rect 20303 18037 20312 18071
rect 20260 18028 20312 18037
rect 20628 18028 20680 18080
rect 7912 17926 7964 17978
rect 7976 17926 8028 17978
rect 8040 17926 8092 17978
rect 8104 17926 8156 17978
rect 14843 17926 14895 17978
rect 14907 17926 14959 17978
rect 14971 17926 15023 17978
rect 15035 17926 15087 17978
rect 4896 17824 4948 17876
rect 6644 17824 6696 17876
rect 7012 17824 7064 17876
rect 7196 17824 7248 17876
rect 9128 17824 9180 17876
rect 9312 17867 9364 17876
rect 9312 17833 9321 17867
rect 9321 17833 9355 17867
rect 9355 17833 9364 17867
rect 9312 17824 9364 17833
rect 13084 17824 13136 17876
rect 13176 17824 13228 17876
rect 6092 17756 6144 17808
rect 6644 17688 6696 17740
rect 7380 17620 7432 17672
rect 7564 17663 7616 17672
rect 7564 17629 7573 17663
rect 7573 17629 7607 17663
rect 7607 17629 7616 17663
rect 7564 17620 7616 17629
rect 8484 17756 8536 17808
rect 10600 17756 10652 17808
rect 8760 17688 8812 17740
rect 9680 17688 9732 17740
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 12440 17756 12492 17808
rect 12532 17756 12584 17808
rect 13636 17756 13688 17808
rect 17500 17824 17552 17876
rect 18972 17867 19024 17876
rect 18972 17833 18981 17867
rect 18981 17833 19015 17867
rect 19015 17833 19024 17867
rect 18972 17824 19024 17833
rect 20260 17824 20312 17876
rect 15200 17756 15252 17808
rect 9588 17620 9640 17672
rect 10968 17620 11020 17672
rect 5816 17484 5868 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 7104 17484 7156 17493
rect 7656 17484 7708 17536
rect 8668 17484 8720 17536
rect 11152 17552 11204 17604
rect 14556 17688 14608 17740
rect 15292 17688 15344 17740
rect 10968 17484 11020 17536
rect 11244 17527 11296 17536
rect 11244 17493 11253 17527
rect 11253 17493 11287 17527
rect 11287 17493 11296 17527
rect 11244 17484 11296 17493
rect 11980 17595 12032 17604
rect 11980 17561 11989 17595
rect 11989 17561 12023 17595
rect 12023 17561 12032 17595
rect 11980 17552 12032 17561
rect 12532 17663 12584 17672
rect 12532 17629 12541 17663
rect 12541 17629 12575 17663
rect 12575 17629 12584 17663
rect 12532 17620 12584 17629
rect 13544 17620 13596 17672
rect 14096 17620 14148 17672
rect 15200 17620 15252 17672
rect 15384 17620 15436 17672
rect 14648 17552 14700 17604
rect 15016 17552 15068 17604
rect 16488 17756 16540 17808
rect 16580 17688 16632 17740
rect 17040 17731 17092 17740
rect 17040 17697 17058 17731
rect 17058 17697 17092 17731
rect 17040 17688 17092 17697
rect 17224 17688 17276 17740
rect 18144 17688 18196 17740
rect 18880 17688 18932 17740
rect 20260 17663 20312 17672
rect 20260 17629 20269 17663
rect 20269 17629 20303 17663
rect 20303 17629 20312 17663
rect 20260 17620 20312 17629
rect 21364 17595 21416 17604
rect 12072 17484 12124 17536
rect 12624 17484 12676 17536
rect 15476 17484 15528 17536
rect 16212 17484 16264 17536
rect 21364 17561 21373 17595
rect 21373 17561 21407 17595
rect 21407 17561 21416 17595
rect 21364 17552 21416 17561
rect 19800 17527 19852 17536
rect 19800 17493 19809 17527
rect 19809 17493 19843 17527
rect 19843 17493 19852 17527
rect 19800 17484 19852 17493
rect 4447 17382 4499 17434
rect 4511 17382 4563 17434
rect 4575 17382 4627 17434
rect 4639 17382 4691 17434
rect 11378 17382 11430 17434
rect 11442 17382 11494 17434
rect 11506 17382 11558 17434
rect 11570 17382 11622 17434
rect 18308 17382 18360 17434
rect 18372 17382 18424 17434
rect 18436 17382 18488 17434
rect 18500 17382 18552 17434
rect 6092 17323 6144 17332
rect 6092 17289 6101 17323
rect 6101 17289 6135 17323
rect 6135 17289 6144 17323
rect 6092 17280 6144 17289
rect 6644 17323 6696 17332
rect 6644 17289 6653 17323
rect 6653 17289 6687 17323
rect 6687 17289 6696 17323
rect 6644 17280 6696 17289
rect 7564 17280 7616 17332
rect 8944 17280 8996 17332
rect 1584 17255 1636 17264
rect 1584 17221 1593 17255
rect 1593 17221 1627 17255
rect 1627 17221 1636 17255
rect 1584 17212 1636 17221
rect 8668 17212 8720 17264
rect 8300 17187 8352 17196
rect 8300 17153 8309 17187
rect 8309 17153 8343 17187
rect 8343 17153 8352 17187
rect 8300 17144 8352 17153
rect 6092 17076 6144 17128
rect 9864 17280 9916 17332
rect 10232 17280 10284 17332
rect 12256 17280 12308 17332
rect 13636 17280 13688 17332
rect 14096 17323 14148 17332
rect 14096 17289 14105 17323
rect 14105 17289 14139 17323
rect 14139 17289 14148 17323
rect 14096 17280 14148 17289
rect 14556 17280 14608 17332
rect 14740 17323 14792 17332
rect 14740 17289 14749 17323
rect 14749 17289 14783 17323
rect 14783 17289 14792 17323
rect 14740 17280 14792 17289
rect 15476 17280 15528 17332
rect 16856 17280 16908 17332
rect 20260 17280 20312 17332
rect 9772 17212 9824 17264
rect 11152 17212 11204 17264
rect 11244 17212 11296 17264
rect 14188 17212 14240 17264
rect 9680 17076 9732 17128
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 12164 17144 12216 17196
rect 12716 17187 12768 17196
rect 12716 17153 12725 17187
rect 12725 17153 12759 17187
rect 12759 17153 12768 17187
rect 12716 17144 12768 17153
rect 14740 17144 14792 17196
rect 15384 17144 15436 17196
rect 17132 17212 17184 17264
rect 16488 17187 16540 17196
rect 16488 17153 16497 17187
rect 16497 17153 16531 17187
rect 16531 17153 16540 17187
rect 16488 17144 16540 17153
rect 17040 17144 17092 17196
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 10968 17076 11020 17128
rect 13544 17076 13596 17128
rect 7380 17008 7432 17060
rect 8944 17008 8996 17060
rect 17408 17076 17460 17128
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 20076 17187 20128 17196
rect 18880 17076 18932 17128
rect 18972 17076 19024 17128
rect 20076 17153 20085 17187
rect 20085 17153 20119 17187
rect 20119 17153 20128 17187
rect 20076 17144 20128 17153
rect 21088 17076 21140 17128
rect 15016 17008 15068 17060
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 5356 16983 5408 16992
rect 5356 16949 5365 16983
rect 5365 16949 5399 16983
rect 5399 16949 5408 16983
rect 5356 16940 5408 16949
rect 5724 16983 5776 16992
rect 5724 16949 5733 16983
rect 5733 16949 5767 16983
rect 5767 16949 5776 16983
rect 5724 16940 5776 16949
rect 9036 16983 9088 16992
rect 9036 16949 9045 16983
rect 9045 16949 9079 16983
rect 9079 16949 9088 16983
rect 9036 16940 9088 16949
rect 9772 16940 9824 16992
rect 13636 16940 13688 16992
rect 15568 17008 15620 17060
rect 16488 16940 16540 16992
rect 17224 17008 17276 17060
rect 20076 17008 20128 17060
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 19432 16940 19484 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 7912 16838 7964 16890
rect 7976 16838 8028 16890
rect 8040 16838 8092 16890
rect 8104 16838 8156 16890
rect 14843 16838 14895 16890
rect 14907 16838 14959 16890
rect 14971 16838 15023 16890
rect 15035 16838 15087 16890
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 8484 16736 8536 16788
rect 8944 16736 8996 16788
rect 9036 16736 9088 16788
rect 10692 16736 10744 16788
rect 10968 16668 11020 16720
rect 5448 16643 5500 16652
rect 5448 16609 5457 16643
rect 5457 16609 5491 16643
rect 5491 16609 5500 16643
rect 5448 16600 5500 16609
rect 7288 16600 7340 16652
rect 8576 16643 8628 16652
rect 8300 16532 8352 16584
rect 8576 16609 8585 16643
rect 8585 16609 8619 16643
rect 8619 16609 8628 16643
rect 8576 16600 8628 16609
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 13728 16736 13780 16788
rect 13912 16736 13964 16788
rect 14280 16736 14332 16788
rect 15292 16779 15344 16788
rect 15292 16745 15301 16779
rect 15301 16745 15335 16779
rect 15335 16745 15344 16779
rect 15292 16736 15344 16745
rect 15568 16779 15620 16788
rect 15568 16745 15577 16779
rect 15577 16745 15611 16779
rect 15611 16745 15620 16779
rect 15568 16736 15620 16745
rect 16212 16779 16264 16788
rect 16212 16745 16221 16779
rect 16221 16745 16255 16779
rect 16255 16745 16264 16779
rect 16212 16736 16264 16745
rect 16488 16779 16540 16788
rect 16488 16745 16497 16779
rect 16497 16745 16531 16779
rect 16531 16745 16540 16779
rect 16488 16736 16540 16745
rect 16856 16736 16908 16788
rect 17500 16779 17552 16788
rect 17500 16745 17509 16779
rect 17509 16745 17543 16779
rect 17543 16745 17552 16779
rect 17500 16736 17552 16745
rect 17684 16736 17736 16788
rect 19892 16736 19944 16788
rect 11704 16668 11756 16720
rect 11980 16668 12032 16720
rect 12532 16668 12584 16720
rect 19524 16668 19576 16720
rect 11244 16600 11296 16652
rect 12164 16643 12216 16652
rect 12164 16609 12173 16643
rect 12173 16609 12207 16643
rect 12207 16609 12216 16643
rect 12164 16600 12216 16609
rect 10232 16532 10284 16584
rect 14280 16600 14332 16652
rect 14556 16600 14608 16652
rect 14924 16600 14976 16652
rect 18696 16643 18748 16652
rect 6552 16507 6604 16516
rect 6552 16473 6561 16507
rect 6561 16473 6595 16507
rect 6595 16473 6604 16507
rect 6552 16464 6604 16473
rect 8576 16464 8628 16516
rect 8944 16464 8996 16516
rect 9312 16464 9364 16516
rect 6000 16396 6052 16448
rect 8300 16396 8352 16448
rect 9680 16396 9732 16448
rect 9772 16396 9824 16448
rect 13360 16532 13412 16584
rect 14740 16575 14792 16584
rect 14740 16541 14749 16575
rect 14749 16541 14783 16575
rect 14783 16541 14792 16575
rect 14740 16532 14792 16541
rect 15016 16532 15068 16584
rect 16212 16532 16264 16584
rect 18696 16609 18705 16643
rect 18705 16609 18739 16643
rect 18739 16609 18748 16643
rect 18696 16600 18748 16609
rect 20628 16643 20680 16652
rect 20628 16609 20637 16643
rect 20637 16609 20671 16643
rect 20671 16609 20680 16643
rect 20628 16600 20680 16609
rect 21364 16643 21416 16652
rect 21364 16609 21373 16643
rect 21373 16609 21407 16643
rect 21407 16609 21416 16643
rect 21364 16600 21416 16609
rect 17040 16575 17092 16584
rect 17040 16541 17049 16575
rect 17049 16541 17083 16575
rect 17083 16541 17092 16575
rect 17040 16532 17092 16541
rect 19432 16532 19484 16584
rect 13544 16507 13596 16516
rect 13544 16473 13553 16507
rect 13553 16473 13587 16507
rect 13587 16473 13596 16507
rect 13544 16464 13596 16473
rect 15476 16464 15528 16516
rect 16304 16464 16356 16516
rect 12072 16396 12124 16448
rect 12440 16396 12492 16448
rect 12808 16396 12860 16448
rect 19800 16396 19852 16448
rect 20260 16439 20312 16448
rect 20260 16405 20269 16439
rect 20269 16405 20303 16439
rect 20303 16405 20312 16439
rect 20260 16396 20312 16405
rect 20812 16439 20864 16448
rect 20812 16405 20821 16439
rect 20821 16405 20855 16439
rect 20855 16405 20864 16439
rect 20812 16396 20864 16405
rect 4447 16294 4499 16346
rect 4511 16294 4563 16346
rect 4575 16294 4627 16346
rect 4639 16294 4691 16346
rect 11378 16294 11430 16346
rect 11442 16294 11494 16346
rect 11506 16294 11558 16346
rect 11570 16294 11622 16346
rect 18308 16294 18360 16346
rect 18372 16294 18424 16346
rect 18436 16294 18488 16346
rect 18500 16294 18552 16346
rect 6000 16235 6052 16244
rect 6000 16201 6009 16235
rect 6009 16201 6043 16235
rect 6043 16201 6052 16235
rect 6000 16192 6052 16201
rect 7012 16192 7064 16244
rect 10232 16192 10284 16244
rect 12348 16192 12400 16244
rect 15476 16192 15528 16244
rect 15752 16235 15804 16244
rect 15752 16201 15761 16235
rect 15761 16201 15795 16235
rect 15795 16201 15804 16235
rect 15752 16192 15804 16201
rect 17132 16192 17184 16244
rect 15568 16124 15620 16176
rect 5356 16031 5408 16040
rect 5356 15997 5365 16031
rect 5365 15997 5399 16031
rect 5399 15997 5408 16031
rect 5356 15988 5408 15997
rect 6460 15988 6512 16040
rect 6552 15988 6604 16040
rect 10232 16099 10284 16108
rect 10232 16065 10241 16099
rect 10241 16065 10275 16099
rect 10275 16065 10284 16099
rect 10232 16056 10284 16065
rect 10324 16099 10376 16108
rect 10324 16065 10333 16099
rect 10333 16065 10367 16099
rect 10367 16065 10376 16099
rect 10324 16056 10376 16065
rect 11244 16056 11296 16108
rect 12348 16056 12400 16108
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14740 16056 14792 16108
rect 15016 16056 15068 16108
rect 8576 15988 8628 16040
rect 9680 15988 9732 16040
rect 11888 15988 11940 16040
rect 12164 15988 12216 16040
rect 5724 15963 5776 15972
rect 5724 15929 5733 15963
rect 5733 15929 5767 15963
rect 5767 15929 5776 15963
rect 5724 15920 5776 15929
rect 5540 15852 5592 15904
rect 6368 15852 6420 15904
rect 8116 15920 8168 15972
rect 8392 15920 8444 15972
rect 8484 15852 8536 15904
rect 8576 15852 8628 15904
rect 12532 15988 12584 16040
rect 13268 15920 13320 15972
rect 14096 15920 14148 15972
rect 15660 15988 15712 16040
rect 20168 16192 20220 16244
rect 20352 16124 20404 16176
rect 17868 16099 17920 16108
rect 17868 16065 17877 16099
rect 17877 16065 17911 16099
rect 17911 16065 17920 16099
rect 17868 16056 17920 16065
rect 17684 16031 17736 16040
rect 17684 15997 17693 16031
rect 17693 15997 17727 16031
rect 17727 15997 17736 16031
rect 17684 15988 17736 15997
rect 18144 15988 18196 16040
rect 20168 16056 20220 16108
rect 19524 15988 19576 16040
rect 17960 15920 18012 15972
rect 19340 15920 19392 15972
rect 21364 15963 21416 15972
rect 21364 15929 21373 15963
rect 21373 15929 21407 15963
rect 21407 15929 21416 15963
rect 21364 15920 21416 15929
rect 11060 15852 11112 15904
rect 11980 15852 12032 15904
rect 14004 15852 14056 15904
rect 15292 15852 15344 15904
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 16120 15895 16172 15904
rect 16120 15861 16129 15895
rect 16129 15861 16163 15895
rect 16163 15861 16172 15895
rect 16120 15852 16172 15861
rect 16212 15852 16264 15904
rect 17040 15852 17092 15904
rect 19616 15852 19668 15904
rect 20260 15852 20312 15904
rect 7912 15750 7964 15802
rect 7976 15750 8028 15802
rect 8040 15750 8092 15802
rect 8104 15750 8156 15802
rect 14843 15750 14895 15802
rect 14907 15750 14959 15802
rect 14971 15750 15023 15802
rect 15035 15750 15087 15802
rect 5724 15691 5776 15700
rect 5724 15657 5733 15691
rect 5733 15657 5767 15691
rect 5767 15657 5776 15691
rect 5724 15648 5776 15657
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 8300 15648 8352 15700
rect 8668 15648 8720 15700
rect 9128 15648 9180 15700
rect 11244 15648 11296 15700
rect 12072 15648 12124 15700
rect 12440 15648 12492 15700
rect 12900 15648 12952 15700
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 14004 15691 14056 15700
rect 14004 15657 14013 15691
rect 14013 15657 14047 15691
rect 14047 15657 14056 15691
rect 14004 15648 14056 15657
rect 15292 15691 15344 15700
rect 15292 15657 15301 15691
rect 15301 15657 15335 15691
rect 15335 15657 15344 15691
rect 15292 15648 15344 15657
rect 16948 15691 17000 15700
rect 8484 15555 8536 15564
rect 8484 15521 8513 15555
rect 8513 15521 8536 15555
rect 8484 15512 8536 15521
rect 8668 15512 8720 15564
rect 10232 15555 10284 15564
rect 10232 15521 10266 15555
rect 10266 15521 10284 15555
rect 10232 15512 10284 15521
rect 9588 15444 9640 15496
rect 12808 15580 12860 15632
rect 16948 15657 16957 15691
rect 16957 15657 16991 15691
rect 16991 15657 17000 15691
rect 16948 15648 17000 15657
rect 17868 15648 17920 15700
rect 18696 15648 18748 15700
rect 19616 15648 19668 15700
rect 12624 15555 12676 15564
rect 12624 15521 12633 15555
rect 12633 15521 12667 15555
rect 12667 15521 12676 15555
rect 12624 15512 12676 15521
rect 13268 15512 13320 15564
rect 14096 15512 14148 15564
rect 5540 15376 5592 15428
rect 6368 15308 6420 15360
rect 6644 15308 6696 15360
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7380 15308 7432 15317
rect 10968 15376 11020 15428
rect 13820 15376 13872 15428
rect 15292 15512 15344 15564
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 15200 15444 15252 15496
rect 16120 15444 16172 15496
rect 16856 15580 16908 15632
rect 19432 15580 19484 15632
rect 16580 15444 16632 15496
rect 15936 15376 15988 15428
rect 19432 15444 19484 15496
rect 20812 15580 20864 15632
rect 12072 15308 12124 15360
rect 12256 15351 12308 15360
rect 12256 15317 12265 15351
rect 12265 15317 12299 15351
rect 12299 15317 12308 15351
rect 12256 15308 12308 15317
rect 14464 15308 14516 15360
rect 15108 15308 15160 15360
rect 15752 15351 15804 15360
rect 15752 15317 15761 15351
rect 15761 15317 15795 15351
rect 15795 15317 15804 15351
rect 15752 15308 15804 15317
rect 16028 15308 16080 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 4447 15206 4499 15258
rect 4511 15206 4563 15258
rect 4575 15206 4627 15258
rect 4639 15206 4691 15258
rect 11378 15206 11430 15258
rect 11442 15206 11494 15258
rect 11506 15206 11558 15258
rect 11570 15206 11622 15258
rect 18308 15206 18360 15258
rect 18372 15206 18424 15258
rect 18436 15206 18488 15258
rect 18500 15206 18552 15258
rect 9680 15104 9732 15156
rect 7840 15079 7892 15088
rect 7840 15045 7849 15079
rect 7849 15045 7883 15079
rect 7883 15045 7892 15079
rect 7840 15036 7892 15045
rect 8576 15011 8628 15020
rect 8576 14977 8585 15011
rect 8585 14977 8619 15011
rect 8619 14977 8628 15011
rect 8576 14968 8628 14977
rect 8668 15011 8720 15020
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 9772 15036 9824 15088
rect 11060 15104 11112 15156
rect 11980 15104 12032 15156
rect 12532 15104 12584 15156
rect 11888 15036 11940 15088
rect 14740 15036 14792 15088
rect 16580 15079 16632 15088
rect 10968 14968 11020 15020
rect 12348 14968 12400 15020
rect 12624 14968 12676 15020
rect 16580 15045 16589 15079
rect 16589 15045 16623 15079
rect 16623 15045 16632 15079
rect 16580 15036 16632 15045
rect 16672 15036 16724 15088
rect 7748 14832 7800 14884
rect 12256 14943 12308 14952
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 8392 14764 8444 14816
rect 9680 14832 9732 14884
rect 9772 14832 9824 14884
rect 9956 14875 10008 14884
rect 9956 14841 9965 14875
rect 9965 14841 9999 14875
rect 9999 14841 10008 14875
rect 9956 14832 10008 14841
rect 10232 14832 10284 14884
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 12256 14909 12265 14943
rect 12265 14909 12299 14943
rect 12299 14909 12308 14943
rect 12256 14900 12308 14909
rect 13636 14900 13688 14952
rect 13820 14943 13872 14952
rect 13820 14909 13854 14943
rect 13854 14909 13872 14943
rect 13820 14900 13872 14909
rect 15108 14900 15160 14952
rect 16212 14968 16264 15020
rect 15844 14900 15896 14952
rect 19340 14968 19392 15020
rect 19616 14968 19668 15020
rect 19248 14900 19300 14952
rect 19432 14900 19484 14952
rect 12164 14832 12216 14884
rect 15568 14832 15620 14884
rect 16212 14832 16264 14884
rect 12256 14764 12308 14816
rect 15752 14764 15804 14816
rect 15844 14764 15896 14816
rect 17960 14764 18012 14816
rect 19524 14832 19576 14884
rect 20352 14943 20404 14952
rect 20352 14909 20370 14943
rect 20370 14909 20404 14943
rect 20352 14900 20404 14909
rect 21364 14875 21416 14884
rect 21364 14841 21373 14875
rect 21373 14841 21407 14875
rect 21407 14841 21416 14875
rect 21364 14832 21416 14841
rect 19248 14807 19300 14816
rect 19248 14773 19257 14807
rect 19257 14773 19291 14807
rect 19291 14773 19300 14807
rect 19248 14764 19300 14773
rect 7912 14662 7964 14714
rect 7976 14662 8028 14714
rect 8040 14662 8092 14714
rect 8104 14662 8156 14714
rect 14843 14662 14895 14714
rect 14907 14662 14959 14714
rect 14971 14662 15023 14714
rect 15035 14662 15087 14714
rect 5540 14560 5592 14612
rect 6184 14560 6236 14612
rect 6460 14603 6512 14612
rect 6460 14569 6469 14603
rect 6469 14569 6503 14603
rect 6503 14569 6512 14603
rect 6460 14560 6512 14569
rect 7288 14560 7340 14612
rect 7656 14560 7708 14612
rect 8392 14603 8444 14612
rect 8392 14569 8401 14603
rect 8401 14569 8435 14603
rect 8435 14569 8444 14603
rect 8392 14560 8444 14569
rect 2688 14492 2740 14544
rect 13544 14560 13596 14612
rect 13912 14560 13964 14612
rect 14280 14560 14332 14612
rect 16672 14560 16724 14612
rect 17316 14560 17368 14612
rect 9220 14492 9272 14544
rect 10968 14492 11020 14544
rect 11704 14492 11756 14544
rect 7656 14467 7708 14476
rect 7656 14433 7665 14467
rect 7665 14433 7699 14467
rect 7699 14433 7708 14467
rect 7656 14424 7708 14433
rect 8300 14467 8352 14476
rect 8300 14433 8309 14467
rect 8309 14433 8343 14467
rect 8343 14433 8352 14467
rect 8300 14424 8352 14433
rect 9588 14424 9640 14476
rect 15384 14492 15436 14544
rect 12164 14467 12216 14476
rect 12164 14433 12173 14467
rect 12173 14433 12207 14467
rect 12207 14433 12216 14467
rect 12164 14424 12216 14433
rect 7380 14356 7432 14408
rect 11244 14356 11296 14408
rect 8852 14288 8904 14340
rect 12072 14356 12124 14408
rect 14188 14424 14240 14476
rect 16120 14424 16172 14476
rect 16488 14424 16540 14476
rect 18144 14467 18196 14476
rect 18144 14433 18153 14467
rect 18153 14433 18187 14467
rect 18187 14433 18196 14467
rect 18144 14424 18196 14433
rect 20352 14492 20404 14544
rect 12808 14399 12860 14408
rect 12808 14365 12817 14399
rect 12817 14365 12851 14399
rect 12851 14365 12860 14399
rect 12808 14356 12860 14365
rect 14464 14356 14516 14408
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 17868 14399 17920 14408
rect 7380 14220 7432 14272
rect 7840 14220 7892 14272
rect 8576 14220 8628 14272
rect 9312 14220 9364 14272
rect 9496 14220 9548 14272
rect 13912 14288 13964 14340
rect 14648 14288 14700 14340
rect 15200 14331 15252 14340
rect 15200 14297 15209 14331
rect 15209 14297 15243 14331
rect 15243 14297 15252 14331
rect 15200 14288 15252 14297
rect 15384 14288 15436 14340
rect 17868 14365 17877 14399
rect 17877 14365 17911 14399
rect 17911 14365 17920 14399
rect 17868 14356 17920 14365
rect 17960 14356 18012 14408
rect 19340 14424 19392 14476
rect 20444 14467 20496 14476
rect 20444 14433 20453 14467
rect 20453 14433 20487 14467
rect 20487 14433 20496 14467
rect 20444 14424 20496 14433
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 21180 14288 21232 14340
rect 21364 14331 21416 14340
rect 21364 14297 21373 14331
rect 21373 14297 21407 14331
rect 21407 14297 21416 14331
rect 21364 14288 21416 14297
rect 11060 14220 11112 14272
rect 11152 14263 11204 14272
rect 11152 14229 11161 14263
rect 11161 14229 11195 14263
rect 11195 14229 11204 14263
rect 18788 14263 18840 14272
rect 11152 14220 11204 14229
rect 18788 14229 18797 14263
rect 18797 14229 18831 14263
rect 18831 14229 18840 14263
rect 18788 14220 18840 14229
rect 19340 14220 19392 14272
rect 20352 14220 20404 14272
rect 4447 14118 4499 14170
rect 4511 14118 4563 14170
rect 4575 14118 4627 14170
rect 4639 14118 4691 14170
rect 11378 14118 11430 14170
rect 11442 14118 11494 14170
rect 11506 14118 11558 14170
rect 11570 14118 11622 14170
rect 18308 14118 18360 14170
rect 18372 14118 18424 14170
rect 18436 14118 18488 14170
rect 18500 14118 18552 14170
rect 6092 14016 6144 14068
rect 7748 14016 7800 14068
rect 8300 14016 8352 14068
rect 8760 14016 8812 14068
rect 10692 14016 10744 14068
rect 12164 14059 12216 14068
rect 12164 14025 12173 14059
rect 12173 14025 12207 14059
rect 12207 14025 12216 14059
rect 12164 14016 12216 14025
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 14096 14059 14148 14068
rect 14096 14025 14105 14059
rect 14105 14025 14139 14059
rect 14139 14025 14148 14059
rect 14096 14016 14148 14025
rect 17868 14016 17920 14068
rect 19892 14059 19944 14068
rect 5172 13948 5224 14000
rect 7840 13991 7892 14000
rect 7840 13957 7849 13991
rect 7849 13957 7883 13991
rect 7883 13957 7892 13991
rect 7840 13948 7892 13957
rect 9496 13948 9548 14000
rect 12440 13948 12492 14000
rect 16028 13948 16080 14000
rect 16488 13948 16540 14000
rect 5448 13880 5500 13932
rect 9956 13880 10008 13932
rect 7656 13812 7708 13864
rect 8852 13855 8904 13864
rect 8852 13821 8861 13855
rect 8861 13821 8895 13855
rect 8895 13821 8904 13855
rect 8852 13812 8904 13821
rect 10416 13812 10468 13864
rect 10324 13744 10376 13796
rect 11612 13812 11664 13864
rect 11888 13812 11940 13864
rect 12440 13855 12492 13864
rect 12440 13821 12449 13855
rect 12449 13821 12483 13855
rect 12483 13821 12492 13855
rect 12440 13812 12492 13821
rect 14464 13812 14516 13864
rect 15384 13880 15436 13932
rect 19892 14025 19901 14059
rect 19901 14025 19935 14059
rect 19935 14025 19944 14059
rect 19892 14016 19944 14025
rect 19248 13948 19300 14000
rect 16304 13855 16356 13864
rect 16304 13821 16313 13855
rect 16313 13821 16347 13855
rect 16347 13821 16356 13855
rect 16304 13812 16356 13821
rect 19432 13880 19484 13932
rect 19616 13880 19668 13932
rect 20352 13923 20404 13932
rect 20352 13889 20361 13923
rect 20361 13889 20395 13923
rect 20395 13889 20404 13923
rect 20352 13880 20404 13889
rect 18788 13812 18840 13864
rect 21364 13855 21416 13864
rect 21364 13821 21373 13855
rect 21373 13821 21407 13855
rect 21407 13821 21416 13855
rect 21364 13812 21416 13821
rect 10692 13787 10744 13796
rect 10692 13753 10710 13787
rect 10710 13753 10744 13787
rect 10692 13744 10744 13753
rect 12808 13744 12860 13796
rect 14556 13787 14608 13796
rect 14556 13753 14565 13787
rect 14565 13753 14599 13787
rect 14599 13753 14608 13787
rect 14556 13744 14608 13753
rect 15200 13744 15252 13796
rect 16212 13787 16264 13796
rect 16212 13753 16221 13787
rect 16221 13753 16255 13787
rect 16255 13753 16264 13787
rect 16212 13744 16264 13753
rect 16396 13744 16448 13796
rect 17868 13744 17920 13796
rect 20260 13787 20312 13796
rect 20260 13753 20269 13787
rect 20269 13753 20303 13787
rect 20303 13753 20312 13787
rect 20260 13744 20312 13753
rect 8944 13676 8996 13728
rect 12532 13676 12584 13728
rect 13360 13676 13412 13728
rect 14188 13676 14240 13728
rect 14740 13676 14792 13728
rect 15844 13719 15896 13728
rect 15844 13685 15853 13719
rect 15853 13685 15887 13719
rect 15887 13685 15896 13719
rect 15844 13676 15896 13685
rect 18880 13719 18932 13728
rect 18880 13685 18889 13719
rect 18889 13685 18923 13719
rect 18923 13685 18932 13719
rect 18880 13676 18932 13685
rect 19248 13719 19300 13728
rect 19248 13685 19257 13719
rect 19257 13685 19291 13719
rect 19291 13685 19300 13719
rect 19248 13676 19300 13685
rect 19708 13676 19760 13728
rect 7912 13574 7964 13626
rect 7976 13574 8028 13626
rect 8040 13574 8092 13626
rect 8104 13574 8156 13626
rect 14843 13574 14895 13626
rect 14907 13574 14959 13626
rect 14971 13574 15023 13626
rect 15035 13574 15087 13626
rect 6736 13515 6788 13524
rect 6736 13481 6745 13515
rect 6745 13481 6779 13515
rect 6779 13481 6788 13515
rect 6736 13472 6788 13481
rect 7748 13404 7800 13456
rect 8944 13404 8996 13456
rect 9864 13404 9916 13456
rect 10784 13404 10836 13456
rect 11060 13404 11112 13456
rect 6736 13336 6788 13388
rect 7104 13336 7156 13388
rect 8300 13379 8352 13388
rect 8300 13345 8309 13379
rect 8309 13345 8343 13379
rect 8343 13345 8352 13379
rect 8300 13336 8352 13345
rect 10048 13336 10100 13388
rect 11612 13379 11664 13388
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 12256 13447 12308 13456
rect 12256 13413 12265 13447
rect 12265 13413 12299 13447
rect 12299 13413 12308 13447
rect 14280 13472 14332 13524
rect 12256 13404 12308 13413
rect 10232 13268 10284 13320
rect 11796 13268 11848 13320
rect 12164 13268 12216 13320
rect 14648 13336 14700 13388
rect 12992 13268 13044 13320
rect 14096 13268 14148 13320
rect 15844 13472 15896 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 16948 13472 17000 13524
rect 19248 13472 19300 13524
rect 17408 13404 17460 13456
rect 17592 13404 17644 13456
rect 20168 13404 20220 13456
rect 21180 13447 21232 13456
rect 21180 13413 21189 13447
rect 21189 13413 21223 13447
rect 21223 13413 21232 13447
rect 21180 13404 21232 13413
rect 17040 13336 17092 13388
rect 17132 13336 17184 13388
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 17776 13311 17828 13320
rect 17776 13277 17785 13311
rect 17785 13277 17819 13311
rect 17819 13277 17828 13311
rect 17776 13268 17828 13277
rect 9680 13243 9732 13252
rect 9680 13209 9689 13243
rect 9689 13209 9723 13243
rect 9723 13209 9732 13243
rect 9680 13200 9732 13209
rect 7380 13132 7432 13184
rect 8392 13132 8444 13184
rect 10692 13132 10744 13184
rect 10876 13132 10928 13184
rect 16580 13200 16632 13252
rect 11888 13175 11940 13184
rect 11888 13141 11897 13175
rect 11897 13141 11931 13175
rect 11931 13141 11940 13175
rect 11888 13132 11940 13141
rect 11980 13132 12032 13184
rect 13268 13175 13320 13184
rect 13268 13141 13277 13175
rect 13277 13141 13311 13175
rect 13311 13141 13320 13175
rect 13268 13132 13320 13141
rect 17960 13200 18012 13252
rect 18144 13268 18196 13320
rect 20076 13268 20128 13320
rect 20628 13200 20680 13252
rect 21364 13243 21416 13252
rect 21364 13209 21373 13243
rect 21373 13209 21407 13243
rect 21407 13209 21416 13243
rect 21364 13200 21416 13209
rect 18052 13175 18104 13184
rect 18052 13141 18061 13175
rect 18061 13141 18095 13175
rect 18095 13141 18104 13175
rect 18052 13132 18104 13141
rect 4447 13030 4499 13082
rect 4511 13030 4563 13082
rect 4575 13030 4627 13082
rect 4639 13030 4691 13082
rect 11378 13030 11430 13082
rect 11442 13030 11494 13082
rect 11506 13030 11558 13082
rect 11570 13030 11622 13082
rect 18308 13030 18360 13082
rect 18372 13030 18424 13082
rect 18436 13030 18488 13082
rect 18500 13030 18552 13082
rect 7748 12928 7800 12980
rect 10876 12928 10928 12980
rect 11244 12928 11296 12980
rect 11980 12928 12032 12980
rect 5080 12860 5132 12912
rect 6828 12860 6880 12912
rect 7656 12860 7708 12912
rect 9864 12903 9916 12912
rect 9864 12869 9873 12903
rect 9873 12869 9907 12903
rect 9907 12869 9916 12903
rect 9864 12860 9916 12869
rect 9956 12860 10008 12912
rect 10232 12860 10284 12912
rect 12164 12860 12216 12912
rect 10784 12835 10836 12844
rect 10784 12801 10793 12835
rect 10793 12801 10827 12835
rect 10827 12801 10836 12835
rect 10784 12792 10836 12801
rect 11888 12792 11940 12844
rect 7288 12724 7340 12776
rect 9404 12724 9456 12776
rect 8392 12656 8444 12708
rect 9588 12724 9640 12776
rect 14464 12860 14516 12912
rect 15292 12928 15344 12980
rect 18880 12928 18932 12980
rect 19708 12928 19760 12980
rect 14096 12835 14148 12844
rect 13268 12724 13320 12776
rect 14096 12801 14105 12835
rect 14105 12801 14139 12835
rect 14139 12801 14148 12835
rect 14096 12792 14148 12801
rect 16212 12792 16264 12844
rect 17132 12792 17184 12844
rect 20628 12792 20680 12844
rect 14464 12724 14516 12776
rect 14740 12724 14792 12776
rect 15016 12724 15068 12776
rect 17408 12724 17460 12776
rect 17684 12767 17736 12776
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 19616 12767 19668 12776
rect 19616 12733 19634 12767
rect 19634 12733 19668 12767
rect 19616 12724 19668 12733
rect 10416 12656 10468 12708
rect 6920 12588 6972 12640
rect 7656 12588 7708 12640
rect 8484 12588 8536 12640
rect 9864 12588 9916 12640
rect 10876 12588 10928 12640
rect 11152 12588 11204 12640
rect 11888 12631 11940 12640
rect 11888 12597 11897 12631
rect 11897 12597 11931 12631
rect 11931 12597 11940 12631
rect 11888 12588 11940 12597
rect 13912 12631 13964 12640
rect 13912 12597 13921 12631
rect 13921 12597 13955 12631
rect 13955 12597 13964 12631
rect 15844 12656 15896 12708
rect 17592 12656 17644 12708
rect 19432 12656 19484 12708
rect 20076 12656 20128 12708
rect 13912 12588 13964 12597
rect 16120 12631 16172 12640
rect 16120 12597 16129 12631
rect 16129 12597 16163 12631
rect 16163 12597 16172 12631
rect 16120 12588 16172 12597
rect 16764 12588 16816 12640
rect 17960 12588 18012 12640
rect 20720 12588 20772 12640
rect 20904 12631 20956 12640
rect 20904 12597 20913 12631
rect 20913 12597 20947 12631
rect 20947 12597 20956 12631
rect 20904 12588 20956 12597
rect 7912 12486 7964 12538
rect 7976 12486 8028 12538
rect 8040 12486 8092 12538
rect 8104 12486 8156 12538
rect 14843 12486 14895 12538
rect 14907 12486 14959 12538
rect 14971 12486 15023 12538
rect 15035 12486 15087 12538
rect 6092 12384 6144 12436
rect 10232 12384 10284 12436
rect 11704 12427 11756 12436
rect 11704 12393 11713 12427
rect 11713 12393 11747 12427
rect 11747 12393 11756 12427
rect 11704 12384 11756 12393
rect 11796 12384 11848 12436
rect 13820 12384 13872 12436
rect 14096 12384 14148 12436
rect 14556 12427 14608 12436
rect 14556 12393 14565 12427
rect 14565 12393 14599 12427
rect 14599 12393 14608 12427
rect 14556 12384 14608 12393
rect 16304 12384 16356 12436
rect 16856 12384 16908 12436
rect 17040 12384 17092 12436
rect 18052 12384 18104 12436
rect 19156 12384 19208 12436
rect 19616 12384 19668 12436
rect 7748 12248 7800 12300
rect 8116 12291 8168 12300
rect 8116 12257 8125 12291
rect 8125 12257 8159 12291
rect 8159 12257 8168 12291
rect 8116 12248 8168 12257
rect 8300 12248 8352 12300
rect 9404 12316 9456 12368
rect 2228 12180 2280 12232
rect 7104 12180 7156 12232
rect 8484 12180 8536 12232
rect 10324 12248 10376 12300
rect 10876 12248 10928 12300
rect 11888 12316 11940 12368
rect 13544 12316 13596 12368
rect 13728 12316 13780 12368
rect 18236 12316 18288 12368
rect 20076 12316 20128 12368
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 13268 12248 13320 12300
rect 14004 12248 14056 12300
rect 10692 12180 10744 12232
rect 10784 12180 10836 12232
rect 11704 12180 11756 12232
rect 12440 12180 12492 12232
rect 8760 12155 8812 12164
rect 8760 12121 8769 12155
rect 8769 12121 8803 12155
rect 8803 12121 8812 12155
rect 8760 12112 8812 12121
rect 9036 12112 9088 12164
rect 9220 12112 9272 12164
rect 6276 12044 6328 12096
rect 6920 12044 6972 12096
rect 11980 12112 12032 12164
rect 10508 12044 10560 12096
rect 14740 12180 14792 12232
rect 16580 12248 16632 12300
rect 17040 12248 17092 12300
rect 17868 12248 17920 12300
rect 18880 12291 18932 12300
rect 16212 12180 16264 12232
rect 17132 12223 17184 12232
rect 17132 12189 17141 12223
rect 17141 12189 17175 12223
rect 17175 12189 17184 12223
rect 17132 12180 17184 12189
rect 17960 12223 18012 12232
rect 17960 12189 17969 12223
rect 17969 12189 18003 12223
rect 18003 12189 18012 12223
rect 17960 12180 18012 12189
rect 18880 12257 18889 12291
rect 18889 12257 18923 12291
rect 18923 12257 18932 12291
rect 18880 12248 18932 12257
rect 20628 12248 20680 12300
rect 18972 12180 19024 12232
rect 13728 12112 13780 12164
rect 14004 12044 14056 12096
rect 18788 12112 18840 12164
rect 16580 12044 16632 12096
rect 4447 11942 4499 11994
rect 4511 11942 4563 11994
rect 4575 11942 4627 11994
rect 4639 11942 4691 11994
rect 11378 11942 11430 11994
rect 11442 11942 11494 11994
rect 11506 11942 11558 11994
rect 11570 11942 11622 11994
rect 18308 11942 18360 11994
rect 18372 11942 18424 11994
rect 18436 11942 18488 11994
rect 18500 11942 18552 11994
rect 7748 11883 7800 11892
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 8760 11840 8812 11892
rect 9312 11840 9364 11892
rect 10048 11883 10100 11892
rect 10048 11849 10057 11883
rect 10057 11849 10091 11883
rect 10091 11849 10100 11883
rect 10048 11840 10100 11849
rect 10232 11840 10284 11892
rect 11796 11840 11848 11892
rect 9772 11815 9824 11824
rect 9772 11781 9781 11815
rect 9781 11781 9815 11815
rect 9815 11781 9824 11815
rect 9772 11772 9824 11781
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 10508 11747 10560 11756
rect 10508 11713 10517 11747
rect 10517 11713 10551 11747
rect 10551 11713 10560 11747
rect 10508 11704 10560 11713
rect 12532 11840 12584 11892
rect 13268 11883 13320 11892
rect 13268 11849 13277 11883
rect 13277 11849 13311 11883
rect 13311 11849 13320 11883
rect 13268 11840 13320 11849
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 14464 11840 14516 11892
rect 16488 11840 16540 11892
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 13820 11772 13872 11824
rect 13268 11704 13320 11756
rect 16304 11772 16356 11824
rect 19892 11840 19944 11892
rect 20628 11840 20680 11892
rect 14556 11704 14608 11756
rect 8484 11636 8536 11688
rect 9220 11636 9272 11688
rect 10232 11636 10284 11688
rect 7380 11568 7432 11620
rect 10968 11636 11020 11688
rect 11980 11636 12032 11688
rect 14280 11636 14332 11688
rect 14372 11636 14424 11688
rect 15752 11704 15804 11756
rect 15476 11636 15528 11688
rect 18604 11636 18656 11688
rect 18972 11679 19024 11688
rect 18972 11645 18990 11679
rect 18990 11645 19024 11679
rect 18972 11636 19024 11645
rect 19340 11636 19392 11688
rect 13084 11568 13136 11620
rect 13820 11568 13872 11620
rect 14096 11568 14148 11620
rect 14648 11568 14700 11620
rect 8208 11500 8260 11552
rect 8852 11500 8904 11552
rect 13636 11500 13688 11552
rect 13728 11500 13780 11552
rect 14556 11500 14608 11552
rect 14740 11500 14792 11552
rect 15752 11500 15804 11552
rect 15844 11500 15896 11552
rect 21180 11568 21232 11620
rect 17868 11543 17920 11552
rect 17868 11509 17877 11543
rect 17877 11509 17911 11543
rect 17911 11509 17920 11543
rect 17868 11500 17920 11509
rect 18144 11500 18196 11552
rect 19156 11500 19208 11552
rect 19524 11543 19576 11552
rect 19524 11509 19533 11543
rect 19533 11509 19567 11543
rect 19567 11509 19576 11543
rect 19524 11500 19576 11509
rect 7912 11398 7964 11450
rect 7976 11398 8028 11450
rect 8040 11398 8092 11450
rect 8104 11398 8156 11450
rect 14843 11398 14895 11450
rect 14907 11398 14959 11450
rect 14971 11398 15023 11450
rect 15035 11398 15087 11450
rect 7380 11296 7432 11348
rect 8208 11296 8260 11348
rect 11612 11296 11664 11348
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 14280 11296 14332 11348
rect 16120 11296 16172 11348
rect 16488 11296 16540 11348
rect 9404 11228 9456 11280
rect 9772 11228 9824 11280
rect 12256 11228 12308 11280
rect 17040 11296 17092 11348
rect 18604 11296 18656 11348
rect 20812 11296 20864 11348
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 10784 11160 10836 11212
rect 10968 11160 11020 11212
rect 12072 11160 12124 11212
rect 12348 11203 12400 11212
rect 12348 11169 12357 11203
rect 12357 11169 12391 11203
rect 12391 11169 12400 11203
rect 12348 11160 12400 11169
rect 13636 11160 13688 11212
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 17868 11160 17920 11212
rect 18788 11160 18840 11212
rect 19708 11160 19760 11212
rect 4804 10956 4856 11008
rect 5632 10956 5684 11008
rect 9036 11092 9088 11144
rect 8392 10956 8444 11008
rect 9220 11024 9272 11076
rect 10324 11024 10376 11076
rect 10600 11024 10652 11076
rect 13084 11135 13136 11144
rect 10876 11024 10928 11076
rect 9956 10956 10008 11008
rect 10692 10999 10744 11008
rect 10692 10965 10701 10999
rect 10701 10965 10735 10999
rect 10735 10965 10744 10999
rect 10692 10956 10744 10965
rect 11704 10956 11756 11008
rect 13084 11101 13093 11135
rect 13093 11101 13127 11135
rect 13127 11101 13136 11135
rect 13084 11092 13136 11101
rect 13268 11135 13320 11144
rect 13268 11101 13277 11135
rect 13277 11101 13311 11135
rect 13311 11101 13320 11135
rect 13268 11092 13320 11101
rect 19064 11135 19116 11144
rect 19064 11101 19073 11135
rect 19073 11101 19107 11135
rect 19107 11101 19116 11135
rect 19064 11092 19116 11101
rect 19340 11092 19392 11144
rect 14372 10956 14424 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 4447 10854 4499 10906
rect 4511 10854 4563 10906
rect 4575 10854 4627 10906
rect 4639 10854 4691 10906
rect 11378 10854 11430 10906
rect 11442 10854 11494 10906
rect 11506 10854 11558 10906
rect 11570 10854 11622 10906
rect 18308 10854 18360 10906
rect 18372 10854 18424 10906
rect 18436 10854 18488 10906
rect 18500 10854 18552 10906
rect 1768 10752 1820 10804
rect 7380 10795 7432 10804
rect 7380 10761 7389 10795
rect 7389 10761 7423 10795
rect 7423 10761 7432 10795
rect 7380 10752 7432 10761
rect 12256 10752 12308 10804
rect 13268 10752 13320 10804
rect 13912 10752 13964 10804
rect 10876 10684 10928 10736
rect 15844 10684 15896 10736
rect 12348 10616 12400 10668
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 8576 10548 8628 10600
rect 8852 10548 8904 10600
rect 9956 10548 10008 10600
rect 10692 10548 10744 10600
rect 11060 10548 11112 10600
rect 14004 10616 14056 10668
rect 17868 10752 17920 10804
rect 18972 10752 19024 10804
rect 20904 10752 20956 10804
rect 18788 10684 18840 10736
rect 17040 10616 17092 10668
rect 17408 10659 17460 10668
rect 13820 10548 13872 10600
rect 14648 10548 14700 10600
rect 16580 10548 16632 10600
rect 17408 10625 17417 10659
rect 17417 10625 17451 10659
rect 17451 10625 17460 10659
rect 17408 10616 17460 10625
rect 18880 10616 18932 10668
rect 21180 10659 21232 10668
rect 21180 10625 21189 10659
rect 21189 10625 21223 10659
rect 21223 10625 21232 10659
rect 21180 10616 21232 10625
rect 17316 10548 17368 10600
rect 15292 10480 15344 10532
rect 19340 10480 19392 10532
rect 20352 10480 20404 10532
rect 4252 10412 4304 10464
rect 8852 10412 8904 10464
rect 9128 10455 9180 10464
rect 9128 10421 9137 10455
rect 9137 10421 9171 10455
rect 9171 10421 9180 10455
rect 9128 10412 9180 10421
rect 9588 10455 9640 10464
rect 9588 10421 9597 10455
rect 9597 10421 9631 10455
rect 9631 10421 9640 10455
rect 9588 10412 9640 10421
rect 9864 10412 9916 10464
rect 11060 10412 11112 10464
rect 11704 10412 11756 10464
rect 12440 10412 12492 10464
rect 12716 10455 12768 10464
rect 12716 10421 12725 10455
rect 12725 10421 12759 10455
rect 12759 10421 12768 10455
rect 12716 10412 12768 10421
rect 12808 10455 12860 10464
rect 12808 10421 12817 10455
rect 12817 10421 12851 10455
rect 12851 10421 12860 10455
rect 12808 10412 12860 10421
rect 14004 10412 14056 10464
rect 14188 10455 14240 10464
rect 14188 10421 14197 10455
rect 14197 10421 14231 10455
rect 14231 10421 14240 10455
rect 14188 10412 14240 10421
rect 14740 10412 14792 10464
rect 16672 10412 16724 10464
rect 18236 10412 18288 10464
rect 20904 10455 20956 10464
rect 20904 10421 20913 10455
rect 20913 10421 20947 10455
rect 20947 10421 20956 10455
rect 20904 10412 20956 10421
rect 21088 10412 21140 10464
rect 7912 10310 7964 10362
rect 7976 10310 8028 10362
rect 8040 10310 8092 10362
rect 8104 10310 8156 10362
rect 14843 10310 14895 10362
rect 14907 10310 14959 10362
rect 14971 10310 15023 10362
rect 15035 10310 15087 10362
rect 8392 10208 8444 10260
rect 8852 10208 8904 10260
rect 10416 10208 10468 10260
rect 9128 10140 9180 10192
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 4804 9868 4856 9920
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 10876 10072 10928 10124
rect 11060 10115 11112 10124
rect 11060 10081 11094 10115
rect 11094 10081 11112 10115
rect 11060 10072 11112 10081
rect 11796 10072 11848 10124
rect 13912 10208 13964 10260
rect 14188 10208 14240 10260
rect 15936 10251 15988 10260
rect 15936 10217 15945 10251
rect 15945 10217 15979 10251
rect 15979 10217 15988 10251
rect 15936 10208 15988 10217
rect 18236 10251 18288 10260
rect 12624 10140 12676 10192
rect 12992 10072 13044 10124
rect 14372 10140 14424 10192
rect 10048 10004 10100 10056
rect 10692 10047 10744 10056
rect 10692 10013 10701 10047
rect 10701 10013 10735 10047
rect 10735 10013 10744 10047
rect 10692 10004 10744 10013
rect 13544 10004 13596 10056
rect 15016 10047 15068 10056
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 18236 10217 18245 10251
rect 18245 10217 18279 10251
rect 18279 10217 18288 10251
rect 18236 10208 18288 10217
rect 18696 10208 18748 10260
rect 19708 10208 19760 10260
rect 20996 10251 21048 10260
rect 20996 10217 21005 10251
rect 21005 10217 21039 10251
rect 21039 10217 21048 10251
rect 20996 10208 21048 10217
rect 20168 10183 20220 10192
rect 20168 10149 20177 10183
rect 20177 10149 20211 10183
rect 20211 10149 20220 10183
rect 20168 10140 20220 10149
rect 17960 10072 18012 10124
rect 18788 10072 18840 10124
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 16028 10004 16080 10056
rect 18144 10004 18196 10056
rect 18604 10004 18656 10056
rect 20260 10047 20312 10056
rect 20260 10013 20269 10047
rect 20269 10013 20303 10047
rect 20303 10013 20312 10047
rect 20260 10004 20312 10013
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 17960 9936 18012 9988
rect 17408 9868 17460 9920
rect 21272 9911 21324 9920
rect 21272 9877 21281 9911
rect 21281 9877 21315 9911
rect 21315 9877 21324 9911
rect 21272 9868 21324 9877
rect 4447 9766 4499 9818
rect 4511 9766 4563 9818
rect 4575 9766 4627 9818
rect 4639 9766 4691 9818
rect 11378 9766 11430 9818
rect 11442 9766 11494 9818
rect 11506 9766 11558 9818
rect 11570 9766 11622 9818
rect 18308 9766 18360 9818
rect 18372 9766 18424 9818
rect 18436 9766 18488 9818
rect 18500 9766 18552 9818
rect 7380 9664 7432 9716
rect 9496 9664 9548 9716
rect 13544 9664 13596 9716
rect 9588 9596 9640 9648
rect 10048 9528 10100 9580
rect 10324 9528 10376 9580
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 9680 9460 9732 9512
rect 9864 9460 9916 9512
rect 13268 9596 13320 9648
rect 14648 9664 14700 9716
rect 16028 9664 16080 9716
rect 15016 9596 15068 9648
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 12624 9528 12676 9580
rect 14556 9571 14608 9580
rect 14556 9537 14565 9571
rect 14565 9537 14599 9571
rect 14599 9537 14608 9571
rect 14556 9528 14608 9537
rect 15384 9528 15436 9580
rect 16672 9528 16724 9580
rect 18604 9664 18656 9716
rect 20352 9664 20404 9716
rect 20996 9571 21048 9580
rect 9404 9392 9456 9444
rect 17040 9460 17092 9512
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 12440 9392 12492 9444
rect 8392 9367 8444 9376
rect 8392 9333 8401 9367
rect 8401 9333 8435 9367
rect 8435 9333 8444 9367
rect 8392 9324 8444 9333
rect 8668 9324 8720 9376
rect 9036 9324 9088 9376
rect 10784 9367 10836 9376
rect 10784 9333 10793 9367
rect 10793 9333 10827 9367
rect 10827 9333 10836 9367
rect 10784 9324 10836 9333
rect 12072 9324 12124 9376
rect 12532 9324 12584 9376
rect 13268 9367 13320 9376
rect 13268 9333 13277 9367
rect 13277 9333 13311 9367
rect 13311 9333 13320 9367
rect 13268 9324 13320 9333
rect 13360 9367 13412 9376
rect 13360 9333 13369 9367
rect 13369 9333 13403 9367
rect 13403 9333 13412 9367
rect 14004 9367 14056 9376
rect 13360 9324 13412 9333
rect 14004 9333 14013 9367
rect 14013 9333 14047 9367
rect 14047 9333 14056 9367
rect 14004 9324 14056 9333
rect 14280 9324 14332 9376
rect 15108 9392 15160 9444
rect 17408 9435 17460 9444
rect 17408 9401 17442 9435
rect 17442 9401 17460 9435
rect 17408 9392 17460 9401
rect 20168 9460 20220 9512
rect 19340 9392 19392 9444
rect 15292 9324 15344 9376
rect 15660 9324 15712 9376
rect 16120 9367 16172 9376
rect 16120 9333 16129 9367
rect 16129 9333 16163 9367
rect 16163 9333 16172 9367
rect 16120 9324 16172 9333
rect 16580 9324 16632 9376
rect 16948 9324 17000 9376
rect 19156 9324 19208 9376
rect 20812 9367 20864 9376
rect 20812 9333 20821 9367
rect 20821 9333 20855 9367
rect 20855 9333 20864 9367
rect 20812 9324 20864 9333
rect 7912 9222 7964 9274
rect 7976 9222 8028 9274
rect 8040 9222 8092 9274
rect 8104 9222 8156 9274
rect 14843 9222 14895 9274
rect 14907 9222 14959 9274
rect 14971 9222 15023 9274
rect 15035 9222 15087 9274
rect 9496 9120 9548 9172
rect 10876 9120 10928 9172
rect 11060 9163 11112 9172
rect 11060 9129 11069 9163
rect 11069 9129 11103 9163
rect 11103 9129 11112 9163
rect 11060 9120 11112 9129
rect 11152 9120 11204 9172
rect 11796 9120 11848 9172
rect 12072 9163 12124 9172
rect 12072 9129 12081 9163
rect 12081 9129 12115 9163
rect 12115 9129 12124 9163
rect 12072 9120 12124 9129
rect 14004 9120 14056 9172
rect 14556 9120 14608 9172
rect 6368 9052 6420 9104
rect 9404 9052 9456 9104
rect 6276 8984 6328 9036
rect 7196 8984 7248 9036
rect 9128 8984 9180 9036
rect 7472 8916 7524 8968
rect 7656 8916 7708 8968
rect 9404 8916 9456 8968
rect 10692 9052 10744 9104
rect 10784 9052 10836 9104
rect 16304 9120 16356 9172
rect 17500 9163 17552 9172
rect 17500 9129 17509 9163
rect 17509 9129 17543 9163
rect 17543 9129 17552 9163
rect 17500 9120 17552 9129
rect 17040 9052 17092 9104
rect 18144 9120 18196 9172
rect 20812 9120 20864 9172
rect 9588 8984 9640 9036
rect 10324 8984 10376 9036
rect 11704 9027 11756 9036
rect 11704 8993 11713 9027
rect 11713 8993 11747 9027
rect 11747 8993 11756 9027
rect 11704 8984 11756 8993
rect 14372 8984 14424 9036
rect 14832 9027 14884 9036
rect 14832 8993 14866 9027
rect 14866 8993 14884 9027
rect 14832 8984 14884 8993
rect 15384 8984 15436 9036
rect 15568 8984 15620 9036
rect 17408 8984 17460 9036
rect 12072 8916 12124 8968
rect 13728 8959 13780 8968
rect 8116 8848 8168 8900
rect 7656 8780 7708 8832
rect 8668 8780 8720 8832
rect 10692 8780 10744 8832
rect 13728 8925 13737 8959
rect 13737 8925 13771 8959
rect 13771 8925 13780 8959
rect 13728 8916 13780 8925
rect 14004 8916 14056 8968
rect 14464 8916 14516 8968
rect 14372 8848 14424 8900
rect 18052 8916 18104 8968
rect 18696 8959 18748 8968
rect 18696 8925 18705 8959
rect 18705 8925 18739 8959
rect 18739 8925 18748 8959
rect 18696 8916 18748 8925
rect 20168 8984 20220 9036
rect 19064 8916 19116 8968
rect 20996 8916 21048 8968
rect 12808 8823 12860 8832
rect 12808 8789 12817 8823
rect 12817 8789 12851 8823
rect 12851 8789 12860 8823
rect 12808 8780 12860 8789
rect 14464 8780 14516 8832
rect 18788 8780 18840 8832
rect 19524 8780 19576 8832
rect 19984 8823 20036 8832
rect 19984 8789 19993 8823
rect 19993 8789 20027 8823
rect 20027 8789 20036 8823
rect 19984 8780 20036 8789
rect 4447 8678 4499 8730
rect 4511 8678 4563 8730
rect 4575 8678 4627 8730
rect 4639 8678 4691 8730
rect 11378 8678 11430 8730
rect 11442 8678 11494 8730
rect 11506 8678 11558 8730
rect 11570 8678 11622 8730
rect 18308 8678 18360 8730
rect 18372 8678 18424 8730
rect 18436 8678 18488 8730
rect 18500 8678 18552 8730
rect 7196 8619 7248 8628
rect 7196 8585 7205 8619
rect 7205 8585 7239 8619
rect 7239 8585 7248 8619
rect 7196 8576 7248 8585
rect 9404 8576 9456 8628
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 9680 8576 9732 8628
rect 9956 8508 10008 8560
rect 10968 8508 11020 8560
rect 11152 8576 11204 8628
rect 13452 8576 13504 8628
rect 13728 8576 13780 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 14280 8619 14332 8628
rect 13820 8576 13872 8585
rect 14280 8585 14289 8619
rect 14289 8585 14323 8619
rect 14323 8585 14332 8619
rect 14280 8576 14332 8585
rect 14372 8576 14424 8628
rect 17960 8576 18012 8628
rect 18696 8576 18748 8628
rect 19248 8576 19300 8628
rect 7748 8372 7800 8424
rect 8116 8372 8168 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 11060 8440 11112 8492
rect 18144 8508 18196 8560
rect 8484 8304 8536 8356
rect 8760 8304 8812 8356
rect 10140 8304 10192 8356
rect 10784 8304 10836 8356
rect 10876 8304 10928 8356
rect 11336 8304 11388 8356
rect 12440 8415 12492 8424
rect 12440 8381 12474 8415
rect 12474 8381 12492 8415
rect 12440 8372 12492 8381
rect 14464 8372 14516 8424
rect 14648 8440 14700 8492
rect 14832 8483 14884 8492
rect 14832 8449 14841 8483
rect 14841 8449 14875 8483
rect 14875 8449 14884 8483
rect 14832 8440 14884 8449
rect 15568 8440 15620 8492
rect 15752 8440 15804 8492
rect 16856 8372 16908 8424
rect 18052 8440 18104 8492
rect 19984 8508 20036 8560
rect 18788 8372 18840 8424
rect 19156 8415 19208 8424
rect 19156 8381 19165 8415
rect 19165 8381 19199 8415
rect 19199 8381 19208 8415
rect 19156 8372 19208 8381
rect 19340 8372 19392 8424
rect 7196 8236 7248 8288
rect 7472 8236 7524 8288
rect 10968 8236 11020 8288
rect 11796 8236 11848 8288
rect 12900 8304 12952 8356
rect 14832 8304 14884 8356
rect 16028 8304 16080 8356
rect 17592 8304 17644 8356
rect 14556 8236 14608 8288
rect 20628 8304 20680 8356
rect 20996 8304 21048 8356
rect 18052 8236 18104 8288
rect 18972 8236 19024 8288
rect 19248 8236 19300 8288
rect 7912 8134 7964 8186
rect 7976 8134 8028 8186
rect 8040 8134 8092 8186
rect 8104 8134 8156 8186
rect 14843 8134 14895 8186
rect 14907 8134 14959 8186
rect 14971 8134 15023 8186
rect 15035 8134 15087 8186
rect 7012 8075 7064 8084
rect 7012 8041 7021 8075
rect 7021 8041 7055 8075
rect 7055 8041 7064 8075
rect 7012 8032 7064 8041
rect 9128 8032 9180 8084
rect 9864 8032 9916 8084
rect 10232 8032 10284 8084
rect 10968 8032 11020 8084
rect 11704 8032 11756 8084
rect 12072 8075 12124 8084
rect 12072 8041 12081 8075
rect 12081 8041 12115 8075
rect 12115 8041 12124 8075
rect 12072 8032 12124 8041
rect 12348 8032 12400 8084
rect 11796 7964 11848 8016
rect 13728 7964 13780 8016
rect 14464 8007 14516 8016
rect 14464 7973 14473 8007
rect 14473 7973 14507 8007
rect 14507 7973 14516 8007
rect 14464 7964 14516 7973
rect 14648 8032 14700 8084
rect 17684 8075 17736 8084
rect 17684 8041 17693 8075
rect 17693 8041 17727 8075
rect 17727 8041 17736 8075
rect 17684 8032 17736 8041
rect 18788 8075 18840 8084
rect 18788 8041 18797 8075
rect 18797 8041 18831 8075
rect 18831 8041 18840 8075
rect 18788 8032 18840 8041
rect 20996 8032 21048 8084
rect 17868 7964 17920 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 8852 7828 8904 7880
rect 9036 7828 9088 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10048 7828 10100 7880
rect 10784 7896 10836 7948
rect 11336 7896 11388 7948
rect 15752 7896 15804 7948
rect 17776 7939 17828 7948
rect 17776 7905 17785 7939
rect 17785 7905 17819 7939
rect 17819 7905 17828 7939
rect 17776 7896 17828 7905
rect 18052 7896 18104 7948
rect 19340 7896 19392 7948
rect 20536 7896 20588 7948
rect 9864 7760 9916 7812
rect 11152 7828 11204 7880
rect 11796 7828 11848 7880
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 16304 7871 16356 7880
rect 16304 7837 16313 7871
rect 16313 7837 16347 7871
rect 16347 7837 16356 7871
rect 16304 7828 16356 7837
rect 16396 7828 16448 7880
rect 17316 7828 17368 7880
rect 12072 7760 12124 7812
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 18972 7692 19024 7744
rect 19156 7735 19208 7744
rect 19156 7701 19165 7735
rect 19165 7701 19199 7735
rect 19199 7701 19208 7735
rect 19156 7692 19208 7701
rect 20996 7692 21048 7744
rect 4447 7590 4499 7642
rect 4511 7590 4563 7642
rect 4575 7590 4627 7642
rect 4639 7590 4691 7642
rect 11378 7590 11430 7642
rect 11442 7590 11494 7642
rect 11506 7590 11558 7642
rect 11570 7590 11622 7642
rect 18308 7590 18360 7642
rect 18372 7590 18424 7642
rect 18436 7590 18488 7642
rect 18500 7590 18552 7642
rect 7656 7488 7708 7540
rect 6828 7420 6880 7472
rect 8116 7420 8168 7472
rect 10048 7488 10100 7540
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 11428 7420 11480 7472
rect 11520 7420 11572 7472
rect 12256 7488 12308 7540
rect 11060 7352 11112 7404
rect 14464 7420 14516 7472
rect 15752 7488 15804 7540
rect 16304 7488 16356 7540
rect 15476 7420 15528 7472
rect 13912 7352 13964 7404
rect 7748 7284 7800 7336
rect 7564 7148 7616 7200
rect 9036 7216 9088 7268
rect 9864 7284 9916 7336
rect 10048 7327 10100 7336
rect 10048 7293 10082 7327
rect 10082 7293 10100 7327
rect 10048 7284 10100 7293
rect 10416 7284 10468 7336
rect 12532 7284 12584 7336
rect 12808 7284 12860 7336
rect 13820 7284 13872 7336
rect 16212 7327 16264 7336
rect 10968 7216 11020 7268
rect 12992 7259 13044 7268
rect 8208 7148 8260 7200
rect 12992 7225 13001 7259
rect 13001 7225 13035 7259
rect 13035 7225 13044 7259
rect 12992 7216 13044 7225
rect 13360 7216 13412 7268
rect 16212 7293 16241 7327
rect 16241 7293 16264 7327
rect 18972 7352 19024 7404
rect 20076 7352 20128 7404
rect 16212 7284 16264 7293
rect 18880 7284 18932 7336
rect 19156 7327 19208 7336
rect 19156 7293 19165 7327
rect 19165 7293 19199 7327
rect 19199 7293 19208 7327
rect 19156 7284 19208 7293
rect 17132 7216 17184 7268
rect 17316 7216 17368 7268
rect 13084 7191 13136 7200
rect 13084 7157 13093 7191
rect 13093 7157 13127 7191
rect 13127 7157 13136 7191
rect 13084 7148 13136 7157
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 14188 7148 14240 7200
rect 17592 7148 17644 7200
rect 19892 7191 19944 7200
rect 19892 7157 19901 7191
rect 19901 7157 19935 7191
rect 19935 7157 19944 7191
rect 19892 7148 19944 7157
rect 20260 7191 20312 7200
rect 20260 7157 20269 7191
rect 20269 7157 20303 7191
rect 20303 7157 20312 7191
rect 20260 7148 20312 7157
rect 20352 7191 20404 7200
rect 20352 7157 20361 7191
rect 20361 7157 20395 7191
rect 20395 7157 20404 7191
rect 20904 7191 20956 7200
rect 20352 7148 20404 7157
rect 20904 7157 20913 7191
rect 20913 7157 20947 7191
rect 20947 7157 20956 7191
rect 20904 7148 20956 7157
rect 7912 7046 7964 7098
rect 7976 7046 8028 7098
rect 8040 7046 8092 7098
rect 8104 7046 8156 7098
rect 14843 7046 14895 7098
rect 14907 7046 14959 7098
rect 14971 7046 15023 7098
rect 15035 7046 15087 7098
rect 9680 6944 9732 6996
rect 10324 6944 10376 6996
rect 11336 6944 11388 6996
rect 11520 6987 11572 6996
rect 11520 6953 11529 6987
rect 11529 6953 11563 6987
rect 11563 6953 11572 6987
rect 11520 6944 11572 6953
rect 11796 6944 11848 6996
rect 12348 6944 12400 6996
rect 8300 6876 8352 6928
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 7656 6851 7708 6860
rect 7656 6817 7665 6851
rect 7665 6817 7699 6851
rect 7699 6817 7708 6851
rect 7656 6808 7708 6817
rect 8116 6851 8168 6860
rect 8116 6817 8125 6851
rect 8125 6817 8159 6851
rect 8159 6817 8168 6851
rect 8116 6808 8168 6817
rect 12440 6876 12492 6928
rect 13176 6876 13228 6928
rect 13544 6944 13596 6996
rect 16396 6987 16448 6996
rect 16396 6953 16405 6987
rect 16405 6953 16439 6987
rect 16439 6953 16448 6987
rect 16396 6944 16448 6953
rect 16488 6944 16540 6996
rect 16120 6876 16172 6928
rect 20904 6944 20956 6996
rect 12624 6851 12676 6860
rect 12624 6817 12642 6851
rect 12642 6817 12676 6851
rect 12624 6808 12676 6817
rect 12808 6808 12860 6860
rect 13820 6808 13872 6860
rect 14740 6808 14792 6860
rect 15200 6808 15252 6860
rect 16212 6808 16264 6860
rect 17500 6851 17552 6860
rect 9036 6740 9088 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10324 6740 10376 6792
rect 10508 6740 10560 6792
rect 10876 6740 10928 6792
rect 13912 6783 13964 6792
rect 13912 6749 13921 6783
rect 13921 6749 13955 6783
rect 13955 6749 13964 6783
rect 13912 6740 13964 6749
rect 14096 6740 14148 6792
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 19064 6876 19116 6928
rect 20076 6919 20128 6928
rect 20076 6885 20110 6919
rect 20110 6885 20128 6919
rect 20076 6876 20128 6885
rect 8760 6672 8812 6724
rect 10692 6672 10744 6724
rect 10784 6672 10836 6724
rect 12900 6672 12952 6724
rect 6276 6647 6328 6656
rect 6276 6613 6285 6647
rect 6285 6613 6319 6647
rect 6319 6613 6328 6647
rect 6276 6604 6328 6613
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 9404 6604 9456 6656
rect 10508 6647 10560 6656
rect 10508 6613 10517 6647
rect 10517 6613 10551 6647
rect 10551 6613 10560 6647
rect 10508 6604 10560 6613
rect 11152 6604 11204 6656
rect 13360 6672 13412 6724
rect 16028 6715 16080 6724
rect 16028 6681 16037 6715
rect 16037 6681 16071 6715
rect 16071 6681 16080 6715
rect 16028 6672 16080 6681
rect 17316 6740 17368 6792
rect 18788 6783 18840 6792
rect 18788 6749 18797 6783
rect 18797 6749 18831 6783
rect 18831 6749 18840 6783
rect 18788 6740 18840 6749
rect 18880 6740 18932 6792
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 13452 6604 13504 6656
rect 17776 6604 17828 6656
rect 17960 6604 18012 6656
rect 19984 6604 20036 6656
rect 20536 6604 20588 6656
rect 4447 6502 4499 6554
rect 4511 6502 4563 6554
rect 4575 6502 4627 6554
rect 4639 6502 4691 6554
rect 11378 6502 11430 6554
rect 11442 6502 11494 6554
rect 11506 6502 11558 6554
rect 11570 6502 11622 6554
rect 18308 6502 18360 6554
rect 18372 6502 18424 6554
rect 18436 6502 18488 6554
rect 18500 6502 18552 6554
rect 6920 6332 6972 6384
rect 7288 6375 7340 6384
rect 7288 6341 7297 6375
rect 7297 6341 7331 6375
rect 7331 6341 7340 6375
rect 9588 6400 9640 6452
rect 7288 6332 7340 6341
rect 8852 6332 8904 6384
rect 13360 6400 13412 6452
rect 12992 6332 13044 6384
rect 13176 6332 13228 6384
rect 7564 6264 7616 6316
rect 2228 6196 2280 6248
rect 7380 6196 7432 6248
rect 10876 6307 10928 6316
rect 10876 6273 10885 6307
rect 10885 6273 10919 6307
rect 10919 6273 10928 6307
rect 10876 6264 10928 6273
rect 13452 6264 13504 6316
rect 5816 6128 5868 6180
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 6276 6060 6328 6112
rect 6920 6060 6972 6112
rect 7748 6128 7800 6180
rect 9404 6196 9456 6248
rect 13728 6196 13780 6248
rect 14372 6196 14424 6248
rect 14832 6400 14884 6452
rect 19708 6400 19760 6452
rect 20076 6400 20128 6452
rect 20260 6400 20312 6452
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 15936 6264 15988 6316
rect 16304 6264 16356 6316
rect 20076 6264 20128 6316
rect 9588 6128 9640 6180
rect 9864 6128 9916 6180
rect 10692 6171 10744 6180
rect 10692 6137 10701 6171
rect 10701 6137 10735 6171
rect 10735 6137 10744 6171
rect 10692 6128 10744 6137
rect 12348 6128 12400 6180
rect 8852 6060 8904 6112
rect 9036 6103 9088 6112
rect 9036 6069 9045 6103
rect 9045 6069 9079 6103
rect 9079 6069 9088 6103
rect 9036 6060 9088 6069
rect 10048 6060 10100 6112
rect 10784 6103 10836 6112
rect 10784 6069 10793 6103
rect 10793 6069 10827 6103
rect 10827 6069 10836 6103
rect 10784 6060 10836 6069
rect 12624 6060 12676 6112
rect 13176 6060 13228 6112
rect 13912 6128 13964 6180
rect 14556 6128 14608 6180
rect 18880 6196 18932 6248
rect 17408 6128 17460 6180
rect 15476 6103 15528 6112
rect 15476 6069 15485 6103
rect 15485 6069 15519 6103
rect 15519 6069 15528 6103
rect 15476 6060 15528 6069
rect 16212 6060 16264 6112
rect 16396 6103 16448 6112
rect 16396 6069 16405 6103
rect 16405 6069 16439 6103
rect 16439 6069 16448 6103
rect 16396 6060 16448 6069
rect 18788 6128 18840 6180
rect 20996 6239 21048 6248
rect 20996 6205 21005 6239
rect 21005 6205 21039 6239
rect 21039 6205 21048 6239
rect 20996 6196 21048 6205
rect 21088 6103 21140 6112
rect 21088 6069 21097 6103
rect 21097 6069 21131 6103
rect 21131 6069 21140 6103
rect 21088 6060 21140 6069
rect 7912 5958 7964 6010
rect 7976 5958 8028 6010
rect 8040 5958 8092 6010
rect 8104 5958 8156 6010
rect 14843 5958 14895 6010
rect 14907 5958 14959 6010
rect 14971 5958 15023 6010
rect 15035 5958 15087 6010
rect 5816 5899 5868 5908
rect 5816 5865 5825 5899
rect 5825 5865 5859 5899
rect 5859 5865 5868 5899
rect 5816 5856 5868 5865
rect 7748 5856 7800 5908
rect 8760 5899 8812 5908
rect 8760 5865 8769 5899
rect 8769 5865 8803 5899
rect 8803 5865 8812 5899
rect 8760 5856 8812 5865
rect 9772 5856 9824 5908
rect 10508 5856 10560 5908
rect 10692 5856 10744 5908
rect 8392 5788 8444 5840
rect 10048 5831 10100 5840
rect 10048 5797 10057 5831
rect 10057 5797 10091 5831
rect 10091 5797 10100 5831
rect 10048 5788 10100 5797
rect 11796 5831 11848 5840
rect 11796 5797 11814 5831
rect 11814 5797 11848 5831
rect 12624 5856 12676 5908
rect 12808 5856 12860 5908
rect 12992 5856 13044 5908
rect 13084 5856 13136 5908
rect 13636 5856 13688 5908
rect 13728 5856 13780 5908
rect 11796 5788 11848 5797
rect 15476 5788 15528 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 7564 5720 7616 5772
rect 7748 5720 7800 5772
rect 8208 5720 8260 5772
rect 9036 5652 9088 5704
rect 10692 5652 10744 5704
rect 6092 5516 6144 5568
rect 7472 5516 7524 5568
rect 10140 5516 10192 5568
rect 10692 5559 10744 5568
rect 10692 5525 10701 5559
rect 10701 5525 10735 5559
rect 10735 5525 10744 5559
rect 10692 5516 10744 5525
rect 12624 5720 12676 5772
rect 12532 5652 12584 5704
rect 12072 5584 12124 5636
rect 12440 5627 12492 5636
rect 12440 5593 12449 5627
rect 12449 5593 12483 5627
rect 12483 5593 12492 5627
rect 13268 5720 13320 5772
rect 14740 5720 14792 5772
rect 15200 5720 15252 5772
rect 15568 5763 15620 5772
rect 13176 5652 13228 5704
rect 15292 5695 15344 5704
rect 15292 5661 15301 5695
rect 15301 5661 15335 5695
rect 15335 5661 15344 5695
rect 15292 5652 15344 5661
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 17868 5856 17920 5908
rect 20352 5856 20404 5908
rect 16212 5788 16264 5840
rect 19800 5788 19852 5840
rect 20076 5788 20128 5840
rect 20628 5788 20680 5840
rect 16488 5652 16540 5704
rect 18880 5652 18932 5704
rect 12440 5584 12492 5593
rect 14188 5584 14240 5636
rect 14740 5559 14792 5568
rect 14740 5525 14749 5559
rect 14749 5525 14783 5559
rect 14783 5525 14792 5559
rect 14740 5516 14792 5525
rect 16120 5584 16172 5636
rect 20996 5627 21048 5636
rect 20996 5593 21005 5627
rect 21005 5593 21039 5627
rect 21039 5593 21048 5627
rect 20996 5584 21048 5593
rect 18696 5516 18748 5568
rect 18972 5559 19024 5568
rect 18972 5525 18981 5559
rect 18981 5525 19015 5559
rect 19015 5525 19024 5559
rect 18972 5516 19024 5525
rect 4447 5414 4499 5466
rect 4511 5414 4563 5466
rect 4575 5414 4627 5466
rect 4639 5414 4691 5466
rect 11378 5414 11430 5466
rect 11442 5414 11494 5466
rect 11506 5414 11558 5466
rect 11570 5414 11622 5466
rect 18308 5414 18360 5466
rect 18372 5414 18424 5466
rect 18436 5414 18488 5466
rect 18500 5414 18552 5466
rect 5724 5312 5776 5364
rect 9220 5312 9272 5364
rect 10324 5355 10376 5364
rect 10324 5321 10333 5355
rect 10333 5321 10367 5355
rect 10367 5321 10376 5355
rect 10324 5312 10376 5321
rect 18604 5312 18656 5364
rect 5816 5244 5868 5296
rect 7564 5244 7616 5296
rect 8300 5244 8352 5296
rect 9036 5244 9088 5296
rect 9312 5244 9364 5296
rect 12808 5244 12860 5296
rect 8576 5108 8628 5160
rect 7288 5040 7340 5092
rect 9312 5108 9364 5160
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 10692 5176 10744 5228
rect 12532 5219 12584 5228
rect 12532 5185 12541 5219
rect 12541 5185 12575 5219
rect 12575 5185 12584 5219
rect 12532 5176 12584 5185
rect 17132 5244 17184 5296
rect 19800 5244 19852 5296
rect 16488 5176 16540 5228
rect 19892 5176 19944 5228
rect 20536 5176 20588 5228
rect 21180 5219 21232 5228
rect 21180 5185 21189 5219
rect 21189 5185 21223 5219
rect 21223 5185 21232 5219
rect 21180 5176 21232 5185
rect 11704 5108 11756 5160
rect 11888 5108 11940 5160
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 14372 5108 14424 5160
rect 14648 5108 14700 5160
rect 8576 4972 8628 5024
rect 11152 5040 11204 5092
rect 11428 5040 11480 5092
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 11244 4972 11296 5024
rect 11704 4972 11756 5024
rect 12072 4972 12124 5024
rect 13452 5040 13504 5092
rect 12624 4972 12676 5024
rect 13084 4972 13136 5024
rect 15292 5108 15344 5160
rect 19984 5151 20036 5160
rect 19984 5117 19993 5151
rect 19993 5117 20027 5151
rect 20027 5117 20036 5151
rect 19984 5108 20036 5117
rect 17592 5083 17644 5092
rect 17592 5049 17601 5083
rect 17601 5049 17635 5083
rect 17635 5049 17644 5083
rect 17592 5040 17644 5049
rect 19248 5040 19300 5092
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 19064 4972 19116 5024
rect 20628 5015 20680 5024
rect 20628 4981 20637 5015
rect 20637 4981 20671 5015
rect 20671 4981 20680 5015
rect 20628 4972 20680 4981
rect 21088 5015 21140 5024
rect 21088 4981 21097 5015
rect 21097 4981 21131 5015
rect 21131 4981 21140 5015
rect 21088 4972 21140 4981
rect 7912 4870 7964 4922
rect 7976 4870 8028 4922
rect 8040 4870 8092 4922
rect 8104 4870 8156 4922
rect 14843 4870 14895 4922
rect 14907 4870 14959 4922
rect 14971 4870 15023 4922
rect 15035 4870 15087 4922
rect 6184 4811 6236 4820
rect 6184 4777 6193 4811
rect 6193 4777 6227 4811
rect 6227 4777 6236 4811
rect 6184 4768 6236 4777
rect 6920 4768 6972 4820
rect 8300 4768 8352 4820
rect 8576 4768 8628 4820
rect 9312 4768 9364 4820
rect 7564 4700 7616 4752
rect 8392 4700 8444 4752
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 6920 4564 6972 4616
rect 9864 4632 9916 4684
rect 10600 4632 10652 4684
rect 14372 4700 14424 4752
rect 14648 4700 14700 4752
rect 14740 4700 14792 4752
rect 16488 4700 16540 4752
rect 17408 4768 17460 4820
rect 18144 4768 18196 4820
rect 18880 4768 18932 4820
rect 21180 4811 21232 4820
rect 21180 4777 21189 4811
rect 21189 4777 21223 4811
rect 21223 4777 21232 4811
rect 21180 4768 21232 4777
rect 17776 4743 17828 4752
rect 17776 4709 17785 4743
rect 17785 4709 17819 4743
rect 17819 4709 17828 4743
rect 17776 4700 17828 4709
rect 22100 4700 22152 4752
rect 12440 4632 12492 4684
rect 13912 4675 13964 4684
rect 13912 4641 13921 4675
rect 13921 4641 13955 4675
rect 13955 4641 13964 4675
rect 13912 4632 13964 4641
rect 18512 4675 18564 4684
rect 11428 4607 11480 4616
rect 8852 4496 8904 4548
rect 9404 4496 9456 4548
rect 7656 4471 7708 4480
rect 7656 4437 7665 4471
rect 7665 4437 7699 4471
rect 7699 4437 7708 4471
rect 7656 4428 7708 4437
rect 8300 4428 8352 4480
rect 8944 4428 8996 4480
rect 9680 4428 9732 4480
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 18512 4641 18521 4675
rect 18521 4641 18555 4675
rect 18555 4641 18564 4675
rect 18512 4632 18564 4641
rect 18788 4632 18840 4684
rect 20076 4675 20128 4684
rect 20076 4641 20110 4675
rect 20110 4641 20128 4675
rect 20076 4632 20128 4641
rect 15936 4607 15988 4616
rect 11152 4539 11204 4548
rect 11152 4505 11161 4539
rect 11161 4505 11195 4539
rect 11195 4505 11204 4539
rect 11152 4496 11204 4505
rect 10968 4428 11020 4480
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 18144 4564 18196 4616
rect 18880 4564 18932 4616
rect 13176 4539 13228 4548
rect 13176 4505 13185 4539
rect 13185 4505 13219 4539
rect 13219 4505 13228 4539
rect 13176 4496 13228 4505
rect 13728 4539 13780 4548
rect 13728 4505 13737 4539
rect 13737 4505 13771 4539
rect 13771 4505 13780 4539
rect 13728 4496 13780 4505
rect 14740 4496 14792 4548
rect 15384 4539 15436 4548
rect 15384 4505 15393 4539
rect 15393 4505 15427 4539
rect 15427 4505 15436 4539
rect 15384 4496 15436 4505
rect 17040 4496 17092 4548
rect 13452 4428 13504 4480
rect 19156 4564 19208 4616
rect 21548 4428 21600 4480
rect 4447 4326 4499 4378
rect 4511 4326 4563 4378
rect 4575 4326 4627 4378
rect 4639 4326 4691 4378
rect 11378 4326 11430 4378
rect 11442 4326 11494 4378
rect 11506 4326 11558 4378
rect 11570 4326 11622 4378
rect 18308 4326 18360 4378
rect 18372 4326 18424 4378
rect 18436 4326 18488 4378
rect 18500 4326 18552 4378
rect 5724 4267 5776 4276
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 9496 4267 9548 4276
rect 9496 4233 9505 4267
rect 9505 4233 9539 4267
rect 9539 4233 9548 4267
rect 9496 4224 9548 4233
rect 10600 4224 10652 4276
rect 18696 4224 18748 4276
rect 21088 4224 21140 4276
rect 8300 4156 8352 4208
rect 9680 4156 9732 4208
rect 10048 4156 10100 4208
rect 10508 4156 10560 4208
rect 6552 4131 6604 4140
rect 6552 4097 6561 4131
rect 6561 4097 6595 4131
rect 6595 4097 6604 4131
rect 6552 4088 6604 4097
rect 10324 4088 10376 4140
rect 11152 4156 11204 4208
rect 12348 4131 12400 4140
rect 8024 4020 8076 4072
rect 8300 4063 8352 4072
rect 8300 4029 8309 4063
rect 8309 4029 8343 4063
rect 8343 4029 8352 4063
rect 8300 4020 8352 4029
rect 4160 3952 4212 4004
rect 9956 4020 10008 4072
rect 10140 4063 10192 4072
rect 10140 4029 10149 4063
rect 10149 4029 10183 4063
rect 10183 4029 10192 4063
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 14556 4131 14608 4140
rect 14556 4097 14565 4131
rect 14565 4097 14599 4131
rect 14599 4097 14608 4131
rect 14556 4088 14608 4097
rect 16212 4131 16264 4140
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 17408 4156 17460 4208
rect 17500 4156 17552 4208
rect 18144 4156 18196 4208
rect 16488 4088 16540 4140
rect 20076 4131 20128 4140
rect 20076 4097 20085 4131
rect 20085 4097 20119 4131
rect 20119 4097 20128 4131
rect 20076 4088 20128 4097
rect 10140 4020 10192 4029
rect 11704 4020 11756 4072
rect 13820 4020 13872 4072
rect 14280 4020 14332 4072
rect 17132 4020 17184 4072
rect 17224 4020 17276 4072
rect 21272 4063 21324 4072
rect 7288 3884 7340 3936
rect 8208 3884 8260 3936
rect 8300 3884 8352 3936
rect 8484 3927 8536 3936
rect 8484 3893 8493 3927
rect 8493 3893 8527 3927
rect 8527 3893 8536 3927
rect 8484 3884 8536 3893
rect 8944 3927 8996 3936
rect 8944 3893 8953 3927
rect 8953 3893 8987 3927
rect 8987 3893 8996 3927
rect 8944 3884 8996 3893
rect 9772 3884 9824 3936
rect 10140 3884 10192 3936
rect 10784 3884 10836 3936
rect 11980 3952 12032 4004
rect 14648 3995 14700 4004
rect 14648 3961 14657 3995
rect 14657 3961 14691 3995
rect 14691 3961 14700 3995
rect 14648 3952 14700 3961
rect 15200 3995 15252 4004
rect 15200 3961 15209 3995
rect 15209 3961 15243 3995
rect 15243 3961 15252 3995
rect 15200 3952 15252 3961
rect 15292 3952 15344 4004
rect 17592 3952 17644 4004
rect 12072 3884 12124 3936
rect 12256 3927 12308 3936
rect 12256 3893 12265 3927
rect 12265 3893 12299 3927
rect 12299 3893 12308 3927
rect 12256 3884 12308 3893
rect 14004 3884 14056 3936
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 16028 3884 16080 3936
rect 21272 4029 21281 4063
rect 21281 4029 21315 4063
rect 21315 4029 21324 4063
rect 21272 4020 21324 4029
rect 18880 3952 18932 4004
rect 20352 3927 20404 3936
rect 20352 3893 20361 3927
rect 20361 3893 20395 3927
rect 20395 3893 20404 3927
rect 20352 3884 20404 3893
rect 7912 3782 7964 3834
rect 7976 3782 8028 3834
rect 8040 3782 8092 3834
rect 8104 3782 8156 3834
rect 14843 3782 14895 3834
rect 14907 3782 14959 3834
rect 14971 3782 15023 3834
rect 15035 3782 15087 3834
rect 7012 3680 7064 3732
rect 7288 3680 7340 3732
rect 7196 3612 7248 3664
rect 10968 3680 11020 3732
rect 11244 3680 11296 3732
rect 11704 3680 11756 3732
rect 14004 3723 14056 3732
rect 14004 3689 14013 3723
rect 14013 3689 14047 3723
rect 14047 3689 14056 3723
rect 14004 3680 14056 3689
rect 15752 3680 15804 3732
rect 15844 3680 15896 3732
rect 16580 3680 16632 3732
rect 18604 3680 18656 3732
rect 18880 3723 18932 3732
rect 18880 3689 18889 3723
rect 18889 3689 18923 3723
rect 18923 3689 18932 3723
rect 18880 3680 18932 3689
rect 19156 3680 19208 3732
rect 20628 3680 20680 3732
rect 7748 3544 7800 3596
rect 7932 3544 7984 3596
rect 14648 3612 14700 3664
rect 8852 3587 8904 3596
rect 8852 3553 8861 3587
rect 8861 3553 8895 3587
rect 8895 3553 8904 3587
rect 8852 3544 8904 3553
rect 9036 3544 9088 3596
rect 10508 3544 10560 3596
rect 10692 3587 10744 3596
rect 10692 3553 10701 3587
rect 10701 3553 10735 3587
rect 10735 3553 10744 3587
rect 10692 3544 10744 3553
rect 5264 3476 5316 3528
rect 7840 3476 7892 3528
rect 10048 3476 10100 3528
rect 10600 3476 10652 3528
rect 12440 3544 12492 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 11152 3476 11204 3528
rect 11612 3476 11664 3528
rect 12348 3476 12400 3528
rect 14372 3544 14424 3596
rect 13268 3476 13320 3528
rect 14096 3476 14148 3528
rect 1308 3408 1360 3460
rect 6552 3408 6604 3460
rect 8116 3408 8168 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 5816 3340 5868 3392
rect 7104 3340 7156 3392
rect 7288 3383 7340 3392
rect 7288 3349 7297 3383
rect 7297 3349 7331 3383
rect 7331 3349 7340 3383
rect 7288 3340 7340 3349
rect 7564 3340 7616 3392
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8024 3340 8076 3392
rect 8392 3340 8444 3392
rect 9404 3408 9456 3460
rect 12624 3451 12676 3460
rect 10048 3340 10100 3392
rect 11796 3340 11848 3392
rect 11980 3340 12032 3392
rect 12624 3417 12633 3451
rect 12633 3417 12667 3451
rect 12667 3417 12676 3451
rect 12624 3408 12676 3417
rect 20444 3612 20496 3664
rect 16396 3544 16448 3596
rect 17592 3544 17644 3596
rect 18144 3544 18196 3596
rect 18696 3544 18748 3596
rect 20904 3612 20956 3664
rect 20720 3587 20772 3596
rect 20720 3553 20729 3587
rect 20729 3553 20763 3587
rect 20763 3553 20772 3587
rect 20720 3544 20772 3553
rect 16580 3476 16632 3528
rect 16948 3519 17000 3528
rect 16948 3485 16957 3519
rect 16957 3485 16991 3519
rect 16991 3485 17000 3519
rect 16948 3476 17000 3485
rect 17132 3476 17184 3528
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 16304 3383 16356 3392
rect 16304 3349 16313 3383
rect 16313 3349 16347 3383
rect 16347 3349 16356 3383
rect 16304 3340 16356 3349
rect 17316 3340 17368 3392
rect 19340 3408 19392 3460
rect 19156 3383 19208 3392
rect 19156 3349 19165 3383
rect 19165 3349 19199 3383
rect 19199 3349 19208 3383
rect 19156 3340 19208 3349
rect 19248 3340 19300 3392
rect 20812 3340 20864 3392
rect 21180 3383 21232 3392
rect 21180 3349 21189 3383
rect 21189 3349 21223 3383
rect 21223 3349 21232 3383
rect 21180 3340 21232 3349
rect 4447 3238 4499 3290
rect 4511 3238 4563 3290
rect 4575 3238 4627 3290
rect 4639 3238 4691 3290
rect 11378 3238 11430 3290
rect 11442 3238 11494 3290
rect 11506 3238 11558 3290
rect 11570 3238 11622 3290
rect 18308 3238 18360 3290
rect 18372 3238 18424 3290
rect 18436 3238 18488 3290
rect 18500 3238 18552 3290
rect 9312 3136 9364 3188
rect 9772 3136 9824 3188
rect 12808 3136 12860 3188
rect 13268 3179 13320 3188
rect 13268 3145 13277 3179
rect 13277 3145 13311 3179
rect 13311 3145 13320 3179
rect 13268 3136 13320 3145
rect 14188 3136 14240 3188
rect 4436 3111 4488 3120
rect 4436 3077 4445 3111
rect 4445 3077 4479 3111
rect 4479 3077 4488 3111
rect 4436 3068 4488 3077
rect 10508 3068 10560 3120
rect 6920 3000 6972 3052
rect 7104 3000 7156 3052
rect 7840 3043 7892 3052
rect 848 2932 900 2984
rect 1308 2932 1360 2984
rect 1492 2932 1544 2984
rect 1952 2932 2004 2984
rect 4712 2975 4764 2984
rect 4712 2941 4721 2975
rect 4721 2941 4755 2975
rect 4755 2941 4764 2975
rect 4712 2932 4764 2941
rect 7012 2975 7064 2984
rect 7012 2941 7021 2975
rect 7021 2941 7055 2975
rect 7055 2941 7064 2975
rect 7012 2932 7064 2941
rect 7288 2932 7340 2984
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8116 3000 8168 3052
rect 7932 2975 7984 2984
rect 2504 2864 2556 2916
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 8024 2932 8076 2984
rect 8484 2932 8536 2984
rect 8760 2932 8812 2984
rect 8944 3000 8996 3052
rect 9312 2975 9364 2984
rect 9312 2941 9321 2975
rect 9321 2941 9355 2975
rect 9355 2941 9364 2975
rect 9312 2932 9364 2941
rect 10140 3000 10192 3052
rect 10048 2932 10100 2984
rect 14648 3136 14700 3188
rect 16948 3068 17000 3120
rect 18144 3136 18196 3188
rect 21180 3136 21232 3188
rect 11704 2932 11756 2984
rect 9220 2864 9272 2916
rect 13084 2932 13136 2984
rect 15108 3000 15160 3052
rect 16672 3000 16724 3052
rect 14372 2932 14424 2984
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 3148 2796 3200 2848
rect 3608 2796 3660 2848
rect 4160 2796 4212 2848
rect 5172 2839 5224 2848
rect 5172 2805 5181 2839
rect 5181 2805 5215 2839
rect 5215 2805 5224 2839
rect 5172 2796 5224 2805
rect 6460 2796 6512 2848
rect 7472 2796 7524 2848
rect 8484 2796 8536 2848
rect 8576 2839 8628 2848
rect 8576 2805 8585 2839
rect 8585 2805 8619 2839
rect 8619 2805 8628 2839
rect 9036 2839 9088 2848
rect 8576 2796 8628 2805
rect 9036 2805 9045 2839
rect 9045 2805 9079 2839
rect 9079 2805 9088 2839
rect 9036 2796 9088 2805
rect 9588 2796 9640 2848
rect 10692 2796 10744 2848
rect 11704 2796 11756 2848
rect 12256 2864 12308 2916
rect 13912 2864 13964 2916
rect 15936 2932 15988 2984
rect 17132 2975 17184 2984
rect 17132 2941 17141 2975
rect 17141 2941 17175 2975
rect 17175 2941 17184 2975
rect 17132 2932 17184 2941
rect 18512 3000 18564 3052
rect 18880 3000 18932 3052
rect 20812 3000 20864 3052
rect 19064 2932 19116 2984
rect 19248 2975 19300 2984
rect 19248 2941 19257 2975
rect 19257 2941 19291 2975
rect 19291 2941 19300 2975
rect 19248 2932 19300 2941
rect 20628 2932 20680 2984
rect 21364 3068 21416 3120
rect 19800 2907 19852 2916
rect 19800 2873 19809 2907
rect 19809 2873 19843 2907
rect 19843 2873 19852 2907
rect 19800 2864 19852 2873
rect 18788 2839 18840 2848
rect 18788 2805 18797 2839
rect 18797 2805 18831 2839
rect 18831 2805 18840 2839
rect 18788 2796 18840 2805
rect 19708 2796 19760 2848
rect 7912 2694 7964 2746
rect 7976 2694 8028 2746
rect 8040 2694 8092 2746
rect 8104 2694 8156 2746
rect 14843 2694 14895 2746
rect 14907 2694 14959 2746
rect 14971 2694 15023 2746
rect 15035 2694 15087 2746
rect 4068 2592 4120 2644
rect 4252 2635 4304 2644
rect 4252 2601 4261 2635
rect 4261 2601 4295 2635
rect 4295 2601 4304 2635
rect 4252 2592 4304 2601
rect 4804 2635 4856 2644
rect 4804 2601 4813 2635
rect 4813 2601 4847 2635
rect 4847 2601 4856 2635
rect 4804 2592 4856 2601
rect 8668 2592 8720 2644
rect 9956 2592 10008 2644
rect 11152 2635 11204 2644
rect 11152 2601 11161 2635
rect 11161 2601 11195 2635
rect 11195 2601 11204 2635
rect 11152 2592 11204 2601
rect 2228 2567 2280 2576
rect 2228 2533 2237 2567
rect 2237 2533 2271 2567
rect 2271 2533 2280 2567
rect 2228 2524 2280 2533
rect 4160 2567 4212 2576
rect 4160 2533 4169 2567
rect 4169 2533 4203 2567
rect 4203 2533 4212 2567
rect 4160 2524 4212 2533
rect 6368 2524 6420 2576
rect 7380 2524 7432 2576
rect 9128 2524 9180 2576
rect 296 2456 348 2508
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1952 2456 2004 2508
rect 2504 2499 2556 2508
rect 2504 2465 2513 2499
rect 2513 2465 2547 2499
rect 2547 2465 2556 2499
rect 2504 2456 2556 2465
rect 3056 2456 3108 2508
rect 5172 2456 5224 2508
rect 5264 2456 5316 2508
rect 5816 2456 5868 2508
rect 6460 2456 6512 2508
rect 7656 2456 7708 2508
rect 8208 2499 8260 2508
rect 8208 2465 8217 2499
rect 8217 2465 8251 2499
rect 8251 2465 8260 2499
rect 8208 2456 8260 2465
rect 8944 2456 8996 2508
rect 4160 2388 4212 2440
rect 10140 2524 10192 2576
rect 10416 2524 10468 2576
rect 11704 2524 11756 2576
rect 14556 2592 14608 2644
rect 15844 2592 15896 2644
rect 16580 2592 16632 2644
rect 18512 2592 18564 2644
rect 18604 2592 18656 2644
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 9772 2456 9824 2508
rect 10324 2456 10376 2508
rect 10600 2499 10652 2508
rect 10600 2465 10609 2499
rect 10609 2465 10643 2499
rect 10643 2465 10652 2499
rect 10600 2456 10652 2465
rect 10876 2456 10928 2508
rect 17592 2524 17644 2576
rect 2688 2295 2740 2304
rect 2688 2261 2697 2295
rect 2697 2261 2731 2295
rect 2731 2261 2740 2295
rect 2688 2252 2740 2261
rect 8484 2320 8536 2372
rect 12072 2363 12124 2372
rect 12072 2329 12081 2363
rect 12081 2329 12115 2363
rect 12115 2329 12124 2363
rect 12072 2320 12124 2329
rect 12256 2388 12308 2440
rect 12716 2320 12768 2372
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 16120 2499 16172 2508
rect 16120 2465 16129 2499
rect 16129 2465 16163 2499
rect 16163 2465 16172 2499
rect 16120 2456 16172 2465
rect 18144 2524 18196 2576
rect 18972 2524 19024 2576
rect 19064 2524 19116 2576
rect 17960 2499 18012 2508
rect 17960 2465 17969 2499
rect 17969 2465 18003 2499
rect 18003 2465 18012 2499
rect 17960 2456 18012 2465
rect 19524 2456 19576 2508
rect 17868 2431 17920 2440
rect 17868 2397 17877 2431
rect 17877 2397 17911 2431
rect 17911 2397 17920 2431
rect 17868 2388 17920 2397
rect 8300 2252 8352 2304
rect 8852 2295 8904 2304
rect 8852 2261 8861 2295
rect 8861 2261 8895 2295
rect 8895 2261 8904 2295
rect 8852 2252 8904 2261
rect 10784 2252 10836 2304
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 13544 2295 13596 2304
rect 12992 2252 13044 2261
rect 13544 2261 13553 2295
rect 13553 2261 13587 2295
rect 13587 2261 13596 2295
rect 13544 2252 13596 2261
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 17776 2320 17828 2372
rect 19156 2320 19208 2372
rect 18144 2252 18196 2304
rect 19248 2252 19300 2304
rect 19432 2320 19484 2372
rect 21088 2363 21140 2372
rect 21088 2329 21097 2363
rect 21097 2329 21131 2363
rect 21131 2329 21140 2363
rect 21088 2320 21140 2329
rect 4447 2150 4499 2202
rect 4511 2150 4563 2202
rect 4575 2150 4627 2202
rect 4639 2150 4691 2202
rect 11378 2150 11430 2202
rect 11442 2150 11494 2202
rect 11506 2150 11558 2202
rect 11570 2150 11622 2202
rect 18308 2150 18360 2202
rect 18372 2150 18424 2202
rect 18436 2150 18488 2202
rect 18500 2150 18552 2202
rect 9036 2048 9088 2100
rect 12256 2048 12308 2100
rect 14096 2048 14148 2100
rect 19892 2048 19944 2100
rect 2044 1980 2096 2032
rect 17960 1980 18012 2032
rect 8668 1912 8720 1964
rect 9496 1912 9548 1964
rect 9864 1912 9916 1964
rect 11428 1912 11480 1964
rect 16764 1912 16816 1964
rect 21088 1912 21140 1964
rect 2688 1844 2740 1896
rect 16120 1844 16172 1896
rect 13544 1776 13596 1828
rect 20444 1776 20496 1828
rect 6184 1708 6236 1760
rect 17868 1708 17920 1760
rect 8852 1640 8904 1692
rect 16856 1640 16908 1692
rect 8944 1572 8996 1624
rect 18052 1572 18104 1624
rect 12992 1504 13044 1556
rect 22652 1504 22704 1556
rect 21916 1436 21968 1488
rect 22008 1411 22060 1420
rect 22008 1377 22017 1411
rect 22017 1377 22051 1411
rect 22051 1377 22060 1411
rect 22008 1368 22060 1377
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 15382 22200 15438 23000
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 17958 22264 18014 22273
rect 308 19310 336 22200
rect 860 20602 888 22200
rect 848 20596 900 20602
rect 848 20538 900 20544
rect 1412 19990 1440 22200
rect 1964 20330 1992 22200
rect 1952 20324 2004 20330
rect 1952 20266 2004 20272
rect 1964 20074 1992 20266
rect 1964 20046 2084 20074
rect 1400 19984 1452 19990
rect 1400 19926 1452 19932
rect 1952 19984 2004 19990
rect 1952 19926 2004 19932
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1688 19310 1716 19858
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 296 19304 348 19310
rect 296 19246 348 19252
rect 1676 19304 1728 19310
rect 1676 19246 1728 19252
rect 1584 17264 1636 17270
rect 1582 17232 1584 17241
rect 1636 17232 1638 17241
rect 1582 17167 1638 17176
rect 1780 10810 1808 19654
rect 1964 19514 1992 19926
rect 2056 19854 2084 20046
rect 2320 20052 2372 20058
rect 2320 19994 2372 20000
rect 2332 19961 2360 19994
rect 2318 19952 2374 19961
rect 2516 19922 2544 22200
rect 3068 20398 3096 22200
rect 3620 20398 3648 22200
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 3608 20392 3660 20398
rect 3608 20334 3660 20340
rect 2688 20256 2740 20262
rect 2688 20198 2740 20204
rect 2318 19887 2374 19896
rect 2504 19916 2556 19922
rect 2504 19858 2556 19864
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 2516 19514 2544 19858
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2240 12238 2268 16934
rect 2700 14550 2728 20198
rect 3068 20058 3096 20334
rect 3620 20058 3648 20334
rect 4172 20262 4200 22200
rect 4724 20890 4752 22200
rect 4724 20862 4844 20890
rect 4421 20700 4717 20720
rect 4477 20698 4501 20700
rect 4557 20698 4581 20700
rect 4637 20698 4661 20700
rect 4499 20646 4501 20698
rect 4563 20646 4575 20698
rect 4637 20646 4639 20698
rect 4477 20644 4501 20646
rect 4557 20644 4581 20646
rect 4637 20644 4661 20646
rect 4421 20624 4717 20644
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 4172 20058 4200 20198
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3608 20052 3660 20058
rect 3608 19994 3660 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4816 19922 4844 20862
rect 5080 20596 5132 20602
rect 5080 20538 5132 20544
rect 4896 20324 4948 20330
rect 4896 20266 4948 20272
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 2778 19816 2834 19825
rect 2778 19751 2780 19760
rect 2832 19751 2834 19760
rect 2780 19722 2832 19728
rect 4421 19612 4717 19632
rect 4477 19610 4501 19612
rect 4557 19610 4581 19612
rect 4637 19610 4661 19612
rect 4499 19558 4501 19610
rect 4563 19558 4575 19610
rect 4637 19558 4639 19610
rect 4477 19556 4501 19558
rect 4557 19556 4581 19558
rect 4637 19556 4661 19558
rect 4421 19536 4717 19556
rect 4816 19514 4844 19858
rect 4804 19508 4856 19514
rect 4804 19450 4856 19456
rect 4421 18524 4717 18544
rect 4477 18522 4501 18524
rect 4557 18522 4581 18524
rect 4637 18522 4661 18524
rect 4499 18470 4501 18522
rect 4563 18470 4575 18522
rect 4637 18470 4639 18522
rect 4477 18468 4501 18470
rect 4557 18468 4581 18470
rect 4637 18468 4661 18470
rect 4421 18448 4717 18468
rect 4908 17882 4936 20266
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4421 17436 4717 17456
rect 4477 17434 4501 17436
rect 4557 17434 4581 17436
rect 4637 17434 4661 17436
rect 4499 17382 4501 17434
rect 4563 17382 4575 17434
rect 4637 17382 4639 17434
rect 4477 17380 4501 17382
rect 4557 17380 4581 17382
rect 4637 17380 4661 17382
rect 4421 17360 4717 17380
rect 4421 16348 4717 16368
rect 4477 16346 4501 16348
rect 4557 16346 4581 16348
rect 4637 16346 4661 16348
rect 4499 16294 4501 16346
rect 4563 16294 4575 16346
rect 4637 16294 4639 16346
rect 4477 16292 4501 16294
rect 4557 16292 4581 16294
rect 4637 16292 4661 16294
rect 4421 16272 4717 16292
rect 4421 15260 4717 15280
rect 4477 15258 4501 15260
rect 4557 15258 4581 15260
rect 4637 15258 4661 15260
rect 4499 15206 4501 15258
rect 4563 15206 4575 15258
rect 4637 15206 4639 15258
rect 4477 15204 4501 15206
rect 4557 15204 4581 15206
rect 4637 15204 4661 15206
rect 4421 15184 4717 15204
rect 2688 14544 2740 14550
rect 2688 14486 2740 14492
rect 4421 14172 4717 14192
rect 4477 14170 4501 14172
rect 4557 14170 4581 14172
rect 4637 14170 4661 14172
rect 4499 14118 4501 14170
rect 4563 14118 4575 14170
rect 4637 14118 4639 14170
rect 4477 14116 4501 14118
rect 4557 14116 4581 14118
rect 4637 14116 4661 14118
rect 4421 14096 4717 14116
rect 4421 13084 4717 13104
rect 4477 13082 4501 13084
rect 4557 13082 4581 13084
rect 4637 13082 4661 13084
rect 4499 13030 4501 13082
rect 4563 13030 4575 13082
rect 4637 13030 4639 13082
rect 4477 13028 4501 13030
rect 4557 13028 4581 13030
rect 4637 13028 4661 13030
rect 4421 13008 4717 13028
rect 5092 12918 5120 20538
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5184 14006 5212 20402
rect 5276 20398 5304 22200
rect 5828 20398 5856 22200
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5276 19310 5304 20334
rect 5264 19304 5316 19310
rect 5264 19246 5316 19252
rect 5828 18970 5856 20334
rect 5908 20256 5960 20262
rect 5908 20198 5960 20204
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5264 18692 5316 18698
rect 5264 18634 5316 18640
rect 5276 17513 5304 18634
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 18148 5500 18154
rect 5448 18090 5500 18096
rect 5262 17504 5318 17513
rect 5262 17439 5318 17448
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16046 5396 16934
rect 5460 16658 5488 18090
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5460 13938 5488 16594
rect 5552 15910 5580 18566
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5552 15434 5580 15846
rect 5540 15428 5592 15434
rect 5540 15370 5592 15376
rect 5552 14618 5580 15370
rect 5540 14612 5592 14618
rect 5540 14554 5592 14560
rect 5448 13932 5500 13938
rect 5448 13874 5500 13880
rect 5080 12912 5132 12918
rect 5080 12854 5132 12860
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 4421 11996 4717 12016
rect 4477 11994 4501 11996
rect 4557 11994 4581 11996
rect 4637 11994 4661 11996
rect 4499 11942 4501 11994
rect 4563 11942 4575 11994
rect 4637 11942 4639 11994
rect 4477 11940 4501 11942
rect 4557 11940 4581 11942
rect 4637 11940 4661 11942
rect 4421 11920 4717 11940
rect 5644 11014 5672 18022
rect 5816 17536 5868 17542
rect 5920 17524 5948 20198
rect 5868 17496 5948 17524
rect 5816 17478 5868 17484
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 5736 16794 5764 16934
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5722 16008 5778 16017
rect 5722 15943 5724 15952
rect 5776 15943 5778 15952
rect 5724 15914 5776 15920
rect 5736 15706 5764 15914
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 4804 11008 4856 11014
rect 4804 10950 4856 10956
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 4421 10908 4717 10928
rect 4477 10906 4501 10908
rect 4557 10906 4581 10908
rect 4637 10906 4661 10908
rect 4499 10854 4501 10906
rect 4563 10854 4575 10906
rect 4637 10854 4639 10906
rect 4477 10852 4501 10854
rect 4557 10852 4581 10854
rect 4637 10852 4661 10854
rect 4421 10832 4717 10852
rect 1768 10804 1820 10810
rect 1768 10746 1820 10752
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 2228 6248 2280 6254
rect 2228 6190 2280 6196
rect 1582 5808 1638 5817
rect 1582 5743 1584 5752
rect 1636 5743 1638 5752
rect 1584 5714 1636 5720
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1320 2990 1348 3402
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 848 2984 900 2990
rect 848 2926 900 2932
rect 1308 2984 1360 2990
rect 1308 2926 1360 2932
rect 296 2508 348 2514
rect 296 2450 348 2456
rect 308 800 336 2450
rect 860 800 888 2926
rect 1412 2514 1440 3334
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1504 2394 1532 2926
rect 1964 2514 1992 2926
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1952 2508 2004 2514
rect 1952 2450 2004 2456
rect 1412 2366 1532 2394
rect 1412 800 1440 2366
rect 1964 800 1992 2450
rect 2056 2038 2084 2790
rect 2240 2582 2268 6190
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 2938 4200 3946
rect 2504 2916 2556 2922
rect 2504 2858 2556 2864
rect 4080 2910 4200 2938
rect 2228 2576 2280 2582
rect 2228 2518 2280 2524
rect 2516 2514 2544 2858
rect 3148 2848 3200 2854
rect 3068 2796 3148 2802
rect 3068 2790 3200 2796
rect 3608 2848 3660 2854
rect 3608 2790 3660 2796
rect 3068 2774 3188 2790
rect 3068 2514 3096 2774
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 3056 2508 3108 2514
rect 3056 2450 3108 2456
rect 2044 2032 2096 2038
rect 2044 1974 2096 1980
rect 2516 800 2544 2450
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 2700 1902 2728 2246
rect 2688 1896 2740 1902
rect 2688 1838 2740 1844
rect 3068 800 3096 2450
rect 3620 800 3648 2790
rect 4080 2650 4108 2910
rect 4160 2848 4212 2854
rect 4160 2790 4212 2796
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4172 2582 4200 2790
rect 4264 2650 4292 10406
rect 4816 9926 4844 10950
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4421 9820 4717 9840
rect 4477 9818 4501 9820
rect 4557 9818 4581 9820
rect 4637 9818 4661 9820
rect 4499 9766 4501 9818
rect 4563 9766 4575 9818
rect 4637 9766 4639 9818
rect 4477 9764 4501 9766
rect 4557 9764 4581 9766
rect 4637 9764 4661 9766
rect 4421 9744 4717 9764
rect 4421 8732 4717 8752
rect 4477 8730 4501 8732
rect 4557 8730 4581 8732
rect 4637 8730 4661 8732
rect 4499 8678 4501 8730
rect 4563 8678 4575 8730
rect 4637 8678 4639 8730
rect 4477 8676 4501 8678
rect 4557 8676 4581 8678
rect 4637 8676 4661 8678
rect 4421 8656 4717 8676
rect 4421 7644 4717 7664
rect 4477 7642 4501 7644
rect 4557 7642 4581 7644
rect 4637 7642 4661 7644
rect 4499 7590 4501 7642
rect 4563 7590 4575 7642
rect 4637 7590 4639 7642
rect 4477 7588 4501 7590
rect 4557 7588 4581 7590
rect 4637 7588 4661 7590
rect 4421 7568 4717 7588
rect 4421 6556 4717 6576
rect 4477 6554 4501 6556
rect 4557 6554 4581 6556
rect 4637 6554 4661 6556
rect 4499 6502 4501 6554
rect 4563 6502 4575 6554
rect 4637 6502 4639 6554
rect 4477 6500 4501 6502
rect 4557 6500 4581 6502
rect 4637 6500 4661 6502
rect 4421 6480 4717 6500
rect 4421 5468 4717 5488
rect 4477 5466 4501 5468
rect 4557 5466 4581 5468
rect 4637 5466 4661 5468
rect 4499 5414 4501 5466
rect 4563 5414 4575 5466
rect 4637 5414 4639 5466
rect 4477 5412 4501 5414
rect 4557 5412 4581 5414
rect 4637 5412 4661 5414
rect 4421 5392 4717 5412
rect 4421 4380 4717 4400
rect 4477 4378 4501 4380
rect 4557 4378 4581 4380
rect 4637 4378 4661 4380
rect 4499 4326 4501 4378
rect 4563 4326 4575 4378
rect 4637 4326 4639 4378
rect 4477 4324 4501 4326
rect 4557 4324 4581 4326
rect 4637 4324 4661 4326
rect 4421 4304 4717 4324
rect 4421 3292 4717 3312
rect 4477 3290 4501 3292
rect 4557 3290 4581 3292
rect 4637 3290 4661 3292
rect 4499 3238 4501 3290
rect 4563 3238 4575 3290
rect 4637 3238 4639 3290
rect 4477 3236 4501 3238
rect 4557 3236 4581 3238
rect 4637 3236 4661 3238
rect 4421 3216 4717 3236
rect 4436 3120 4488 3126
rect 4434 3088 4436 3097
rect 4488 3088 4490 3097
rect 4434 3023 4490 3032
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4160 2576 4212 2582
rect 4160 2518 4212 2524
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4172 800 4200 2382
rect 4724 2292 4752 2926
rect 4816 2650 4844 9862
rect 5828 6186 5856 17478
rect 6012 16454 6040 20470
rect 6472 20398 6500 22200
rect 6920 20460 6972 20466
rect 6920 20402 6972 20408
rect 6460 20392 6512 20398
rect 6460 20334 6512 20340
rect 6092 19916 6144 19922
rect 6092 19858 6144 19864
rect 6104 18834 6132 19858
rect 6472 19514 6500 20334
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 6460 19508 6512 19514
rect 6460 19450 6512 19456
rect 6182 19272 6238 19281
rect 6564 19242 6592 19858
rect 6644 19848 6696 19854
rect 6828 19848 6880 19854
rect 6696 19808 6828 19836
rect 6644 19790 6696 19796
rect 6828 19790 6880 19796
rect 6644 19712 6696 19718
rect 6828 19712 6880 19718
rect 6644 19654 6696 19660
rect 6826 19680 6828 19689
rect 6880 19680 6882 19689
rect 6656 19514 6684 19654
rect 6826 19615 6882 19624
rect 6734 19544 6790 19553
rect 6644 19508 6696 19514
rect 6734 19479 6790 19488
rect 6644 19450 6696 19456
rect 6182 19207 6238 19216
rect 6552 19236 6604 19242
rect 6196 19174 6224 19207
rect 6552 19178 6604 19184
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6276 19168 6328 19174
rect 6276 19110 6328 19116
rect 6184 18896 6236 18902
rect 6184 18838 6236 18844
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6092 17808 6144 17814
rect 6196 17796 6224 18838
rect 6288 18766 6316 19110
rect 6276 18760 6328 18766
rect 6276 18702 6328 18708
rect 6144 17768 6224 17796
rect 6092 17750 6144 17756
rect 6104 17338 6132 17750
rect 6092 17332 6144 17338
rect 6092 17274 6144 17280
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 6012 16250 6040 16390
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6104 14074 6132 17070
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6092 14068 6144 14074
rect 6092 14010 6144 14016
rect 6104 12442 6132 14010
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 5816 6180 5868 6186
rect 5816 6122 5868 6128
rect 5828 5914 5856 6122
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 5816 5908 5868 5914
rect 5816 5850 5868 5856
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5736 4282 5764 5306
rect 5828 5302 5856 5850
rect 6104 5574 6132 6054
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6196 4826 6224 14554
rect 6288 12102 6316 18702
rect 6748 18290 6776 19479
rect 6826 18456 6882 18465
rect 6826 18391 6882 18400
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6642 18184 6698 18193
rect 6642 18119 6698 18128
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6380 17241 6408 18022
rect 6656 17882 6684 18119
rect 6644 17876 6696 17882
rect 6644 17818 6696 17824
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6656 17338 6684 17682
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6366 17232 6422 17241
rect 6366 17167 6422 17176
rect 6552 16516 6604 16522
rect 6552 16458 6604 16464
rect 6564 16046 6592 16458
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6368 15904 6420 15910
rect 6368 15846 6420 15852
rect 6380 15366 6408 15846
rect 6472 15609 6500 15982
rect 6656 15706 6684 17274
rect 6748 16130 6776 18226
rect 6840 18154 6868 18391
rect 6828 18148 6880 18154
rect 6828 18090 6880 18096
rect 6932 16232 6960 20402
rect 7024 19922 7052 22200
rect 7576 20534 7604 22200
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 7564 20528 7616 20534
rect 7564 20470 7616 20476
rect 7116 20058 7144 20470
rect 7576 20398 7604 20470
rect 8128 20398 8156 22200
rect 8208 20528 8260 20534
rect 8680 20516 8708 22200
rect 8944 20596 8996 20602
rect 8944 20538 8996 20544
rect 8680 20488 8800 20516
rect 8208 20470 8260 20476
rect 7564 20392 7616 20398
rect 7564 20334 7616 20340
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 7288 20324 7340 20330
rect 7288 20266 7340 20272
rect 7472 20324 7524 20330
rect 7472 20266 7524 20272
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7102 19952 7158 19961
rect 7012 19916 7064 19922
rect 7102 19887 7158 19896
rect 7012 19858 7064 19864
rect 7024 18970 7052 19858
rect 7116 19718 7144 19887
rect 7196 19780 7248 19786
rect 7196 19722 7248 19728
rect 7104 19712 7156 19718
rect 7104 19654 7156 19660
rect 7104 19304 7156 19310
rect 7104 19246 7156 19252
rect 7012 18964 7064 18970
rect 7012 18906 7064 18912
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 7024 17882 7052 18294
rect 7116 18086 7144 19246
rect 7104 18080 7156 18086
rect 7104 18022 7156 18028
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7024 17377 7052 17818
rect 7116 17762 7144 18022
rect 7208 17882 7236 19722
rect 7300 19378 7328 20266
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7392 19553 7420 20198
rect 7378 19544 7434 19553
rect 7378 19479 7434 19488
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7116 17734 7236 17762
rect 7104 17536 7156 17542
rect 7104 17478 7156 17484
rect 7010 17368 7066 17377
rect 7010 17303 7066 17312
rect 7012 16244 7064 16250
rect 6932 16204 7012 16232
rect 7012 16186 7064 16192
rect 6748 16102 6960 16130
rect 6734 16008 6790 16017
rect 6734 15943 6790 15952
rect 6644 15700 6696 15706
rect 6564 15660 6644 15688
rect 6458 15600 6514 15609
rect 6458 15535 6514 15544
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 6472 14618 6500 15535
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6564 12434 6592 15660
rect 6644 15642 6696 15648
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6472 12406 6592 12434
rect 6276 12096 6328 12102
rect 6276 12038 6328 12044
rect 6472 9674 6500 12406
rect 6656 12322 6684 15302
rect 6748 13530 6776 15943
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6380 9646 6500 9674
rect 6564 12294 6684 12322
rect 6380 9110 6408 9646
rect 6368 9104 6420 9110
rect 6368 9046 6420 9052
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6288 6662 6316 8978
rect 6276 6656 6328 6662
rect 6276 6598 6328 6604
rect 6288 6118 6316 6598
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5184 2514 5212 2790
rect 5276 2514 5304 3470
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5828 2514 5856 3334
rect 5172 2508 5224 2514
rect 5172 2450 5224 2456
rect 5264 2508 5316 2514
rect 5264 2450 5316 2456
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 4724 2264 4844 2292
rect 4421 2204 4717 2224
rect 4477 2202 4501 2204
rect 4557 2202 4581 2204
rect 4637 2202 4661 2204
rect 4499 2150 4501 2202
rect 4563 2150 4575 2202
rect 4637 2150 4639 2202
rect 4477 2148 4501 2150
rect 4557 2148 4581 2150
rect 4637 2148 4661 2150
rect 4421 2128 4717 2148
rect 4816 1442 4844 2264
rect 4724 1414 4844 1442
rect 4724 800 4752 1414
rect 5276 800 5304 2450
rect 5828 800 5856 2450
rect 6196 1766 6224 4762
rect 6380 2582 6408 9046
rect 6564 7313 6592 12294
rect 6550 7304 6606 7313
rect 6550 7239 6606 7248
rect 6564 6866 6592 7239
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 6564 4146 6592 6802
rect 6748 4434 6776 13330
rect 6828 12912 6880 12918
rect 6828 12854 6880 12860
rect 6840 12220 6868 12854
rect 6932 12646 6960 16102
rect 7024 14822 7052 16186
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 7024 12322 7052 14758
rect 7116 13394 7144 17478
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 7208 12434 7236 17734
rect 7300 16833 7328 19314
rect 7380 19304 7432 19310
rect 7378 19272 7380 19281
rect 7432 19272 7434 19281
rect 7378 19207 7434 19216
rect 7380 19168 7432 19174
rect 7380 19110 7432 19116
rect 7392 18290 7420 19110
rect 7484 18970 7512 20266
rect 7886 20156 8182 20176
rect 7942 20154 7966 20156
rect 8022 20154 8046 20156
rect 8102 20154 8126 20156
rect 7964 20102 7966 20154
rect 8028 20102 8040 20154
rect 8102 20102 8104 20154
rect 7942 20100 7966 20102
rect 8022 20100 8046 20102
rect 8102 20100 8126 20102
rect 7886 20080 8182 20100
rect 8220 20058 8248 20470
rect 8772 20398 8800 20488
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8850 20360 8906 20369
rect 8392 20324 8444 20330
rect 8850 20295 8906 20304
rect 8392 20266 8444 20272
rect 8404 20233 8432 20266
rect 8864 20262 8892 20295
rect 8668 20256 8720 20262
rect 8390 20224 8446 20233
rect 8668 20198 8720 20204
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8390 20159 8446 20168
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7656 19916 7708 19922
rect 7656 19858 7708 19864
rect 8116 19916 8168 19922
rect 8392 19916 8444 19922
rect 8168 19876 8248 19904
rect 8116 19858 8168 19864
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7484 18426 7512 18634
rect 7472 18420 7524 18426
rect 7472 18362 7524 18368
rect 7576 18358 7604 19314
rect 7564 18352 7616 18358
rect 7470 18320 7526 18329
rect 7380 18284 7432 18290
rect 7564 18294 7616 18300
rect 7470 18255 7526 18264
rect 7668 18272 7696 19858
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 8128 19689 8156 19722
rect 8114 19680 8170 19689
rect 8114 19615 8170 19624
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7760 18737 7788 19110
rect 7886 19068 8182 19088
rect 7942 19066 7966 19068
rect 8022 19066 8046 19068
rect 8102 19066 8126 19068
rect 7964 19014 7966 19066
rect 8028 19014 8040 19066
rect 8102 19014 8104 19066
rect 7942 19012 7966 19014
rect 8022 19012 8046 19014
rect 8102 19012 8126 19014
rect 7886 18992 8182 19012
rect 7852 18822 8064 18850
rect 7746 18728 7802 18737
rect 7852 18698 7880 18822
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 7746 18663 7802 18672
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7840 18420 7892 18426
rect 7760 18380 7840 18408
rect 7380 18226 7432 18232
rect 7484 18086 7512 18255
rect 7668 18244 7716 18272
rect 7472 18080 7524 18086
rect 7688 18068 7716 18244
rect 7472 18022 7524 18028
rect 7668 18040 7716 18068
rect 7378 17776 7434 17785
rect 7378 17711 7434 17720
rect 7392 17678 7420 17711
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7286 16824 7342 16833
rect 7286 16759 7342 16768
rect 7288 16652 7340 16658
rect 7288 16594 7340 16600
rect 7300 14618 7328 16594
rect 7392 15366 7420 17002
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7288 14612 7340 14618
rect 7288 14554 7340 14560
rect 7300 12782 7328 14554
rect 7392 14414 7420 15302
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7380 14272 7432 14278
rect 7380 14214 7432 14220
rect 7392 13190 7420 14214
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7208 12406 7328 12434
rect 7024 12294 7236 12322
rect 7104 12232 7156 12238
rect 6840 12192 7052 12220
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6840 5692 6868 7414
rect 6932 6390 6960 12038
rect 7024 8090 7052 12192
rect 7104 12174 7156 12180
rect 7116 8922 7144 12174
rect 7208 9042 7236 12294
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7194 8936 7250 8945
rect 7116 8894 7194 8922
rect 7194 8871 7250 8880
rect 7208 8634 7236 8871
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 8514 7328 12406
rect 7392 11626 7420 13126
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7392 11354 7420 11562
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7392 9722 7420 10746
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7116 8486 7328 8514
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6932 5817 6960 6054
rect 6918 5808 6974 5817
rect 6918 5743 6974 5752
rect 6840 5664 6960 5692
rect 6932 4826 6960 5664
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6932 4622 6960 4762
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6748 4406 6960 4434
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6564 3466 6592 4082
rect 6552 3460 6604 3466
rect 6552 3402 6604 3408
rect 6932 3233 6960 4406
rect 7024 3738 7052 8026
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7024 3369 7052 3674
rect 7116 3505 7144 8486
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7208 7449 7236 8230
rect 7194 7440 7250 7449
rect 7194 7375 7250 7384
rect 7208 3670 7236 7375
rect 7392 7154 7420 9658
rect 7484 9081 7512 18022
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7576 17338 7604 17614
rect 7668 17542 7696 18040
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7564 17332 7616 17338
rect 7564 17274 7616 17280
rect 7760 15552 7788 18380
rect 7840 18362 7892 18368
rect 7944 18329 7972 18702
rect 8036 18426 8064 18822
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 7930 18320 7986 18329
rect 7930 18255 7986 18264
rect 7886 17980 8182 18000
rect 7942 17978 7966 17980
rect 8022 17978 8046 17980
rect 8102 17978 8126 17980
rect 7964 17926 7966 17978
rect 8028 17926 8040 17978
rect 8102 17926 8104 17978
rect 7942 17924 7966 17926
rect 8022 17924 8046 17926
rect 8102 17924 8126 17926
rect 7886 17904 8182 17924
rect 8220 17241 8248 19876
rect 8392 19858 8444 19864
rect 8576 19916 8628 19922
rect 8576 19858 8628 19864
rect 8298 19272 8354 19281
rect 8298 19207 8354 19216
rect 8312 19174 8340 19207
rect 8300 19168 8352 19174
rect 8300 19110 8352 19116
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8206 17232 8262 17241
rect 8312 17202 8340 18022
rect 8206 17167 8262 17176
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7886 16892 8182 16912
rect 7942 16890 7966 16892
rect 8022 16890 8046 16892
rect 8102 16890 8126 16892
rect 7964 16838 7966 16890
rect 8028 16838 8040 16890
rect 8102 16838 8104 16890
rect 7942 16836 7966 16838
rect 8022 16836 8046 16838
rect 8102 16836 8126 16838
rect 7886 16816 8182 16836
rect 8114 16688 8170 16697
rect 8114 16623 8170 16632
rect 8128 15978 8156 16623
rect 8312 16590 8340 17138
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8300 16448 8352 16454
rect 8300 16390 8352 16396
rect 8116 15972 8168 15978
rect 8116 15914 8168 15920
rect 8312 15858 8340 16390
rect 8404 15978 8432 19858
rect 8484 18828 8536 18834
rect 8484 18770 8536 18776
rect 8496 17814 8524 18770
rect 8588 18630 8616 19858
rect 8576 18624 8628 18630
rect 8576 18566 8628 18572
rect 8574 18184 8630 18193
rect 8574 18119 8630 18128
rect 8484 17808 8536 17814
rect 8484 17750 8536 17756
rect 8496 16794 8524 17750
rect 8588 16810 8616 18119
rect 8680 18057 8708 20198
rect 8956 20058 8984 20538
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 9232 19310 9260 22200
rect 9784 20312 9812 22200
rect 10048 20460 10100 20466
rect 10048 20402 10100 20408
rect 9864 20324 9916 20330
rect 9784 20284 9864 20312
rect 9864 20266 9916 20272
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9312 19916 9364 19922
rect 9364 19876 9444 19904
rect 9312 19858 9364 19864
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 9220 19304 9272 19310
rect 9220 19246 9272 19252
rect 8760 19168 8812 19174
rect 8760 19110 8812 19116
rect 8772 18329 8800 19110
rect 8864 19009 8892 19246
rect 8850 19000 8906 19009
rect 8850 18935 8906 18944
rect 8758 18320 8814 18329
rect 8758 18255 8814 18264
rect 8852 18148 8904 18154
rect 8852 18090 8904 18096
rect 8666 18048 8722 18057
rect 8864 18034 8892 18090
rect 8864 18006 8984 18034
rect 8666 17983 8722 17992
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8680 17270 8708 17478
rect 8668 17264 8720 17270
rect 8668 17206 8720 17212
rect 8484 16788 8536 16794
rect 8588 16782 8708 16810
rect 8484 16730 8536 16736
rect 8574 16688 8630 16697
rect 8574 16623 8576 16632
rect 8628 16623 8630 16632
rect 8576 16594 8628 16600
rect 8576 16516 8628 16522
rect 8576 16458 8628 16464
rect 8588 16046 8616 16458
rect 8576 16040 8628 16046
rect 8576 15982 8628 15988
rect 8392 15972 8444 15978
rect 8392 15914 8444 15920
rect 8484 15904 8536 15910
rect 8312 15830 8432 15858
rect 8484 15846 8536 15852
rect 8576 15904 8628 15910
rect 8576 15846 8628 15852
rect 7886 15804 8182 15824
rect 7942 15802 7966 15804
rect 8022 15802 8046 15804
rect 8102 15802 8126 15804
rect 7964 15750 7966 15802
rect 8028 15750 8040 15802
rect 8102 15750 8104 15802
rect 7942 15748 7966 15750
rect 8022 15748 8046 15750
rect 8102 15748 8126 15750
rect 7886 15728 8182 15748
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 7576 15524 7788 15552
rect 7470 9072 7526 9081
rect 7470 9007 7526 9016
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7484 8294 7512 8910
rect 7472 8288 7524 8294
rect 7472 8230 7524 8236
rect 7576 7426 7604 15524
rect 7840 15088 7892 15094
rect 7840 15030 7892 15036
rect 7656 14952 7708 14958
rect 7852 14929 7880 15030
rect 7656 14894 7708 14900
rect 7838 14920 7894 14929
rect 7668 14618 7696 14894
rect 7748 14884 7800 14890
rect 7838 14855 7894 14864
rect 7748 14826 7800 14832
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7656 14476 7708 14482
rect 7656 14418 7708 14424
rect 7668 13870 7696 14418
rect 7760 14074 7788 14826
rect 7886 14716 8182 14736
rect 7942 14714 7966 14716
rect 8022 14714 8046 14716
rect 8102 14714 8126 14716
rect 7964 14662 7966 14714
rect 8028 14662 8040 14714
rect 8102 14662 8104 14714
rect 7942 14660 7966 14662
rect 8022 14660 8046 14662
rect 8102 14660 8126 14662
rect 7886 14640 8182 14660
rect 8312 14482 8340 15642
rect 8404 14906 8432 15830
rect 8496 15570 8524 15846
rect 8484 15564 8536 15570
rect 8484 15506 8536 15512
rect 8588 15026 8616 15846
rect 8680 15706 8708 16782
rect 8668 15700 8720 15706
rect 8668 15642 8720 15648
rect 8668 15564 8720 15570
rect 8668 15506 8720 15512
rect 8680 15026 8708 15506
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8404 14878 8524 14906
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8404 14618 8432 14758
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7760 13462 7788 14010
rect 7852 14006 7880 14214
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 7840 14000 7892 14006
rect 7840 13942 7892 13948
rect 7886 13628 8182 13648
rect 7942 13626 7966 13628
rect 8022 13626 8046 13628
rect 8102 13626 8126 13628
rect 7964 13574 7966 13626
rect 8028 13574 8040 13626
rect 8102 13574 8104 13626
rect 7942 13572 7966 13574
rect 8022 13572 8046 13574
rect 8102 13572 8126 13574
rect 7886 13552 8182 13572
rect 7748 13456 7800 13462
rect 7654 13424 7710 13433
rect 7748 13398 7800 13404
rect 7654 13359 7710 13368
rect 7668 12918 7696 13359
rect 7760 12986 7788 13398
rect 8312 13394 8340 14010
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8496 13274 8524 14878
rect 8576 14272 8628 14278
rect 8574 14240 8576 14249
rect 8628 14240 8630 14249
rect 8574 14175 8630 14184
rect 8220 13246 8524 13274
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 8974 7696 12582
rect 7886 12540 8182 12560
rect 7942 12538 7966 12540
rect 8022 12538 8046 12540
rect 8102 12538 8126 12540
rect 7964 12486 7966 12538
rect 8028 12486 8040 12538
rect 8102 12486 8104 12538
rect 7942 12484 7966 12486
rect 8022 12484 8046 12486
rect 8102 12484 8126 12486
rect 7886 12464 8182 12484
rect 8114 12336 8170 12345
rect 7748 12300 7800 12306
rect 8114 12271 8116 12280
rect 7748 12242 7800 12248
rect 8168 12271 8170 12280
rect 8116 12242 8168 12248
rect 7760 11898 7788 12242
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7760 11801 7788 11834
rect 7746 11792 7802 11801
rect 7746 11727 7802 11736
rect 8220 11642 8248 13246
rect 8392 13184 8444 13190
rect 8392 13126 8444 13132
rect 8404 12714 8432 13126
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8298 12472 8354 12481
rect 8298 12407 8354 12416
rect 8312 12306 8340 12407
rect 8300 12300 8352 12306
rect 8300 12242 8352 12248
rect 8404 11762 8432 12650
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12238 8524 12582
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8496 11694 8524 12174
rect 8484 11688 8536 11694
rect 8220 11614 8340 11642
rect 8484 11630 8536 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 7886 11452 8182 11472
rect 7942 11450 7966 11452
rect 8022 11450 8046 11452
rect 8102 11450 8126 11452
rect 7964 11398 7966 11450
rect 8028 11398 8040 11450
rect 8102 11398 8104 11450
rect 7942 11396 7966 11398
rect 8022 11396 8046 11398
rect 8102 11396 8126 11398
rect 7886 11376 8182 11396
rect 8220 11354 8248 11494
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11234 8340 11614
rect 8220 11206 8340 11234
rect 7886 10364 8182 10384
rect 7942 10362 7966 10364
rect 8022 10362 8046 10364
rect 8102 10362 8126 10364
rect 7964 10310 7966 10362
rect 8028 10310 8040 10362
rect 8102 10310 8104 10362
rect 7942 10308 7966 10310
rect 8022 10308 8046 10310
rect 8102 10308 8126 10310
rect 7746 10296 7802 10305
rect 7886 10288 8182 10308
rect 7746 10231 7802 10240
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7656 8832 7708 8838
rect 7760 8820 7788 10231
rect 8220 9330 8248 11206
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8404 10266 8432 10950
rect 8588 10690 8616 14175
rect 8772 14074 8800 17682
rect 8956 17338 8984 18006
rect 9048 17649 9076 19246
rect 9312 19168 9364 19174
rect 9232 19128 9312 19156
rect 9232 18766 9260 19128
rect 9312 19110 9364 19116
rect 9312 18896 9364 18902
rect 9416 18873 9444 19876
rect 9312 18838 9364 18844
rect 9402 18864 9458 18873
rect 9220 18760 9272 18766
rect 9140 18720 9220 18748
rect 9140 18086 9168 18720
rect 9220 18702 9272 18708
rect 9324 18290 9352 18838
rect 9402 18799 9458 18808
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9128 18080 9180 18086
rect 9128 18022 9180 18028
rect 9140 17882 9168 18022
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 9034 17640 9090 17649
rect 9034 17575 9090 17584
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9048 17184 9076 17575
rect 9232 17513 9260 18090
rect 9324 17882 9352 18226
rect 9508 18170 9536 20198
rect 9770 20088 9826 20097
rect 9770 20023 9826 20032
rect 9784 19990 9812 20023
rect 9772 19984 9824 19990
rect 9772 19926 9824 19932
rect 9588 19916 9640 19922
rect 9588 19858 9640 19864
rect 9416 18142 9536 18170
rect 9416 17921 9444 18142
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9402 17912 9458 17921
rect 9312 17876 9364 17882
rect 9402 17847 9458 17856
rect 9312 17818 9364 17824
rect 9218 17504 9274 17513
rect 9218 17439 9274 17448
rect 9048 17156 9168 17184
rect 9034 17096 9090 17105
rect 8944 17060 8996 17066
rect 9034 17031 9090 17040
rect 8944 17002 8996 17008
rect 8956 16794 8984 17002
rect 9048 16998 9076 17031
rect 9036 16992 9088 16998
rect 9036 16934 9088 16940
rect 9140 16810 9168 17156
rect 9048 16794 9168 16810
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 9036 16788 9168 16794
rect 9088 16782 9168 16788
rect 9036 16730 9088 16736
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8850 14376 8906 14385
rect 8850 14311 8852 14320
rect 8904 14311 8906 14320
rect 8852 14282 8904 14288
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 8956 13954 8984 16458
rect 8772 13926 8984 13954
rect 8772 12434 8800 13926
rect 8852 13864 8904 13870
rect 8852 13806 8904 13812
rect 8496 10662 8616 10690
rect 8680 12406 8800 12434
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8392 9376 8444 9382
rect 8220 9302 8340 9330
rect 8496 9364 8524 10662
rect 8576 10600 8628 10606
rect 8574 10568 8576 10577
rect 8628 10568 8630 10577
rect 8574 10503 8630 10512
rect 8444 9336 8524 9364
rect 8392 9318 8444 9324
rect 7886 9276 8182 9296
rect 7942 9274 7966 9276
rect 8022 9274 8046 9276
rect 8102 9274 8126 9276
rect 7964 9222 7966 9274
rect 8028 9222 8040 9274
rect 8102 9222 8104 9274
rect 7942 9220 7966 9222
rect 8022 9220 8046 9222
rect 8102 9220 8126 9222
rect 7886 9200 8182 9220
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 7708 8792 7788 8820
rect 7656 8774 7708 8780
rect 7668 7546 7696 8774
rect 8128 8430 8156 8842
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7576 7398 7696 7426
rect 7564 7200 7616 7206
rect 7392 7126 7512 7154
rect 7564 7142 7616 7148
rect 7668 7154 7696 7398
rect 7760 7342 7788 8366
rect 7886 8188 8182 8208
rect 7942 8186 7966 8188
rect 8022 8186 8046 8188
rect 8102 8186 8126 8188
rect 7964 8134 7966 8186
rect 8028 8134 8040 8186
rect 8102 8134 8104 8186
rect 7942 8132 7966 8134
rect 8022 8132 8046 8134
rect 8102 8132 8126 8134
rect 7886 8112 8182 8132
rect 8312 7834 8340 9302
rect 8128 7806 8340 7834
rect 8128 7478 8156 7806
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 8208 7200 8260 7206
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7300 5522 7328 6326
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5681 7420 6190
rect 7378 5672 7434 5681
rect 7378 5607 7434 5616
rect 7484 5574 7512 7126
rect 7576 6322 7604 7142
rect 7668 7126 7788 7154
rect 8208 7142 8260 7148
rect 7654 6896 7710 6905
rect 7654 6831 7656 6840
rect 7708 6831 7710 6840
rect 7656 6802 7708 6808
rect 7760 6746 7788 7126
rect 7886 7100 8182 7120
rect 7942 7098 7966 7100
rect 8022 7098 8046 7100
rect 8102 7098 8126 7100
rect 7964 7046 7966 7098
rect 8028 7046 8040 7098
rect 8102 7046 8104 7098
rect 7942 7044 7966 7046
rect 8022 7044 8046 7046
rect 8102 7044 8126 7046
rect 7886 7024 8182 7044
rect 8116 6860 8168 6866
rect 8116 6802 8168 6808
rect 7668 6718 7788 6746
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7576 5778 7604 6258
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 7472 5568 7524 5574
rect 7300 5494 7420 5522
rect 7472 5510 7524 5516
rect 7288 5092 7340 5098
rect 7288 5034 7340 5040
rect 7300 4593 7328 5034
rect 7286 4584 7342 4593
rect 7286 4519 7342 4528
rect 7300 3942 7328 4519
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7300 3738 7328 3878
rect 7288 3732 7340 3738
rect 7288 3674 7340 3680
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7102 3496 7158 3505
rect 7102 3431 7158 3440
rect 7104 3392 7156 3398
rect 7010 3360 7066 3369
rect 7104 3334 7156 3340
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7010 3295 7066 3304
rect 6918 3224 6974 3233
rect 6918 3159 6974 3168
rect 7116 3058 7144 3334
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 6932 2961 6960 2994
rect 7300 2990 7328 3334
rect 7012 2984 7064 2990
rect 6918 2952 6974 2961
rect 7012 2926 7064 2932
rect 7288 2984 7340 2990
rect 7288 2926 7340 2932
rect 6918 2887 6974 2896
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6368 2576 6420 2582
rect 6368 2518 6420 2524
rect 6472 2514 6500 2790
rect 6460 2508 6512 2514
rect 6460 2450 6512 2456
rect 6184 1760 6236 1766
rect 6184 1702 6236 1708
rect 6472 800 6500 2450
rect 7024 800 7052 2926
rect 7392 2582 7420 5494
rect 7576 5302 7604 5607
rect 7564 5296 7616 5302
rect 7564 5238 7616 5244
rect 7576 4758 7604 5238
rect 7668 5137 7696 6718
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6225 7880 6598
rect 8128 6361 8156 6802
rect 8114 6352 8170 6361
rect 8114 6287 8170 6296
rect 7838 6216 7894 6225
rect 7748 6180 7800 6186
rect 7838 6151 7894 6160
rect 7748 6122 7800 6128
rect 7760 5914 7788 6122
rect 7886 6012 8182 6032
rect 7942 6010 7966 6012
rect 8022 6010 8046 6012
rect 8102 6010 8126 6012
rect 7964 5958 7966 6010
rect 8028 5958 8040 6010
rect 8102 5958 8104 6010
rect 7942 5956 7966 5958
rect 8022 5956 8046 5958
rect 8102 5956 8126 5958
rect 7886 5936 8182 5956
rect 7748 5908 7800 5914
rect 7748 5850 7800 5856
rect 8220 5778 8248 7142
rect 8312 6934 8340 7686
rect 8404 7041 8432 9318
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8390 7032 8446 7041
rect 8390 6967 8446 6976
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8404 5846 8432 6967
rect 8392 5840 8444 5846
rect 8392 5782 8444 5788
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 7654 5128 7710 5137
rect 7654 5063 7710 5072
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7656 4480 7708 4486
rect 7656 4422 7708 4428
rect 7470 3632 7526 3641
rect 7470 3567 7526 3576
rect 7484 2854 7512 3567
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7380 2576 7432 2582
rect 7380 2518 7432 2524
rect 7576 2496 7604 3334
rect 7668 2961 7696 4422
rect 7760 3720 7788 5714
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 7886 4924 8182 4944
rect 7942 4922 7966 4924
rect 8022 4922 8046 4924
rect 8102 4922 8126 4924
rect 7964 4870 7966 4922
rect 8028 4870 8040 4922
rect 8102 4870 8104 4922
rect 7942 4868 7966 4870
rect 8022 4868 8046 4870
rect 8102 4868 8126 4870
rect 7886 4848 8182 4868
rect 8312 4826 8340 5238
rect 8300 4820 8352 4826
rect 8300 4762 8352 4768
rect 8392 4752 8444 4758
rect 8392 4694 8444 4700
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8022 4312 8078 4321
rect 8022 4247 8078 4256
rect 8036 4078 8064 4247
rect 8312 4214 8340 4422
rect 8300 4208 8352 4214
rect 8300 4150 8352 4156
rect 8312 4078 8340 4150
rect 8024 4072 8076 4078
rect 8024 4014 8076 4020
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3936 8260 3942
rect 8300 3936 8352 3942
rect 8208 3878 8260 3884
rect 8298 3904 8300 3913
rect 8352 3904 8354 3913
rect 7886 3836 8182 3856
rect 7942 3834 7966 3836
rect 8022 3834 8046 3836
rect 8102 3834 8126 3836
rect 7964 3782 7966 3834
rect 8028 3782 8040 3834
rect 8102 3782 8104 3834
rect 7942 3780 7966 3782
rect 8022 3780 8046 3782
rect 8102 3780 8126 3782
rect 7886 3760 8182 3780
rect 7760 3692 7972 3720
rect 7944 3602 7972 3692
rect 7748 3596 7800 3602
rect 7748 3538 7800 3544
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7654 2952 7710 2961
rect 7654 2887 7710 2896
rect 7760 2553 7788 3538
rect 7840 3528 7892 3534
rect 7840 3470 7892 3476
rect 7852 3058 7880 3470
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7944 2990 7972 3334
rect 8036 2990 8064 3334
rect 8128 3058 8156 3402
rect 8116 3052 8168 3058
rect 8116 2994 8168 3000
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7886 2748 8182 2768
rect 7942 2746 7966 2748
rect 8022 2746 8046 2748
rect 8102 2746 8126 2748
rect 7964 2694 7966 2746
rect 8028 2694 8040 2746
rect 8102 2694 8104 2746
rect 7942 2692 7966 2694
rect 8022 2692 8046 2694
rect 8102 2692 8126 2694
rect 7886 2672 8182 2692
rect 7746 2544 7802 2553
rect 7656 2508 7708 2514
rect 7576 2468 7656 2496
rect 7576 800 7604 2468
rect 8220 2514 8248 3878
rect 8298 3839 8354 3848
rect 8404 3398 8432 4694
rect 8496 4321 8524 8298
rect 8588 5166 8616 10503
rect 8680 9382 8708 12406
rect 8758 12200 8814 12209
rect 8758 12135 8760 12144
rect 8812 12135 8814 12144
rect 8760 12106 8812 12112
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8680 8430 8708 8774
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8772 8362 8800 11834
rect 8864 11558 8892 13806
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8956 13462 8984 13670
rect 8944 13456 8996 13462
rect 8944 13398 8996 13404
rect 9048 12434 9076 16730
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8956 12406 9076 12434
rect 8852 11552 8904 11558
rect 8852 11494 8904 11500
rect 8864 10606 8892 11494
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8852 10464 8904 10470
rect 8850 10432 8852 10441
rect 8904 10432 8906 10441
rect 8850 10367 8906 10376
rect 8852 10260 8904 10266
rect 8852 10202 8904 10208
rect 8760 8356 8812 8362
rect 8760 8298 8812 8304
rect 8864 7886 8892 10202
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8956 7698 8984 12406
rect 9036 12164 9088 12170
rect 9036 12106 9088 12112
rect 9048 11393 9076 12106
rect 9034 11384 9090 11393
rect 9034 11319 9090 11328
rect 9048 11150 9076 11319
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9140 10554 9168 15642
rect 9232 14550 9260 17439
rect 9310 17368 9366 17377
rect 9310 17303 9366 17312
rect 9324 16522 9352 17303
rect 9416 16833 9444 17847
rect 9402 16824 9458 16833
rect 9402 16759 9458 16768
rect 9508 16658 9536 18022
rect 9600 17678 9628 19858
rect 9876 19854 9904 20266
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 9678 19408 9734 19417
rect 9678 19343 9734 19352
rect 9692 19310 9720 19343
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9692 18465 9720 19246
rect 9678 18456 9734 18465
rect 9678 18391 9734 18400
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9692 17746 9720 18294
rect 9772 18080 9824 18086
rect 9772 18022 9824 18028
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9600 16946 9628 17614
rect 9692 17134 9720 17682
rect 9784 17270 9812 18022
rect 9876 17338 9904 18022
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9862 17232 9918 17241
rect 9862 17167 9918 17176
rect 9680 17128 9732 17134
rect 9680 17070 9732 17076
rect 9772 16992 9824 16998
rect 9600 16940 9772 16946
rect 9600 16934 9824 16940
rect 9600 16918 9812 16934
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9600 16538 9628 16918
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9416 16510 9628 16538
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9416 14396 9444 16510
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9692 16046 9720 16390
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9588 15496 9640 15502
rect 9588 15438 9640 15444
rect 9678 15464 9734 15473
rect 9600 14482 9628 15438
rect 9678 15399 9734 15408
rect 9692 15162 9720 15399
rect 9680 15156 9732 15162
rect 9680 15098 9732 15104
rect 9784 15094 9812 16390
rect 9772 15088 9824 15094
rect 9772 15030 9824 15036
rect 9680 14884 9732 14890
rect 9680 14826 9732 14832
rect 9772 14884 9824 14890
rect 9772 14826 9824 14832
rect 9692 14793 9720 14826
rect 9678 14784 9734 14793
rect 9678 14719 9734 14728
rect 9784 14657 9812 14826
rect 9770 14648 9826 14657
rect 9770 14583 9826 14592
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9232 14368 9444 14396
rect 9232 12170 9260 14368
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9324 14113 9352 14214
rect 9310 14104 9366 14113
rect 9310 14039 9366 14048
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9324 11898 9352 14039
rect 9508 14006 9536 14214
rect 9496 14000 9548 14006
rect 9416 13960 9496 13988
rect 9416 12782 9444 13960
rect 9496 13942 9548 13948
rect 9494 13832 9550 13841
rect 9494 13767 9550 13776
rect 9404 12776 9456 12782
rect 9404 12718 9456 12724
rect 9402 12472 9458 12481
rect 9402 12407 9458 12416
rect 9416 12374 9444 12407
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9220 11688 9272 11694
rect 9220 11630 9272 11636
rect 9232 11082 9260 11630
rect 9508 11370 9536 13767
rect 9600 13716 9628 14418
rect 9876 13818 9904 17167
rect 9968 15065 9996 20198
rect 10060 19990 10088 20402
rect 10336 20398 10364 22200
rect 10598 20496 10654 20505
rect 10888 20482 10916 22200
rect 11440 20890 11468 22200
rect 11256 20862 11468 20890
rect 10888 20454 11008 20482
rect 10598 20431 10654 20440
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10416 20324 10468 20330
rect 10416 20266 10468 20272
rect 10508 20324 10560 20330
rect 10508 20266 10560 20272
rect 10048 19984 10100 19990
rect 10048 19926 10100 19932
rect 10324 19916 10376 19922
rect 10152 19876 10324 19904
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 19689 10088 19790
rect 10152 19786 10180 19876
rect 10324 19858 10376 19864
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 10046 19680 10102 19689
rect 10046 19615 10102 19624
rect 10048 19168 10100 19174
rect 10244 19156 10272 19722
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 10100 19128 10272 19156
rect 10048 19110 10100 19116
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 9954 15056 10010 15065
rect 9954 14991 10010 15000
rect 10152 15008 10180 18158
rect 10230 17368 10286 17377
rect 10230 17303 10232 17312
rect 10284 17303 10286 17312
rect 10232 17274 10284 17280
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 16250 10272 16526
rect 10232 16244 10284 16250
rect 10232 16186 10284 16192
rect 10336 16114 10364 19654
rect 10232 16108 10284 16114
rect 10232 16050 10284 16056
rect 10324 16108 10376 16114
rect 10324 16050 10376 16056
rect 10244 15570 10272 16050
rect 10232 15564 10284 15570
rect 10232 15506 10284 15512
rect 10428 15473 10456 20266
rect 10520 18034 10548 20266
rect 10612 19310 10640 20431
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10690 19680 10746 19689
rect 10690 19615 10746 19624
rect 10600 19304 10652 19310
rect 10600 19246 10652 19252
rect 10704 19242 10732 19615
rect 10692 19236 10744 19242
rect 10692 19178 10744 19184
rect 10704 18970 10732 19178
rect 10796 19145 10824 20334
rect 10782 19136 10838 19145
rect 10782 19071 10838 19080
rect 10692 18964 10744 18970
rect 10692 18906 10744 18912
rect 10782 18592 10838 18601
rect 10782 18527 10838 18536
rect 10796 18170 10824 18527
rect 10888 18358 10916 20334
rect 10980 20312 11008 20454
rect 11060 20324 11112 20330
rect 10980 20284 11060 20312
rect 11060 20266 11112 20272
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19961 11192 20198
rect 11150 19952 11206 19961
rect 11060 19916 11112 19922
rect 11150 19887 11206 19896
rect 11060 19858 11112 19864
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10980 19378 11008 19790
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10796 18142 10916 18170
rect 10520 18006 10824 18034
rect 10600 17808 10652 17814
rect 10600 17750 10652 17756
rect 10612 16153 10640 17750
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10704 16794 10732 17070
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10598 16144 10654 16153
rect 10520 16102 10598 16130
rect 10414 15464 10470 15473
rect 10414 15399 10470 15408
rect 10152 14980 10364 15008
rect 9956 14884 10008 14890
rect 10232 14884 10284 14890
rect 10008 14844 10232 14872
rect 9956 14826 10008 14832
rect 10232 14826 10284 14832
rect 9954 13968 10010 13977
rect 10336 13954 10364 14980
rect 9954 13903 9956 13912
rect 10008 13903 10010 13912
rect 10152 13926 10364 13954
rect 9956 13874 10008 13880
rect 9876 13790 9996 13818
rect 9600 13705 9720 13716
rect 9600 13696 9734 13705
rect 9600 13688 9678 13696
rect 9600 12782 9628 13688
rect 9968 13682 9996 13790
rect 9678 13631 9734 13640
rect 9876 13654 9996 13682
rect 9876 13546 9904 13654
rect 9784 13518 9904 13546
rect 9678 13288 9734 13297
rect 9678 13223 9680 13232
rect 9732 13223 9734 13232
rect 9680 13194 9732 13200
rect 9784 12889 9812 13518
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9876 12918 9904 13398
rect 10048 13388 10100 13394
rect 10048 13330 10100 13336
rect 9954 13016 10010 13025
rect 9954 12951 10010 12960
rect 9968 12918 9996 12951
rect 9864 12912 9916 12918
rect 9770 12880 9826 12889
rect 9864 12854 9916 12860
rect 9956 12912 10008 12918
rect 9956 12854 10008 12860
rect 9770 12815 9826 12824
rect 9588 12776 9640 12782
rect 9588 12718 9640 12724
rect 9784 11914 9812 12815
rect 9876 12646 9904 12854
rect 9864 12640 9916 12646
rect 9864 12582 9916 12588
rect 9784 11886 9904 11914
rect 10060 11898 10088 13330
rect 9772 11824 9824 11830
rect 9772 11766 9824 11772
rect 9324 11342 9536 11370
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 9140 10526 9260 10554
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 9140 10198 9168 10406
rect 9128 10192 9180 10198
rect 9128 10134 9180 10140
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9048 7970 9076 9318
rect 9140 9042 9168 10134
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9140 8090 9168 8366
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9048 7942 9168 7970
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8680 7670 8984 7698
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8576 5024 8628 5030
rect 8576 4966 8628 4972
rect 8588 4826 8616 4966
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8574 4720 8630 4729
rect 8574 4655 8630 4664
rect 8482 4312 8538 4321
rect 8482 4247 8538 4256
rect 8482 4040 8538 4049
rect 8482 3975 8538 3984
rect 8496 3942 8524 3975
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8484 2984 8536 2990
rect 8404 2932 8484 2938
rect 8404 2926 8536 2932
rect 8404 2910 8524 2926
rect 8404 2774 8432 2910
rect 8588 2854 8616 4655
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8312 2746 8432 2774
rect 7746 2479 7802 2488
rect 8208 2508 8260 2514
rect 7656 2450 7708 2456
rect 8208 2450 8260 2456
rect 8220 2122 8248 2450
rect 8312 2310 8340 2746
rect 8496 2378 8524 2790
rect 8680 2650 8708 7670
rect 9048 7562 9076 7822
rect 8956 7534 9076 7562
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8772 5914 8800 6666
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8864 6118 8892 6326
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8956 4842 8984 7534
rect 9036 7268 9088 7274
rect 9036 7210 9088 7216
rect 9048 6798 9076 7210
rect 9036 6792 9088 6798
rect 9036 6734 9088 6740
rect 9048 6118 9076 6734
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 9048 5710 9076 6054
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 9048 4865 9076 5238
rect 8772 4814 8984 4842
rect 9034 4856 9090 4865
rect 8772 2990 8800 4814
rect 9034 4791 9090 4800
rect 8852 4548 8904 4554
rect 8852 4490 8904 4496
rect 8864 3602 8892 4490
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8956 4185 8984 4422
rect 8942 4176 8998 4185
rect 8942 4111 8998 4120
rect 8944 3936 8996 3942
rect 8944 3878 8996 3884
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8850 3496 8906 3505
rect 8850 3431 8906 3440
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8864 2825 8892 3431
rect 8956 3058 8984 3878
rect 9048 3602 9076 4791
rect 9036 3596 9088 3602
rect 9036 3538 9088 3544
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 9036 2848 9088 2854
rect 8850 2816 8906 2825
rect 9036 2790 9088 2796
rect 8850 2751 8906 2760
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8128 2094 8248 2122
rect 8128 800 8156 2094
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8680 800 8708 1906
rect 8864 1698 8892 2246
rect 8852 1692 8904 1698
rect 8852 1634 8904 1640
rect 8956 1630 8984 2450
rect 9048 2106 9076 2790
rect 9140 2582 9168 7942
rect 9232 5370 9260 10526
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 5001 9260 5306
rect 9324 5302 9352 11342
rect 9784 11286 9812 11766
rect 9404 11280 9456 11286
rect 9772 11280 9824 11286
rect 9456 11228 9720 11234
rect 9404 11222 9720 11228
rect 9772 11222 9824 11228
rect 9416 11206 9720 11222
rect 9588 10464 9640 10470
rect 9588 10406 9640 10412
rect 9600 10169 9628 10406
rect 9586 10160 9642 10169
rect 9586 10095 9642 10104
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9508 9722 9536 9862
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9404 9444 9456 9450
rect 9404 9386 9456 9392
rect 9416 9110 9444 9386
rect 9508 9178 9536 9454
rect 9600 9194 9628 9590
rect 9692 9518 9720 11206
rect 9876 11132 9904 11886
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9784 11104 9904 11132
rect 9680 9512 9732 9518
rect 9680 9454 9732 9460
rect 9496 9172 9548 9178
rect 9600 9166 9720 9194
rect 9496 9114 9548 9120
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9416 8634 9444 8910
rect 9494 8800 9550 8809
rect 9494 8735 9550 8744
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 6254 9444 6598
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9402 6080 9458 6089
rect 9402 6015 9458 6024
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9312 5160 9364 5166
rect 9312 5102 9364 5108
rect 9218 4992 9274 5001
rect 9218 4927 9274 4936
rect 9232 3074 9260 4927
rect 9324 4826 9352 5102
rect 9312 4820 9364 4826
rect 9312 4762 9364 4768
rect 9312 4684 9364 4690
rect 9312 4626 9364 4632
rect 9324 4457 9352 4626
rect 9416 4554 9444 6015
rect 9404 4548 9456 4554
rect 9404 4490 9456 4496
rect 9310 4448 9366 4457
rect 9310 4383 9366 4392
rect 9508 4282 9536 8735
rect 9600 8634 9628 8978
rect 9692 8634 9720 9166
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9784 7993 9812 11104
rect 9956 11008 10008 11014
rect 9956 10950 10008 10956
rect 9968 10606 9996 10950
rect 9956 10600 10008 10606
rect 10008 10560 10088 10588
rect 9956 10542 10008 10548
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10062 9904 10406
rect 10060 10062 10088 10560
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 10048 10056 10100 10062
rect 10048 9998 10100 10004
rect 10046 9616 10102 9625
rect 10046 9551 10048 9560
rect 10100 9551 10102 9560
rect 10048 9522 10100 9528
rect 9864 9512 9916 9518
rect 9864 9454 9916 9460
rect 9876 8090 9904 9454
rect 10152 8650 10180 13926
rect 10416 13864 10468 13870
rect 10416 13806 10468 13812
rect 10324 13796 10376 13802
rect 10324 13738 10376 13744
rect 10336 13705 10364 13738
rect 10322 13696 10378 13705
rect 10322 13631 10378 13640
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 10244 12918 10272 13262
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10428 12714 10456 13806
rect 10416 12708 10468 12714
rect 10416 12650 10468 12656
rect 10232 12436 10284 12442
rect 10520 12434 10548 16102
rect 10598 16079 10654 16088
rect 10796 15314 10824 18006
rect 10612 15286 10824 15314
rect 10612 14521 10640 15286
rect 10690 15056 10746 15065
rect 10690 14991 10746 15000
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10232 12378 10284 12384
rect 10428 12406 10548 12434
rect 10244 11898 10272 12378
rect 10324 12300 10376 12306
rect 10324 12242 10376 12248
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 9968 8622 10180 8650
rect 9968 8566 9996 8622
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 10138 8392 10194 8401
rect 10244 8378 10272 11630
rect 10336 11082 10364 12242
rect 10324 11076 10376 11082
rect 10324 11018 10376 11024
rect 10428 10266 10456 12406
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11762 10548 12038
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10612 11234 10640 14447
rect 10704 14074 10732 14991
rect 10888 14906 10916 18142
rect 10980 17678 11008 19314
rect 11072 18766 11100 19858
rect 11256 19802 11284 20862
rect 11352 20700 11648 20720
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11430 20646 11432 20698
rect 11494 20646 11506 20698
rect 11568 20646 11570 20698
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11352 20624 11648 20644
rect 12084 20534 12112 22200
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 11428 20528 11480 20534
rect 11428 20470 11480 20476
rect 12072 20528 12124 20534
rect 12268 20505 12296 20538
rect 12636 20534 12664 22200
rect 13188 20534 13216 22200
rect 13740 20534 13768 22200
rect 12624 20528 12676 20534
rect 12072 20470 12124 20476
rect 12254 20496 12310 20505
rect 11440 20058 11468 20470
rect 12624 20470 12676 20476
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 12254 20431 12310 20440
rect 11704 20324 11756 20330
rect 11704 20266 11756 20272
rect 12808 20324 12860 20330
rect 12808 20266 12860 20272
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 11428 20052 11480 20058
rect 11428 19994 11480 20000
rect 11164 19774 11284 19802
rect 11164 18850 11192 19774
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11256 18970 11284 19654
rect 11352 19612 11648 19632
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11430 19558 11432 19610
rect 11494 19558 11506 19610
rect 11568 19558 11570 19610
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11352 19536 11648 19556
rect 11428 19168 11480 19174
rect 11428 19110 11480 19116
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11164 18834 11284 18850
rect 11164 18828 11296 18834
rect 11164 18822 11244 18828
rect 11244 18770 11296 18776
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11060 18760 11112 18766
rect 11348 18714 11376 18770
rect 11440 18766 11468 19110
rect 11060 18702 11112 18708
rect 11256 18686 11376 18714
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11152 18216 11204 18222
rect 11152 18158 11204 18164
rect 11164 17785 11192 18158
rect 11256 18154 11284 18686
rect 11352 18524 11648 18544
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11430 18470 11432 18522
rect 11494 18470 11506 18522
rect 11568 18470 11570 18522
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11352 18448 11648 18468
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11150 17776 11206 17785
rect 11060 17740 11112 17746
rect 11150 17711 11206 17720
rect 11060 17682 11112 17688
rect 10968 17672 11020 17678
rect 10968 17614 11020 17620
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10980 17134 11008 17478
rect 11072 17241 11100 17682
rect 11164 17610 11192 17711
rect 11152 17604 11204 17610
rect 11152 17546 11204 17552
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 11256 17270 11284 17478
rect 11352 17436 11648 17456
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11430 17382 11432 17434
rect 11494 17382 11506 17434
rect 11568 17382 11570 17434
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11352 17360 11648 17380
rect 11152 17264 11204 17270
rect 11058 17232 11114 17241
rect 11152 17206 11204 17212
rect 11244 17264 11296 17270
rect 11244 17206 11296 17212
rect 11058 17167 11114 17176
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 10968 16720 11020 16726
rect 10968 16662 11020 16668
rect 10980 16561 11008 16662
rect 10966 16552 11022 16561
rect 10966 16487 11022 16496
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 10968 15428 11020 15434
rect 10968 15370 11020 15376
rect 10980 15026 11008 15370
rect 11072 15162 11100 15846
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10796 14878 10916 14906
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10692 13796 10744 13802
rect 10692 13738 10744 13744
rect 10704 13190 10732 13738
rect 10796 13462 10824 14878
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14550 11008 14758
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10692 13184 10744 13190
rect 10876 13184 10928 13190
rect 10744 13132 10824 13138
rect 10692 13126 10824 13132
rect 10876 13126 10928 13132
rect 10704 13110 10824 13126
rect 10796 12850 10824 13110
rect 10888 12986 10916 13126
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10784 12844 10836 12850
rect 10784 12786 10836 12792
rect 10690 12472 10746 12481
rect 10690 12407 10746 12416
rect 10704 12238 10732 12407
rect 10796 12238 10824 12786
rect 10876 12640 10928 12646
rect 10874 12608 10876 12617
rect 10928 12608 10930 12617
rect 10874 12543 10930 12552
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10692 12232 10744 12238
rect 10692 12174 10744 12180
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10520 11206 10640 11234
rect 10784 11212 10836 11218
rect 10416 10260 10468 10266
rect 10416 10202 10468 10208
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 9042 10364 9522
rect 10324 9036 10376 9042
rect 10324 8978 10376 8984
rect 10244 8350 10364 8378
rect 10138 8327 10140 8336
rect 10192 8327 10194 8336
rect 10140 8298 10192 8304
rect 9954 8256 10010 8265
rect 9954 8191 10010 8200
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9770 7984 9826 7993
rect 9680 7948 9732 7954
rect 9770 7919 9826 7928
rect 9680 7890 9732 7896
rect 9692 7002 9720 7890
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9862 7848 9918 7857
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9678 6760 9734 6769
rect 9600 6458 9628 6734
rect 9678 6695 9734 6704
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9692 6202 9720 6695
rect 9600 6186 9720 6202
rect 9588 6180 9720 6186
rect 9640 6174 9720 6180
rect 9588 6122 9640 6128
rect 9600 5545 9628 6122
rect 9784 5914 9812 7822
rect 9862 7783 9864 7792
rect 9916 7783 9918 7792
rect 9864 7754 9916 7760
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 9876 7177 9904 7278
rect 9862 7168 9918 7177
rect 9862 7103 9918 7112
rect 9864 6180 9916 6186
rect 9864 6122 9916 6128
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9876 5794 9904 6122
rect 9692 5766 9904 5794
rect 9586 5536 9642 5545
rect 9586 5471 9642 5480
rect 9692 4486 9720 5766
rect 9862 5400 9918 5409
rect 9862 5335 9918 5344
rect 9876 4690 9904 5335
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9680 4208 9732 4214
rect 9680 4150 9732 4156
rect 9692 4026 9720 4150
rect 9968 4078 9996 8191
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10060 7546 10088 7822
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10060 7342 10088 7482
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 10060 5846 10088 6054
rect 10048 5840 10100 5846
rect 10048 5782 10100 5788
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5166 10180 5510
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10138 4312 10194 4321
rect 10138 4247 10194 4256
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9956 4072 10008 4078
rect 9692 3998 9904 4026
rect 9956 4014 10008 4020
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9310 3632 9366 3641
rect 9310 3567 9366 3576
rect 9324 3194 9352 3567
rect 9494 3496 9550 3505
rect 9404 3460 9456 3466
rect 9456 3440 9494 3448
rect 9456 3431 9550 3440
rect 9456 3420 9536 3431
rect 9404 3402 9456 3408
rect 9784 3194 9812 3878
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9232 3046 9352 3074
rect 9324 2990 9352 3046
rect 9312 2984 9364 2990
rect 9312 2926 9364 2932
rect 9220 2916 9272 2922
rect 9220 2858 9272 2864
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 8944 1624 8996 1630
rect 8944 1566 8996 1572
rect 9232 800 9260 2858
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9508 2514 9536 2615
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 9508 1970 9536 2450
rect 9600 2417 9628 2790
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9586 2408 9642 2417
rect 9586 2343 9642 2352
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9784 800 9812 2450
rect 9876 1970 9904 3998
rect 10060 3534 10088 4150
rect 10152 4078 10180 4247
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10048 3392 10100 3398
rect 10048 3334 10100 3340
rect 10060 2990 10088 3334
rect 10152 3058 10180 3878
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10048 2984 10100 2990
rect 10048 2926 10100 2932
rect 9954 2680 10010 2689
rect 9954 2615 9956 2624
rect 10008 2615 10010 2624
rect 9956 2586 10008 2592
rect 10140 2576 10192 2582
rect 10244 2564 10272 8026
rect 10336 7002 10364 8350
rect 10428 7342 10456 10202
rect 10416 7336 10468 7342
rect 10416 7278 10468 7284
rect 10324 6996 10376 7002
rect 10324 6938 10376 6944
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 5681 10364 6734
rect 10322 5672 10378 5681
rect 10322 5607 10378 5616
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10336 5273 10364 5306
rect 10322 5264 10378 5273
rect 10322 5199 10378 5208
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10192 2536 10272 2564
rect 10140 2518 10192 2524
rect 10336 2514 10364 4082
rect 10428 2582 10456 7278
rect 10520 6798 10548 11206
rect 10784 11154 10836 11160
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 5914 10548 6598
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10612 4808 10640 11018
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10606 10732 10950
rect 10796 10713 10824 11154
rect 10888 11082 10916 12242
rect 10980 11694 11008 14486
rect 11164 14278 11192 17206
rect 11716 17202 11744 20266
rect 12070 20224 12126 20233
rect 12070 20159 12126 20168
rect 12084 19990 12112 20159
rect 12072 19984 12124 19990
rect 11794 19952 11850 19961
rect 12072 19926 12124 19932
rect 11794 19887 11850 19896
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11256 16114 11284 16594
rect 11352 16348 11648 16368
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11430 16294 11432 16346
rect 11494 16294 11506 16346
rect 11568 16294 11570 16346
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11352 16272 11648 16292
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15706 11284 16050
rect 11244 15700 11296 15706
rect 11244 15642 11296 15648
rect 11352 15260 11648 15280
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11430 15206 11432 15258
rect 11494 15206 11506 15258
rect 11568 15206 11570 15258
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11352 15184 11648 15204
rect 11716 14793 11744 16662
rect 11702 14784 11758 14793
rect 11702 14719 11758 14728
rect 11704 14544 11756 14550
rect 11704 14486 11756 14492
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 11060 14272 11112 14278
rect 11060 14214 11112 14220
rect 11152 14272 11204 14278
rect 11152 14214 11204 14220
rect 11072 13462 11100 14214
rect 11060 13456 11112 13462
rect 11060 13398 11112 13404
rect 11256 12986 11284 14350
rect 11352 14172 11648 14192
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11430 14118 11432 14170
rect 11494 14118 11506 14170
rect 11568 14118 11570 14170
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11352 14096 11648 14116
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11624 13394 11652 13806
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11352 13084 11648 13104
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11430 13030 11432 13082
rect 11494 13030 11506 13082
rect 11568 13030 11570 13082
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11352 13008 11648 13028
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11242 12608 11298 12617
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11218 11008 11630
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 10980 11121 11008 11154
rect 10966 11112 11022 11121
rect 10876 11076 10928 11082
rect 10966 11047 11022 11056
rect 10876 11018 10928 11024
rect 10876 10736 10928 10742
rect 10782 10704 10838 10713
rect 10876 10678 10928 10684
rect 10782 10639 10838 10648
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10888 10130 10916 10678
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 11072 10470 11100 10542
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 11060 10124 11112 10130
rect 11060 10066 11112 10072
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10704 9110 10732 9998
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 9110 10824 9318
rect 11072 9178 11100 10066
rect 11164 9178 11192 12582
rect 11242 12543 11298 12552
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 11060 9172 11112 9178
rect 11060 9114 11112 9120
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10784 9104 10836 9110
rect 10784 9046 10836 9052
rect 10888 9058 10916 9114
rect 10704 8922 10732 9046
rect 10888 9030 11192 9058
rect 10704 8894 11008 8922
rect 10692 8832 10744 8838
rect 10690 8800 10692 8809
rect 10744 8800 10746 8809
rect 10690 8735 10746 8744
rect 10980 8566 11008 8894
rect 11164 8634 11192 9030
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 10968 8560 11020 8566
rect 10690 8528 10746 8537
rect 10968 8502 11020 8508
rect 10690 8463 10746 8472
rect 11060 8492 11112 8498
rect 10704 6730 10732 8463
rect 11060 8434 11112 8440
rect 10784 8356 10836 8362
rect 10784 8298 10836 8304
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10796 7954 10824 8298
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 10888 7018 10916 8298
rect 10968 8288 11020 8294
rect 10968 8230 11020 8236
rect 10980 8090 11008 8230
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 10966 7984 11022 7993
rect 10966 7919 11022 7928
rect 10980 7274 11008 7919
rect 11072 7410 11100 8434
rect 11152 7880 11204 7886
rect 11152 7822 11204 7828
rect 11164 7546 11192 7822
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 10968 7268 11020 7274
rect 11256 7256 11284 12543
rect 11716 12442 11744 14486
rect 11808 13326 11836 19887
rect 12348 19712 12400 19718
rect 12348 19654 12400 19660
rect 12360 19242 12388 19654
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12440 19236 12492 19242
rect 12440 19178 12492 19184
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 11980 18624 12032 18630
rect 11886 18592 11942 18601
rect 11980 18566 12032 18572
rect 11886 18527 11942 18536
rect 11900 18290 11928 18527
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11992 18086 12020 18566
rect 12084 18290 12112 18770
rect 12176 18358 12204 19178
rect 12346 19000 12402 19009
rect 12256 18964 12308 18970
rect 12346 18935 12402 18944
rect 12256 18906 12308 18912
rect 12164 18352 12216 18358
rect 12164 18294 12216 18300
rect 12072 18284 12124 18290
rect 12072 18226 12124 18232
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11900 16046 11928 18022
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 16726 12020 17546
rect 12072 17536 12124 17542
rect 12268 17513 12296 18906
rect 12360 18850 12388 18935
rect 12452 18850 12480 19178
rect 12716 19168 12768 19174
rect 12716 19110 12768 19116
rect 12360 18822 12480 18850
rect 12346 18184 12402 18193
rect 12346 18119 12402 18128
rect 12360 17785 12388 18119
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12622 18048 12678 18057
rect 12452 17814 12480 18022
rect 12622 17983 12678 17992
rect 12440 17808 12492 17814
rect 12346 17776 12402 17785
rect 12532 17808 12584 17814
rect 12440 17750 12492 17756
rect 12530 17776 12532 17785
rect 12584 17776 12586 17785
rect 12346 17711 12402 17720
rect 12530 17711 12586 17720
rect 12532 17672 12584 17678
rect 12360 17620 12532 17626
rect 12360 17614 12584 17620
rect 12360 17598 12572 17614
rect 12072 17478 12124 17484
rect 12254 17504 12310 17513
rect 11980 16720 12032 16726
rect 11980 16662 12032 16668
rect 12084 16538 12112 17478
rect 12254 17439 12310 17448
rect 12254 17368 12310 17377
rect 12254 17303 12256 17312
rect 12308 17303 12310 17312
rect 12256 17274 12308 17280
rect 12164 17196 12216 17202
rect 12164 17138 12216 17144
rect 12176 16658 12204 17138
rect 12164 16652 12216 16658
rect 12164 16594 12216 16600
rect 12084 16510 12204 16538
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 11888 16040 11940 16046
rect 11888 15982 11940 15988
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15162 12020 15846
rect 12084 15706 12112 16390
rect 12176 16130 12204 16510
rect 12360 16250 12388 17598
rect 12636 17542 12664 17983
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12728 17202 12756 19110
rect 12820 18970 12848 20266
rect 13740 20058 13768 20266
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 12912 19514 12940 19858
rect 13268 19848 13320 19854
rect 13082 19816 13138 19825
rect 13268 19790 13320 19796
rect 13082 19751 13138 19760
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12806 18864 12862 18873
rect 12806 18799 12862 18808
rect 12820 18193 12848 18799
rect 12806 18184 12862 18193
rect 13096 18170 13124 19751
rect 13280 19514 13308 19790
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13542 19136 13598 19145
rect 13542 19071 13598 19080
rect 13556 18970 13584 19071
rect 13544 18964 13596 18970
rect 13544 18906 13596 18912
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13096 18142 13216 18170
rect 12806 18119 12862 18128
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12820 17082 12848 18119
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 12912 17785 12940 18022
rect 13096 17882 13124 18022
rect 13188 17882 13216 18142
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13176 17876 13228 17882
rect 13176 17818 13228 17824
rect 12898 17776 12954 17785
rect 12898 17711 12954 17720
rect 12728 17054 12848 17082
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12348 16244 12400 16250
rect 12348 16186 12400 16192
rect 12176 16102 12296 16130
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12072 15700 12124 15706
rect 12072 15642 12124 15648
rect 12176 15586 12204 15982
rect 12084 15558 12204 15586
rect 12084 15366 12112 15558
rect 12268 15450 12296 16102
rect 12348 16108 12400 16114
rect 12348 16050 12400 16056
rect 12176 15422 12296 15450
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11888 15088 11940 15094
rect 11888 15030 11940 15036
rect 11900 13870 11928 15030
rect 12176 15008 12204 15422
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 11992 14980 12204 15008
rect 11888 13864 11940 13870
rect 11888 13806 11940 13812
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 11992 13190 12020 14980
rect 12268 14958 12296 15302
rect 12360 15026 12388 16050
rect 12452 15994 12480 16390
rect 12544 16153 12572 16662
rect 12530 16144 12586 16153
rect 12530 16079 12586 16088
rect 12532 16040 12584 16046
rect 12452 15988 12532 15994
rect 12452 15982 12584 15988
rect 12452 15966 12572 15982
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12348 15020 12400 15026
rect 12348 14962 12400 14968
rect 12256 14952 12308 14958
rect 12256 14894 12308 14900
rect 12164 14884 12216 14890
rect 12164 14826 12216 14832
rect 12176 14482 12204 14826
rect 12256 14816 12308 14822
rect 12256 14758 12308 14764
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 12072 14408 12124 14414
rect 12070 14376 12072 14385
rect 12124 14376 12126 14385
rect 12070 14311 12126 14320
rect 12162 14104 12218 14113
rect 12162 14039 12164 14048
rect 12216 14039 12218 14048
rect 12164 14010 12216 14016
rect 12268 13462 12296 14758
rect 12452 14006 12480 15642
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12532 15156 12584 15162
rect 12532 15098 12584 15104
rect 12544 14657 12572 15098
rect 12636 15026 12664 15506
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12530 14648 12586 14657
rect 12530 14583 12586 14592
rect 12440 14000 12492 14006
rect 12492 13948 12664 13954
rect 12440 13942 12664 13948
rect 12452 13926 12664 13942
rect 12440 13864 12492 13870
rect 12440 13806 12492 13812
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 11888 13184 11940 13190
rect 11888 13126 11940 13132
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11900 12850 11928 13126
rect 11992 12986 12020 13126
rect 11980 12980 12032 12986
rect 11980 12922 12032 12928
rect 12176 12918 12204 13262
rect 12268 13161 12296 13398
rect 12254 13152 12310 13161
rect 12254 13087 12310 13096
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11704 12232 11756 12238
rect 11704 12174 11756 12180
rect 11352 11996 11648 12016
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11430 11942 11432 11994
rect 11494 11942 11506 11994
rect 11568 11942 11570 11994
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11352 11920 11648 11940
rect 11610 11656 11666 11665
rect 11610 11591 11666 11600
rect 11624 11354 11652 11591
rect 11612 11348 11664 11354
rect 11612 11290 11664 11296
rect 11716 11098 11744 12174
rect 11808 11898 11836 12378
rect 11900 12374 11928 12582
rect 12176 12434 12204 12854
rect 12452 12628 12480 13806
rect 12532 13728 12584 13734
rect 12532 13670 12584 13676
rect 12544 13025 12572 13670
rect 12530 13016 12586 13025
rect 12530 12951 12586 12960
rect 12452 12600 12572 12628
rect 12084 12406 12204 12434
rect 11888 12368 11940 12374
rect 11888 12310 11940 12316
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11992 11694 12020 12106
rect 11980 11688 12032 11694
rect 11980 11630 12032 11636
rect 12084 11336 12112 12406
rect 12162 12336 12218 12345
rect 12544 12306 12572 12600
rect 12162 12271 12218 12280
rect 12532 12300 12584 12306
rect 12176 11801 12204 12271
rect 12532 12242 12584 12248
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12162 11792 12218 11801
rect 12162 11727 12218 11736
rect 12452 11370 12480 12174
rect 12544 11898 12572 12242
rect 12532 11892 12584 11898
rect 12532 11834 12584 11840
rect 12636 11642 12664 13926
rect 12728 12434 12756 17054
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 15638 12848 16390
rect 12912 15706 12940 17711
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13268 15972 13320 15978
rect 13268 15914 13320 15920
rect 12900 15700 12952 15706
rect 12900 15642 12952 15648
rect 12808 15632 12860 15638
rect 12808 15574 12860 15580
rect 13280 15570 13308 15914
rect 13268 15564 13320 15570
rect 13268 15506 13320 15512
rect 12808 14408 12860 14414
rect 12808 14350 12860 14356
rect 12820 13802 12848 14350
rect 13372 13977 13400 16526
rect 13358 13968 13414 13977
rect 13358 13903 13414 13912
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 13372 13734 13400 13903
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 12728 12406 12848 12434
rect 12636 11614 12756 11642
rect 12268 11342 12480 11370
rect 12084 11308 12204 11336
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 11716 11070 12020 11098
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11352 10908 11648 10928
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11430 10854 11432 10906
rect 11494 10854 11506 10906
rect 11568 10854 11570 10906
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11352 10832 11648 10852
rect 11716 10470 11744 10950
rect 11704 10464 11756 10470
rect 11756 10424 11928 10452
rect 11704 10406 11756 10412
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11352 9820 11648 9840
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11430 9766 11432 9818
rect 11494 9766 11506 9818
rect 11568 9766 11570 9818
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11352 9744 11648 9764
rect 11808 9489 11836 10066
rect 11794 9480 11850 9489
rect 11794 9415 11850 9424
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11352 8732 11648 8752
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11430 8678 11432 8730
rect 11494 8678 11506 8730
rect 11568 8678 11570 8730
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11352 8656 11648 8676
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7954 11376 8298
rect 11716 8090 11744 8978
rect 11808 8294 11836 9114
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11796 8016 11848 8022
rect 11794 7984 11796 7993
rect 11848 7984 11850 7993
rect 11336 7948 11388 7954
rect 11794 7919 11850 7928
rect 11336 7890 11388 7896
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11352 7644 11648 7664
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11430 7590 11432 7642
rect 11494 7590 11506 7642
rect 11568 7590 11570 7642
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11352 7568 11648 7588
rect 11428 7472 11480 7478
rect 11428 7414 11480 7420
rect 11520 7472 11572 7478
rect 11808 7426 11836 7822
rect 11520 7414 11572 7420
rect 10968 7210 11020 7216
rect 11164 7228 11284 7256
rect 11164 7018 11192 7228
rect 10888 6990 11008 7018
rect 10876 6792 10928 6798
rect 10876 6734 10928 6740
rect 10692 6724 10744 6730
rect 10692 6666 10744 6672
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10704 5914 10732 6122
rect 10796 6118 10824 6666
rect 10888 6322 10916 6734
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 6112 10836 6118
rect 10784 6054 10836 6060
rect 10692 5908 10744 5914
rect 10692 5850 10744 5856
rect 10692 5704 10744 5710
rect 10796 5692 10824 6054
rect 10874 5944 10930 5953
rect 10874 5879 10930 5888
rect 10744 5664 10824 5692
rect 10692 5646 10744 5652
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 5234 10732 5510
rect 10888 5409 10916 5879
rect 10874 5400 10930 5409
rect 10874 5335 10930 5344
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10520 4780 10640 4808
rect 10520 4214 10548 4780
rect 10600 4684 10652 4690
rect 10704 4672 10732 5170
rect 10652 4644 10732 4672
rect 10600 4626 10652 4632
rect 10598 4448 10654 4457
rect 10598 4383 10654 4392
rect 10612 4282 10640 4383
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10888 4026 10916 5335
rect 10980 5030 11008 6990
rect 11072 6990 11192 7018
rect 11336 6996 11388 7002
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 10520 3998 10916 4026
rect 10520 3602 10548 3998
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 10692 3596 10744 3602
rect 10692 3538 10744 3544
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10508 3120 10560 3126
rect 10508 3062 10560 3068
rect 10520 2904 10548 3062
rect 10612 2972 10640 3470
rect 10704 3369 10732 3538
rect 10690 3360 10746 3369
rect 10690 3295 10746 3304
rect 10612 2944 10732 2972
rect 10520 2876 10640 2904
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 10612 2514 10640 2876
rect 10704 2854 10732 2944
rect 10692 2848 10744 2854
rect 10692 2790 10744 2796
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10600 2508 10652 2514
rect 10600 2450 10652 2456
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 10612 1850 10640 2450
rect 10796 2310 10824 3878
rect 10980 3738 11008 4422
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11072 3380 11100 6990
rect 11440 6984 11468 7414
rect 11532 7002 11560 7414
rect 11716 7398 11836 7426
rect 11388 6956 11468 6984
rect 11520 6996 11572 7002
rect 11336 6938 11388 6944
rect 11520 6938 11572 6944
rect 11152 6656 11204 6662
rect 11152 6598 11204 6604
rect 11164 5098 11192 6598
rect 11352 6556 11648 6576
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11430 6502 11432 6554
rect 11494 6502 11506 6554
rect 11568 6502 11570 6554
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11352 6480 11648 6500
rect 11352 5468 11648 5488
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11430 5414 11432 5466
rect 11494 5414 11506 5466
rect 11568 5414 11570 5466
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11352 5392 11648 5412
rect 11716 5166 11744 7398
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11808 5846 11836 6938
rect 11796 5840 11848 5846
rect 11796 5782 11848 5788
rect 11900 5692 11928 10424
rect 11808 5664 11928 5692
rect 11704 5160 11756 5166
rect 11704 5102 11756 5108
rect 11152 5092 11204 5098
rect 11152 5034 11204 5040
rect 11428 5092 11480 5098
rect 11428 5034 11480 5040
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11164 4214 11192 4490
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11164 3534 11192 4150
rect 11256 3738 11284 4966
rect 11440 4622 11468 5034
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11352 4380 11648 4400
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11430 4326 11432 4378
rect 11494 4326 11506 4378
rect 11568 4326 11570 4378
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11352 4304 11648 4324
rect 11716 4162 11744 4966
rect 11624 4134 11744 4162
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11624 3534 11652 4134
rect 11704 4072 11756 4078
rect 11704 4014 11756 4020
rect 11716 3738 11744 4014
rect 11704 3732 11756 3738
rect 11704 3674 11756 3680
rect 11808 3618 11836 5664
rect 11888 5160 11940 5166
rect 11888 5102 11940 5108
rect 11900 5001 11928 5102
rect 11886 4992 11942 5001
rect 11886 4927 11942 4936
rect 11992 4842 12020 11070
rect 12084 9674 12112 11154
rect 12176 9738 12204 11308
rect 12268 11286 12296 11342
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12348 11212 12400 11218
rect 12348 11154 12400 11160
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12268 10713 12296 10746
rect 12254 10704 12310 10713
rect 12360 10674 12388 11154
rect 12254 10639 12310 10648
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12440 10464 12492 10470
rect 12438 10432 12440 10441
rect 12492 10432 12494 10441
rect 12438 10367 12494 10376
rect 12636 10198 12664 10610
rect 12728 10470 12756 11614
rect 12820 10470 12848 12406
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12624 10192 12676 10198
rect 12624 10134 12676 10140
rect 12176 9710 12388 9738
rect 12084 9646 12204 9674
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 9178 12112 9318
rect 12072 9172 12124 9178
rect 12072 9114 12124 9120
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 8090 12112 8910
rect 12072 8084 12124 8090
rect 12072 8026 12124 8032
rect 12072 7812 12124 7818
rect 12072 7754 12124 7760
rect 12084 5642 12112 7754
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12072 5024 12124 5030
rect 12070 4992 12072 5001
rect 12124 4992 12126 5001
rect 12070 4927 12126 4936
rect 11992 4814 12112 4842
rect 12084 4049 12112 4814
rect 12070 4040 12126 4049
rect 11980 4004 12032 4010
rect 12070 3975 12126 3984
rect 11980 3946 12032 3952
rect 11716 3590 11836 3618
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11612 3528 11664 3534
rect 11612 3470 11664 3476
rect 11072 3352 11192 3380
rect 11164 2650 11192 3352
rect 11352 3292 11648 3312
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11430 3238 11432 3290
rect 11494 3238 11506 3290
rect 11568 3238 11570 3290
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11352 3216 11648 3236
rect 11716 2990 11744 3590
rect 11992 3398 12020 3946
rect 12072 3936 12124 3942
rect 12070 3904 12072 3913
rect 12124 3904 12126 3913
rect 12070 3839 12126 3848
rect 12176 3777 12204 9646
rect 12254 9072 12310 9081
rect 12254 9007 12310 9016
rect 12268 7546 12296 9007
rect 12360 8090 12388 9710
rect 12636 9586 12664 10134
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12544 9489 12572 9522
rect 12530 9480 12586 9489
rect 12440 9444 12492 9450
rect 12530 9415 12586 9424
rect 12440 9386 12492 9392
rect 12452 8430 12480 9386
rect 12532 9376 12584 9382
rect 12532 9318 12584 9324
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12544 8242 12572 9318
rect 12820 8838 12848 10406
rect 13004 10130 13032 13262
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13280 12782 13308 13126
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13464 12434 13492 18770
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13542 18456 13598 18465
rect 13542 18391 13544 18400
rect 13596 18391 13598 18400
rect 13544 18362 13596 18368
rect 13740 18290 13768 18702
rect 13728 18284 13780 18290
rect 13728 18226 13780 18232
rect 13832 17898 13860 19858
rect 13740 17870 13860 17898
rect 13636 17808 13688 17814
rect 13636 17750 13688 17756
rect 13544 17672 13596 17678
rect 13544 17614 13596 17620
rect 13556 17134 13584 17614
rect 13648 17338 13676 17750
rect 13636 17332 13688 17338
rect 13636 17274 13688 17280
rect 13544 17128 13596 17134
rect 13740 17082 13768 17870
rect 13544 17070 13596 17076
rect 13556 16522 13584 17070
rect 13648 17054 13768 17082
rect 13648 16998 13676 17054
rect 13636 16992 13688 16998
rect 13636 16934 13688 16940
rect 13924 16794 13952 20266
rect 14292 19990 14320 22200
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14476 20058 14504 20538
rect 14844 20346 14872 22200
rect 14752 20318 14872 20346
rect 14752 20058 14780 20318
rect 14817 20156 15113 20176
rect 14873 20154 14897 20156
rect 14953 20154 14977 20156
rect 15033 20154 15057 20156
rect 14895 20102 14897 20154
rect 14959 20102 14971 20154
rect 15033 20102 15035 20154
rect 14873 20100 14897 20102
rect 14953 20100 14977 20102
rect 15033 20100 15057 20102
rect 14817 20080 15113 20100
rect 15212 20058 15332 20074
rect 14464 20052 14516 20058
rect 14464 19994 14516 20000
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 15200 20052 15332 20058
rect 15252 20046 15332 20052
rect 15200 19994 15252 20000
rect 14280 19984 14332 19990
rect 14280 19926 14332 19932
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 15200 19916 15252 19922
rect 15200 19858 15252 19864
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14188 19168 14240 19174
rect 14188 19110 14240 19116
rect 14200 18970 14228 19110
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14004 18896 14056 18902
rect 14002 18864 14004 18873
rect 14056 18864 14058 18873
rect 14002 18799 14058 18808
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 13728 16788 13780 16794
rect 13728 16730 13780 16736
rect 13912 16788 13964 16794
rect 13912 16730 13964 16736
rect 13634 16552 13690 16561
rect 13544 16516 13596 16522
rect 13634 16487 13690 16496
rect 13544 16458 13596 16464
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13556 14618 13584 15642
rect 13648 14958 13676 16487
rect 13740 16425 13768 16730
rect 13726 16416 13782 16425
rect 13726 16351 13782 16360
rect 14016 15994 14044 18566
rect 14108 17678 14136 18702
rect 14200 18290 14228 18906
rect 14292 18698 14320 19246
rect 14280 18692 14332 18698
rect 14280 18634 14332 18640
rect 14384 18290 14412 19654
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14476 18170 14504 19858
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 14384 18142 14504 18170
rect 14278 18048 14334 18057
rect 14278 17983 14334 17992
rect 14096 17672 14148 17678
rect 14096 17614 14148 17620
rect 14108 17338 14136 17614
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 13924 15966 14044 15994
rect 14108 15978 14136 17274
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14096 15972 14148 15978
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 14958 13860 15370
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13832 14074 13860 14894
rect 13924 14618 13952 15966
rect 14096 15914 14148 15920
rect 14004 15904 14056 15910
rect 14004 15846 14056 15852
rect 14016 15706 14044 15846
rect 14004 15700 14056 15706
rect 14004 15642 14056 15648
rect 14096 15564 14148 15570
rect 14096 15506 14148 15512
rect 13912 14612 13964 14618
rect 13912 14554 13964 14560
rect 13910 14376 13966 14385
rect 13910 14311 13912 14320
rect 13964 14311 13966 14320
rect 13912 14282 13964 14288
rect 14108 14074 14136 15506
rect 14200 14482 14228 17206
rect 14292 16794 14320 17983
rect 14280 16788 14332 16794
rect 14280 16730 14332 16736
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 14292 14618 14320 16594
rect 14280 14612 14332 14618
rect 14280 14554 14332 14560
rect 14188 14476 14240 14482
rect 14188 14418 14240 14424
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14188 13728 14240 13734
rect 14188 13670 14240 13676
rect 14096 13320 14148 13326
rect 14096 13262 14148 13268
rect 14108 12850 14136 13262
rect 14096 12844 14148 12850
rect 14096 12786 14148 12792
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13372 12406 13492 12434
rect 13820 12436 13872 12442
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 13280 11898 13308 12242
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13280 11762 13308 11834
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11150 13124 11562
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 13268 11144 13320 11150
rect 13268 11086 13320 11092
rect 13280 10810 13308 11086
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13268 9648 13320 9654
rect 13372 9625 13400 12406
rect 13820 12378 13872 12384
rect 13544 12368 13596 12374
rect 13728 12368 13780 12374
rect 13544 12310 13596 12316
rect 13726 12336 13728 12345
rect 13780 12336 13782 12345
rect 13556 11898 13584 12310
rect 13726 12271 13782 12280
rect 13726 12200 13782 12209
rect 13726 12135 13728 12144
rect 13780 12135 13782 12144
rect 13728 12106 13780 12112
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13832 11830 13860 12378
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 13820 11620 13872 11626
rect 13820 11562 13872 11568
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13648 11218 13676 11494
rect 13740 11354 13768 11494
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13832 10690 13860 11562
rect 13924 10810 13952 12582
rect 14108 12442 14136 12786
rect 14096 12436 14148 12442
rect 14096 12378 14148 12384
rect 14004 12300 14056 12306
rect 14004 12242 14056 12248
rect 14016 12102 14044 12242
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13832 10662 13952 10690
rect 14016 10674 14044 12038
rect 14200 11937 14228 13670
rect 14292 13530 14320 14554
rect 14280 13524 14332 13530
rect 14280 13466 14332 13472
rect 14292 12209 14320 13466
rect 14278 12200 14334 12209
rect 14278 12135 14334 12144
rect 14186 11928 14242 11937
rect 14186 11863 14242 11872
rect 14292 11778 14320 12135
rect 14384 12073 14412 18142
rect 14464 18080 14516 18086
rect 14462 18048 14464 18057
rect 14516 18048 14518 18057
rect 14462 17983 14518 17992
rect 14568 17746 14596 19654
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14752 19417 14780 19450
rect 14738 19408 14794 19417
rect 14738 19343 14794 19352
rect 14752 19122 14780 19343
rect 14660 19094 14780 19122
rect 14556 17740 14608 17746
rect 14556 17682 14608 17688
rect 14660 17610 14688 19094
rect 14817 19068 15113 19088
rect 14873 19066 14897 19068
rect 14953 19066 14977 19068
rect 15033 19066 15057 19068
rect 14895 19014 14897 19066
rect 14959 19014 14971 19066
rect 15033 19014 15035 19066
rect 14873 19012 14897 19014
rect 14953 19012 14977 19014
rect 15033 19012 15057 19014
rect 14817 18992 15113 19012
rect 15212 18834 15240 19858
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 15200 18352 15252 18358
rect 15304 18340 15332 20046
rect 15396 19990 15424 22200
rect 15948 19990 15976 22200
rect 16396 20528 16448 20534
rect 16396 20470 16448 20476
rect 16120 20324 16172 20330
rect 16120 20266 16172 20272
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15936 19984 15988 19990
rect 15936 19926 15988 19932
rect 16132 19446 16160 20266
rect 16408 19990 16436 20470
rect 16500 20074 16528 22200
rect 16672 20324 16724 20330
rect 16672 20266 16724 20272
rect 16500 20046 16620 20074
rect 16592 19990 16620 20046
rect 16396 19984 16448 19990
rect 16396 19926 16448 19932
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16684 19786 16712 20266
rect 17052 19990 17080 22200
rect 17696 20534 17724 22200
rect 17958 22199 18014 22208
rect 18234 22200 18290 23000
rect 18786 22200 18842 23000
rect 19246 22672 19302 22681
rect 19246 22607 19302 22616
rect 17972 20534 18000 22199
rect 18248 20890 18276 22200
rect 18602 21720 18658 21729
rect 18602 21655 18658 21664
rect 18156 20862 18276 20890
rect 18156 20602 18184 20862
rect 18282 20700 18578 20720
rect 18338 20698 18362 20700
rect 18418 20698 18442 20700
rect 18498 20698 18522 20700
rect 18360 20646 18362 20698
rect 18424 20646 18436 20698
rect 18498 20646 18500 20698
rect 18338 20644 18362 20646
rect 18418 20644 18442 20646
rect 18498 20644 18522 20646
rect 18282 20624 18578 20644
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18616 20534 18644 21655
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17960 20528 18012 20534
rect 17960 20470 18012 20476
rect 18604 20528 18656 20534
rect 18604 20470 18656 20476
rect 18800 20466 18828 22200
rect 18970 21312 19026 21321
rect 18970 21247 19026 21256
rect 18984 20534 19012 21247
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17960 20324 18012 20330
rect 17960 20266 18012 20272
rect 18788 20324 18840 20330
rect 18788 20266 18840 20272
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17040 19984 17092 19990
rect 17040 19926 17092 19932
rect 16948 19916 17000 19922
rect 16948 19858 17000 19864
rect 16672 19780 16724 19786
rect 16672 19722 16724 19728
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16580 19168 16632 19174
rect 16580 19110 16632 19116
rect 16592 18970 16620 19110
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16672 18964 16724 18970
rect 16672 18906 16724 18912
rect 15384 18896 15436 18902
rect 16684 18850 16712 18906
rect 15384 18838 15436 18844
rect 15252 18312 15332 18340
rect 15200 18294 15252 18300
rect 15292 18216 15344 18222
rect 15396 18204 15424 18838
rect 16132 18822 16712 18850
rect 15936 18692 15988 18698
rect 15936 18634 15988 18640
rect 15948 18222 15976 18634
rect 15344 18176 15424 18204
rect 15292 18158 15344 18164
rect 14740 18148 14792 18154
rect 14740 18090 14792 18096
rect 14648 17604 14700 17610
rect 14648 17546 14700 17552
rect 14554 17504 14610 17513
rect 14554 17439 14610 17448
rect 14568 17338 14596 17439
rect 14752 17338 14780 18090
rect 14817 17980 15113 18000
rect 14873 17978 14897 17980
rect 14953 17978 14977 17980
rect 15033 17978 15057 17980
rect 14895 17926 14897 17978
rect 14959 17926 14971 17978
rect 15033 17926 15035 17978
rect 14873 17924 14897 17926
rect 14953 17924 14977 17926
rect 15033 17924 15057 17926
rect 14817 17904 15113 17924
rect 15200 17808 15252 17814
rect 15198 17776 15200 17785
rect 15396 17785 15424 18176
rect 15936 18216 15988 18222
rect 16028 18216 16080 18222
rect 15936 18158 15988 18164
rect 16026 18184 16028 18193
rect 16080 18184 16082 18193
rect 15752 18148 15804 18154
rect 16026 18119 16082 18128
rect 15752 18090 15804 18096
rect 15252 17776 15254 17785
rect 15382 17776 15438 17785
rect 15198 17711 15254 17720
rect 15292 17740 15344 17746
rect 15382 17711 15438 17720
rect 15292 17682 15344 17688
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14740 17332 14792 17338
rect 14740 17274 14792 17280
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14556 16652 14608 16658
rect 14556 16594 14608 16600
rect 14462 16552 14518 16561
rect 14462 16487 14518 16496
rect 14476 16114 14504 16487
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14476 15366 14504 16050
rect 14464 15360 14516 15366
rect 14464 15302 14516 15308
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14476 13870 14504 14350
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14476 12918 14504 13806
rect 14568 13802 14596 16594
rect 14752 16590 14780 17138
rect 15028 17066 15056 17546
rect 15016 17060 15068 17066
rect 15016 17002 15068 17008
rect 14817 16892 15113 16912
rect 14873 16890 14897 16892
rect 14953 16890 14977 16892
rect 15033 16890 15057 16892
rect 14895 16838 14897 16890
rect 14959 16838 14971 16890
rect 15033 16838 15035 16890
rect 14873 16836 14897 16838
rect 14953 16836 14977 16838
rect 15033 16836 15057 16838
rect 14817 16816 15113 16836
rect 14924 16652 14976 16658
rect 14844 16612 14924 16640
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14844 16232 14872 16612
rect 14924 16594 14976 16600
rect 15016 16584 15068 16590
rect 15212 16561 15240 17614
rect 15304 16794 15332 17682
rect 15396 17678 15424 17711
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15382 17368 15438 17377
rect 15488 17338 15516 17478
rect 15382 17303 15438 17312
rect 15476 17332 15528 17338
rect 15396 17202 15424 17303
rect 15476 17274 15528 17280
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15568 17060 15620 17066
rect 15568 17002 15620 17008
rect 15580 16794 15608 17002
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15016 16526 15068 16532
rect 15198 16552 15254 16561
rect 14660 16204 14872 16232
rect 14660 14346 14688 16204
rect 15028 16114 15056 16526
rect 15198 16487 15254 16496
rect 15476 16516 15528 16522
rect 15476 16458 15528 16464
rect 15488 16250 15516 16458
rect 15764 16250 15792 18090
rect 15842 16416 15898 16425
rect 15842 16351 15898 16360
rect 15476 16244 15528 16250
rect 15476 16186 15528 16192
rect 15752 16244 15804 16250
rect 15752 16186 15804 16192
rect 15568 16176 15620 16182
rect 15568 16118 15620 16124
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 14752 15094 14780 16050
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 14817 15804 15113 15824
rect 14873 15802 14897 15804
rect 14953 15802 14977 15804
rect 15033 15802 15057 15804
rect 14895 15750 14897 15802
rect 14959 15750 14971 15802
rect 15033 15750 15035 15802
rect 14873 15748 14897 15750
rect 14953 15748 14977 15750
rect 15033 15748 15057 15750
rect 14817 15728 15113 15748
rect 15304 15706 15332 15846
rect 15292 15700 15344 15706
rect 15292 15642 15344 15648
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 15120 14958 15148 15302
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 14817 14716 15113 14736
rect 14873 14714 14897 14716
rect 14953 14714 14977 14716
rect 15033 14714 15057 14716
rect 14895 14662 14897 14714
rect 14959 14662 14971 14714
rect 15033 14662 15035 14714
rect 14873 14660 14897 14662
rect 14953 14660 14977 14662
rect 15033 14660 15057 14662
rect 14817 14640 15113 14660
rect 15212 14346 15240 15438
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 14556 13796 14608 13802
rect 14556 13738 14608 13744
rect 15200 13796 15252 13802
rect 15200 13738 15252 13744
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14464 12912 14516 12918
rect 14464 12854 14516 12860
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14370 12064 14426 12073
rect 14370 11999 14426 12008
rect 14476 11898 14504 12718
rect 14556 12436 14608 12442
rect 14556 12378 14608 12384
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14200 11750 14320 11778
rect 14462 11792 14518 11801
rect 14096 11620 14148 11626
rect 14096 11562 14148 11568
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13556 9722 13584 9998
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13268 9590 13320 9596
rect 13358 9616 13414 9625
rect 13280 9382 13308 9590
rect 13358 9551 13414 9560
rect 13450 9480 13506 9489
rect 13450 9415 13506 9424
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 12808 8832 12860 8838
rect 12808 8774 12860 8780
rect 12452 8214 12572 8242
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12360 7585 12388 8026
rect 12346 7576 12402 7585
rect 12256 7540 12308 7546
rect 12346 7511 12402 7520
rect 12256 7482 12308 7488
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12254 6760 12310 6769
rect 12254 6695 12310 6704
rect 12268 5817 12296 6695
rect 12360 6186 12388 6938
rect 12452 6934 12480 8214
rect 12530 8120 12586 8129
rect 12820 8106 12848 8774
rect 12898 8392 12954 8401
rect 12898 8327 12900 8336
rect 12952 8327 12954 8336
rect 12900 8298 12952 8304
rect 12530 8055 12586 8064
rect 12728 8078 12848 8106
rect 12544 7886 12572 8055
rect 12532 7880 12584 7886
rect 12532 7822 12584 7828
rect 12544 7342 12572 7822
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12530 6488 12586 6497
rect 12530 6423 12586 6432
rect 12544 6225 12572 6423
rect 12530 6216 12586 6225
rect 12348 6180 12400 6186
rect 12530 6151 12586 6160
rect 12348 6122 12400 6128
rect 12254 5808 12310 5817
rect 12254 5743 12310 5752
rect 12360 5692 12388 6122
rect 12636 6118 12664 6802
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12636 5778 12664 5850
rect 12624 5772 12676 5778
rect 12624 5714 12676 5720
rect 12268 5664 12388 5692
rect 12532 5704 12584 5710
rect 12268 3942 12296 5664
rect 12532 5646 12584 5652
rect 12440 5636 12492 5642
rect 12440 5578 12492 5584
rect 12452 5545 12480 5578
rect 12438 5536 12494 5545
rect 12438 5471 12494 5480
rect 12544 5386 12572 5646
rect 12360 5358 12572 5386
rect 12360 4146 12388 5358
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12256 3936 12308 3942
rect 12256 3878 12308 3884
rect 12162 3768 12218 3777
rect 12162 3703 12218 3712
rect 12346 3632 12402 3641
rect 12452 3602 12480 4626
rect 12544 4146 12572 5170
rect 12636 5030 12664 5714
rect 12624 5024 12676 5030
rect 12624 4966 12676 4972
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12346 3567 12402 3576
rect 12440 3596 12492 3602
rect 12360 3534 12388 3567
rect 12440 3538 12492 3544
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 12624 3460 12676 3466
rect 12624 3402 12676 3408
rect 11796 3392 11848 3398
rect 11980 3392 12032 3398
rect 11848 3340 11928 3346
rect 11796 3334 11928 3340
rect 11980 3334 12032 3340
rect 12070 3360 12126 3369
rect 11808 3318 11928 3334
rect 11794 3224 11850 3233
rect 11794 3159 11850 3168
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11716 2582 11744 2790
rect 11808 2689 11836 3159
rect 11900 2904 11928 3318
rect 12070 3295 12126 3304
rect 12084 3097 12112 3295
rect 12070 3088 12126 3097
rect 12070 3023 12126 3032
rect 12530 2952 12586 2961
rect 12256 2916 12308 2922
rect 11900 2876 12256 2904
rect 12530 2887 12586 2896
rect 12256 2858 12308 2864
rect 12544 2774 12572 2887
rect 12452 2746 12572 2774
rect 11794 2680 11850 2689
rect 11794 2615 11850 2624
rect 11704 2576 11756 2582
rect 12452 2553 12480 2746
rect 11704 2518 11756 2524
rect 12438 2544 12494 2553
rect 10876 2508 10928 2514
rect 12438 2479 12494 2488
rect 10876 2450 10928 2456
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10336 1822 10640 1850
rect 10336 800 10364 1822
rect 10888 800 10916 2450
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12072 2372 12124 2378
rect 12072 2314 12124 2320
rect 11352 2204 11648 2224
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11430 2150 11432 2202
rect 11494 2150 11506 2202
rect 11568 2150 11570 2202
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11352 2128 11648 2148
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11440 800 11468 1906
rect 12084 800 12112 2314
rect 12268 2106 12296 2382
rect 12256 2100 12308 2106
rect 12256 2042 12308 2048
rect 12636 800 12664 3402
rect 12728 2378 12756 8078
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12820 6866 12848 7278
rect 13372 7274 13400 9318
rect 13464 8634 13492 9415
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13740 8634 13768 8910
rect 13832 8634 13860 10542
rect 13924 10266 13952 10662
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 14004 10464 14056 10470
rect 14108 10452 14136 11562
rect 14200 11234 14228 11750
rect 14568 11762 14596 12378
rect 14462 11727 14518 11736
rect 14556 11756 14608 11762
rect 14280 11688 14332 11694
rect 14280 11630 14332 11636
rect 14372 11688 14424 11694
rect 14372 11630 14424 11636
rect 14292 11354 14320 11630
rect 14280 11348 14332 11354
rect 14280 11290 14332 11296
rect 14200 11206 14320 11234
rect 14056 10424 14136 10452
rect 14004 10406 14056 10412
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14004 9376 14056 9382
rect 14004 9318 14056 9324
rect 14016 9178 14044 9318
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14004 8968 14056 8974
rect 14004 8910 14056 8916
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13740 8022 13768 8570
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13726 7712 13782 7721
rect 13726 7647 13782 7656
rect 13542 7304 13598 7313
rect 12992 7268 13044 7274
rect 12992 7210 13044 7216
rect 13360 7268 13412 7274
rect 13542 7239 13598 7248
rect 13360 7210 13412 7216
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12820 5914 12848 6802
rect 12900 6724 12952 6730
rect 12900 6666 12952 6672
rect 12912 5953 12940 6666
rect 13004 6390 13032 7210
rect 13084 7200 13136 7206
rect 13084 7142 13136 7148
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12990 6216 13046 6225
rect 12990 6151 13046 6160
rect 12898 5944 12954 5953
rect 12808 5908 12860 5914
rect 13004 5914 13032 6151
rect 13096 5914 13124 7142
rect 13176 6928 13228 6934
rect 13176 6870 13228 6876
rect 13188 6390 13216 6870
rect 13372 6730 13400 7210
rect 13556 7002 13584 7239
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13176 6384 13228 6390
rect 13176 6326 13228 6332
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12898 5879 12954 5888
rect 12992 5908 13044 5914
rect 12808 5850 12860 5856
rect 12992 5850 13044 5856
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13188 5710 13216 6054
rect 13280 5778 13308 6598
rect 13360 6452 13412 6458
rect 13360 6394 13412 6400
rect 13372 5794 13400 6394
rect 13464 6322 13492 6598
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13648 5914 13676 7142
rect 13740 6254 13768 7647
rect 13832 7342 13860 8570
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13924 7410 13952 7686
rect 13912 7404 13964 7410
rect 13912 7346 13964 7352
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13818 7032 13874 7041
rect 13818 6967 13874 6976
rect 13832 6866 13860 6967
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13924 6798 13952 7346
rect 13912 6792 13964 6798
rect 13912 6734 13964 6740
rect 13728 6248 13780 6254
rect 13728 6190 13780 6196
rect 13924 6186 13952 6734
rect 13912 6180 13964 6186
rect 13912 6122 13964 6128
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13728 5908 13780 5914
rect 13728 5850 13780 5856
rect 13740 5794 13768 5850
rect 13268 5772 13320 5778
rect 13372 5766 13768 5794
rect 13268 5714 13320 5720
rect 13176 5704 13228 5710
rect 13176 5646 13228 5652
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12820 4049 12848 5238
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 5030 13124 5102
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12806 4040 12862 4049
rect 12806 3975 12862 3984
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12820 3194 12848 3538
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 13096 2990 13124 4966
rect 13176 4548 13228 4554
rect 13176 4490 13228 4496
rect 13084 2984 13136 2990
rect 13084 2926 13136 2932
rect 12716 2372 12768 2378
rect 12716 2314 12768 2320
rect 12992 2304 13044 2310
rect 12992 2246 13044 2252
rect 13004 1562 13032 2246
rect 12992 1556 13044 1562
rect 12992 1498 13044 1504
rect 13188 800 13216 4490
rect 13464 4486 13492 5034
rect 13912 4684 13964 4690
rect 13912 4626 13964 4632
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13464 4146 13492 4422
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13280 3194 13308 3470
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 1834 13584 2246
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13740 800 13768 4490
rect 13820 4072 13872 4078
rect 13820 4014 13872 4020
rect 13832 3913 13860 4014
rect 13818 3904 13874 3913
rect 13818 3839 13874 3848
rect 13924 2922 13952 4626
rect 14016 4026 14044 8910
rect 14108 6798 14136 10424
rect 14188 10464 14240 10470
rect 14188 10406 14240 10412
rect 14200 10266 14228 10406
rect 14188 10260 14240 10266
rect 14188 10202 14240 10208
rect 14292 10146 14320 11206
rect 14384 11014 14412 11630
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10713 14412 10950
rect 14370 10704 14426 10713
rect 14370 10639 14426 10648
rect 14384 10198 14412 10639
rect 14200 10118 14320 10146
rect 14372 10192 14424 10198
rect 14372 10134 14424 10140
rect 14200 8514 14228 10118
rect 14280 9376 14332 9382
rect 14280 9318 14332 9324
rect 14292 8634 14320 9318
rect 14384 9042 14412 10134
rect 14372 9036 14424 9042
rect 14372 8978 14424 8984
rect 14476 8974 14504 11727
rect 14556 11698 14608 11704
rect 14660 11626 14688 13330
rect 14752 12782 14780 13670
rect 14817 13628 15113 13648
rect 14873 13626 14897 13628
rect 14953 13626 14977 13628
rect 15033 13626 15057 13628
rect 14895 13574 14897 13626
rect 14959 13574 14971 13626
rect 15033 13574 15035 13626
rect 14873 13572 14897 13574
rect 14953 13572 14977 13574
rect 15033 13572 15057 13574
rect 14817 13552 15113 13572
rect 15014 12880 15070 12889
rect 15014 12815 15070 12824
rect 15028 12782 15056 12815
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14817 12540 15113 12560
rect 14873 12538 14897 12540
rect 14953 12538 14977 12540
rect 15033 12538 15057 12540
rect 14895 12486 14897 12538
rect 14959 12486 14971 12538
rect 15033 12486 15035 12538
rect 14873 12484 14897 12486
rect 14953 12484 14977 12486
rect 15033 12484 15057 12486
rect 14817 12464 15113 12484
rect 15212 12345 15240 13738
rect 15304 12986 15332 15506
rect 15382 14784 15438 14793
rect 15382 14719 15438 14728
rect 15396 14550 15424 14719
rect 15384 14544 15436 14550
rect 15384 14486 15436 14492
rect 15384 14340 15436 14346
rect 15384 14282 15436 14288
rect 15396 13938 15424 14282
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15198 12336 15254 12345
rect 15198 12271 15254 12280
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14648 11620 14700 11626
rect 14648 11562 14700 11568
rect 14752 11558 14780 12174
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14568 9994 14596 11494
rect 14817 11452 15113 11472
rect 14873 11450 14897 11452
rect 14953 11450 14977 11452
rect 15033 11450 15057 11452
rect 14895 11398 14897 11450
rect 14959 11398 14971 11450
rect 15033 11398 15035 11450
rect 14873 11396 14897 11398
rect 14953 11396 14977 11398
rect 15033 11396 15057 11398
rect 14817 11376 15113 11396
rect 14648 10600 14700 10606
rect 14648 10542 14700 10548
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14660 9722 14688 10542
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14556 9580 14608 9586
rect 14556 9522 14608 9528
rect 14568 9178 14596 9522
rect 14752 9432 14780 10406
rect 14817 10364 15113 10384
rect 14873 10362 14897 10364
rect 14953 10362 14977 10364
rect 15033 10362 15057 10364
rect 14895 10310 14897 10362
rect 14959 10310 14971 10362
rect 15033 10310 15035 10362
rect 14873 10308 14897 10310
rect 14953 10308 14977 10310
rect 15033 10308 15057 10310
rect 14817 10288 15113 10308
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15028 9654 15056 9998
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15108 9444 15160 9450
rect 14752 9404 15108 9432
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14464 8968 14516 8974
rect 14464 8910 14516 8916
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 14384 8634 14412 8842
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14200 8486 14320 8514
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14200 5642 14228 7142
rect 14292 6633 14320 8486
rect 14476 8430 14504 8774
rect 14752 8537 14780 9404
rect 15108 9386 15160 9392
rect 14817 9276 15113 9296
rect 14873 9274 14897 9276
rect 14953 9274 14977 9276
rect 15033 9274 15057 9276
rect 14895 9222 14897 9274
rect 14959 9222 14971 9274
rect 15033 9222 15035 9274
rect 14873 9220 14897 9222
rect 14953 9220 14977 9222
rect 15033 9220 15057 9222
rect 14817 9200 15113 9220
rect 14832 9036 14884 9042
rect 14832 8978 14884 8984
rect 14738 8528 14794 8537
rect 14648 8492 14700 8498
rect 14844 8498 14872 8978
rect 14738 8463 14794 8472
rect 14832 8492 14884 8498
rect 14648 8434 14700 8440
rect 14832 8434 14884 8440
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 14476 8022 14504 8366
rect 14556 8288 14608 8294
rect 14554 8256 14556 8265
rect 14608 8256 14610 8265
rect 14554 8191 14610 8200
rect 14660 8090 14688 8434
rect 14832 8356 14884 8362
rect 14752 8316 14832 8344
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14464 7472 14516 7478
rect 14464 7414 14516 7420
rect 14476 6633 14504 7414
rect 14752 6866 14780 8316
rect 14832 8298 14884 8304
rect 14817 8188 15113 8208
rect 14873 8186 14897 8188
rect 14953 8186 14977 8188
rect 15033 8186 15057 8188
rect 14895 8134 14897 8186
rect 14959 8134 14971 8186
rect 15033 8134 15035 8186
rect 14873 8132 14897 8134
rect 14953 8132 14977 8134
rect 15033 8132 15057 8134
rect 14817 8112 15113 8132
rect 15212 8072 15240 12271
rect 15488 11694 15516 15846
rect 15580 14890 15608 16118
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15672 15609 15700 15982
rect 15658 15600 15714 15609
rect 15658 15535 15714 15544
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15672 14414 15700 15535
rect 15752 15360 15804 15366
rect 15752 15302 15804 15308
rect 15764 14822 15792 15302
rect 15856 14958 15884 16351
rect 16132 15910 16160 18822
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 16304 18624 16356 18630
rect 16304 18566 16356 18572
rect 16212 17536 16264 17542
rect 16212 17478 16264 17484
rect 16224 16794 16252 17478
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16212 16584 16264 16590
rect 16212 16526 16264 16532
rect 16224 16017 16252 16526
rect 16316 16522 16344 18566
rect 16684 18426 16712 18702
rect 16672 18420 16724 18426
rect 16672 18362 16724 18368
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16488 17808 16540 17814
rect 16488 17750 16540 17756
rect 16500 17202 16528 17750
rect 16592 17746 16620 18022
rect 16580 17740 16632 17746
rect 16580 17682 16632 17688
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16488 17196 16540 17202
rect 16488 17138 16540 17144
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16794 16528 16934
rect 16868 16794 16896 17274
rect 16488 16788 16540 16794
rect 16488 16730 16540 16736
rect 16856 16788 16908 16794
rect 16856 16730 16908 16736
rect 16304 16516 16356 16522
rect 16304 16458 16356 16464
rect 16210 16008 16266 16017
rect 16210 15943 16266 15952
rect 16224 15910 16252 15943
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 16132 15502 16160 15846
rect 16224 15570 16252 15846
rect 16960 15706 16988 19858
rect 17236 19514 17264 20198
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17224 19508 17276 19514
rect 17224 19450 17276 19456
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 17052 18465 17080 19246
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17038 18456 17094 18465
rect 17038 18391 17094 18400
rect 17224 18284 17276 18290
rect 17224 18226 17276 18232
rect 17236 17785 17264 18226
rect 17222 17776 17278 17785
rect 17040 17740 17092 17746
rect 17222 17711 17224 17720
rect 17040 17682 17092 17688
rect 17276 17711 17278 17720
rect 17224 17682 17276 17688
rect 17052 17202 17080 17682
rect 17222 17504 17278 17513
rect 17222 17439 17278 17448
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 17196 17092 17202
rect 17040 17138 17092 17144
rect 17052 16590 17080 17138
rect 17040 16584 17092 16590
rect 17040 16526 17092 16532
rect 17144 16250 17172 17206
rect 17236 17066 17264 17439
rect 17224 17060 17276 17066
rect 17224 17002 17276 17008
rect 17132 16244 17184 16250
rect 17132 16186 17184 16192
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 16948 15700 17000 15706
rect 16948 15642 17000 15648
rect 16856 15632 16908 15638
rect 16856 15574 16908 15580
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16120 15496 16172 15502
rect 16026 15464 16082 15473
rect 15936 15428 15988 15434
rect 16580 15496 16632 15502
rect 16172 15444 16252 15450
rect 16120 15438 16252 15444
rect 16580 15438 16632 15444
rect 16026 15399 16082 15408
rect 16132 15422 16252 15438
rect 15936 15370 15988 15376
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15752 14816 15804 14822
rect 15752 14758 15804 14764
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15660 14408 15712 14414
rect 15856 14385 15884 14758
rect 15660 14350 15712 14356
rect 15842 14376 15898 14385
rect 15842 14311 15898 14320
rect 15844 13728 15896 13734
rect 15844 13670 15896 13676
rect 15856 13530 15884 13670
rect 15844 13524 15896 13530
rect 15844 13466 15896 13472
rect 15844 12708 15896 12714
rect 15844 12650 15896 12656
rect 15856 12434 15884 12650
rect 15672 12406 15884 12434
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15304 10441 15332 10474
rect 15290 10432 15346 10441
rect 15290 10367 15346 10376
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9081 15332 9318
rect 15290 9072 15346 9081
rect 15396 9042 15424 9522
rect 15672 9382 15700 12406
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15764 11558 15792 11698
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 10742 15884 11494
rect 15844 10736 15896 10742
rect 15844 10678 15896 10684
rect 15948 10266 15976 15370
rect 16040 15366 16068 15399
rect 16132 15373 16160 15422
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16224 15026 16252 15422
rect 16592 15094 16620 15438
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16672 15088 16724 15094
rect 16672 15030 16724 15036
rect 16212 15020 16264 15026
rect 16132 14980 16212 15008
rect 16132 14482 16160 14980
rect 16212 14962 16264 14968
rect 16212 14884 16264 14890
rect 16212 14826 16264 14832
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 16028 14000 16080 14006
rect 16028 13942 16080 13948
rect 16040 13326 16068 13942
rect 16224 13802 16252 14826
rect 16684 14618 16712 15030
rect 16672 14612 16724 14618
rect 16672 14554 16724 14560
rect 16488 14476 16540 14482
rect 16488 14418 16540 14424
rect 16500 14006 16528 14418
rect 16488 14000 16540 14006
rect 16488 13942 16540 13948
rect 16304 13864 16356 13870
rect 16304 13806 16356 13812
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16212 12844 16264 12850
rect 16212 12786 16264 12792
rect 16120 12640 16172 12646
rect 16120 12582 16172 12588
rect 16132 11354 16160 12582
rect 16224 12238 16252 12786
rect 16316 12442 16344 13806
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16408 13530 16436 13738
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16580 13252 16632 13258
rect 16580 13194 16632 13200
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16592 12345 16620 13194
rect 16762 13152 16818 13161
rect 16762 13087 16818 13096
rect 16776 12646 16804 13087
rect 16764 12640 16816 12646
rect 16764 12582 16816 12588
rect 16578 12336 16634 12345
rect 16578 12271 16580 12280
rect 16632 12271 16634 12280
rect 16580 12242 16632 12248
rect 16212 12232 16264 12238
rect 16592 12211 16620 12242
rect 16212 12174 16264 12180
rect 16580 12096 16632 12102
rect 16580 12038 16632 12044
rect 16488 11892 16540 11898
rect 16488 11834 16540 11840
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16132 11234 16160 11290
rect 16132 11206 16252 11234
rect 16316 11218 16344 11766
rect 16500 11354 16528 11834
rect 16488 11348 16540 11354
rect 16488 11290 16540 11296
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9722 16068 9998
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 15660 9376 15712 9382
rect 15660 9318 15712 9324
rect 16120 9376 16172 9382
rect 16120 9318 16172 9324
rect 15474 9072 15530 9081
rect 15290 9007 15346 9016
rect 15384 9036 15436 9042
rect 15474 9007 15530 9016
rect 15568 9036 15620 9042
rect 15384 8978 15436 8984
rect 15212 8044 15424 8072
rect 15198 7984 15254 7993
rect 15198 7919 15254 7928
rect 15212 7177 15240 7919
rect 15198 7168 15254 7177
rect 14817 7100 15113 7120
rect 15198 7103 15254 7112
rect 14873 7098 14897 7100
rect 14953 7098 14977 7100
rect 15033 7098 15057 7100
rect 14895 7046 14897 7098
rect 14959 7046 14971 7098
rect 15033 7046 15035 7098
rect 14873 7044 14897 7046
rect 14953 7044 14977 7046
rect 15033 7044 15057 7046
rect 14817 7024 15113 7044
rect 14740 6860 14792 6866
rect 14740 6802 14792 6808
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 14462 6624 14518 6633
rect 14462 6559 14518 6568
rect 14372 6248 14424 6254
rect 14372 6190 14424 6196
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 14384 5166 14412 6190
rect 14556 6180 14608 6186
rect 14556 6122 14608 6128
rect 14568 6089 14596 6122
rect 14554 6080 14610 6089
rect 14554 6015 14610 6024
rect 14752 5778 14780 6802
rect 15106 6760 15162 6769
rect 15212 6746 15240 6802
rect 15162 6718 15240 6746
rect 15106 6695 15162 6704
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14844 6225 14872 6394
rect 14830 6216 14886 6225
rect 14830 6151 14886 6160
rect 15120 6168 15148 6695
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15120 6140 15240 6168
rect 14817 6012 15113 6032
rect 14873 6010 14897 6012
rect 14953 6010 14977 6012
rect 15033 6010 15057 6012
rect 14895 5958 14897 6010
rect 14959 5958 14971 6010
rect 15033 5958 15035 6010
rect 14873 5956 14897 5958
rect 14953 5956 14977 5958
rect 15033 5956 15057 5958
rect 14817 5936 15113 5956
rect 15212 5778 15240 6140
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 15200 5772 15252 5778
rect 15200 5714 15252 5720
rect 15304 5710 15332 6258
rect 15292 5704 15344 5710
rect 15396 5692 15424 8044
rect 15488 7478 15516 9007
rect 15568 8978 15620 8984
rect 15580 8498 15608 8978
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15764 7954 15792 8434
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15752 7948 15804 7954
rect 15752 7890 15804 7896
rect 15764 7546 15792 7890
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15476 7472 15528 7478
rect 15476 7414 15528 7420
rect 16040 6730 16068 8298
rect 16132 6934 16160 9318
rect 16224 9160 16252 11206
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16592 10606 16620 12038
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 9586 16712 10406
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16304 9172 16356 9178
rect 16224 9132 16304 9160
rect 16304 9114 16356 9120
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16316 7546 16344 7822
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 16120 6928 16172 6934
rect 16120 6870 16172 6876
rect 16224 6866 16252 7278
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16028 6724 16080 6730
rect 16028 6666 16080 6672
rect 16316 6322 16344 7482
rect 16408 7002 16436 7822
rect 16486 7304 16542 7313
rect 16486 7239 16542 7248
rect 16500 7002 16528 7239
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16488 6996 16540 7002
rect 16488 6938 16540 6944
rect 15936 6316 15988 6322
rect 15936 6258 15988 6264
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15476 6112 15528 6118
rect 15476 6054 15528 6060
rect 15488 5846 15516 6054
rect 15476 5840 15528 5846
rect 15476 5782 15528 5788
rect 15566 5808 15622 5817
rect 15566 5743 15568 5752
rect 15620 5743 15622 5752
rect 15568 5714 15620 5720
rect 15396 5664 15516 5692
rect 15292 5646 15344 5652
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14372 5160 14424 5166
rect 14372 5102 14424 5108
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14660 4758 14688 5102
rect 14752 4758 14780 5510
rect 15304 5166 15332 5646
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 14817 4924 15113 4944
rect 14873 4922 14897 4924
rect 14953 4922 14977 4924
rect 15033 4922 15057 4924
rect 14895 4870 14897 4922
rect 14959 4870 14971 4922
rect 15033 4870 15035 4922
rect 14873 4868 14897 4870
rect 14953 4868 14977 4870
rect 15033 4868 15057 4870
rect 14817 4848 15113 4868
rect 14372 4752 14424 4758
rect 14372 4694 14424 4700
rect 14648 4752 14700 4758
rect 14648 4694 14700 4700
rect 14740 4752 14792 4758
rect 14740 4694 14792 4700
rect 14280 4072 14332 4078
rect 14016 3998 14136 4026
rect 14280 4014 14332 4020
rect 14004 3936 14056 3942
rect 14004 3878 14056 3884
rect 14016 3738 14044 3878
rect 14004 3732 14056 3738
rect 14004 3674 14056 3680
rect 14108 3534 14136 3998
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 3210 14136 3470
rect 14108 3194 14228 3210
rect 14108 3188 14240 3194
rect 14108 3182 14188 3188
rect 14108 2961 14136 3182
rect 14188 3130 14240 3136
rect 14094 2952 14150 2961
rect 13912 2916 13964 2922
rect 14094 2887 14150 2896
rect 13912 2858 13964 2864
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 2106 14136 2246
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 14292 800 14320 4014
rect 14384 3602 14412 4694
rect 14660 4593 14688 4694
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 14556 4140 14608 4146
rect 14556 4082 14608 4088
rect 14372 3596 14424 3602
rect 14372 3538 14424 3544
rect 14384 2990 14412 3538
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14568 2650 14596 4082
rect 14648 4004 14700 4010
rect 14648 3946 14700 3952
rect 14660 3670 14688 3946
rect 14648 3664 14700 3670
rect 14648 3606 14700 3612
rect 14660 3194 14688 3606
rect 14648 3188 14700 3194
rect 14648 3130 14700 3136
rect 14556 2644 14608 2650
rect 14556 2586 14608 2592
rect 14752 898 14780 4490
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 14817 3836 15113 3856
rect 14873 3834 14897 3836
rect 14953 3834 14977 3836
rect 15033 3834 15057 3836
rect 14895 3782 14897 3834
rect 14959 3782 14971 3834
rect 15033 3782 15035 3834
rect 14873 3780 14897 3782
rect 14953 3780 14977 3782
rect 15033 3780 15057 3782
rect 14817 3760 15113 3780
rect 15212 3074 15240 3946
rect 15120 3058 15240 3074
rect 15108 3052 15240 3058
rect 15160 3046 15240 3052
rect 15108 2994 15160 3000
rect 14817 2748 15113 2768
rect 14873 2746 14897 2748
rect 14953 2746 14977 2748
rect 15033 2746 15057 2748
rect 14895 2694 14897 2746
rect 14959 2694 14971 2746
rect 15033 2694 15035 2746
rect 14873 2692 14897 2694
rect 14953 2692 14977 2694
rect 15033 2692 15057 2694
rect 14817 2672 15113 2692
rect 15304 2417 15332 3946
rect 15290 2408 15346 2417
rect 15290 2343 15346 2352
rect 14752 870 14872 898
rect 14844 800 14872 870
rect 15396 800 15424 4490
rect 15488 3641 15516 5664
rect 15948 4622 15976 6258
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16224 5846 16252 6054
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15936 4616 15988 4622
rect 15934 4584 15936 4593
rect 15988 4584 15990 4593
rect 15934 4519 15990 4528
rect 16132 4128 16160 5578
rect 16212 4140 16264 4146
rect 16132 4100 16212 4128
rect 16212 4082 16264 4088
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15764 3738 15792 3878
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 15474 3632 15530 3641
rect 15474 3567 15530 3576
rect 15856 3369 15884 3674
rect 15936 3392 15988 3398
rect 15842 3360 15898 3369
rect 15936 3334 15988 3340
rect 15842 3295 15898 3304
rect 15856 2650 15884 3295
rect 15948 2990 15976 3334
rect 15936 2984 15988 2990
rect 15936 2926 15988 2932
rect 15844 2644 15896 2650
rect 15844 2586 15896 2592
rect 15948 2446 15976 2926
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 16040 1442 16068 3878
rect 16408 3602 16436 6054
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16500 5234 16528 5646
rect 16488 5228 16540 5234
rect 16488 5170 16540 5176
rect 16500 4758 16528 5170
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16316 3233 16344 3334
rect 16302 3224 16358 3233
rect 16302 3159 16358 3168
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16132 1902 16160 2450
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 15948 1414 16068 1442
rect 15948 800 15976 1414
rect 16500 800 16528 4082
rect 16592 3738 16620 9318
rect 16580 3732 16632 3738
rect 16580 3674 16632 3680
rect 16592 3618 16620 3674
rect 16592 3590 16712 3618
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16592 2650 16620 3470
rect 16684 3058 16712 3590
rect 16672 3052 16724 3058
rect 16672 2994 16724 3000
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16776 1970 16804 12582
rect 16868 12442 16896 15574
rect 17052 14770 17080 15846
rect 17328 15065 17356 18770
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17420 17134 17448 18158
rect 17512 17882 17540 19858
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17604 18601 17632 19246
rect 17696 18970 17724 20266
rect 17972 19174 18000 20266
rect 18800 20058 18828 20266
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18510 19952 18566 19961
rect 18510 19887 18512 19896
rect 18564 19887 18566 19896
rect 18604 19916 18656 19922
rect 18512 19858 18564 19864
rect 18604 19858 18656 19864
rect 18282 19612 18578 19632
rect 18338 19610 18362 19612
rect 18418 19610 18442 19612
rect 18498 19610 18522 19612
rect 18360 19558 18362 19610
rect 18424 19558 18436 19610
rect 18498 19558 18500 19610
rect 18338 19556 18362 19558
rect 18418 19556 18442 19558
rect 18498 19556 18522 19558
rect 18282 19536 18578 19556
rect 18616 19378 18644 19858
rect 18604 19372 18656 19378
rect 18604 19314 18656 19320
rect 19260 19310 19288 22607
rect 19338 22200 19394 23000
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
rect 19352 19990 19380 22200
rect 19522 20768 19578 20777
rect 19522 20703 19578 20712
rect 19536 20534 19564 20703
rect 19524 20528 19576 20534
rect 19524 20470 19576 20476
rect 19432 20324 19484 20330
rect 19432 20266 19484 20272
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 18420 19304 18472 19310
rect 18420 19246 18472 19252
rect 19064 19304 19116 19310
rect 19064 19246 19116 19252
rect 19248 19304 19300 19310
rect 19248 19246 19300 19252
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17684 18964 17736 18970
rect 17684 18906 17736 18912
rect 18432 18873 18460 19246
rect 18418 18864 18474 18873
rect 18052 18828 18104 18834
rect 18418 18799 18474 18808
rect 18052 18770 18104 18776
rect 17960 18760 18012 18766
rect 17960 18702 18012 18708
rect 17590 18592 17646 18601
rect 17590 18527 17646 18536
rect 17500 17876 17552 17882
rect 17500 17818 17552 17824
rect 17408 17128 17460 17134
rect 17408 17070 17460 17076
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16794 17540 16934
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17696 16046 17724 16730
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17684 16040 17736 16046
rect 17684 15982 17736 15988
rect 17880 15706 17908 16050
rect 17972 15978 18000 18702
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17314 15056 17370 15065
rect 17314 14991 17370 15000
rect 16960 14742 17080 14770
rect 17960 14816 18012 14822
rect 18064 14804 18092 18770
rect 18282 18524 18578 18544
rect 18338 18522 18362 18524
rect 18418 18522 18442 18524
rect 18498 18522 18522 18524
rect 18360 18470 18362 18522
rect 18424 18470 18436 18522
rect 18498 18470 18500 18522
rect 18338 18468 18362 18470
rect 18418 18468 18442 18470
rect 18498 18468 18522 18470
rect 18282 18448 18578 18468
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18892 17746 18920 18022
rect 18984 17882 19012 18090
rect 18972 17876 19024 17882
rect 18972 17818 19024 17824
rect 18144 17740 18196 17746
rect 18144 17682 18196 17688
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18156 17202 18184 17682
rect 18282 17436 18578 17456
rect 18338 17434 18362 17436
rect 18418 17434 18442 17436
rect 18498 17434 18522 17436
rect 18360 17382 18362 17434
rect 18424 17382 18436 17434
rect 18498 17382 18500 17434
rect 18338 17380 18362 17382
rect 18418 17380 18442 17382
rect 18498 17380 18522 17382
rect 18282 17360 18578 17380
rect 18602 17232 18658 17241
rect 18144 17196 18196 17202
rect 18602 17167 18658 17176
rect 18144 17138 18196 17144
rect 18156 16046 18184 17138
rect 18282 16348 18578 16368
rect 18338 16346 18362 16348
rect 18418 16346 18442 16348
rect 18498 16346 18522 16348
rect 18360 16294 18362 16346
rect 18424 16294 18436 16346
rect 18498 16294 18500 16346
rect 18338 16292 18362 16294
rect 18418 16292 18442 16294
rect 18498 16292 18522 16294
rect 18282 16272 18578 16292
rect 18144 16040 18196 16046
rect 18144 15982 18196 15988
rect 18616 15586 18644 17167
rect 18892 17134 18920 17682
rect 18984 17134 19012 17818
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18708 15706 18736 16594
rect 18696 15700 18748 15706
rect 18696 15642 18748 15648
rect 18616 15558 18736 15586
rect 18282 15260 18578 15280
rect 18338 15258 18362 15260
rect 18418 15258 18442 15260
rect 18498 15258 18522 15260
rect 18360 15206 18362 15258
rect 18424 15206 18436 15258
rect 18498 15206 18500 15258
rect 18338 15204 18362 15206
rect 18418 15204 18442 15206
rect 18498 15204 18522 15206
rect 18282 15184 18578 15204
rect 18012 14776 18092 14804
rect 17960 14758 18012 14764
rect 16960 13530 16988 14742
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 16868 8514 16896 12378
rect 16960 9382 16988 13466
rect 17040 13388 17092 13394
rect 17040 13330 17092 13336
rect 17132 13388 17184 13394
rect 17132 13330 17184 13336
rect 17052 12442 17080 13330
rect 17144 12850 17172 13330
rect 17132 12844 17184 12850
rect 17132 12786 17184 12792
rect 17040 12436 17092 12442
rect 17040 12378 17092 12384
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 17052 12209 17080 12242
rect 17144 12238 17172 12786
rect 17132 12232 17184 12238
rect 17038 12200 17094 12209
rect 17132 12174 17184 12180
rect 17038 12135 17094 12144
rect 17328 11898 17356 14554
rect 18144 14476 18196 14482
rect 18144 14418 18196 14424
rect 17868 14408 17920 14414
rect 17868 14350 17920 14356
rect 17960 14408 18012 14414
rect 17960 14350 18012 14356
rect 17880 14074 17908 14350
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17880 13954 17908 14010
rect 17788 13926 17908 13954
rect 17408 13456 17460 13462
rect 17592 13456 17644 13462
rect 17460 13404 17540 13410
rect 17408 13398 17540 13404
rect 17592 13398 17644 13404
rect 17682 13424 17738 13433
rect 17420 13382 17540 13398
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17052 10674 17080 11290
rect 17420 10674 17448 12718
rect 17040 10668 17092 10674
rect 17040 10610 17092 10616
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17328 10010 17356 10542
rect 17328 9982 17448 10010
rect 17420 9926 17448 9982
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 17052 9110 17080 9454
rect 17420 9450 17448 9862
rect 17408 9444 17460 9450
rect 17408 9386 17460 9392
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17420 9042 17448 9386
rect 17512 9178 17540 13382
rect 17604 12714 17632 13398
rect 17682 13359 17738 13368
rect 17696 12782 17724 13359
rect 17788 13326 17816 13926
rect 17868 13796 17920 13802
rect 17868 13738 17920 13744
rect 17776 13320 17828 13326
rect 17776 13262 17828 13268
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17592 12708 17644 12714
rect 17592 12650 17644 12656
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17408 9036 17460 9042
rect 17408 8978 17460 8984
rect 16868 8486 17080 8514
rect 16856 8424 16908 8430
rect 16856 8366 16908 8372
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 16868 1698 16896 8366
rect 17052 5114 17080 8486
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17328 7274 17356 7822
rect 17132 7268 17184 7274
rect 17132 7210 17184 7216
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17144 5302 17172 7210
rect 17328 6798 17356 7210
rect 17512 6866 17540 9114
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17604 7206 17632 8298
rect 17696 8090 17724 12718
rect 17788 12345 17816 13262
rect 17774 12336 17830 12345
rect 17880 12306 17908 13738
rect 17972 13258 18000 14350
rect 18156 14113 18184 14418
rect 18282 14172 18578 14192
rect 18338 14170 18362 14172
rect 18418 14170 18442 14172
rect 18498 14170 18522 14172
rect 18360 14118 18362 14170
rect 18424 14118 18436 14170
rect 18498 14118 18500 14170
rect 18338 14116 18362 14118
rect 18418 14116 18442 14118
rect 18498 14116 18522 14118
rect 18142 14104 18198 14113
rect 18282 14096 18578 14116
rect 18142 14039 18198 14048
rect 18144 13320 18196 13326
rect 18144 13262 18196 13268
rect 17960 13252 18012 13258
rect 17960 13194 18012 13200
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 12640 18012 12646
rect 17960 12582 18012 12588
rect 17774 12271 17830 12280
rect 17868 12300 17920 12306
rect 17868 12242 17920 12248
rect 17972 12238 18000 12582
rect 18064 12442 18092 13126
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18156 11558 18184 13262
rect 18282 13084 18578 13104
rect 18338 13082 18362 13084
rect 18418 13082 18442 13084
rect 18498 13082 18522 13084
rect 18360 13030 18362 13082
rect 18424 13030 18436 13082
rect 18498 13030 18500 13082
rect 18338 13028 18362 13030
rect 18418 13028 18442 13030
rect 18498 13028 18522 13030
rect 18282 13008 18578 13028
rect 18236 12368 18288 12374
rect 18234 12336 18236 12345
rect 18288 12336 18290 12345
rect 18234 12271 18290 12280
rect 18282 11996 18578 12016
rect 18338 11994 18362 11996
rect 18418 11994 18442 11996
rect 18498 11994 18522 11996
rect 18360 11942 18362 11994
rect 18424 11942 18436 11994
rect 18498 11942 18500 11994
rect 18338 11940 18362 11942
rect 18418 11940 18442 11942
rect 18498 11940 18522 11942
rect 18282 11920 18578 11940
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17880 11218 17908 11494
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17880 10810 17908 11154
rect 18156 11121 18184 11494
rect 18616 11354 18644 11630
rect 18604 11348 18656 11354
rect 18604 11290 18656 11296
rect 18142 11112 18198 11121
rect 18142 11047 18198 11056
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17972 10146 18000 10950
rect 18282 10908 18578 10928
rect 18338 10906 18362 10908
rect 18418 10906 18442 10908
rect 18498 10906 18522 10908
rect 18360 10854 18362 10906
rect 18424 10854 18436 10906
rect 18498 10854 18500 10906
rect 18338 10852 18362 10854
rect 18418 10852 18442 10854
rect 18498 10852 18522 10854
rect 18282 10832 18578 10852
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18248 10266 18276 10406
rect 18708 10266 18736 15558
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 18800 13870 18828 14214
rect 18788 13864 18840 13870
rect 18788 13806 18840 13812
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18892 12986 18920 13670
rect 19076 13297 19104 19246
rect 19260 18970 19288 19246
rect 19352 19174 19380 19790
rect 19444 19446 19472 20266
rect 19904 19990 19932 22200
rect 20456 20466 20484 22200
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20168 20392 20220 20398
rect 20168 20334 20220 20340
rect 20442 20360 20498 20369
rect 19892 19984 19944 19990
rect 19892 19926 19944 19932
rect 19616 19916 19668 19922
rect 19616 19858 19668 19864
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19248 18964 19300 18970
rect 19248 18906 19300 18912
rect 19156 18624 19208 18630
rect 19156 18566 19208 18572
rect 19524 18624 19576 18630
rect 19524 18566 19576 18572
rect 19168 18154 19196 18566
rect 19156 18148 19208 18154
rect 19156 18090 19208 18096
rect 19432 16992 19484 16998
rect 19432 16934 19484 16940
rect 19444 16590 19472 16934
rect 19536 16726 19564 18566
rect 19628 18329 19656 19858
rect 19708 19236 19760 19242
rect 19708 19178 19760 19184
rect 19984 19236 20036 19242
rect 19984 19178 20036 19184
rect 19614 18320 19670 18329
rect 19614 18255 19670 18264
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19432 16584 19484 16590
rect 19432 16526 19484 16532
rect 19340 15972 19392 15978
rect 19340 15914 19392 15920
rect 19352 15026 19380 15914
rect 19444 15638 19472 16526
rect 19524 16040 19576 16046
rect 19524 15982 19576 15988
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19444 14958 19472 15438
rect 19248 14952 19300 14958
rect 19432 14952 19484 14958
rect 19300 14900 19380 14906
rect 19248 14894 19380 14900
rect 19432 14894 19484 14900
rect 19260 14878 19380 14894
rect 19248 14816 19300 14822
rect 19246 14784 19248 14793
rect 19300 14784 19302 14793
rect 19246 14719 19302 14728
rect 19260 14006 19288 14719
rect 19352 14482 19380 14878
rect 19340 14476 19392 14482
rect 19340 14418 19392 14424
rect 19340 14272 19392 14278
rect 19340 14214 19392 14220
rect 19248 14000 19300 14006
rect 19248 13942 19300 13948
rect 19248 13728 19300 13734
rect 19248 13670 19300 13676
rect 19260 13530 19288 13670
rect 19248 13524 19300 13530
rect 19248 13466 19300 13472
rect 19062 13288 19118 13297
rect 19062 13223 19118 13232
rect 18880 12980 18932 12986
rect 18880 12922 18932 12928
rect 19154 12744 19210 12753
rect 19352 12730 19380 14214
rect 19444 13938 19472 14894
rect 19536 14890 19564 15982
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 19628 15706 19656 15846
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19616 15020 19668 15026
rect 19720 15008 19748 19178
rect 19892 18080 19944 18086
rect 19892 18022 19944 18028
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19812 16454 19840 17478
rect 19904 16794 19932 18022
rect 19892 16788 19944 16794
rect 19892 16730 19944 16736
rect 19890 16688 19946 16697
rect 19890 16623 19946 16632
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19668 14980 19748 15008
rect 19616 14962 19668 14968
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19904 14074 19932 16623
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19432 13932 19484 13938
rect 19432 13874 19484 13880
rect 19616 13932 19668 13938
rect 19616 13874 19668 13880
rect 19210 12702 19380 12730
rect 19444 12714 19472 13874
rect 19628 12782 19656 13874
rect 19708 13728 19760 13734
rect 19708 13670 19760 13676
rect 19720 12986 19748 13670
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19616 12776 19668 12782
rect 19616 12718 19668 12724
rect 19432 12708 19484 12714
rect 19154 12679 19210 12688
rect 19168 12442 19196 12679
rect 19432 12650 19484 12656
rect 19628 12442 19656 12718
rect 19156 12436 19208 12442
rect 19156 12378 19208 12384
rect 19616 12436 19668 12442
rect 19996 12434 20024 19178
rect 20076 18828 20128 18834
rect 20076 18770 20128 18776
rect 20088 18737 20116 18770
rect 20074 18728 20130 18737
rect 20074 18663 20130 18672
rect 20074 17640 20130 17649
rect 20074 17575 20130 17584
rect 20088 17202 20116 17575
rect 20076 17196 20128 17202
rect 20076 17138 20128 17144
rect 20180 17105 20208 20334
rect 20810 20360 20866 20369
rect 20442 20295 20498 20304
rect 20628 20324 20680 20330
rect 20456 18902 20484 20295
rect 20810 20295 20812 20304
rect 20628 20266 20680 20272
rect 20864 20295 20866 20304
rect 20812 20266 20864 20272
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 19281 20576 19858
rect 20640 19514 20668 20266
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20534 19272 20590 19281
rect 20534 19207 20590 19216
rect 21008 18902 21036 22200
rect 21180 20324 21232 20330
rect 21180 20266 21232 20272
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 21100 19310 21128 20198
rect 21088 19304 21140 19310
rect 21088 19246 21140 19252
rect 21088 19168 21140 19174
rect 21088 19110 21140 19116
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20996 18896 21048 18902
rect 20996 18838 21048 18844
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20272 18426 20300 18770
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20260 18420 20312 18426
rect 20260 18362 20312 18368
rect 20640 18222 20668 18634
rect 20628 18216 20680 18222
rect 20628 18158 20680 18164
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20628 18080 20680 18086
rect 20628 18022 20680 18028
rect 20272 17882 20300 18022
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20272 17338 20300 17614
rect 20640 17513 20668 18022
rect 20626 17504 20682 17513
rect 20626 17439 20682 17448
rect 20260 17332 20312 17338
rect 20260 17274 20312 17280
rect 21100 17134 21128 19110
rect 21088 17128 21140 17134
rect 20166 17096 20222 17105
rect 20076 17060 20128 17066
rect 21088 17070 21140 17076
rect 20166 17031 20222 17040
rect 20076 17002 20128 17008
rect 20088 13326 20116 17002
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16250 20208 16934
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 20168 16108 20220 16114
rect 20272 16096 20300 16390
rect 20352 16176 20404 16182
rect 20352 16118 20404 16124
rect 20220 16068 20300 16096
rect 20168 16050 20220 16056
rect 20180 13462 20208 16050
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 20272 13802 20300 15846
rect 20364 14958 20392 16118
rect 20352 14952 20404 14958
rect 20640 14929 20668 16594
rect 20812 16448 20864 16454
rect 21192 16402 21220 20266
rect 21468 19825 21496 20266
rect 21560 20058 21588 22200
rect 21548 20052 21600 20058
rect 21548 19994 21600 20000
rect 21454 19816 21510 19825
rect 21364 19780 21416 19786
rect 21454 19751 21510 19760
rect 21364 19722 21416 19728
rect 21376 19417 21404 19722
rect 22112 19718 22140 22200
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21364 19236 21416 19242
rect 21364 19178 21416 19184
rect 21376 18873 21404 19178
rect 22664 18970 22692 22200
rect 22652 18964 22704 18970
rect 22652 18906 22704 18912
rect 21362 18864 21418 18873
rect 21362 18799 21418 18808
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21376 18465 21404 18634
rect 21362 18456 21418 18465
rect 21362 18391 21418 18400
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21376 18057 21404 18090
rect 21362 18048 21418 18057
rect 21362 17983 21418 17992
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21376 17105 21404 17546
rect 21362 17096 21418 17105
rect 21362 17031 21418 17040
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21284 16561 21312 16934
rect 21364 16652 21416 16658
rect 21364 16594 21416 16600
rect 21270 16552 21326 16561
rect 21270 16487 21326 16496
rect 20812 16390 20864 16396
rect 20824 15638 20852 16390
rect 21008 16374 21220 16402
rect 20812 15632 20864 15638
rect 20812 15574 20864 15580
rect 20352 14894 20404 14900
rect 20626 14920 20682 14929
rect 20364 14550 20392 14894
rect 20626 14855 20682 14864
rect 20352 14544 20404 14550
rect 20352 14486 20404 14492
rect 20534 14512 20590 14521
rect 20444 14476 20496 14482
rect 20534 14447 20590 14456
rect 20444 14418 20496 14424
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 13938 20392 14214
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20260 13796 20312 13802
rect 20260 13738 20312 13744
rect 20168 13456 20220 13462
rect 20168 13398 20220 13404
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20076 12708 20128 12714
rect 20076 12650 20128 12656
rect 19616 12378 19668 12384
rect 19904 12406 20024 12434
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18800 11937 18828 12106
rect 18786 11928 18842 11937
rect 18786 11863 18842 11872
rect 18786 11248 18842 11257
rect 18786 11183 18788 11192
rect 18840 11183 18842 11192
rect 18788 11154 18840 11160
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18236 10260 18288 10266
rect 18236 10202 18288 10208
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 17972 10130 18092 10146
rect 18800 10130 18828 10678
rect 18892 10674 18920 12242
rect 18972 12232 19024 12238
rect 18972 12174 19024 12180
rect 18984 11694 19012 12174
rect 19904 11898 19932 12406
rect 20088 12374 20116 12650
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 18972 11688 19024 11694
rect 18972 11630 19024 11636
rect 19340 11688 19392 11694
rect 19340 11630 19392 11636
rect 18984 11132 19012 11630
rect 19156 11552 19208 11558
rect 19156 11494 19208 11500
rect 19064 11144 19116 11150
rect 18984 11104 19064 11132
rect 18984 10810 19012 11104
rect 19064 11086 19116 11092
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 19168 10690 19196 11494
rect 19352 11150 19380 11630
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18984 10662 19196 10690
rect 18878 10160 18934 10169
rect 17960 10124 18092 10130
rect 18012 10118 18092 10124
rect 17960 10066 18012 10072
rect 17958 10024 18014 10033
rect 17958 9959 17960 9968
rect 18012 9959 18014 9968
rect 17960 9930 18012 9936
rect 18064 8974 18092 10118
rect 18788 10124 18840 10130
rect 18878 10095 18934 10104
rect 18788 10066 18840 10072
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18604 10056 18656 10062
rect 18604 9998 18656 10004
rect 18156 9178 18184 9998
rect 18282 9820 18578 9840
rect 18338 9818 18362 9820
rect 18418 9818 18442 9820
rect 18498 9818 18522 9820
rect 18360 9766 18362 9818
rect 18424 9766 18436 9818
rect 18498 9766 18500 9818
rect 18338 9764 18362 9766
rect 18418 9764 18442 9766
rect 18498 9764 18522 9766
rect 18282 9744 18578 9764
rect 18616 9722 18644 9998
rect 18892 9761 18920 10095
rect 18878 9752 18934 9761
rect 18604 9716 18656 9722
rect 18878 9687 18934 9696
rect 18604 9658 18656 9664
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 18696 8968 18748 8974
rect 18696 8910 18748 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17972 8129 18000 8570
rect 18064 8498 18092 8910
rect 18282 8732 18578 8752
rect 18338 8730 18362 8732
rect 18418 8730 18442 8732
rect 18498 8730 18522 8732
rect 18360 8678 18362 8730
rect 18424 8678 18436 8730
rect 18498 8678 18500 8730
rect 18338 8676 18362 8678
rect 18418 8676 18442 8678
rect 18498 8676 18522 8678
rect 18282 8656 18578 8676
rect 18708 8634 18736 8910
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18800 8673 18828 8774
rect 18786 8664 18842 8673
rect 18696 8628 18748 8634
rect 18786 8599 18842 8608
rect 18696 8570 18748 8576
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17958 8120 18014 8129
rect 17684 8084 17736 8090
rect 17958 8055 18014 8064
rect 17684 8026 17736 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17788 7449 17816 7890
rect 17774 7440 17830 7449
rect 17774 7375 17830 7384
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17328 5914 17356 6734
rect 17776 6656 17828 6662
rect 17590 6624 17646 6633
rect 17776 6598 17828 6604
rect 17590 6559 17646 6568
rect 17408 6180 17460 6186
rect 17408 6122 17460 6128
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17314 5536 17370 5545
rect 17314 5471 17370 5480
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17052 5086 17264 5114
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16960 3126 16988 3470
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16856 1692 16908 1698
rect 16856 1634 16908 1640
rect 17052 800 17080 4490
rect 17144 4078 17172 4966
rect 17236 4078 17264 5086
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17144 2990 17172 3470
rect 17328 3398 17356 5471
rect 17420 4826 17448 6122
rect 17604 5098 17632 6559
rect 17592 5092 17644 5098
rect 17592 5034 17644 5040
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17420 4214 17448 4762
rect 17788 4758 17816 6598
rect 17880 5914 17908 7958
rect 18064 7954 18092 8230
rect 18052 7948 18104 7954
rect 18052 7890 18104 7896
rect 18064 7721 18092 7890
rect 18050 7712 18106 7721
rect 18050 7647 18106 7656
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17868 5908 17920 5914
rect 17868 5850 17920 5856
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17512 3534 17540 4150
rect 17592 4004 17644 4010
rect 17592 3946 17644 3952
rect 17604 3602 17632 3946
rect 17592 3596 17644 3602
rect 17592 3538 17644 3544
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17316 3392 17368 3398
rect 17316 3334 17368 3340
rect 17132 2984 17184 2990
rect 17132 2926 17184 2932
rect 17972 2666 18000 6598
rect 18156 5522 18184 8502
rect 18788 8424 18840 8430
rect 18788 8366 18840 8372
rect 18800 8090 18828 8366
rect 18788 8084 18840 8090
rect 18788 8026 18840 8032
rect 18892 7970 18920 9687
rect 18984 8294 19012 10662
rect 19352 10538 19380 11086
rect 19536 10577 19564 11494
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19522 10568 19578 10577
rect 19340 10532 19392 10538
rect 19522 10503 19578 10512
rect 19340 10474 19392 10480
rect 19352 9450 19380 10474
rect 19720 10266 19748 11154
rect 20352 10532 20404 10538
rect 20352 10474 20404 10480
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 20168 10192 20220 10198
rect 20168 10134 20220 10140
rect 20180 9518 20208 10134
rect 20364 10062 20392 10474
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20168 9512 20220 9518
rect 20168 9454 20220 9460
rect 19340 9444 19392 9450
rect 19340 9386 19392 9392
rect 19156 9376 19208 9382
rect 19156 9318 19208 9324
rect 19064 8968 19116 8974
rect 19064 8910 19116 8916
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18800 7942 18920 7970
rect 18282 7644 18578 7664
rect 18338 7642 18362 7644
rect 18418 7642 18442 7644
rect 18498 7642 18522 7644
rect 18360 7590 18362 7642
rect 18424 7590 18436 7642
rect 18498 7590 18500 7642
rect 18338 7588 18362 7590
rect 18418 7588 18442 7590
rect 18498 7588 18522 7590
rect 18282 7568 18578 7588
rect 18800 6798 18828 7942
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18984 7410 19012 7686
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18892 6798 18920 7278
rect 19076 6934 19104 8910
rect 19168 8430 19196 9318
rect 19246 8936 19302 8945
rect 19246 8871 19302 8880
rect 19260 8634 19288 8871
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19352 8430 19380 9386
rect 20272 9058 20300 9998
rect 20364 9722 20392 9998
rect 20352 9716 20404 9722
rect 20352 9658 20404 9664
rect 20180 9042 20300 9058
rect 20168 9036 20300 9042
rect 20220 9030 20300 9036
rect 20168 8978 20220 8984
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19248 8288 19300 8294
rect 19248 8230 19300 8236
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19168 7342 19196 7686
rect 19156 7336 19208 7342
rect 19156 7278 19208 7284
rect 19260 7154 19288 8230
rect 19352 7954 19380 8366
rect 19340 7948 19392 7954
rect 19340 7890 19392 7896
rect 19168 7126 19288 7154
rect 19064 6928 19116 6934
rect 19064 6870 19116 6876
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18282 6556 18578 6576
rect 18338 6554 18362 6556
rect 18418 6554 18442 6556
rect 18498 6554 18522 6556
rect 18360 6502 18362 6554
rect 18424 6502 18436 6554
rect 18498 6502 18500 6554
rect 18338 6500 18362 6502
rect 18418 6500 18442 6502
rect 18498 6500 18522 6502
rect 18282 6480 18578 6500
rect 18892 6254 18920 6734
rect 18880 6248 18932 6254
rect 18880 6190 18932 6196
rect 18788 6180 18840 6186
rect 18788 6122 18840 6128
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18708 5574 18736 5743
rect 17604 2638 18000 2666
rect 18064 5494 18184 5522
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 17604 2582 17632 2638
rect 17592 2576 17644 2582
rect 17592 2518 17644 2524
rect 17960 2508 18012 2514
rect 17960 2450 18012 2456
rect 17868 2440 17920 2446
rect 17868 2382 17920 2388
rect 17776 2372 17828 2378
rect 17776 2314 17828 2320
rect 17788 1170 17816 2314
rect 17880 1766 17908 2382
rect 17972 2038 18000 2450
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 17868 1760 17920 1766
rect 17868 1702 17920 1708
rect 18064 1630 18092 5494
rect 18282 5468 18578 5488
rect 18338 5466 18362 5468
rect 18418 5466 18442 5468
rect 18498 5466 18522 5468
rect 18360 5414 18362 5466
rect 18424 5414 18436 5466
rect 18498 5414 18500 5466
rect 18338 5412 18362 5414
rect 18418 5412 18442 5414
rect 18498 5412 18522 5414
rect 18282 5392 18578 5412
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18142 5264 18198 5273
rect 18142 5199 18198 5208
rect 18156 4826 18184 5199
rect 18616 4865 18644 5306
rect 18602 4856 18658 4865
rect 18144 4820 18196 4826
rect 18800 4842 18828 6122
rect 18892 5710 18920 6190
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18602 4791 18658 4800
rect 18708 4814 18828 4842
rect 18892 4826 18920 5646
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18880 4820 18932 4826
rect 18144 4762 18196 4768
rect 18510 4720 18566 4729
rect 18510 4655 18512 4664
rect 18564 4655 18566 4664
rect 18512 4626 18564 4632
rect 18144 4616 18196 4622
rect 18708 4570 18736 4814
rect 18880 4762 18932 4768
rect 18788 4684 18840 4690
rect 18788 4626 18840 4632
rect 18144 4558 18196 4564
rect 18156 4214 18184 4558
rect 18616 4542 18736 4570
rect 18282 4380 18578 4400
rect 18338 4378 18362 4380
rect 18418 4378 18442 4380
rect 18498 4378 18522 4380
rect 18360 4326 18362 4378
rect 18424 4326 18436 4378
rect 18498 4326 18500 4378
rect 18338 4324 18362 4326
rect 18418 4324 18442 4326
rect 18498 4324 18522 4326
rect 18282 4304 18578 4324
rect 18144 4208 18196 4214
rect 18144 4150 18196 4156
rect 18616 3890 18644 4542
rect 18694 4448 18750 4457
rect 18694 4383 18750 4392
rect 18708 4282 18736 4383
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18616 3862 18736 3890
rect 18604 3732 18656 3738
rect 18604 3674 18656 3680
rect 18144 3596 18196 3602
rect 18144 3538 18196 3544
rect 18156 3194 18184 3538
rect 18282 3292 18578 3312
rect 18338 3290 18362 3292
rect 18418 3290 18442 3292
rect 18498 3290 18522 3292
rect 18360 3238 18362 3290
rect 18424 3238 18436 3290
rect 18498 3238 18500 3290
rect 18338 3236 18362 3238
rect 18418 3236 18442 3238
rect 18498 3236 18522 3238
rect 18282 3216 18578 3236
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18156 2582 18184 3130
rect 18512 3052 18564 3058
rect 18512 2994 18564 3000
rect 18524 2650 18552 2994
rect 18616 2650 18644 3674
rect 18708 3602 18736 3862
rect 18696 3596 18748 3602
rect 18696 3538 18748 3544
rect 18800 3505 18828 4626
rect 18892 4622 18920 4762
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18880 4004 18932 4010
rect 18880 3946 18932 3952
rect 18892 3738 18920 3946
rect 18880 3732 18932 3738
rect 18880 3674 18932 3680
rect 18786 3496 18842 3505
rect 18786 3431 18842 3440
rect 18892 3058 18920 3674
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18878 2952 18934 2961
rect 18878 2887 18934 2896
rect 18788 2848 18840 2854
rect 18786 2816 18788 2825
rect 18840 2816 18842 2825
rect 18786 2751 18842 2760
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18604 2644 18656 2650
rect 18604 2586 18656 2592
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 18052 1624 18104 1630
rect 18052 1566 18104 1572
rect 17696 1142 17816 1170
rect 18156 1170 18184 2246
rect 18282 2204 18578 2224
rect 18338 2202 18362 2204
rect 18418 2202 18442 2204
rect 18498 2202 18522 2204
rect 18360 2150 18362 2202
rect 18424 2150 18436 2202
rect 18498 2150 18500 2202
rect 18338 2148 18362 2150
rect 18418 2148 18442 2150
rect 18498 2148 18522 2150
rect 18282 2128 18578 2148
rect 18156 1142 18276 1170
rect 17696 800 17724 1142
rect 18248 800 18276 1142
rect 18892 898 18920 2887
rect 18984 2582 19012 5510
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 2990 19104 4966
rect 19168 4729 19196 7126
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19154 4720 19210 4729
rect 19154 4655 19210 4664
rect 19156 4616 19208 4622
rect 19156 4558 19208 4564
rect 19168 3738 19196 4558
rect 19156 3732 19208 3738
rect 19156 3674 19208 3680
rect 19154 3632 19210 3641
rect 19260 3618 19288 5034
rect 19260 3590 19472 3618
rect 19154 3567 19210 3576
rect 19168 3516 19196 3567
rect 19168 3488 19288 3516
rect 19260 3398 19288 3488
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19248 3392 19300 3398
rect 19248 3334 19300 3340
rect 19064 2984 19116 2990
rect 19064 2926 19116 2932
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 19076 2582 19104 2751
rect 18972 2576 19024 2582
rect 18972 2518 19024 2524
rect 19064 2576 19116 2582
rect 19064 2518 19116 2524
rect 19168 2378 19196 3334
rect 19248 2984 19300 2990
rect 19248 2926 19300 2932
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 19260 2310 19288 2926
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 18800 870 18920 898
rect 18800 800 18828 870
rect 19352 800 19380 3402
rect 19444 2378 19472 3590
rect 19536 2553 19564 8774
rect 19996 8566 20024 8774
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19720 2854 19748 6394
rect 19800 5840 19852 5846
rect 19800 5782 19852 5788
rect 19812 5302 19840 5782
rect 19800 5296 19852 5302
rect 19800 5238 19852 5244
rect 19904 5234 19932 7142
rect 20088 6934 20116 7346
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19996 5166 20024 6598
rect 20088 6458 20116 6870
rect 20076 6452 20128 6458
rect 20076 6394 20128 6400
rect 20180 6361 20208 8978
rect 20260 7200 20312 7206
rect 20260 7142 20312 7148
rect 20352 7200 20404 7206
rect 20352 7142 20404 7148
rect 20272 6458 20300 7142
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20166 6352 20222 6361
rect 20076 6316 20128 6322
rect 20166 6287 20222 6296
rect 20076 6258 20128 6264
rect 20088 5846 20116 6258
rect 20364 5914 20392 7142
rect 20352 5908 20404 5914
rect 20352 5850 20404 5856
rect 20076 5840 20128 5846
rect 20076 5782 20128 5788
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20088 4146 20116 4626
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20352 3936 20404 3942
rect 20352 3878 20404 3884
rect 20364 3097 20392 3878
rect 20456 3670 20484 14418
rect 20548 14414 20576 14447
rect 20536 14408 20588 14414
rect 20536 14350 20588 14356
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 20640 12850 20668 13194
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20640 12306 20668 12786
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20640 11898 20668 12242
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20732 9761 20760 12582
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20824 10130 20852 11290
rect 20916 10810 20944 12582
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20718 9752 20774 9761
rect 20718 9687 20774 9696
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20824 9178 20852 9318
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20628 8356 20680 8362
rect 20628 8298 20680 8304
rect 20536 7948 20588 7954
rect 20536 7890 20588 7896
rect 20548 6662 20576 7890
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20548 5234 20576 6598
rect 20640 5846 20668 8298
rect 20916 7970 20944 10406
rect 21008 10266 21036 16374
rect 21376 16153 21404 16594
rect 21362 16144 21418 16153
rect 21362 16079 21418 16088
rect 21364 15972 21416 15978
rect 21364 15914 21416 15920
rect 21376 15609 21404 15914
rect 21362 15600 21418 15609
rect 21362 15535 21418 15544
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21284 15201 21312 15302
rect 21270 15192 21326 15201
rect 21270 15127 21326 15136
rect 21364 14884 21416 14890
rect 21364 14826 21416 14832
rect 21376 14657 21404 14826
rect 21362 14648 21418 14657
rect 21362 14583 21418 14592
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21192 13462 21220 14282
rect 21376 14249 21404 14282
rect 21362 14240 21418 14249
rect 21362 14175 21418 14184
rect 21364 13864 21416 13870
rect 21362 13832 21364 13841
rect 21416 13832 21418 13841
rect 21362 13767 21418 13776
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21362 13288 21418 13297
rect 21362 13223 21364 13232
rect 21416 13223 21418 13232
rect 21364 13194 21416 13200
rect 21180 11620 21232 11626
rect 21180 11562 21232 11568
rect 21192 11354 21220 11562
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21192 10674 21220 11290
rect 21180 10668 21232 10674
rect 21180 10610 21232 10616
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 8974 21036 9522
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21008 8362 21036 8910
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 21008 8090 21036 8298
rect 20996 8084 21048 8090
rect 20996 8026 21048 8032
rect 20916 7942 21036 7970
rect 21008 7750 21036 7942
rect 20996 7744 21048 7750
rect 20996 7686 21048 7692
rect 20904 7200 20956 7206
rect 20904 7142 20956 7148
rect 20916 7002 20944 7142
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 21008 6254 21036 7686
rect 20996 6248 21048 6254
rect 20996 6190 21048 6196
rect 21100 6118 21128 10406
rect 21272 9920 21324 9926
rect 21272 9862 21324 9868
rect 21088 6112 21140 6118
rect 21088 6054 21140 6060
rect 20628 5840 20680 5846
rect 20628 5782 20680 5788
rect 20996 5636 21048 5642
rect 20996 5578 21048 5584
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20626 5128 20682 5137
rect 20626 5063 20682 5072
rect 20640 5030 20668 5063
rect 20628 5024 20680 5030
rect 20628 4966 20680 4972
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20444 3664 20496 3670
rect 20444 3606 20496 3612
rect 20350 3088 20406 3097
rect 20350 3023 20406 3032
rect 20640 2990 20668 3674
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20732 3505 20760 3538
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20812 3392 20864 3398
rect 20812 3334 20864 3340
rect 20824 3058 20852 3334
rect 20812 3052 20864 3058
rect 20812 2994 20864 3000
rect 20628 2984 20680 2990
rect 19798 2952 19854 2961
rect 20628 2926 20680 2932
rect 19798 2887 19800 2896
rect 19852 2887 19854 2896
rect 19800 2858 19852 2864
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 20640 2774 20668 2926
rect 20640 2746 20760 2774
rect 19522 2544 19578 2553
rect 19522 2479 19524 2488
rect 19576 2479 19578 2488
rect 19524 2450 19576 2456
rect 19536 2419 19564 2450
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 19892 2100 19944 2106
rect 19892 2042 19944 2048
rect 19904 800 19932 2042
rect 20732 2009 20760 2746
rect 20718 2000 20774 2009
rect 20718 1935 20774 1944
rect 20444 1828 20496 1834
rect 20444 1770 20496 1776
rect 20456 800 20484 1770
rect 20916 1601 20944 3606
rect 20902 1592 20958 1601
rect 20902 1527 20958 1536
rect 21008 800 21036 5578
rect 21100 5545 21128 6054
rect 21086 5536 21142 5545
rect 21086 5471 21142 5480
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21088 5024 21140 5030
rect 21088 4966 21140 4972
rect 21100 4282 21128 4966
rect 21192 4826 21220 5170
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21088 4276 21140 4282
rect 21088 4218 21140 4224
rect 21284 4078 21312 9862
rect 22100 4752 22152 4758
rect 22100 4694 22152 4700
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21180 3392 21232 3398
rect 21180 3334 21232 3340
rect 21192 3194 21220 3334
rect 21180 3188 21232 3194
rect 21180 3130 21232 3136
rect 21284 2961 21312 4014
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21270 2952 21326 2961
rect 21270 2887 21326 2896
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21100 1970 21128 2314
rect 21088 1964 21140 1970
rect 21088 1906 21140 1912
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2502 0 2558 800
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17038 0 17094 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21376 649 21404 3062
rect 21560 800 21588 4422
rect 21916 1488 21968 1494
rect 21916 1430 21968 1436
rect 21362 640 21418 649
rect 21362 575 21418 584
rect 21546 0 21602 800
rect 21928 241 21956 1430
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 22020 1057 22048 1362
rect 22006 1048 22062 1057
rect 22006 983 22062 992
rect 22112 800 22140 4694
rect 22652 1556 22704 1562
rect 22652 1498 22704 1504
rect 22664 800 22692 1498
rect 21914 232 21970 241
rect 21914 167 21970 176
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 17958 22208 18014 22264
rect 1582 17212 1584 17232
rect 1584 17212 1636 17232
rect 1636 17212 1638 17232
rect 1582 17176 1638 17212
rect 2318 19896 2374 19952
rect 4421 20698 4477 20700
rect 4501 20698 4557 20700
rect 4581 20698 4637 20700
rect 4661 20698 4717 20700
rect 4421 20646 4447 20698
rect 4447 20646 4477 20698
rect 4501 20646 4511 20698
rect 4511 20646 4557 20698
rect 4581 20646 4627 20698
rect 4627 20646 4637 20698
rect 4661 20646 4691 20698
rect 4691 20646 4717 20698
rect 4421 20644 4477 20646
rect 4501 20644 4557 20646
rect 4581 20644 4637 20646
rect 4661 20644 4717 20646
rect 2778 19780 2834 19816
rect 2778 19760 2780 19780
rect 2780 19760 2832 19780
rect 2832 19760 2834 19780
rect 4421 19610 4477 19612
rect 4501 19610 4557 19612
rect 4581 19610 4637 19612
rect 4661 19610 4717 19612
rect 4421 19558 4447 19610
rect 4447 19558 4477 19610
rect 4501 19558 4511 19610
rect 4511 19558 4557 19610
rect 4581 19558 4627 19610
rect 4627 19558 4637 19610
rect 4661 19558 4691 19610
rect 4691 19558 4717 19610
rect 4421 19556 4477 19558
rect 4501 19556 4557 19558
rect 4581 19556 4637 19558
rect 4661 19556 4717 19558
rect 4421 18522 4477 18524
rect 4501 18522 4557 18524
rect 4581 18522 4637 18524
rect 4661 18522 4717 18524
rect 4421 18470 4447 18522
rect 4447 18470 4477 18522
rect 4501 18470 4511 18522
rect 4511 18470 4557 18522
rect 4581 18470 4627 18522
rect 4627 18470 4637 18522
rect 4661 18470 4691 18522
rect 4691 18470 4717 18522
rect 4421 18468 4477 18470
rect 4501 18468 4557 18470
rect 4581 18468 4637 18470
rect 4661 18468 4717 18470
rect 4421 17434 4477 17436
rect 4501 17434 4557 17436
rect 4581 17434 4637 17436
rect 4661 17434 4717 17436
rect 4421 17382 4447 17434
rect 4447 17382 4477 17434
rect 4501 17382 4511 17434
rect 4511 17382 4557 17434
rect 4581 17382 4627 17434
rect 4627 17382 4637 17434
rect 4661 17382 4691 17434
rect 4691 17382 4717 17434
rect 4421 17380 4477 17382
rect 4501 17380 4557 17382
rect 4581 17380 4637 17382
rect 4661 17380 4717 17382
rect 4421 16346 4477 16348
rect 4501 16346 4557 16348
rect 4581 16346 4637 16348
rect 4661 16346 4717 16348
rect 4421 16294 4447 16346
rect 4447 16294 4477 16346
rect 4501 16294 4511 16346
rect 4511 16294 4557 16346
rect 4581 16294 4627 16346
rect 4627 16294 4637 16346
rect 4661 16294 4691 16346
rect 4691 16294 4717 16346
rect 4421 16292 4477 16294
rect 4501 16292 4557 16294
rect 4581 16292 4637 16294
rect 4661 16292 4717 16294
rect 4421 15258 4477 15260
rect 4501 15258 4557 15260
rect 4581 15258 4637 15260
rect 4661 15258 4717 15260
rect 4421 15206 4447 15258
rect 4447 15206 4477 15258
rect 4501 15206 4511 15258
rect 4511 15206 4557 15258
rect 4581 15206 4627 15258
rect 4627 15206 4637 15258
rect 4661 15206 4691 15258
rect 4691 15206 4717 15258
rect 4421 15204 4477 15206
rect 4501 15204 4557 15206
rect 4581 15204 4637 15206
rect 4661 15204 4717 15206
rect 4421 14170 4477 14172
rect 4501 14170 4557 14172
rect 4581 14170 4637 14172
rect 4661 14170 4717 14172
rect 4421 14118 4447 14170
rect 4447 14118 4477 14170
rect 4501 14118 4511 14170
rect 4511 14118 4557 14170
rect 4581 14118 4627 14170
rect 4627 14118 4637 14170
rect 4661 14118 4691 14170
rect 4691 14118 4717 14170
rect 4421 14116 4477 14118
rect 4501 14116 4557 14118
rect 4581 14116 4637 14118
rect 4661 14116 4717 14118
rect 4421 13082 4477 13084
rect 4501 13082 4557 13084
rect 4581 13082 4637 13084
rect 4661 13082 4717 13084
rect 4421 13030 4447 13082
rect 4447 13030 4477 13082
rect 4501 13030 4511 13082
rect 4511 13030 4557 13082
rect 4581 13030 4627 13082
rect 4627 13030 4637 13082
rect 4661 13030 4691 13082
rect 4691 13030 4717 13082
rect 4421 13028 4477 13030
rect 4501 13028 4557 13030
rect 4581 13028 4637 13030
rect 4661 13028 4717 13030
rect 5262 17448 5318 17504
rect 4421 11994 4477 11996
rect 4501 11994 4557 11996
rect 4581 11994 4637 11996
rect 4661 11994 4717 11996
rect 4421 11942 4447 11994
rect 4447 11942 4477 11994
rect 4501 11942 4511 11994
rect 4511 11942 4557 11994
rect 4581 11942 4627 11994
rect 4627 11942 4637 11994
rect 4661 11942 4691 11994
rect 4691 11942 4717 11994
rect 4421 11940 4477 11942
rect 4501 11940 4557 11942
rect 4581 11940 4637 11942
rect 4661 11940 4717 11942
rect 5722 15972 5778 16008
rect 5722 15952 5724 15972
rect 5724 15952 5776 15972
rect 5776 15952 5778 15972
rect 4421 10906 4477 10908
rect 4501 10906 4557 10908
rect 4581 10906 4637 10908
rect 4661 10906 4717 10908
rect 4421 10854 4447 10906
rect 4447 10854 4477 10906
rect 4501 10854 4511 10906
rect 4511 10854 4557 10906
rect 4581 10854 4627 10906
rect 4627 10854 4637 10906
rect 4661 10854 4691 10906
rect 4691 10854 4717 10906
rect 4421 10852 4477 10854
rect 4501 10852 4557 10854
rect 4581 10852 4637 10854
rect 4661 10852 4717 10854
rect 1582 5772 1638 5808
rect 1582 5752 1584 5772
rect 1584 5752 1636 5772
rect 1636 5752 1638 5772
rect 4421 9818 4477 9820
rect 4501 9818 4557 9820
rect 4581 9818 4637 9820
rect 4661 9818 4717 9820
rect 4421 9766 4447 9818
rect 4447 9766 4477 9818
rect 4501 9766 4511 9818
rect 4511 9766 4557 9818
rect 4581 9766 4627 9818
rect 4627 9766 4637 9818
rect 4661 9766 4691 9818
rect 4691 9766 4717 9818
rect 4421 9764 4477 9766
rect 4501 9764 4557 9766
rect 4581 9764 4637 9766
rect 4661 9764 4717 9766
rect 4421 8730 4477 8732
rect 4501 8730 4557 8732
rect 4581 8730 4637 8732
rect 4661 8730 4717 8732
rect 4421 8678 4447 8730
rect 4447 8678 4477 8730
rect 4501 8678 4511 8730
rect 4511 8678 4557 8730
rect 4581 8678 4627 8730
rect 4627 8678 4637 8730
rect 4661 8678 4691 8730
rect 4691 8678 4717 8730
rect 4421 8676 4477 8678
rect 4501 8676 4557 8678
rect 4581 8676 4637 8678
rect 4661 8676 4717 8678
rect 4421 7642 4477 7644
rect 4501 7642 4557 7644
rect 4581 7642 4637 7644
rect 4661 7642 4717 7644
rect 4421 7590 4447 7642
rect 4447 7590 4477 7642
rect 4501 7590 4511 7642
rect 4511 7590 4557 7642
rect 4581 7590 4627 7642
rect 4627 7590 4637 7642
rect 4661 7590 4691 7642
rect 4691 7590 4717 7642
rect 4421 7588 4477 7590
rect 4501 7588 4557 7590
rect 4581 7588 4637 7590
rect 4661 7588 4717 7590
rect 4421 6554 4477 6556
rect 4501 6554 4557 6556
rect 4581 6554 4637 6556
rect 4661 6554 4717 6556
rect 4421 6502 4447 6554
rect 4447 6502 4477 6554
rect 4501 6502 4511 6554
rect 4511 6502 4557 6554
rect 4581 6502 4627 6554
rect 4627 6502 4637 6554
rect 4661 6502 4691 6554
rect 4691 6502 4717 6554
rect 4421 6500 4477 6502
rect 4501 6500 4557 6502
rect 4581 6500 4637 6502
rect 4661 6500 4717 6502
rect 4421 5466 4477 5468
rect 4501 5466 4557 5468
rect 4581 5466 4637 5468
rect 4661 5466 4717 5468
rect 4421 5414 4447 5466
rect 4447 5414 4477 5466
rect 4501 5414 4511 5466
rect 4511 5414 4557 5466
rect 4581 5414 4627 5466
rect 4627 5414 4637 5466
rect 4661 5414 4691 5466
rect 4691 5414 4717 5466
rect 4421 5412 4477 5414
rect 4501 5412 4557 5414
rect 4581 5412 4637 5414
rect 4661 5412 4717 5414
rect 4421 4378 4477 4380
rect 4501 4378 4557 4380
rect 4581 4378 4637 4380
rect 4661 4378 4717 4380
rect 4421 4326 4447 4378
rect 4447 4326 4477 4378
rect 4501 4326 4511 4378
rect 4511 4326 4557 4378
rect 4581 4326 4627 4378
rect 4627 4326 4637 4378
rect 4661 4326 4691 4378
rect 4691 4326 4717 4378
rect 4421 4324 4477 4326
rect 4501 4324 4557 4326
rect 4581 4324 4637 4326
rect 4661 4324 4717 4326
rect 4421 3290 4477 3292
rect 4501 3290 4557 3292
rect 4581 3290 4637 3292
rect 4661 3290 4717 3292
rect 4421 3238 4447 3290
rect 4447 3238 4477 3290
rect 4501 3238 4511 3290
rect 4511 3238 4557 3290
rect 4581 3238 4627 3290
rect 4627 3238 4637 3290
rect 4661 3238 4691 3290
rect 4691 3238 4717 3290
rect 4421 3236 4477 3238
rect 4501 3236 4557 3238
rect 4581 3236 4637 3238
rect 4661 3236 4717 3238
rect 4434 3068 4436 3088
rect 4436 3068 4488 3088
rect 4488 3068 4490 3088
rect 4434 3032 4490 3068
rect 6182 19216 6238 19272
rect 6826 19660 6828 19680
rect 6828 19660 6880 19680
rect 6880 19660 6882 19680
rect 6826 19624 6882 19660
rect 6734 19488 6790 19544
rect 6826 18400 6882 18456
rect 6642 18128 6698 18184
rect 6366 17176 6422 17232
rect 7102 19896 7158 19952
rect 7378 19488 7434 19544
rect 7010 17312 7066 17368
rect 6734 15952 6790 16008
rect 6458 15544 6514 15600
rect 4421 2202 4477 2204
rect 4501 2202 4557 2204
rect 4581 2202 4637 2204
rect 4661 2202 4717 2204
rect 4421 2150 4447 2202
rect 4447 2150 4477 2202
rect 4501 2150 4511 2202
rect 4511 2150 4557 2202
rect 4581 2150 4627 2202
rect 4627 2150 4637 2202
rect 4661 2150 4691 2202
rect 4691 2150 4717 2202
rect 4421 2148 4477 2150
rect 4501 2148 4557 2150
rect 4581 2148 4637 2150
rect 4661 2148 4717 2150
rect 6550 7248 6606 7304
rect 7378 19252 7380 19272
rect 7380 19252 7432 19272
rect 7432 19252 7434 19272
rect 7378 19216 7434 19252
rect 7886 20154 7942 20156
rect 7966 20154 8022 20156
rect 8046 20154 8102 20156
rect 8126 20154 8182 20156
rect 7886 20102 7912 20154
rect 7912 20102 7942 20154
rect 7966 20102 7976 20154
rect 7976 20102 8022 20154
rect 8046 20102 8092 20154
rect 8092 20102 8102 20154
rect 8126 20102 8156 20154
rect 8156 20102 8182 20154
rect 7886 20100 7942 20102
rect 7966 20100 8022 20102
rect 8046 20100 8102 20102
rect 8126 20100 8182 20102
rect 8850 20304 8906 20360
rect 8390 20168 8446 20224
rect 7470 18264 7526 18320
rect 8114 19624 8170 19680
rect 7886 19066 7942 19068
rect 7966 19066 8022 19068
rect 8046 19066 8102 19068
rect 8126 19066 8182 19068
rect 7886 19014 7912 19066
rect 7912 19014 7942 19066
rect 7966 19014 7976 19066
rect 7976 19014 8022 19066
rect 8046 19014 8092 19066
rect 8092 19014 8102 19066
rect 8126 19014 8156 19066
rect 8156 19014 8182 19066
rect 7886 19012 7942 19014
rect 7966 19012 8022 19014
rect 8046 19012 8102 19014
rect 8126 19012 8182 19014
rect 7746 18672 7802 18728
rect 7378 17720 7434 17776
rect 7286 16768 7342 16824
rect 7194 8880 7250 8936
rect 6918 5752 6974 5808
rect 7194 7384 7250 7440
rect 7930 18264 7986 18320
rect 7886 17978 7942 17980
rect 7966 17978 8022 17980
rect 8046 17978 8102 17980
rect 8126 17978 8182 17980
rect 7886 17926 7912 17978
rect 7912 17926 7942 17978
rect 7966 17926 7976 17978
rect 7976 17926 8022 17978
rect 8046 17926 8092 17978
rect 8092 17926 8102 17978
rect 8126 17926 8156 17978
rect 8156 17926 8182 17978
rect 7886 17924 7942 17926
rect 7966 17924 8022 17926
rect 8046 17924 8102 17926
rect 8126 17924 8182 17926
rect 8298 19216 8354 19272
rect 8206 17176 8262 17232
rect 7886 16890 7942 16892
rect 7966 16890 8022 16892
rect 8046 16890 8102 16892
rect 8126 16890 8182 16892
rect 7886 16838 7912 16890
rect 7912 16838 7942 16890
rect 7966 16838 7976 16890
rect 7976 16838 8022 16890
rect 8046 16838 8092 16890
rect 8092 16838 8102 16890
rect 8126 16838 8156 16890
rect 8156 16838 8182 16890
rect 7886 16836 7942 16838
rect 7966 16836 8022 16838
rect 8046 16836 8102 16838
rect 8126 16836 8182 16838
rect 8114 16632 8170 16688
rect 8574 18128 8630 18184
rect 8850 18944 8906 19000
rect 8758 18264 8814 18320
rect 8666 17992 8722 18048
rect 8574 16652 8630 16688
rect 8574 16632 8576 16652
rect 8576 16632 8628 16652
rect 8628 16632 8630 16652
rect 7886 15802 7942 15804
rect 7966 15802 8022 15804
rect 8046 15802 8102 15804
rect 8126 15802 8182 15804
rect 7886 15750 7912 15802
rect 7912 15750 7942 15802
rect 7966 15750 7976 15802
rect 7976 15750 8022 15802
rect 8046 15750 8092 15802
rect 8092 15750 8102 15802
rect 8126 15750 8156 15802
rect 8156 15750 8182 15802
rect 7886 15748 7942 15750
rect 7966 15748 8022 15750
rect 8046 15748 8102 15750
rect 8126 15748 8182 15750
rect 7470 9016 7526 9072
rect 7838 14864 7894 14920
rect 7886 14714 7942 14716
rect 7966 14714 8022 14716
rect 8046 14714 8102 14716
rect 8126 14714 8182 14716
rect 7886 14662 7912 14714
rect 7912 14662 7942 14714
rect 7966 14662 7976 14714
rect 7976 14662 8022 14714
rect 8046 14662 8092 14714
rect 8092 14662 8102 14714
rect 8126 14662 8156 14714
rect 8156 14662 8182 14714
rect 7886 14660 7942 14662
rect 7966 14660 8022 14662
rect 8046 14660 8102 14662
rect 8126 14660 8182 14662
rect 7886 13626 7942 13628
rect 7966 13626 8022 13628
rect 8046 13626 8102 13628
rect 8126 13626 8182 13628
rect 7886 13574 7912 13626
rect 7912 13574 7942 13626
rect 7966 13574 7976 13626
rect 7976 13574 8022 13626
rect 8046 13574 8092 13626
rect 8092 13574 8102 13626
rect 8126 13574 8156 13626
rect 8156 13574 8182 13626
rect 7886 13572 7942 13574
rect 7966 13572 8022 13574
rect 8046 13572 8102 13574
rect 8126 13572 8182 13574
rect 7654 13368 7710 13424
rect 8574 14220 8576 14240
rect 8576 14220 8628 14240
rect 8628 14220 8630 14240
rect 8574 14184 8630 14220
rect 7886 12538 7942 12540
rect 7966 12538 8022 12540
rect 8046 12538 8102 12540
rect 8126 12538 8182 12540
rect 7886 12486 7912 12538
rect 7912 12486 7942 12538
rect 7966 12486 7976 12538
rect 7976 12486 8022 12538
rect 8046 12486 8092 12538
rect 8092 12486 8102 12538
rect 8126 12486 8156 12538
rect 8156 12486 8182 12538
rect 7886 12484 7942 12486
rect 7966 12484 8022 12486
rect 8046 12484 8102 12486
rect 8126 12484 8182 12486
rect 8114 12300 8170 12336
rect 8114 12280 8116 12300
rect 8116 12280 8168 12300
rect 8168 12280 8170 12300
rect 7746 11736 7802 11792
rect 8298 12416 8354 12472
rect 7886 11450 7942 11452
rect 7966 11450 8022 11452
rect 8046 11450 8102 11452
rect 8126 11450 8182 11452
rect 7886 11398 7912 11450
rect 7912 11398 7942 11450
rect 7966 11398 7976 11450
rect 7976 11398 8022 11450
rect 8046 11398 8092 11450
rect 8092 11398 8102 11450
rect 8126 11398 8156 11450
rect 8156 11398 8182 11450
rect 7886 11396 7942 11398
rect 7966 11396 8022 11398
rect 8046 11396 8102 11398
rect 8126 11396 8182 11398
rect 7886 10362 7942 10364
rect 7966 10362 8022 10364
rect 8046 10362 8102 10364
rect 8126 10362 8182 10364
rect 7886 10310 7912 10362
rect 7912 10310 7942 10362
rect 7966 10310 7976 10362
rect 7976 10310 8022 10362
rect 8046 10310 8092 10362
rect 8092 10310 8102 10362
rect 8126 10310 8156 10362
rect 8156 10310 8182 10362
rect 7886 10308 7942 10310
rect 7966 10308 8022 10310
rect 8046 10308 8102 10310
rect 8126 10308 8182 10310
rect 7746 10240 7802 10296
rect 9402 18808 9458 18864
rect 9034 17584 9090 17640
rect 9770 20032 9826 20088
rect 9402 17856 9458 17912
rect 9218 17448 9274 17504
rect 9034 17040 9090 17096
rect 8850 14340 8906 14376
rect 8850 14320 8852 14340
rect 8852 14320 8904 14340
rect 8904 14320 8906 14340
rect 8574 10548 8576 10568
rect 8576 10548 8628 10568
rect 8628 10548 8630 10568
rect 8574 10512 8630 10548
rect 7886 9274 7942 9276
rect 7966 9274 8022 9276
rect 8046 9274 8102 9276
rect 8126 9274 8182 9276
rect 7886 9222 7912 9274
rect 7912 9222 7942 9274
rect 7966 9222 7976 9274
rect 7976 9222 8022 9274
rect 8046 9222 8092 9274
rect 8092 9222 8102 9274
rect 8126 9222 8156 9274
rect 8156 9222 8182 9274
rect 7886 9220 7942 9222
rect 7966 9220 8022 9222
rect 8046 9220 8102 9222
rect 8126 9220 8182 9222
rect 7886 8186 7942 8188
rect 7966 8186 8022 8188
rect 8046 8186 8102 8188
rect 8126 8186 8182 8188
rect 7886 8134 7912 8186
rect 7912 8134 7942 8186
rect 7966 8134 7976 8186
rect 7976 8134 8022 8186
rect 8046 8134 8092 8186
rect 8092 8134 8102 8186
rect 8126 8134 8156 8186
rect 8156 8134 8182 8186
rect 7886 8132 7942 8134
rect 7966 8132 8022 8134
rect 8046 8132 8102 8134
rect 8126 8132 8182 8134
rect 7378 5616 7434 5672
rect 7654 6860 7710 6896
rect 7654 6840 7656 6860
rect 7656 6840 7708 6860
rect 7708 6840 7710 6860
rect 7886 7098 7942 7100
rect 7966 7098 8022 7100
rect 8046 7098 8102 7100
rect 8126 7098 8182 7100
rect 7886 7046 7912 7098
rect 7912 7046 7942 7098
rect 7966 7046 7976 7098
rect 7976 7046 8022 7098
rect 8046 7046 8092 7098
rect 8092 7046 8102 7098
rect 8126 7046 8156 7098
rect 8156 7046 8182 7098
rect 7886 7044 7942 7046
rect 7966 7044 8022 7046
rect 8046 7044 8102 7046
rect 8126 7044 8182 7046
rect 7562 5616 7618 5672
rect 7286 4528 7342 4584
rect 7102 3440 7158 3496
rect 7010 3304 7066 3360
rect 6918 3168 6974 3224
rect 6918 2896 6974 2952
rect 8114 6296 8170 6352
rect 7838 6160 7894 6216
rect 7886 6010 7942 6012
rect 7966 6010 8022 6012
rect 8046 6010 8102 6012
rect 8126 6010 8182 6012
rect 7886 5958 7912 6010
rect 7912 5958 7942 6010
rect 7966 5958 7976 6010
rect 7976 5958 8022 6010
rect 8046 5958 8092 6010
rect 8092 5958 8102 6010
rect 8126 5958 8156 6010
rect 8156 5958 8182 6010
rect 7886 5956 7942 5958
rect 7966 5956 8022 5958
rect 8046 5956 8102 5958
rect 8126 5956 8182 5958
rect 8390 6976 8446 7032
rect 7654 5072 7710 5128
rect 7470 3576 7526 3632
rect 7886 4922 7942 4924
rect 7966 4922 8022 4924
rect 8046 4922 8102 4924
rect 8126 4922 8182 4924
rect 7886 4870 7912 4922
rect 7912 4870 7942 4922
rect 7966 4870 7976 4922
rect 7976 4870 8022 4922
rect 8046 4870 8092 4922
rect 8092 4870 8102 4922
rect 8126 4870 8156 4922
rect 8156 4870 8182 4922
rect 7886 4868 7942 4870
rect 7966 4868 8022 4870
rect 8046 4868 8102 4870
rect 8126 4868 8182 4870
rect 8022 4256 8078 4312
rect 8298 3884 8300 3904
rect 8300 3884 8352 3904
rect 8352 3884 8354 3904
rect 7886 3834 7942 3836
rect 7966 3834 8022 3836
rect 8046 3834 8102 3836
rect 8126 3834 8182 3836
rect 7886 3782 7912 3834
rect 7912 3782 7942 3834
rect 7966 3782 7976 3834
rect 7976 3782 8022 3834
rect 8046 3782 8092 3834
rect 8092 3782 8102 3834
rect 8126 3782 8156 3834
rect 8156 3782 8182 3834
rect 7886 3780 7942 3782
rect 7966 3780 8022 3782
rect 8046 3780 8102 3782
rect 8126 3780 8182 3782
rect 7654 2896 7710 2952
rect 7886 2746 7942 2748
rect 7966 2746 8022 2748
rect 8046 2746 8102 2748
rect 8126 2746 8182 2748
rect 7886 2694 7912 2746
rect 7912 2694 7942 2746
rect 7966 2694 7976 2746
rect 7976 2694 8022 2746
rect 8046 2694 8092 2746
rect 8092 2694 8102 2746
rect 8126 2694 8156 2746
rect 8156 2694 8182 2746
rect 7886 2692 7942 2694
rect 7966 2692 8022 2694
rect 8046 2692 8102 2694
rect 8126 2692 8182 2694
rect 7746 2488 7802 2544
rect 8298 3848 8354 3884
rect 8758 12164 8814 12200
rect 8758 12144 8760 12164
rect 8760 12144 8812 12164
rect 8812 12144 8814 12164
rect 8850 10412 8852 10432
rect 8852 10412 8904 10432
rect 8904 10412 8906 10432
rect 8850 10376 8906 10412
rect 9034 11328 9090 11384
rect 9310 17312 9366 17368
rect 9402 16768 9458 16824
rect 9678 19352 9734 19408
rect 9678 18400 9734 18456
rect 9862 17176 9918 17232
rect 9678 15408 9734 15464
rect 9678 14728 9734 14784
rect 9770 14592 9826 14648
rect 9310 14048 9366 14104
rect 9494 13776 9550 13832
rect 9402 12416 9458 12472
rect 10598 20440 10654 20496
rect 10046 19624 10102 19680
rect 9954 15000 10010 15056
rect 10230 17332 10286 17368
rect 10230 17312 10232 17332
rect 10232 17312 10284 17332
rect 10284 17312 10286 17332
rect 10690 19624 10746 19680
rect 10782 19080 10838 19136
rect 10782 18536 10838 18592
rect 11150 19896 11206 19952
rect 10414 15408 10470 15464
rect 9954 13932 10010 13968
rect 9954 13912 9956 13932
rect 9956 13912 10008 13932
rect 10008 13912 10010 13932
rect 9678 13640 9734 13696
rect 9678 13252 9734 13288
rect 9678 13232 9680 13252
rect 9680 13232 9732 13252
rect 9732 13232 9734 13252
rect 9954 12960 10010 13016
rect 9770 12824 9826 12880
rect 8574 4664 8630 4720
rect 8482 4256 8538 4312
rect 8482 3984 8538 4040
rect 9034 4800 9090 4856
rect 8942 4120 8998 4176
rect 8850 3440 8906 3496
rect 8850 2760 8906 2816
rect 9586 10104 9642 10160
rect 9494 8744 9550 8800
rect 9402 6024 9458 6080
rect 9218 4936 9274 4992
rect 9310 4392 9366 4448
rect 10046 9580 10102 9616
rect 10046 9560 10048 9580
rect 10048 9560 10100 9580
rect 10100 9560 10102 9580
rect 10322 13640 10378 13696
rect 10598 16088 10654 16144
rect 10690 15000 10746 15056
rect 10598 14456 10654 14512
rect 10138 8356 10194 8392
rect 10138 8336 10140 8356
rect 10140 8336 10192 8356
rect 10192 8336 10194 8356
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11378 20698
rect 11378 20646 11408 20698
rect 11432 20646 11442 20698
rect 11442 20646 11488 20698
rect 11512 20646 11558 20698
rect 11558 20646 11568 20698
rect 11592 20646 11622 20698
rect 11622 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 12254 20440 12310 20496
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11378 19610
rect 11378 19558 11408 19610
rect 11432 19558 11442 19610
rect 11442 19558 11488 19610
rect 11512 19558 11558 19610
rect 11558 19558 11568 19610
rect 11592 19558 11622 19610
rect 11622 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11378 18522
rect 11378 18470 11408 18522
rect 11432 18470 11442 18522
rect 11442 18470 11488 18522
rect 11512 18470 11558 18522
rect 11558 18470 11568 18522
rect 11592 18470 11622 18522
rect 11622 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11150 17720 11206 17776
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11378 17434
rect 11378 17382 11408 17434
rect 11432 17382 11442 17434
rect 11442 17382 11488 17434
rect 11512 17382 11558 17434
rect 11558 17382 11568 17434
rect 11592 17382 11622 17434
rect 11622 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11058 17176 11114 17232
rect 10966 16496 11022 16552
rect 10690 12416 10746 12472
rect 10874 12588 10876 12608
rect 10876 12588 10928 12608
rect 10928 12588 10930 12608
rect 10874 12552 10930 12588
rect 9954 8200 10010 8256
rect 9770 7928 9826 7984
rect 9678 6704 9734 6760
rect 9862 7812 9918 7848
rect 9862 7792 9864 7812
rect 9864 7792 9916 7812
rect 9916 7792 9918 7812
rect 9862 7112 9918 7168
rect 9586 5480 9642 5536
rect 9862 5344 9918 5400
rect 10138 4256 10194 4312
rect 9310 3576 9366 3632
rect 9494 3440 9550 3496
rect 9494 2624 9550 2680
rect 9586 2352 9642 2408
rect 9954 2644 10010 2680
rect 9954 2624 9956 2644
rect 9956 2624 10008 2644
rect 10008 2624 10010 2644
rect 10322 5616 10378 5672
rect 10322 5208 10378 5264
rect 12070 20168 12126 20224
rect 11794 19896 11850 19952
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11378 16346
rect 11378 16294 11408 16346
rect 11432 16294 11442 16346
rect 11442 16294 11488 16346
rect 11512 16294 11558 16346
rect 11558 16294 11568 16346
rect 11592 16294 11622 16346
rect 11622 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11378 15258
rect 11378 15206 11408 15258
rect 11432 15206 11442 15258
rect 11442 15206 11488 15258
rect 11512 15206 11558 15258
rect 11558 15206 11568 15258
rect 11592 15206 11622 15258
rect 11622 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11702 14728 11758 14784
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11378 14170
rect 11378 14118 11408 14170
rect 11432 14118 11442 14170
rect 11442 14118 11488 14170
rect 11512 14118 11558 14170
rect 11558 14118 11568 14170
rect 11592 14118 11622 14170
rect 11622 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11378 13082
rect 11378 13030 11408 13082
rect 11432 13030 11442 13082
rect 11442 13030 11488 13082
rect 11512 13030 11558 13082
rect 11558 13030 11568 13082
rect 11592 13030 11622 13082
rect 11622 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10966 11056 11022 11112
rect 10782 10648 10838 10704
rect 11242 12552 11298 12608
rect 10690 8780 10692 8800
rect 10692 8780 10744 8800
rect 10744 8780 10746 8800
rect 10690 8744 10746 8780
rect 10690 8472 10746 8528
rect 10966 7928 11022 7984
rect 11886 18536 11942 18592
rect 12346 18944 12402 19000
rect 12346 18128 12402 18184
rect 12622 17992 12678 18048
rect 12346 17720 12402 17776
rect 12530 17756 12532 17776
rect 12532 17756 12584 17776
rect 12584 17756 12586 17776
rect 12530 17720 12586 17756
rect 12254 17448 12310 17504
rect 12254 17332 12310 17368
rect 12254 17312 12256 17332
rect 12256 17312 12308 17332
rect 12308 17312 12310 17332
rect 13082 19760 13138 19816
rect 12806 18808 12862 18864
rect 12806 18128 12862 18184
rect 13542 19080 13598 19136
rect 12898 17720 12954 17776
rect 12530 16088 12586 16144
rect 12070 14356 12072 14376
rect 12072 14356 12124 14376
rect 12124 14356 12126 14376
rect 12070 14320 12126 14356
rect 12162 14068 12218 14104
rect 12162 14048 12164 14068
rect 12164 14048 12216 14068
rect 12216 14048 12218 14068
rect 12530 14592 12586 14648
rect 12254 13096 12310 13152
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11378 11994
rect 11378 11942 11408 11994
rect 11432 11942 11442 11994
rect 11442 11942 11488 11994
rect 11512 11942 11558 11994
rect 11558 11942 11568 11994
rect 11592 11942 11622 11994
rect 11622 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11610 11600 11666 11656
rect 12530 12960 12586 13016
rect 12162 12280 12218 12336
rect 12162 11736 12218 11792
rect 13358 13912 13414 13968
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11378 10906
rect 11378 10854 11408 10906
rect 11432 10854 11442 10906
rect 11442 10854 11488 10906
rect 11512 10854 11558 10906
rect 11558 10854 11568 10906
rect 11592 10854 11622 10906
rect 11622 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11378 9818
rect 11378 9766 11408 9818
rect 11432 9766 11442 9818
rect 11442 9766 11488 9818
rect 11512 9766 11558 9818
rect 11558 9766 11568 9818
rect 11592 9766 11622 9818
rect 11622 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11794 9424 11850 9480
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11378 8730
rect 11378 8678 11408 8730
rect 11432 8678 11442 8730
rect 11442 8678 11488 8730
rect 11512 8678 11558 8730
rect 11558 8678 11568 8730
rect 11592 8678 11622 8730
rect 11622 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11794 7964 11796 7984
rect 11796 7964 11848 7984
rect 11848 7964 11850 7984
rect 11794 7928 11850 7964
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11378 7642
rect 11378 7590 11408 7642
rect 11432 7590 11442 7642
rect 11442 7590 11488 7642
rect 11512 7590 11558 7642
rect 11558 7590 11568 7642
rect 11592 7590 11622 7642
rect 11622 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 10874 5888 10930 5944
rect 10874 5344 10930 5400
rect 10598 4392 10654 4448
rect 10690 3304 10746 3360
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11378 6554
rect 11378 6502 11408 6554
rect 11432 6502 11442 6554
rect 11442 6502 11488 6554
rect 11512 6502 11558 6554
rect 11558 6502 11568 6554
rect 11592 6502 11622 6554
rect 11622 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11378 5466
rect 11378 5414 11408 5466
rect 11432 5414 11442 5466
rect 11442 5414 11488 5466
rect 11512 5414 11558 5466
rect 11558 5414 11568 5466
rect 11592 5414 11622 5466
rect 11622 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11378 4378
rect 11378 4326 11408 4378
rect 11432 4326 11442 4378
rect 11442 4326 11488 4378
rect 11512 4326 11558 4378
rect 11558 4326 11568 4378
rect 11592 4326 11622 4378
rect 11622 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11886 4936 11942 4992
rect 12254 10648 12310 10704
rect 12438 10412 12440 10432
rect 12440 10412 12492 10432
rect 12492 10412 12494 10432
rect 12438 10376 12494 10412
rect 12070 4972 12072 4992
rect 12072 4972 12124 4992
rect 12124 4972 12126 4992
rect 12070 4936 12126 4972
rect 12070 3984 12126 4040
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11378 3290
rect 11378 3238 11408 3290
rect 11432 3238 11442 3290
rect 11442 3238 11488 3290
rect 11512 3238 11558 3290
rect 11558 3238 11568 3290
rect 11592 3238 11622 3290
rect 11622 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12070 3884 12072 3904
rect 12072 3884 12124 3904
rect 12124 3884 12126 3904
rect 12070 3848 12126 3884
rect 12254 9016 12310 9072
rect 12530 9424 12586 9480
rect 13542 18420 13598 18456
rect 13542 18400 13544 18420
rect 13544 18400 13596 18420
rect 13596 18400 13598 18420
rect 14817 20154 14873 20156
rect 14897 20154 14953 20156
rect 14977 20154 15033 20156
rect 15057 20154 15113 20156
rect 14817 20102 14843 20154
rect 14843 20102 14873 20154
rect 14897 20102 14907 20154
rect 14907 20102 14953 20154
rect 14977 20102 15023 20154
rect 15023 20102 15033 20154
rect 15057 20102 15087 20154
rect 15087 20102 15113 20154
rect 14817 20100 14873 20102
rect 14897 20100 14953 20102
rect 14977 20100 15033 20102
rect 15057 20100 15113 20102
rect 14002 18844 14004 18864
rect 14004 18844 14056 18864
rect 14056 18844 14058 18864
rect 14002 18808 14058 18844
rect 13634 16496 13690 16552
rect 13726 16360 13782 16416
rect 14278 17992 14334 18048
rect 13910 14340 13966 14376
rect 13910 14320 13912 14340
rect 13912 14320 13964 14340
rect 13964 14320 13966 14340
rect 13726 12316 13728 12336
rect 13728 12316 13780 12336
rect 13780 12316 13782 12336
rect 13726 12280 13782 12316
rect 13726 12164 13782 12200
rect 13726 12144 13728 12164
rect 13728 12144 13780 12164
rect 13780 12144 13782 12164
rect 14278 12144 14334 12200
rect 14186 11872 14242 11928
rect 14462 18028 14464 18048
rect 14464 18028 14516 18048
rect 14516 18028 14518 18048
rect 14462 17992 14518 18028
rect 14738 19352 14794 19408
rect 14817 19066 14873 19068
rect 14897 19066 14953 19068
rect 14977 19066 15033 19068
rect 15057 19066 15113 19068
rect 14817 19014 14843 19066
rect 14843 19014 14873 19066
rect 14897 19014 14907 19066
rect 14907 19014 14953 19066
rect 14977 19014 15023 19066
rect 15023 19014 15033 19066
rect 15057 19014 15087 19066
rect 15087 19014 15113 19066
rect 14817 19012 14873 19014
rect 14897 19012 14953 19014
rect 14977 19012 15033 19014
rect 15057 19012 15113 19014
rect 19246 22616 19302 22672
rect 18602 21664 18658 21720
rect 18282 20698 18338 20700
rect 18362 20698 18418 20700
rect 18442 20698 18498 20700
rect 18522 20698 18578 20700
rect 18282 20646 18308 20698
rect 18308 20646 18338 20698
rect 18362 20646 18372 20698
rect 18372 20646 18418 20698
rect 18442 20646 18488 20698
rect 18488 20646 18498 20698
rect 18522 20646 18552 20698
rect 18552 20646 18578 20698
rect 18282 20644 18338 20646
rect 18362 20644 18418 20646
rect 18442 20644 18498 20646
rect 18522 20644 18578 20646
rect 18970 21256 19026 21312
rect 14554 17448 14610 17504
rect 14817 17978 14873 17980
rect 14897 17978 14953 17980
rect 14977 17978 15033 17980
rect 15057 17978 15113 17980
rect 14817 17926 14843 17978
rect 14843 17926 14873 17978
rect 14897 17926 14907 17978
rect 14907 17926 14953 17978
rect 14977 17926 15023 17978
rect 15023 17926 15033 17978
rect 15057 17926 15087 17978
rect 15087 17926 15113 17978
rect 14817 17924 14873 17926
rect 14897 17924 14953 17926
rect 14977 17924 15033 17926
rect 15057 17924 15113 17926
rect 16026 18164 16028 18184
rect 16028 18164 16080 18184
rect 16080 18164 16082 18184
rect 16026 18128 16082 18164
rect 15198 17756 15200 17776
rect 15200 17756 15252 17776
rect 15252 17756 15254 17776
rect 15198 17720 15254 17756
rect 15382 17720 15438 17776
rect 14462 16496 14518 16552
rect 14817 16890 14873 16892
rect 14897 16890 14953 16892
rect 14977 16890 15033 16892
rect 15057 16890 15113 16892
rect 14817 16838 14843 16890
rect 14843 16838 14873 16890
rect 14897 16838 14907 16890
rect 14907 16838 14953 16890
rect 14977 16838 15023 16890
rect 15023 16838 15033 16890
rect 15057 16838 15087 16890
rect 15087 16838 15113 16890
rect 14817 16836 14873 16838
rect 14897 16836 14953 16838
rect 14977 16836 15033 16838
rect 15057 16836 15113 16838
rect 15382 17312 15438 17368
rect 15198 16496 15254 16552
rect 15842 16360 15898 16416
rect 14817 15802 14873 15804
rect 14897 15802 14953 15804
rect 14977 15802 15033 15804
rect 15057 15802 15113 15804
rect 14817 15750 14843 15802
rect 14843 15750 14873 15802
rect 14897 15750 14907 15802
rect 14907 15750 14953 15802
rect 14977 15750 15023 15802
rect 15023 15750 15033 15802
rect 15057 15750 15087 15802
rect 15087 15750 15113 15802
rect 14817 15748 14873 15750
rect 14897 15748 14953 15750
rect 14977 15748 15033 15750
rect 15057 15748 15113 15750
rect 14817 14714 14873 14716
rect 14897 14714 14953 14716
rect 14977 14714 15033 14716
rect 15057 14714 15113 14716
rect 14817 14662 14843 14714
rect 14843 14662 14873 14714
rect 14897 14662 14907 14714
rect 14907 14662 14953 14714
rect 14977 14662 15023 14714
rect 15023 14662 15033 14714
rect 15057 14662 15087 14714
rect 15087 14662 15113 14714
rect 14817 14660 14873 14662
rect 14897 14660 14953 14662
rect 14977 14660 15033 14662
rect 15057 14660 15113 14662
rect 14370 12008 14426 12064
rect 13358 9560 13414 9616
rect 13450 9424 13506 9480
rect 12346 7520 12402 7576
rect 12254 6704 12310 6760
rect 12530 8064 12586 8120
rect 12898 8356 12954 8392
rect 12898 8336 12900 8356
rect 12900 8336 12952 8356
rect 12952 8336 12954 8356
rect 12530 6432 12586 6488
rect 12530 6160 12586 6216
rect 12254 5752 12310 5808
rect 12438 5480 12494 5536
rect 12162 3712 12218 3768
rect 12346 3576 12402 3632
rect 11794 3168 11850 3224
rect 12070 3304 12126 3360
rect 12070 3032 12126 3088
rect 12530 2896 12586 2952
rect 11794 2624 11850 2680
rect 12438 2488 12494 2544
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11378 2202
rect 11378 2150 11408 2202
rect 11432 2150 11442 2202
rect 11442 2150 11488 2202
rect 11512 2150 11558 2202
rect 11558 2150 11568 2202
rect 11592 2150 11622 2202
rect 11622 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 14462 11736 14518 11792
rect 13726 7656 13782 7712
rect 13542 7248 13598 7304
rect 12990 6160 13046 6216
rect 12898 5888 12954 5944
rect 13818 6976 13874 7032
rect 12806 3984 12862 4040
rect 13818 3848 13874 3904
rect 14370 10648 14426 10704
rect 14817 13626 14873 13628
rect 14897 13626 14953 13628
rect 14977 13626 15033 13628
rect 15057 13626 15113 13628
rect 14817 13574 14843 13626
rect 14843 13574 14873 13626
rect 14897 13574 14907 13626
rect 14907 13574 14953 13626
rect 14977 13574 15023 13626
rect 15023 13574 15033 13626
rect 15057 13574 15087 13626
rect 15087 13574 15113 13626
rect 14817 13572 14873 13574
rect 14897 13572 14953 13574
rect 14977 13572 15033 13574
rect 15057 13572 15113 13574
rect 15014 12824 15070 12880
rect 14817 12538 14873 12540
rect 14897 12538 14953 12540
rect 14977 12538 15033 12540
rect 15057 12538 15113 12540
rect 14817 12486 14843 12538
rect 14843 12486 14873 12538
rect 14897 12486 14907 12538
rect 14907 12486 14953 12538
rect 14977 12486 15023 12538
rect 15023 12486 15033 12538
rect 15057 12486 15087 12538
rect 15087 12486 15113 12538
rect 14817 12484 14873 12486
rect 14897 12484 14953 12486
rect 14977 12484 15033 12486
rect 15057 12484 15113 12486
rect 15382 14728 15438 14784
rect 15198 12280 15254 12336
rect 14817 11450 14873 11452
rect 14897 11450 14953 11452
rect 14977 11450 15033 11452
rect 15057 11450 15113 11452
rect 14817 11398 14843 11450
rect 14843 11398 14873 11450
rect 14897 11398 14907 11450
rect 14907 11398 14953 11450
rect 14977 11398 15023 11450
rect 15023 11398 15033 11450
rect 15057 11398 15087 11450
rect 15087 11398 15113 11450
rect 14817 11396 14873 11398
rect 14897 11396 14953 11398
rect 14977 11396 15033 11398
rect 15057 11396 15113 11398
rect 14817 10362 14873 10364
rect 14897 10362 14953 10364
rect 14977 10362 15033 10364
rect 15057 10362 15113 10364
rect 14817 10310 14843 10362
rect 14843 10310 14873 10362
rect 14897 10310 14907 10362
rect 14907 10310 14953 10362
rect 14977 10310 15023 10362
rect 15023 10310 15033 10362
rect 15057 10310 15087 10362
rect 15087 10310 15113 10362
rect 14817 10308 14873 10310
rect 14897 10308 14953 10310
rect 14977 10308 15033 10310
rect 15057 10308 15113 10310
rect 14817 9274 14873 9276
rect 14897 9274 14953 9276
rect 14977 9274 15033 9276
rect 15057 9274 15113 9276
rect 14817 9222 14843 9274
rect 14843 9222 14873 9274
rect 14897 9222 14907 9274
rect 14907 9222 14953 9274
rect 14977 9222 15023 9274
rect 15023 9222 15033 9274
rect 15057 9222 15087 9274
rect 15087 9222 15113 9274
rect 14817 9220 14873 9222
rect 14897 9220 14953 9222
rect 14977 9220 15033 9222
rect 15057 9220 15113 9222
rect 14738 8472 14794 8528
rect 14554 8236 14556 8256
rect 14556 8236 14608 8256
rect 14608 8236 14610 8256
rect 14554 8200 14610 8236
rect 14817 8186 14873 8188
rect 14897 8186 14953 8188
rect 14977 8186 15033 8188
rect 15057 8186 15113 8188
rect 14817 8134 14843 8186
rect 14843 8134 14873 8186
rect 14897 8134 14907 8186
rect 14907 8134 14953 8186
rect 14977 8134 15023 8186
rect 15023 8134 15033 8186
rect 15057 8134 15087 8186
rect 15087 8134 15113 8186
rect 14817 8132 14873 8134
rect 14897 8132 14953 8134
rect 14977 8132 15033 8134
rect 15057 8132 15113 8134
rect 15658 15544 15714 15600
rect 16210 15952 16266 16008
rect 17038 18400 17094 18456
rect 17222 17740 17278 17776
rect 17222 17720 17224 17740
rect 17224 17720 17276 17740
rect 17276 17720 17278 17740
rect 17222 17448 17278 17504
rect 16026 15408 16082 15464
rect 15842 14320 15898 14376
rect 15290 10376 15346 10432
rect 15290 9016 15346 9072
rect 16762 13096 16818 13152
rect 16578 12300 16634 12336
rect 16578 12280 16580 12300
rect 16580 12280 16632 12300
rect 16632 12280 16634 12300
rect 15474 9016 15530 9072
rect 15198 7928 15254 7984
rect 15198 7112 15254 7168
rect 14817 7098 14873 7100
rect 14897 7098 14953 7100
rect 14977 7098 15033 7100
rect 15057 7098 15113 7100
rect 14817 7046 14843 7098
rect 14843 7046 14873 7098
rect 14897 7046 14907 7098
rect 14907 7046 14953 7098
rect 14977 7046 15023 7098
rect 15023 7046 15033 7098
rect 15057 7046 15087 7098
rect 15087 7046 15113 7098
rect 14817 7044 14873 7046
rect 14897 7044 14953 7046
rect 14977 7044 15033 7046
rect 15057 7044 15113 7046
rect 14278 6568 14334 6624
rect 14462 6568 14518 6624
rect 14554 6024 14610 6080
rect 15106 6704 15162 6760
rect 14830 6160 14886 6216
rect 14817 6010 14873 6012
rect 14897 6010 14953 6012
rect 14977 6010 15033 6012
rect 15057 6010 15113 6012
rect 14817 5958 14843 6010
rect 14843 5958 14873 6010
rect 14897 5958 14907 6010
rect 14907 5958 14953 6010
rect 14977 5958 15023 6010
rect 15023 5958 15033 6010
rect 15057 5958 15087 6010
rect 15087 5958 15113 6010
rect 14817 5956 14873 5958
rect 14897 5956 14953 5958
rect 14977 5956 15033 5958
rect 15057 5956 15113 5958
rect 16486 7248 16542 7304
rect 15566 5772 15622 5808
rect 15566 5752 15568 5772
rect 15568 5752 15620 5772
rect 15620 5752 15622 5772
rect 14817 4922 14873 4924
rect 14897 4922 14953 4924
rect 14977 4922 15033 4924
rect 15057 4922 15113 4924
rect 14817 4870 14843 4922
rect 14843 4870 14873 4922
rect 14897 4870 14907 4922
rect 14907 4870 14953 4922
rect 14977 4870 15023 4922
rect 15023 4870 15033 4922
rect 15057 4870 15087 4922
rect 15087 4870 15113 4922
rect 14817 4868 14873 4870
rect 14897 4868 14953 4870
rect 14977 4868 15033 4870
rect 15057 4868 15113 4870
rect 14094 2896 14150 2952
rect 14646 4528 14702 4584
rect 14817 3834 14873 3836
rect 14897 3834 14953 3836
rect 14977 3834 15033 3836
rect 15057 3834 15113 3836
rect 14817 3782 14843 3834
rect 14843 3782 14873 3834
rect 14897 3782 14907 3834
rect 14907 3782 14953 3834
rect 14977 3782 15023 3834
rect 15023 3782 15033 3834
rect 15057 3782 15087 3834
rect 15087 3782 15113 3834
rect 14817 3780 14873 3782
rect 14897 3780 14953 3782
rect 14977 3780 15033 3782
rect 15057 3780 15113 3782
rect 14817 2746 14873 2748
rect 14897 2746 14953 2748
rect 14977 2746 15033 2748
rect 15057 2746 15113 2748
rect 14817 2694 14843 2746
rect 14843 2694 14873 2746
rect 14897 2694 14907 2746
rect 14907 2694 14953 2746
rect 14977 2694 15023 2746
rect 15023 2694 15033 2746
rect 15057 2694 15087 2746
rect 15087 2694 15113 2746
rect 14817 2692 14873 2694
rect 14897 2692 14953 2694
rect 14977 2692 15033 2694
rect 15057 2692 15113 2694
rect 15290 2352 15346 2408
rect 15934 4564 15936 4584
rect 15936 4564 15988 4584
rect 15988 4564 15990 4584
rect 15934 4528 15990 4564
rect 15474 3576 15530 3632
rect 15842 3304 15898 3360
rect 16302 3168 16358 3224
rect 18510 19916 18566 19952
rect 18510 19896 18512 19916
rect 18512 19896 18564 19916
rect 18564 19896 18566 19916
rect 18282 19610 18338 19612
rect 18362 19610 18418 19612
rect 18442 19610 18498 19612
rect 18522 19610 18578 19612
rect 18282 19558 18308 19610
rect 18308 19558 18338 19610
rect 18362 19558 18372 19610
rect 18372 19558 18418 19610
rect 18442 19558 18488 19610
rect 18488 19558 18498 19610
rect 18522 19558 18552 19610
rect 18552 19558 18578 19610
rect 18282 19556 18338 19558
rect 18362 19556 18418 19558
rect 18442 19556 18498 19558
rect 18522 19556 18578 19558
rect 19522 20712 19578 20768
rect 18418 18808 18474 18864
rect 17590 18536 17646 18592
rect 17314 15000 17370 15056
rect 18282 18522 18338 18524
rect 18362 18522 18418 18524
rect 18442 18522 18498 18524
rect 18522 18522 18578 18524
rect 18282 18470 18308 18522
rect 18308 18470 18338 18522
rect 18362 18470 18372 18522
rect 18372 18470 18418 18522
rect 18442 18470 18488 18522
rect 18488 18470 18498 18522
rect 18522 18470 18552 18522
rect 18552 18470 18578 18522
rect 18282 18468 18338 18470
rect 18362 18468 18418 18470
rect 18442 18468 18498 18470
rect 18522 18468 18578 18470
rect 18282 17434 18338 17436
rect 18362 17434 18418 17436
rect 18442 17434 18498 17436
rect 18522 17434 18578 17436
rect 18282 17382 18308 17434
rect 18308 17382 18338 17434
rect 18362 17382 18372 17434
rect 18372 17382 18418 17434
rect 18442 17382 18488 17434
rect 18488 17382 18498 17434
rect 18522 17382 18552 17434
rect 18552 17382 18578 17434
rect 18282 17380 18338 17382
rect 18362 17380 18418 17382
rect 18442 17380 18498 17382
rect 18522 17380 18578 17382
rect 18602 17176 18658 17232
rect 18282 16346 18338 16348
rect 18362 16346 18418 16348
rect 18442 16346 18498 16348
rect 18522 16346 18578 16348
rect 18282 16294 18308 16346
rect 18308 16294 18338 16346
rect 18362 16294 18372 16346
rect 18372 16294 18418 16346
rect 18442 16294 18488 16346
rect 18488 16294 18498 16346
rect 18522 16294 18552 16346
rect 18552 16294 18578 16346
rect 18282 16292 18338 16294
rect 18362 16292 18418 16294
rect 18442 16292 18498 16294
rect 18522 16292 18578 16294
rect 18282 15258 18338 15260
rect 18362 15258 18418 15260
rect 18442 15258 18498 15260
rect 18522 15258 18578 15260
rect 18282 15206 18308 15258
rect 18308 15206 18338 15258
rect 18362 15206 18372 15258
rect 18372 15206 18418 15258
rect 18442 15206 18488 15258
rect 18488 15206 18498 15258
rect 18522 15206 18552 15258
rect 18552 15206 18578 15258
rect 18282 15204 18338 15206
rect 18362 15204 18418 15206
rect 18442 15204 18498 15206
rect 18522 15204 18578 15206
rect 17038 12144 17094 12200
rect 17682 13368 17738 13424
rect 17774 12280 17830 12336
rect 18282 14170 18338 14172
rect 18362 14170 18418 14172
rect 18442 14170 18498 14172
rect 18522 14170 18578 14172
rect 18282 14118 18308 14170
rect 18308 14118 18338 14170
rect 18362 14118 18372 14170
rect 18372 14118 18418 14170
rect 18442 14118 18488 14170
rect 18488 14118 18498 14170
rect 18522 14118 18552 14170
rect 18552 14118 18578 14170
rect 18282 14116 18338 14118
rect 18362 14116 18418 14118
rect 18442 14116 18498 14118
rect 18522 14116 18578 14118
rect 18142 14048 18198 14104
rect 18282 13082 18338 13084
rect 18362 13082 18418 13084
rect 18442 13082 18498 13084
rect 18522 13082 18578 13084
rect 18282 13030 18308 13082
rect 18308 13030 18338 13082
rect 18362 13030 18372 13082
rect 18372 13030 18418 13082
rect 18442 13030 18488 13082
rect 18488 13030 18498 13082
rect 18522 13030 18552 13082
rect 18552 13030 18578 13082
rect 18282 13028 18338 13030
rect 18362 13028 18418 13030
rect 18442 13028 18498 13030
rect 18522 13028 18578 13030
rect 18234 12316 18236 12336
rect 18236 12316 18288 12336
rect 18288 12316 18290 12336
rect 18234 12280 18290 12316
rect 18282 11994 18338 11996
rect 18362 11994 18418 11996
rect 18442 11994 18498 11996
rect 18522 11994 18578 11996
rect 18282 11942 18308 11994
rect 18308 11942 18338 11994
rect 18362 11942 18372 11994
rect 18372 11942 18418 11994
rect 18442 11942 18488 11994
rect 18488 11942 18498 11994
rect 18522 11942 18552 11994
rect 18552 11942 18578 11994
rect 18282 11940 18338 11942
rect 18362 11940 18418 11942
rect 18442 11940 18498 11942
rect 18522 11940 18578 11942
rect 18142 11056 18198 11112
rect 18282 10906 18338 10908
rect 18362 10906 18418 10908
rect 18442 10906 18498 10908
rect 18522 10906 18578 10908
rect 18282 10854 18308 10906
rect 18308 10854 18338 10906
rect 18362 10854 18372 10906
rect 18372 10854 18418 10906
rect 18442 10854 18488 10906
rect 18488 10854 18498 10906
rect 18522 10854 18552 10906
rect 18552 10854 18578 10906
rect 18282 10852 18338 10854
rect 18362 10852 18418 10854
rect 18442 10852 18498 10854
rect 18522 10852 18578 10854
rect 19614 18264 19670 18320
rect 19246 14764 19248 14784
rect 19248 14764 19300 14784
rect 19300 14764 19302 14784
rect 19246 14728 19302 14764
rect 19062 13232 19118 13288
rect 19154 12688 19210 12744
rect 19890 16632 19946 16688
rect 20074 18672 20130 18728
rect 20074 17584 20130 17640
rect 20442 20304 20498 20360
rect 20810 20324 20866 20360
rect 20810 20304 20812 20324
rect 20812 20304 20864 20324
rect 20864 20304 20866 20324
rect 20534 19216 20590 19272
rect 20626 17448 20682 17504
rect 20166 17040 20222 17096
rect 21454 19760 21510 19816
rect 21362 19352 21418 19408
rect 21362 18808 21418 18864
rect 21362 18400 21418 18456
rect 21362 17992 21418 18048
rect 21362 17040 21418 17096
rect 21270 16496 21326 16552
rect 20626 14864 20682 14920
rect 20534 14456 20590 14512
rect 18786 11872 18842 11928
rect 18786 11212 18842 11248
rect 18786 11192 18788 11212
rect 18788 11192 18840 11212
rect 18840 11192 18842 11212
rect 17958 9988 18014 10024
rect 17958 9968 17960 9988
rect 17960 9968 18012 9988
rect 18012 9968 18014 9988
rect 18878 10104 18934 10160
rect 18282 9818 18338 9820
rect 18362 9818 18418 9820
rect 18442 9818 18498 9820
rect 18522 9818 18578 9820
rect 18282 9766 18308 9818
rect 18308 9766 18338 9818
rect 18362 9766 18372 9818
rect 18372 9766 18418 9818
rect 18442 9766 18488 9818
rect 18488 9766 18498 9818
rect 18522 9766 18552 9818
rect 18552 9766 18578 9818
rect 18282 9764 18338 9766
rect 18362 9764 18418 9766
rect 18442 9764 18498 9766
rect 18522 9764 18578 9766
rect 18878 9696 18934 9752
rect 18282 8730 18338 8732
rect 18362 8730 18418 8732
rect 18442 8730 18498 8732
rect 18522 8730 18578 8732
rect 18282 8678 18308 8730
rect 18308 8678 18338 8730
rect 18362 8678 18372 8730
rect 18372 8678 18418 8730
rect 18442 8678 18488 8730
rect 18488 8678 18498 8730
rect 18522 8678 18552 8730
rect 18552 8678 18578 8730
rect 18282 8676 18338 8678
rect 18362 8676 18418 8678
rect 18442 8676 18498 8678
rect 18522 8676 18578 8678
rect 18786 8608 18842 8664
rect 17958 8064 18014 8120
rect 17774 7384 17830 7440
rect 17590 6568 17646 6624
rect 17314 5480 17370 5536
rect 18050 7656 18106 7712
rect 19522 10512 19578 10568
rect 18282 7642 18338 7644
rect 18362 7642 18418 7644
rect 18442 7642 18498 7644
rect 18522 7642 18578 7644
rect 18282 7590 18308 7642
rect 18308 7590 18338 7642
rect 18362 7590 18372 7642
rect 18372 7590 18418 7642
rect 18442 7590 18488 7642
rect 18488 7590 18498 7642
rect 18522 7590 18552 7642
rect 18552 7590 18578 7642
rect 18282 7588 18338 7590
rect 18362 7588 18418 7590
rect 18442 7588 18498 7590
rect 18522 7588 18578 7590
rect 19246 8880 19302 8936
rect 18282 6554 18338 6556
rect 18362 6554 18418 6556
rect 18442 6554 18498 6556
rect 18522 6554 18578 6556
rect 18282 6502 18308 6554
rect 18308 6502 18338 6554
rect 18362 6502 18372 6554
rect 18372 6502 18418 6554
rect 18442 6502 18488 6554
rect 18488 6502 18498 6554
rect 18522 6502 18552 6554
rect 18552 6502 18578 6554
rect 18282 6500 18338 6502
rect 18362 6500 18418 6502
rect 18442 6500 18498 6502
rect 18522 6500 18578 6502
rect 18694 5752 18750 5808
rect 18282 5466 18338 5468
rect 18362 5466 18418 5468
rect 18442 5466 18498 5468
rect 18522 5466 18578 5468
rect 18282 5414 18308 5466
rect 18308 5414 18338 5466
rect 18362 5414 18372 5466
rect 18372 5414 18418 5466
rect 18442 5414 18488 5466
rect 18488 5414 18498 5466
rect 18522 5414 18552 5466
rect 18552 5414 18578 5466
rect 18282 5412 18338 5414
rect 18362 5412 18418 5414
rect 18442 5412 18498 5414
rect 18522 5412 18578 5414
rect 18142 5208 18198 5264
rect 18602 4800 18658 4856
rect 18510 4684 18566 4720
rect 18510 4664 18512 4684
rect 18512 4664 18564 4684
rect 18564 4664 18566 4684
rect 18282 4378 18338 4380
rect 18362 4378 18418 4380
rect 18442 4378 18498 4380
rect 18522 4378 18578 4380
rect 18282 4326 18308 4378
rect 18308 4326 18338 4378
rect 18362 4326 18372 4378
rect 18372 4326 18418 4378
rect 18442 4326 18488 4378
rect 18488 4326 18498 4378
rect 18522 4326 18552 4378
rect 18552 4326 18578 4378
rect 18282 4324 18338 4326
rect 18362 4324 18418 4326
rect 18442 4324 18498 4326
rect 18522 4324 18578 4326
rect 18694 4392 18750 4448
rect 18282 3290 18338 3292
rect 18362 3290 18418 3292
rect 18442 3290 18498 3292
rect 18522 3290 18578 3292
rect 18282 3238 18308 3290
rect 18308 3238 18338 3290
rect 18362 3238 18372 3290
rect 18372 3238 18418 3290
rect 18442 3238 18488 3290
rect 18488 3238 18498 3290
rect 18522 3238 18552 3290
rect 18552 3238 18578 3290
rect 18282 3236 18338 3238
rect 18362 3236 18418 3238
rect 18442 3236 18498 3238
rect 18522 3236 18578 3238
rect 18786 3440 18842 3496
rect 18878 2896 18934 2952
rect 18786 2796 18788 2816
rect 18788 2796 18840 2816
rect 18840 2796 18842 2816
rect 18786 2760 18842 2796
rect 18282 2202 18338 2204
rect 18362 2202 18418 2204
rect 18442 2202 18498 2204
rect 18522 2202 18578 2204
rect 18282 2150 18308 2202
rect 18308 2150 18338 2202
rect 18362 2150 18372 2202
rect 18372 2150 18418 2202
rect 18442 2150 18488 2202
rect 18488 2150 18498 2202
rect 18522 2150 18552 2202
rect 18552 2150 18578 2202
rect 18282 2148 18338 2150
rect 18362 2148 18418 2150
rect 18442 2148 18498 2150
rect 18522 2148 18578 2150
rect 19154 4664 19210 4720
rect 19154 3576 19210 3632
rect 19062 2760 19118 2816
rect 20166 6296 20222 6352
rect 20718 9696 20774 9752
rect 21362 16088 21418 16144
rect 21362 15544 21418 15600
rect 21270 15136 21326 15192
rect 21362 14592 21418 14648
rect 21362 14184 21418 14240
rect 21362 13812 21364 13832
rect 21364 13812 21416 13832
rect 21416 13812 21418 13832
rect 21362 13776 21418 13812
rect 21362 13252 21418 13288
rect 21362 13232 21364 13252
rect 21364 13232 21416 13252
rect 21416 13232 21418 13252
rect 20626 5072 20682 5128
rect 20350 3032 20406 3088
rect 20718 3440 20774 3496
rect 19798 2916 19854 2952
rect 19798 2896 19800 2916
rect 19800 2896 19852 2916
rect 19852 2896 19854 2916
rect 19522 2508 19578 2544
rect 19522 2488 19524 2508
rect 19524 2488 19576 2508
rect 19576 2488 19578 2508
rect 20718 1944 20774 2000
rect 20902 1536 20958 1592
rect 21086 5480 21142 5536
rect 21270 2896 21326 2952
rect 21362 584 21418 640
rect 22006 992 22062 1048
rect 21914 176 21970 232
<< metal3 >>
rect 19241 22674 19307 22677
rect 22200 22674 23000 22704
rect 19241 22672 23000 22674
rect 19241 22616 19246 22672
rect 19302 22616 23000 22672
rect 19241 22614 23000 22616
rect 19241 22611 19307 22614
rect 22200 22584 23000 22614
rect 17953 22266 18019 22269
rect 22200 22266 23000 22296
rect 17953 22264 23000 22266
rect 17953 22208 17958 22264
rect 18014 22208 23000 22264
rect 17953 22206 23000 22208
rect 17953 22203 18019 22206
rect 22200 22176 23000 22206
rect 18597 21722 18663 21725
rect 22200 21722 23000 21752
rect 18597 21720 23000 21722
rect 18597 21664 18602 21720
rect 18658 21664 23000 21720
rect 18597 21662 23000 21664
rect 18597 21659 18663 21662
rect 22200 21632 23000 21662
rect 18965 21314 19031 21317
rect 22200 21314 23000 21344
rect 18965 21312 23000 21314
rect 18965 21256 18970 21312
rect 19026 21256 23000 21312
rect 18965 21254 23000 21256
rect 18965 21251 19031 21254
rect 22200 21224 23000 21254
rect 19517 20770 19583 20773
rect 22200 20770 23000 20800
rect 19517 20768 23000 20770
rect 19517 20712 19522 20768
rect 19578 20712 23000 20768
rect 19517 20710 23000 20712
rect 19517 20707 19583 20710
rect 4409 20704 4729 20705
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 20639 4729 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 18270 20704 18590 20705
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18590 20704
rect 22200 20680 23000 20710
rect 18270 20639 18590 20640
rect 10593 20498 10659 20501
rect 12249 20498 12315 20501
rect 10593 20496 12315 20498
rect 10593 20440 10598 20496
rect 10654 20440 12254 20496
rect 12310 20440 12315 20496
rect 10593 20438 12315 20440
rect 10593 20435 10659 20438
rect 12249 20435 12315 20438
rect 8845 20362 8911 20365
rect 20437 20362 20503 20365
rect 8845 20360 20503 20362
rect 8845 20304 8850 20360
rect 8906 20304 20442 20360
rect 20498 20304 20503 20360
rect 8845 20302 20503 20304
rect 8845 20299 8911 20302
rect 20437 20299 20503 20302
rect 20805 20362 20871 20365
rect 22200 20362 23000 20392
rect 20805 20360 23000 20362
rect 20805 20304 20810 20360
rect 20866 20304 23000 20360
rect 20805 20302 23000 20304
rect 20805 20299 20871 20302
rect 22200 20272 23000 20302
rect 8385 20226 8451 20229
rect 12065 20226 12131 20229
rect 8385 20224 12131 20226
rect 8385 20168 8390 20224
rect 8446 20168 12070 20224
rect 12126 20168 12131 20224
rect 8385 20166 12131 20168
rect 8385 20163 8451 20166
rect 12065 20163 12131 20166
rect 7874 20160 8194 20161
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8194 20160
rect 7874 20095 8194 20096
rect 14805 20160 15125 20161
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 20095 15125 20096
rect 9765 20090 9831 20093
rect 9765 20088 14106 20090
rect 9765 20032 9770 20088
rect 9826 20032 14106 20088
rect 9765 20030 14106 20032
rect 9765 20027 9831 20030
rect 2313 19954 2379 19957
rect 7097 19954 7163 19957
rect 2313 19952 7163 19954
rect 2313 19896 2318 19952
rect 2374 19896 7102 19952
rect 7158 19896 7163 19952
rect 2313 19894 7163 19896
rect 2313 19891 2379 19894
rect 7097 19891 7163 19894
rect 11145 19954 11211 19957
rect 11789 19954 11855 19957
rect 11145 19952 11855 19954
rect 11145 19896 11150 19952
rect 11206 19896 11794 19952
rect 11850 19896 11855 19952
rect 11145 19894 11855 19896
rect 14046 19954 14106 20030
rect 18505 19954 18571 19957
rect 14046 19952 18571 19954
rect 14046 19896 18510 19952
rect 18566 19896 18571 19952
rect 14046 19894 18571 19896
rect 11145 19891 11211 19894
rect 11789 19891 11855 19894
rect 18505 19891 18571 19894
rect 2773 19818 2839 19821
rect 13077 19818 13143 19821
rect 2773 19816 13143 19818
rect 2773 19760 2778 19816
rect 2834 19760 13082 19816
rect 13138 19760 13143 19816
rect 2773 19758 13143 19760
rect 2773 19755 2839 19758
rect 13077 19755 13143 19758
rect 21449 19818 21515 19821
rect 22200 19818 23000 19848
rect 21449 19816 23000 19818
rect 21449 19760 21454 19816
rect 21510 19760 23000 19816
rect 21449 19758 23000 19760
rect 21449 19755 21515 19758
rect 22200 19728 23000 19758
rect 6821 19682 6887 19685
rect 8109 19682 8175 19685
rect 6821 19680 8175 19682
rect 6821 19624 6826 19680
rect 6882 19624 8114 19680
rect 8170 19624 8175 19680
rect 6821 19622 8175 19624
rect 6821 19619 6887 19622
rect 8109 19619 8175 19622
rect 10041 19682 10107 19685
rect 10685 19682 10751 19685
rect 10041 19680 10751 19682
rect 10041 19624 10046 19680
rect 10102 19624 10690 19680
rect 10746 19624 10751 19680
rect 10041 19622 10751 19624
rect 10041 19619 10107 19622
rect 10685 19619 10751 19622
rect 4409 19616 4729 19617
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 19551 4729 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 18270 19616 18590 19617
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18590 19616
rect 18270 19551 18590 19552
rect 6729 19546 6795 19549
rect 7373 19546 7439 19549
rect 6729 19544 7439 19546
rect 6729 19488 6734 19544
rect 6790 19488 7378 19544
rect 7434 19488 7439 19544
rect 6729 19486 7439 19488
rect 6729 19483 6795 19486
rect 7373 19483 7439 19486
rect 9673 19410 9739 19413
rect 14733 19410 14799 19413
rect 9673 19408 14799 19410
rect 9673 19352 9678 19408
rect 9734 19352 14738 19408
rect 14794 19352 14799 19408
rect 9673 19350 14799 19352
rect 9673 19347 9739 19350
rect 14733 19347 14799 19350
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 6177 19274 6243 19277
rect 7373 19274 7439 19277
rect 8293 19274 8359 19277
rect 20529 19274 20595 19277
rect 6177 19272 7666 19274
rect 6177 19216 6182 19272
rect 6238 19216 7378 19272
rect 7434 19216 7666 19272
rect 6177 19214 7666 19216
rect 6177 19211 6243 19214
rect 7373 19211 7439 19214
rect 7606 18594 7666 19214
rect 8293 19272 20595 19274
rect 8293 19216 8298 19272
rect 8354 19216 20534 19272
rect 20590 19216 20595 19272
rect 8293 19214 20595 19216
rect 8293 19211 8359 19214
rect 20529 19211 20595 19214
rect 10777 19138 10843 19141
rect 13537 19138 13603 19141
rect 10777 19136 13603 19138
rect 10777 19080 10782 19136
rect 10838 19080 13542 19136
rect 13598 19080 13603 19136
rect 10777 19078 13603 19080
rect 10777 19075 10843 19078
rect 13537 19075 13603 19078
rect 7874 19072 8194 19073
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8194 19072
rect 7874 19007 8194 19008
rect 14805 19072 15125 19073
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 19007 15125 19008
rect 8845 19002 8911 19005
rect 12341 19002 12407 19005
rect 8845 19000 12407 19002
rect 8845 18944 8850 19000
rect 8906 18944 12346 19000
rect 12402 18944 12407 19000
rect 8845 18942 12407 18944
rect 8845 18939 8911 18942
rect 12341 18939 12407 18942
rect 9397 18866 9463 18869
rect 12801 18866 12867 18869
rect 9397 18864 12867 18866
rect 9397 18808 9402 18864
rect 9458 18808 12806 18864
rect 12862 18808 12867 18864
rect 9397 18806 12867 18808
rect 9397 18803 9463 18806
rect 12801 18803 12867 18806
rect 13997 18866 14063 18869
rect 18413 18866 18479 18869
rect 13997 18864 18479 18866
rect 13997 18808 14002 18864
rect 14058 18808 18418 18864
rect 18474 18808 18479 18864
rect 13997 18806 18479 18808
rect 13997 18803 14063 18806
rect 18413 18803 18479 18806
rect 21357 18866 21423 18869
rect 22200 18866 23000 18896
rect 21357 18864 23000 18866
rect 21357 18808 21362 18864
rect 21418 18808 23000 18864
rect 21357 18806 23000 18808
rect 21357 18803 21423 18806
rect 22200 18776 23000 18806
rect 7741 18730 7807 18733
rect 20069 18730 20135 18733
rect 7741 18728 20135 18730
rect 7741 18672 7746 18728
rect 7802 18672 20074 18728
rect 20130 18672 20135 18728
rect 7741 18670 20135 18672
rect 7741 18667 7807 18670
rect 20069 18667 20135 18670
rect 10777 18594 10843 18597
rect 7606 18592 10843 18594
rect 7606 18536 10782 18592
rect 10838 18536 10843 18592
rect 7606 18534 10843 18536
rect 10777 18531 10843 18534
rect 11881 18594 11947 18597
rect 17585 18594 17651 18597
rect 11881 18592 17651 18594
rect 11881 18536 11886 18592
rect 11942 18536 17590 18592
rect 17646 18536 17651 18592
rect 11881 18534 17651 18536
rect 11881 18531 11947 18534
rect 17585 18531 17651 18534
rect 4409 18528 4729 18529
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 18463 4729 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 18270 18528 18590 18529
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18590 18528
rect 18270 18463 18590 18464
rect 6821 18458 6887 18461
rect 9673 18458 9739 18461
rect 6821 18456 9739 18458
rect 6821 18400 6826 18456
rect 6882 18400 9678 18456
rect 9734 18400 9739 18456
rect 6821 18398 9739 18400
rect 6821 18395 6887 18398
rect 9673 18395 9739 18398
rect 13537 18458 13603 18461
rect 17033 18458 17099 18461
rect 13537 18456 17099 18458
rect 13537 18400 13542 18456
rect 13598 18400 17038 18456
rect 17094 18400 17099 18456
rect 13537 18398 17099 18400
rect 13537 18395 13603 18398
rect 17033 18395 17099 18398
rect 21357 18458 21423 18461
rect 22200 18458 23000 18488
rect 21357 18456 23000 18458
rect 21357 18400 21362 18456
rect 21418 18400 23000 18456
rect 21357 18398 23000 18400
rect 21357 18395 21423 18398
rect 22200 18368 23000 18398
rect 7465 18322 7531 18325
rect 7925 18322 7991 18325
rect 7465 18320 7991 18322
rect 7465 18264 7470 18320
rect 7526 18264 7930 18320
rect 7986 18264 7991 18320
rect 7465 18262 7991 18264
rect 7465 18259 7531 18262
rect 7925 18259 7991 18262
rect 8753 18322 8819 18325
rect 19609 18322 19675 18325
rect 8753 18320 19675 18322
rect 8753 18264 8758 18320
rect 8814 18264 19614 18320
rect 19670 18264 19675 18320
rect 8753 18262 19675 18264
rect 8753 18259 8819 18262
rect 19609 18259 19675 18262
rect 6637 18186 6703 18189
rect 8569 18186 8635 18189
rect 12341 18186 12407 18189
rect 6637 18184 12407 18186
rect 6637 18128 6642 18184
rect 6698 18128 8574 18184
rect 8630 18128 12346 18184
rect 12402 18128 12407 18184
rect 6637 18126 12407 18128
rect 6637 18123 6703 18126
rect 8569 18123 8635 18126
rect 12341 18123 12407 18126
rect 12801 18186 12867 18189
rect 16021 18186 16087 18189
rect 12801 18184 16087 18186
rect 12801 18128 12806 18184
rect 12862 18128 16026 18184
rect 16082 18128 16087 18184
rect 12801 18126 16087 18128
rect 12801 18123 12867 18126
rect 16021 18123 16087 18126
rect 8661 18050 8727 18053
rect 9622 18050 9628 18052
rect 8661 18048 9628 18050
rect 8661 17992 8666 18048
rect 8722 17992 9628 18048
rect 8661 17990 9628 17992
rect 8661 17987 8727 17990
rect 9622 17988 9628 17990
rect 9692 18050 9698 18052
rect 12617 18050 12683 18053
rect 9692 18048 12683 18050
rect 9692 17992 12622 18048
rect 12678 17992 12683 18048
rect 9692 17990 12683 17992
rect 9692 17988 9698 17990
rect 12617 17987 12683 17990
rect 14273 18050 14339 18053
rect 14457 18050 14523 18053
rect 14273 18048 14523 18050
rect 14273 17992 14278 18048
rect 14334 17992 14462 18048
rect 14518 17992 14523 18048
rect 14273 17990 14523 17992
rect 14273 17987 14339 17990
rect 14457 17987 14523 17990
rect 21357 18050 21423 18053
rect 22200 18050 23000 18080
rect 21357 18048 23000 18050
rect 21357 17992 21362 18048
rect 21418 17992 23000 18048
rect 21357 17990 23000 17992
rect 21357 17987 21423 17990
rect 7874 17984 8194 17985
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8194 17984
rect 7874 17919 8194 17920
rect 14805 17984 15125 17985
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 22200 17960 23000 17990
rect 14805 17919 15125 17920
rect 9397 17914 9463 17917
rect 9397 17912 12266 17914
rect 9397 17856 9402 17912
rect 9458 17856 12266 17912
rect 9397 17854 12266 17856
rect 9397 17851 9463 17854
rect 7373 17778 7439 17781
rect 11145 17778 11211 17781
rect 7373 17776 11211 17778
rect 7373 17720 7378 17776
rect 7434 17720 11150 17776
rect 11206 17720 11211 17776
rect 7373 17718 11211 17720
rect 7373 17715 7439 17718
rect 11145 17715 11211 17718
rect 9029 17642 9095 17645
rect 12206 17642 12266 17854
rect 12341 17778 12407 17781
rect 12525 17778 12591 17781
rect 12341 17776 12591 17778
rect 12341 17720 12346 17776
rect 12402 17720 12530 17776
rect 12586 17720 12591 17776
rect 12341 17718 12591 17720
rect 12341 17715 12407 17718
rect 12525 17715 12591 17718
rect 12893 17778 12959 17781
rect 15193 17778 15259 17781
rect 12893 17776 15259 17778
rect 12893 17720 12898 17776
rect 12954 17720 15198 17776
rect 15254 17720 15259 17776
rect 12893 17718 15259 17720
rect 12893 17715 12959 17718
rect 15193 17715 15259 17718
rect 15377 17778 15443 17781
rect 17217 17778 17283 17781
rect 15377 17776 17283 17778
rect 15377 17720 15382 17776
rect 15438 17720 17222 17776
rect 17278 17720 17283 17776
rect 15377 17718 17283 17720
rect 15377 17715 15443 17718
rect 17217 17715 17283 17718
rect 20069 17642 20135 17645
rect 9029 17640 12128 17642
rect 9029 17584 9034 17640
rect 9090 17584 12128 17640
rect 9029 17582 12128 17584
rect 12206 17640 20135 17642
rect 12206 17584 20074 17640
rect 20130 17584 20135 17640
rect 12206 17582 20135 17584
rect 9029 17579 9095 17582
rect 5257 17506 5323 17509
rect 9213 17506 9279 17509
rect 5257 17504 9279 17506
rect 5257 17448 5262 17504
rect 5318 17448 9218 17504
rect 9274 17448 9279 17504
rect 5257 17446 9279 17448
rect 12068 17506 12128 17582
rect 20069 17579 20135 17582
rect 12249 17506 12315 17509
rect 14549 17506 14615 17509
rect 17217 17506 17283 17509
rect 12068 17504 17283 17506
rect 12068 17448 12254 17504
rect 12310 17448 14554 17504
rect 14610 17448 17222 17504
rect 17278 17448 17283 17504
rect 12068 17446 17283 17448
rect 5257 17443 5323 17446
rect 9213 17443 9279 17446
rect 12249 17443 12315 17446
rect 14549 17443 14615 17446
rect 17217 17443 17283 17446
rect 20621 17506 20687 17509
rect 22200 17506 23000 17536
rect 20621 17504 23000 17506
rect 20621 17448 20626 17504
rect 20682 17448 23000 17504
rect 20621 17446 23000 17448
rect 20621 17443 20687 17446
rect 4409 17440 4729 17441
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 17375 4729 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 18270 17440 18590 17441
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18590 17440
rect 22200 17416 23000 17446
rect 18270 17375 18590 17376
rect 7005 17370 7071 17373
rect 9305 17370 9371 17373
rect 10225 17370 10291 17373
rect 7005 17368 10291 17370
rect 7005 17312 7010 17368
rect 7066 17312 9310 17368
rect 9366 17312 10230 17368
rect 10286 17312 10291 17368
rect 7005 17310 10291 17312
rect 7005 17307 7071 17310
rect 9305 17307 9371 17310
rect 10225 17307 10291 17310
rect 12249 17370 12315 17373
rect 15377 17370 15443 17373
rect 12249 17368 15443 17370
rect 12249 17312 12254 17368
rect 12310 17312 15382 17368
rect 15438 17312 15443 17368
rect 12249 17310 15443 17312
rect 12249 17307 12315 17310
rect 15377 17307 15443 17310
rect 0 17234 800 17264
rect 1577 17234 1643 17237
rect 0 17232 1643 17234
rect 0 17176 1582 17232
rect 1638 17176 1643 17232
rect 0 17174 1643 17176
rect 0 17144 800 17174
rect 1577 17171 1643 17174
rect 6361 17234 6427 17237
rect 8201 17234 8267 17237
rect 9857 17234 9923 17237
rect 6361 17232 9923 17234
rect 6361 17176 6366 17232
rect 6422 17176 8206 17232
rect 8262 17176 9862 17232
rect 9918 17176 9923 17232
rect 6361 17174 9923 17176
rect 6361 17171 6427 17174
rect 8201 17171 8267 17174
rect 9857 17171 9923 17174
rect 11053 17234 11119 17237
rect 18597 17234 18663 17237
rect 11053 17232 18663 17234
rect 11053 17176 11058 17232
rect 11114 17176 18602 17232
rect 18658 17176 18663 17232
rect 11053 17174 18663 17176
rect 11053 17171 11119 17174
rect 18597 17171 18663 17174
rect 9029 17098 9095 17101
rect 20161 17098 20227 17101
rect 9029 17096 20227 17098
rect 9029 17040 9034 17096
rect 9090 17040 20166 17096
rect 20222 17040 20227 17096
rect 9029 17038 20227 17040
rect 9029 17035 9095 17038
rect 20161 17035 20227 17038
rect 21357 17098 21423 17101
rect 22200 17098 23000 17128
rect 21357 17096 23000 17098
rect 21357 17040 21362 17096
rect 21418 17040 23000 17096
rect 21357 17038 23000 17040
rect 21357 17035 21423 17038
rect 22200 17008 23000 17038
rect 7874 16896 8194 16897
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8194 16896
rect 7874 16831 8194 16832
rect 14805 16896 15125 16897
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 16831 15125 16832
rect 7281 16826 7347 16829
rect 7598 16826 7604 16828
rect 7281 16824 7604 16826
rect 7281 16768 7286 16824
rect 7342 16768 7604 16824
rect 7281 16766 7604 16768
rect 7281 16763 7347 16766
rect 7598 16764 7604 16766
rect 7668 16764 7674 16828
rect 9397 16826 9463 16829
rect 8342 16824 9463 16826
rect 8342 16768 9402 16824
rect 9458 16768 9463 16824
rect 8342 16766 9463 16768
rect 8109 16690 8175 16693
rect 8342 16690 8402 16766
rect 9397 16763 9463 16766
rect 8109 16688 8402 16690
rect 8109 16632 8114 16688
rect 8170 16632 8402 16688
rect 8109 16630 8402 16632
rect 8569 16690 8635 16693
rect 19885 16690 19951 16693
rect 8569 16688 19951 16690
rect 8569 16632 8574 16688
rect 8630 16632 19890 16688
rect 19946 16632 19951 16688
rect 8569 16630 19951 16632
rect 8109 16627 8175 16630
rect 8569 16627 8635 16630
rect 19885 16627 19951 16630
rect 10961 16554 11027 16557
rect 13629 16554 13695 16557
rect 14457 16554 14523 16557
rect 15193 16554 15259 16557
rect 10961 16552 15259 16554
rect 10961 16496 10966 16552
rect 11022 16496 13634 16552
rect 13690 16496 14462 16552
rect 14518 16496 15198 16552
rect 15254 16496 15259 16552
rect 10961 16494 15259 16496
rect 10961 16491 11027 16494
rect 13629 16491 13695 16494
rect 14457 16491 14523 16494
rect 15193 16491 15259 16494
rect 21265 16554 21331 16557
rect 22200 16554 23000 16584
rect 21265 16552 23000 16554
rect 21265 16496 21270 16552
rect 21326 16496 23000 16552
rect 21265 16494 23000 16496
rect 21265 16491 21331 16494
rect 22200 16464 23000 16494
rect 13721 16418 13787 16421
rect 15837 16418 15903 16421
rect 13721 16416 15903 16418
rect 13721 16360 13726 16416
rect 13782 16360 15842 16416
rect 15898 16360 15903 16416
rect 13721 16358 15903 16360
rect 13721 16355 13787 16358
rect 15837 16355 15903 16358
rect 4409 16352 4729 16353
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 16287 4729 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 18270 16352 18590 16353
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18590 16352
rect 18270 16287 18590 16288
rect 10593 16146 10659 16149
rect 12525 16146 12591 16149
rect 10593 16144 12591 16146
rect 10593 16088 10598 16144
rect 10654 16088 12530 16144
rect 12586 16088 12591 16144
rect 10593 16086 12591 16088
rect 10593 16083 10659 16086
rect 12525 16083 12591 16086
rect 21357 16146 21423 16149
rect 22200 16146 23000 16176
rect 21357 16144 23000 16146
rect 21357 16088 21362 16144
rect 21418 16088 23000 16144
rect 21357 16086 23000 16088
rect 21357 16083 21423 16086
rect 22200 16056 23000 16086
rect 5717 16010 5783 16013
rect 6729 16010 6795 16013
rect 16205 16010 16271 16013
rect 5717 16008 16271 16010
rect 5717 15952 5722 16008
rect 5778 15952 6734 16008
rect 6790 15952 16210 16008
rect 16266 15952 16271 16008
rect 5717 15950 16271 15952
rect 5717 15947 5783 15950
rect 6729 15947 6795 15950
rect 16205 15947 16271 15950
rect 7874 15808 8194 15809
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8194 15808
rect 7874 15743 8194 15744
rect 14805 15808 15125 15809
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 15743 15125 15744
rect 6453 15602 6519 15605
rect 15653 15602 15719 15605
rect 6453 15600 15719 15602
rect 6453 15544 6458 15600
rect 6514 15544 15658 15600
rect 15714 15544 15719 15600
rect 6453 15542 15719 15544
rect 6453 15539 6519 15542
rect 15653 15539 15719 15542
rect 21357 15602 21423 15605
rect 22200 15602 23000 15632
rect 21357 15600 23000 15602
rect 21357 15544 21362 15600
rect 21418 15544 23000 15600
rect 21357 15542 23000 15544
rect 21357 15539 21423 15542
rect 22200 15512 23000 15542
rect 9673 15466 9739 15469
rect 9806 15466 9812 15468
rect 9673 15464 9812 15466
rect 9673 15408 9678 15464
rect 9734 15408 9812 15464
rect 9673 15406 9812 15408
rect 9673 15403 9739 15406
rect 9806 15404 9812 15406
rect 9876 15466 9882 15468
rect 10409 15466 10475 15469
rect 16021 15466 16087 15469
rect 9876 15464 16087 15466
rect 9876 15408 10414 15464
rect 10470 15408 16026 15464
rect 16082 15408 16087 15464
rect 9876 15406 16087 15408
rect 9876 15404 9882 15406
rect 10409 15403 10475 15406
rect 16021 15403 16087 15406
rect 4409 15264 4729 15265
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 15199 4729 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 18270 15264 18590 15265
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18590 15264
rect 18270 15199 18590 15200
rect 21265 15194 21331 15197
rect 22200 15194 23000 15224
rect 21265 15192 23000 15194
rect 21265 15136 21270 15192
rect 21326 15136 23000 15192
rect 21265 15134 23000 15136
rect 21265 15131 21331 15134
rect 22200 15104 23000 15134
rect 9949 15060 10015 15061
rect 9949 15056 9996 15060
rect 10060 15058 10066 15060
rect 10685 15058 10751 15061
rect 17309 15058 17375 15061
rect 9949 15000 9954 15056
rect 9949 14996 9996 15000
rect 10060 14998 10106 15058
rect 10685 15056 17375 15058
rect 10685 15000 10690 15056
rect 10746 15000 17314 15056
rect 17370 15000 17375 15056
rect 10685 14998 17375 15000
rect 10060 14996 10066 14998
rect 9949 14995 10015 14996
rect 10685 14995 10751 14998
rect 17309 14995 17375 14998
rect 7833 14922 7899 14925
rect 20621 14922 20687 14925
rect 7833 14920 20687 14922
rect 7833 14864 7838 14920
rect 7894 14864 20626 14920
rect 20682 14864 20687 14920
rect 7833 14862 20687 14864
rect 7833 14859 7899 14862
rect 20621 14859 20687 14862
rect 9673 14786 9739 14789
rect 11697 14786 11763 14789
rect 9673 14784 11763 14786
rect 9673 14728 9678 14784
rect 9734 14728 11702 14784
rect 11758 14728 11763 14784
rect 9673 14726 11763 14728
rect 9673 14723 9739 14726
rect 11697 14723 11763 14726
rect 15377 14786 15443 14789
rect 19241 14786 19307 14789
rect 15377 14784 19307 14786
rect 15377 14728 15382 14784
rect 15438 14728 19246 14784
rect 19302 14728 19307 14784
rect 15377 14726 19307 14728
rect 15377 14723 15443 14726
rect 19241 14723 19307 14726
rect 7874 14720 8194 14721
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8194 14720
rect 7874 14655 8194 14656
rect 14805 14720 15125 14721
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 14655 15125 14656
rect 9765 14650 9831 14653
rect 12525 14650 12591 14653
rect 9765 14648 12591 14650
rect 9765 14592 9770 14648
rect 9826 14592 12530 14648
rect 12586 14592 12591 14648
rect 9765 14590 12591 14592
rect 9765 14587 9831 14590
rect 12525 14587 12591 14590
rect 21357 14650 21423 14653
rect 22200 14650 23000 14680
rect 21357 14648 23000 14650
rect 21357 14592 21362 14648
rect 21418 14592 23000 14648
rect 21357 14590 23000 14592
rect 21357 14587 21423 14590
rect 22200 14560 23000 14590
rect 10593 14514 10659 14517
rect 20529 14514 20595 14517
rect 10182 14512 20595 14514
rect 10182 14456 10598 14512
rect 10654 14456 20534 14512
rect 20590 14456 20595 14512
rect 10182 14454 20595 14456
rect 8845 14378 8911 14381
rect 10182 14378 10242 14454
rect 10593 14451 10659 14454
rect 20529 14451 20595 14454
rect 12065 14378 12131 14381
rect 8845 14376 10242 14378
rect 8845 14320 8850 14376
rect 8906 14320 10242 14376
rect 8845 14318 10242 14320
rect 11102 14376 12131 14378
rect 11102 14320 12070 14376
rect 12126 14320 12131 14376
rect 11102 14318 12131 14320
rect 8845 14315 8911 14318
rect 8569 14242 8635 14245
rect 11102 14242 11162 14318
rect 12065 14315 12131 14318
rect 13905 14378 13971 14381
rect 15837 14378 15903 14381
rect 13905 14376 15903 14378
rect 13905 14320 13910 14376
rect 13966 14320 15842 14376
rect 15898 14320 15903 14376
rect 13905 14318 15903 14320
rect 13905 14315 13971 14318
rect 15837 14315 15903 14318
rect 8569 14240 11162 14242
rect 8569 14184 8574 14240
rect 8630 14184 11162 14240
rect 8569 14182 11162 14184
rect 21357 14242 21423 14245
rect 22200 14242 23000 14272
rect 21357 14240 23000 14242
rect 21357 14184 21362 14240
rect 21418 14184 23000 14240
rect 21357 14182 23000 14184
rect 8569 14179 8635 14182
rect 21357 14179 21423 14182
rect 4409 14176 4729 14177
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 14111 4729 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 18270 14176 18590 14177
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18590 14176
rect 22200 14152 23000 14182
rect 18270 14111 18590 14112
rect 9305 14106 9371 14109
rect 9622 14106 9628 14108
rect 9305 14104 9628 14106
rect 9305 14048 9310 14104
rect 9366 14048 9628 14104
rect 9305 14046 9628 14048
rect 9305 14043 9371 14046
rect 9622 14044 9628 14046
rect 9692 14044 9698 14108
rect 12157 14106 12223 14109
rect 18137 14106 18203 14109
rect 12157 14104 18203 14106
rect 12157 14048 12162 14104
rect 12218 14048 18142 14104
rect 18198 14048 18203 14104
rect 12157 14046 18203 14048
rect 12157 14043 12223 14046
rect 18137 14043 18203 14046
rect 9949 13970 10015 13973
rect 13353 13970 13419 13973
rect 9949 13968 13419 13970
rect 9949 13912 9954 13968
rect 10010 13912 13358 13968
rect 13414 13912 13419 13968
rect 9949 13910 13419 13912
rect 9949 13907 10015 13910
rect 13353 13907 13419 13910
rect 9489 13834 9555 13837
rect 9806 13834 9812 13836
rect 9489 13832 9812 13834
rect 9489 13776 9494 13832
rect 9550 13776 9812 13832
rect 9489 13774 9812 13776
rect 9489 13771 9555 13774
rect 9806 13772 9812 13774
rect 9876 13772 9882 13836
rect 21357 13834 21423 13837
rect 22200 13834 23000 13864
rect 21357 13832 23000 13834
rect 21357 13776 21362 13832
rect 21418 13776 23000 13832
rect 21357 13774 23000 13776
rect 21357 13771 21423 13774
rect 22200 13744 23000 13774
rect 9673 13698 9739 13701
rect 10317 13698 10383 13701
rect 9673 13696 10383 13698
rect 9673 13640 9678 13696
rect 9734 13640 10322 13696
rect 10378 13640 10383 13696
rect 9673 13638 10383 13640
rect 9673 13635 9739 13638
rect 10317 13635 10383 13638
rect 7874 13632 8194 13633
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8194 13632
rect 7874 13567 8194 13568
rect 14805 13632 15125 13633
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 13567 15125 13568
rect 7649 13426 7715 13429
rect 17677 13426 17743 13429
rect 7649 13424 17743 13426
rect 7649 13368 7654 13424
rect 7710 13368 17682 13424
rect 17738 13368 17743 13424
rect 7649 13366 17743 13368
rect 7649 13363 7715 13366
rect 17677 13363 17743 13366
rect 9673 13290 9739 13293
rect 19057 13290 19123 13293
rect 9673 13288 19123 13290
rect 9673 13232 9678 13288
rect 9734 13232 19062 13288
rect 19118 13232 19123 13288
rect 9673 13230 19123 13232
rect 9673 13227 9739 13230
rect 19057 13227 19123 13230
rect 21357 13290 21423 13293
rect 22200 13290 23000 13320
rect 21357 13288 23000 13290
rect 21357 13232 21362 13288
rect 21418 13232 23000 13288
rect 21357 13230 23000 13232
rect 21357 13227 21423 13230
rect 22200 13200 23000 13230
rect 12249 13154 12315 13157
rect 16757 13154 16823 13157
rect 12249 13152 16823 13154
rect 12249 13096 12254 13152
rect 12310 13096 16762 13152
rect 16818 13096 16823 13152
rect 12249 13094 16823 13096
rect 12249 13091 12315 13094
rect 16757 13091 16823 13094
rect 4409 13088 4729 13089
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 13023 4729 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 18270 13088 18590 13089
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18590 13088
rect 18270 13023 18590 13024
rect 9949 13020 10015 13021
rect 9949 13018 9996 13020
rect 9904 13016 9996 13018
rect 9904 12960 9954 13016
rect 9904 12958 9996 12960
rect 9949 12956 9996 12958
rect 10060 12956 10066 13020
rect 12525 13018 12591 13021
rect 12525 13016 15210 13018
rect 12525 12960 12530 13016
rect 12586 12960 15210 13016
rect 12525 12958 15210 12960
rect 9949 12955 10015 12956
rect 12525 12955 12591 12958
rect 9765 12882 9831 12885
rect 15009 12882 15075 12885
rect 9765 12880 15075 12882
rect 9765 12824 9770 12880
rect 9826 12824 15014 12880
rect 15070 12824 15075 12880
rect 9765 12822 15075 12824
rect 15150 12882 15210 12958
rect 22200 12882 23000 12912
rect 15150 12822 23000 12882
rect 9765 12819 9831 12822
rect 15009 12819 15075 12822
rect 22200 12792 23000 12822
rect 19149 12746 19215 12749
rect 12390 12744 19215 12746
rect 12390 12688 19154 12744
rect 19210 12688 19215 12744
rect 12390 12686 19215 12688
rect 10869 12610 10935 12613
rect 11237 12610 11303 12613
rect 12390 12610 12450 12686
rect 19149 12683 19215 12686
rect 10869 12608 12450 12610
rect 10869 12552 10874 12608
rect 10930 12552 11242 12608
rect 11298 12552 12450 12608
rect 10869 12550 12450 12552
rect 10869 12547 10935 12550
rect 11237 12547 11303 12550
rect 7874 12544 8194 12545
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8194 12544
rect 7874 12479 8194 12480
rect 14805 12544 15125 12545
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 12479 15125 12480
rect 8293 12474 8359 12477
rect 9397 12474 9463 12477
rect 8293 12472 9463 12474
rect 8293 12416 8298 12472
rect 8354 12416 9402 12472
rect 9458 12416 9463 12472
rect 8293 12414 9463 12416
rect 8293 12411 8359 12414
rect 9397 12411 9463 12414
rect 10685 12474 10751 12477
rect 10685 12472 13922 12474
rect 10685 12416 10690 12472
rect 10746 12416 13922 12472
rect 10685 12414 13922 12416
rect 10685 12411 10751 12414
rect 8109 12338 8175 12341
rect 12157 12338 12223 12341
rect 13721 12338 13787 12341
rect 8109 12336 12082 12338
rect 8109 12280 8114 12336
rect 8170 12280 12082 12336
rect 8109 12278 12082 12280
rect 8109 12275 8175 12278
rect 8753 12202 8819 12205
rect 12022 12202 12082 12278
rect 12157 12336 13787 12338
rect 12157 12280 12162 12336
rect 12218 12280 13726 12336
rect 13782 12280 13787 12336
rect 12157 12278 13787 12280
rect 13862 12338 13922 12414
rect 15193 12338 15259 12341
rect 13862 12336 15259 12338
rect 13862 12280 15198 12336
rect 15254 12280 15259 12336
rect 13862 12278 15259 12280
rect 12157 12275 12223 12278
rect 13721 12275 13787 12278
rect 15193 12275 15259 12278
rect 16573 12338 16639 12341
rect 17769 12338 17835 12341
rect 16573 12336 17835 12338
rect 16573 12280 16578 12336
rect 16634 12280 17774 12336
rect 17830 12280 17835 12336
rect 16573 12278 17835 12280
rect 16573 12275 16639 12278
rect 17769 12275 17835 12278
rect 18229 12338 18295 12341
rect 22200 12338 23000 12368
rect 18229 12336 23000 12338
rect 18229 12280 18234 12336
rect 18290 12280 23000 12336
rect 18229 12278 23000 12280
rect 18229 12275 18295 12278
rect 22200 12248 23000 12278
rect 13721 12202 13787 12205
rect 8753 12200 11898 12202
rect 8753 12144 8758 12200
rect 8814 12144 11898 12200
rect 8753 12142 11898 12144
rect 12022 12200 13787 12202
rect 12022 12144 13726 12200
rect 13782 12144 13787 12200
rect 12022 12142 13787 12144
rect 8753 12139 8819 12142
rect 11838 12066 11898 12142
rect 13721 12139 13787 12142
rect 14273 12202 14339 12205
rect 17033 12202 17099 12205
rect 14273 12200 17099 12202
rect 14273 12144 14278 12200
rect 14334 12144 17038 12200
rect 17094 12144 17099 12200
rect 14273 12142 17099 12144
rect 14273 12139 14339 12142
rect 17033 12139 17099 12142
rect 14365 12066 14431 12069
rect 11838 12064 14431 12066
rect 11838 12008 14370 12064
rect 14426 12008 14431 12064
rect 11838 12006 14431 12008
rect 14365 12003 14431 12006
rect 4409 12000 4729 12001
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 11935 4729 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 18270 12000 18590 12001
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18590 12000
rect 18270 11935 18590 11936
rect 14181 11928 14247 11933
rect 14181 11872 14186 11928
rect 14242 11872 14247 11928
rect 14181 11867 14247 11872
rect 18781 11930 18847 11933
rect 22200 11930 23000 11960
rect 18781 11928 23000 11930
rect 18781 11872 18786 11928
rect 18842 11872 23000 11928
rect 18781 11870 23000 11872
rect 18781 11867 18847 11870
rect 7741 11794 7807 11797
rect 12157 11794 12223 11797
rect 7741 11792 12223 11794
rect 7741 11736 7746 11792
rect 7802 11736 12162 11792
rect 12218 11736 12223 11792
rect 7741 11734 12223 11736
rect 14184 11794 14244 11867
rect 22200 11840 23000 11870
rect 14457 11794 14523 11797
rect 14184 11792 14523 11794
rect 14184 11736 14462 11792
rect 14518 11736 14523 11792
rect 14184 11734 14523 11736
rect 7741 11731 7807 11734
rect 12157 11731 12223 11734
rect 14457 11731 14523 11734
rect 11605 11658 11671 11661
rect 11605 11656 19350 11658
rect 11605 11600 11610 11656
rect 11666 11600 19350 11656
rect 11605 11598 19350 11600
rect 11605 11595 11671 11598
rect 7874 11456 8194 11457
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8194 11456
rect 7874 11391 8194 11392
rect 14805 11456 15125 11457
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 11391 15125 11392
rect 9029 11386 9095 11389
rect 19290 11386 19350 11598
rect 22200 11386 23000 11416
rect 9029 11384 9690 11386
rect 9029 11328 9034 11384
rect 9090 11328 9690 11384
rect 9029 11326 9690 11328
rect 19290 11326 23000 11386
rect 9029 11323 9095 11326
rect 9630 11250 9690 11326
rect 22200 11296 23000 11326
rect 18781 11250 18847 11253
rect 9630 11248 18847 11250
rect 9630 11192 18786 11248
rect 18842 11192 18847 11248
rect 9630 11190 18847 11192
rect 18781 11187 18847 11190
rect 10961 11114 11027 11117
rect 18137 11114 18203 11117
rect 10961 11112 18203 11114
rect 10961 11056 10966 11112
rect 11022 11056 18142 11112
rect 18198 11056 18203 11112
rect 10961 11054 18203 11056
rect 10961 11051 11027 11054
rect 18137 11051 18203 11054
rect 22200 10978 23000 11008
rect 19290 10918 23000 10978
rect 4409 10912 4729 10913
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 10847 4729 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 18270 10912 18590 10913
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18590 10912
rect 18270 10847 18590 10848
rect 11792 10782 14658 10842
rect 10777 10706 10843 10709
rect 11792 10706 11852 10782
rect 10777 10704 11852 10706
rect 10777 10648 10782 10704
rect 10838 10648 11852 10704
rect 10777 10646 11852 10648
rect 12249 10706 12315 10709
rect 14365 10706 14431 10709
rect 12249 10704 14431 10706
rect 12249 10648 12254 10704
rect 12310 10648 14370 10704
rect 14426 10648 14431 10704
rect 12249 10646 14431 10648
rect 14598 10706 14658 10782
rect 19290 10706 19350 10918
rect 22200 10888 23000 10918
rect 14598 10646 19350 10706
rect 10777 10643 10843 10646
rect 12249 10643 12315 10646
rect 14365 10643 14431 10646
rect 8569 10570 8635 10573
rect 19517 10570 19583 10573
rect 8569 10568 19583 10570
rect 8569 10512 8574 10568
rect 8630 10512 19522 10568
rect 19578 10512 19583 10568
rect 8569 10510 19583 10512
rect 8569 10507 8635 10510
rect 19517 10507 19583 10510
rect 8845 10434 8911 10437
rect 12433 10434 12499 10437
rect 8845 10432 12499 10434
rect 8845 10376 8850 10432
rect 8906 10376 12438 10432
rect 12494 10376 12499 10432
rect 8845 10374 12499 10376
rect 8845 10371 8911 10374
rect 12433 10371 12499 10374
rect 15285 10434 15351 10437
rect 22200 10434 23000 10464
rect 15285 10432 23000 10434
rect 15285 10376 15290 10432
rect 15346 10376 23000 10432
rect 15285 10374 23000 10376
rect 15285 10371 15351 10374
rect 7874 10368 8194 10369
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8194 10368
rect 7874 10303 8194 10304
rect 14805 10368 15125 10369
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 22200 10344 23000 10374
rect 14805 10303 15125 10304
rect 7598 10236 7604 10300
rect 7668 10298 7674 10300
rect 7741 10298 7807 10301
rect 7668 10296 7807 10298
rect 7668 10240 7746 10296
rect 7802 10240 7807 10296
rect 7668 10238 7807 10240
rect 7668 10236 7674 10238
rect 7741 10235 7807 10238
rect 9581 10162 9647 10165
rect 18873 10162 18939 10165
rect 9581 10160 18939 10162
rect 9581 10104 9586 10160
rect 9642 10104 18878 10160
rect 18934 10104 18939 10160
rect 9581 10102 18939 10104
rect 9581 10099 9647 10102
rect 18873 10099 18939 10102
rect 17953 10026 18019 10029
rect 22200 10026 23000 10056
rect 17953 10024 23000 10026
rect 17953 9968 17958 10024
rect 18014 9968 23000 10024
rect 17953 9966 23000 9968
rect 17953 9963 18019 9966
rect 22200 9936 23000 9966
rect 4409 9824 4729 9825
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 9759 4729 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 18270 9824 18590 9825
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18590 9824
rect 18270 9759 18590 9760
rect 18873 9754 18939 9757
rect 20713 9754 20779 9757
rect 18873 9752 20779 9754
rect 18873 9696 18878 9752
rect 18934 9696 20718 9752
rect 20774 9696 20779 9752
rect 18873 9694 20779 9696
rect 18873 9691 18939 9694
rect 20713 9691 20779 9694
rect 10041 9618 10107 9621
rect 13353 9618 13419 9621
rect 10041 9616 13419 9618
rect 10041 9560 10046 9616
rect 10102 9560 13358 9616
rect 13414 9560 13419 9616
rect 10041 9558 13419 9560
rect 10041 9555 10107 9558
rect 13353 9555 13419 9558
rect 11789 9482 11855 9485
rect 12525 9482 12591 9485
rect 11789 9480 12591 9482
rect 11789 9424 11794 9480
rect 11850 9424 12530 9480
rect 12586 9424 12591 9480
rect 11789 9422 12591 9424
rect 11789 9419 11855 9422
rect 12525 9419 12591 9422
rect 13445 9482 13511 9485
rect 22200 9482 23000 9512
rect 13445 9480 23000 9482
rect 13445 9424 13450 9480
rect 13506 9424 23000 9480
rect 13445 9422 23000 9424
rect 13445 9419 13511 9422
rect 22200 9392 23000 9422
rect 7874 9280 8194 9281
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8194 9280
rect 7874 9215 8194 9216
rect 14805 9280 15125 9281
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 9215 15125 9216
rect 7465 9074 7531 9077
rect 9622 9074 9628 9076
rect 7465 9072 9628 9074
rect 7465 9016 7470 9072
rect 7526 9016 9628 9072
rect 7465 9014 9628 9016
rect 7465 9011 7531 9014
rect 9622 9012 9628 9014
rect 9692 9012 9698 9076
rect 12249 9074 12315 9077
rect 15285 9074 15351 9077
rect 12249 9072 15351 9074
rect 12249 9016 12254 9072
rect 12310 9016 15290 9072
rect 15346 9016 15351 9072
rect 12249 9014 15351 9016
rect 12249 9011 12315 9014
rect 15285 9011 15351 9014
rect 15469 9074 15535 9077
rect 22200 9074 23000 9104
rect 15469 9072 23000 9074
rect 15469 9016 15474 9072
rect 15530 9016 23000 9072
rect 15469 9014 23000 9016
rect 15469 9011 15535 9014
rect 22200 8984 23000 9014
rect 7189 8938 7255 8941
rect 19241 8938 19307 8941
rect 7189 8936 19307 8938
rect 7189 8880 7194 8936
rect 7250 8880 19246 8936
rect 19302 8880 19307 8936
rect 7189 8878 19307 8880
rect 7189 8875 7255 8878
rect 19241 8875 19307 8878
rect 9489 8802 9555 8805
rect 10685 8802 10751 8805
rect 9489 8800 10751 8802
rect 9489 8744 9494 8800
rect 9550 8744 10690 8800
rect 10746 8744 10751 8800
rect 9489 8742 10751 8744
rect 9489 8739 9555 8742
rect 10685 8739 10751 8742
rect 4409 8736 4729 8737
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 8671 4729 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 18270 8736 18590 8737
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18590 8736
rect 18270 8671 18590 8672
rect 18781 8666 18847 8669
rect 22200 8666 23000 8696
rect 18781 8664 23000 8666
rect 18781 8608 18786 8664
rect 18842 8608 23000 8664
rect 18781 8606 23000 8608
rect 18781 8603 18847 8606
rect 22200 8576 23000 8606
rect 10685 8530 10751 8533
rect 14733 8530 14799 8533
rect 10685 8528 14799 8530
rect 10685 8472 10690 8528
rect 10746 8472 14738 8528
rect 14794 8472 14799 8528
rect 10685 8470 14799 8472
rect 10685 8467 10751 8470
rect 14733 8467 14799 8470
rect 10133 8394 10199 8397
rect 12893 8394 12959 8397
rect 10133 8392 12959 8394
rect 10133 8336 10138 8392
rect 10194 8336 12898 8392
rect 12954 8336 12959 8392
rect 10133 8334 12959 8336
rect 10133 8331 10199 8334
rect 12893 8331 12959 8334
rect 9949 8258 10015 8261
rect 14549 8258 14615 8261
rect 9949 8256 14615 8258
rect 9949 8200 9954 8256
rect 10010 8200 14554 8256
rect 14610 8200 14615 8256
rect 9949 8198 14615 8200
rect 9949 8195 10015 8198
rect 14549 8195 14615 8198
rect 7874 8192 8194 8193
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8194 8192
rect 7874 8127 8194 8128
rect 14805 8192 15125 8193
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 14805 8127 15125 8128
rect 12525 8122 12591 8125
rect 10964 8120 12591 8122
rect 10964 8064 12530 8120
rect 12586 8064 12591 8120
rect 10964 8062 12591 8064
rect 10964 7989 11024 8062
rect 12525 8059 12591 8062
rect 17953 8122 18019 8125
rect 22200 8122 23000 8152
rect 17953 8120 23000 8122
rect 17953 8064 17958 8120
rect 18014 8064 23000 8120
rect 17953 8062 23000 8064
rect 17953 8059 18019 8062
rect 22200 8032 23000 8062
rect 9765 7988 9831 7989
rect 9765 7986 9812 7988
rect 9720 7984 9812 7986
rect 9720 7928 9770 7984
rect 9720 7926 9812 7928
rect 9765 7924 9812 7926
rect 9876 7924 9882 7988
rect 10961 7984 11027 7989
rect 10961 7928 10966 7984
rect 11022 7928 11027 7984
rect 9765 7923 9831 7924
rect 10961 7923 11027 7928
rect 11789 7986 11855 7989
rect 15193 7986 15259 7989
rect 11789 7984 15259 7986
rect 11789 7928 11794 7984
rect 11850 7928 15198 7984
rect 15254 7928 15259 7984
rect 11789 7926 15259 7928
rect 11789 7923 11855 7926
rect 15193 7923 15259 7926
rect 9857 7850 9923 7853
rect 9857 7848 19350 7850
rect 9857 7792 9862 7848
rect 9918 7792 19350 7848
rect 9857 7790 19350 7792
rect 9857 7787 9923 7790
rect 13721 7714 13787 7717
rect 18045 7714 18111 7717
rect 13721 7712 18111 7714
rect 13721 7656 13726 7712
rect 13782 7656 18050 7712
rect 18106 7656 18111 7712
rect 13721 7654 18111 7656
rect 19290 7714 19350 7790
rect 22200 7714 23000 7744
rect 19290 7654 23000 7714
rect 13721 7651 13787 7654
rect 18045 7651 18111 7654
rect 4409 7648 4729 7649
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 7583 4729 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 18270 7648 18590 7649
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18590 7648
rect 22200 7624 23000 7654
rect 18270 7583 18590 7584
rect 12198 7516 12204 7580
rect 12268 7578 12274 7580
rect 12341 7578 12407 7581
rect 12268 7576 12407 7578
rect 12268 7520 12346 7576
rect 12402 7520 12407 7576
rect 12268 7518 12407 7520
rect 12268 7516 12274 7518
rect 12341 7515 12407 7518
rect 7189 7442 7255 7445
rect 17769 7442 17835 7445
rect 7189 7440 17835 7442
rect 7189 7384 7194 7440
rect 7250 7384 17774 7440
rect 17830 7384 17835 7440
rect 7189 7382 17835 7384
rect 7189 7379 7255 7382
rect 17769 7379 17835 7382
rect 6545 7306 6611 7309
rect 13537 7306 13603 7309
rect 16481 7306 16547 7309
rect 6545 7304 13603 7306
rect 6545 7248 6550 7304
rect 6606 7248 13542 7304
rect 13598 7248 13603 7304
rect 6545 7246 13603 7248
rect 6545 7243 6611 7246
rect 13537 7243 13603 7246
rect 14046 7304 16547 7306
rect 14046 7248 16486 7304
rect 16542 7248 16547 7304
rect 14046 7246 16547 7248
rect 9857 7170 9923 7173
rect 14046 7170 14106 7246
rect 16481 7243 16547 7246
rect 9857 7168 14106 7170
rect 9857 7112 9862 7168
rect 9918 7112 14106 7168
rect 9857 7110 14106 7112
rect 15193 7170 15259 7173
rect 22200 7170 23000 7200
rect 15193 7168 23000 7170
rect 15193 7112 15198 7168
rect 15254 7112 23000 7168
rect 15193 7110 23000 7112
rect 9857 7107 9923 7110
rect 15193 7107 15259 7110
rect 7874 7104 8194 7105
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8194 7104
rect 7874 7039 8194 7040
rect 14805 7104 15125 7105
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 22200 7080 23000 7110
rect 14805 7039 15125 7040
rect 8385 7034 8451 7037
rect 13813 7034 13879 7037
rect 8385 7032 13879 7034
rect 8385 6976 8390 7032
rect 8446 6976 13818 7032
rect 13874 6976 13879 7032
rect 8385 6974 13879 6976
rect 8385 6971 8451 6974
rect 13813 6971 13879 6974
rect 7649 6898 7715 6901
rect 7649 6896 17418 6898
rect 7649 6840 7654 6896
rect 7710 6840 17418 6896
rect 7649 6838 17418 6840
rect 7649 6835 7715 6838
rect 9673 6762 9739 6765
rect 12249 6762 12315 6765
rect 15101 6762 15167 6765
rect 9673 6760 11852 6762
rect 9673 6704 9678 6760
rect 9734 6704 11852 6760
rect 9673 6702 11852 6704
rect 9673 6699 9739 6702
rect 11792 6626 11852 6702
rect 12249 6760 15167 6762
rect 12249 6704 12254 6760
rect 12310 6704 15106 6760
rect 15162 6704 15167 6760
rect 12249 6702 15167 6704
rect 17358 6762 17418 6838
rect 22200 6762 23000 6792
rect 17358 6702 23000 6762
rect 12249 6699 12315 6702
rect 15101 6699 15167 6702
rect 22200 6672 23000 6702
rect 14273 6626 14339 6629
rect 11792 6624 14339 6626
rect 11792 6568 14278 6624
rect 14334 6568 14339 6624
rect 11792 6566 14339 6568
rect 14273 6563 14339 6566
rect 14457 6626 14523 6629
rect 17585 6626 17651 6629
rect 14457 6624 17651 6626
rect 14457 6568 14462 6624
rect 14518 6568 17590 6624
rect 17646 6568 17651 6624
rect 14457 6566 17651 6568
rect 14457 6563 14523 6566
rect 17585 6563 17651 6566
rect 4409 6560 4729 6561
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 6495 4729 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 18270 6560 18590 6561
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18590 6560
rect 18270 6495 18590 6496
rect 12525 6490 12591 6493
rect 12525 6488 17970 6490
rect 12525 6432 12530 6488
rect 12586 6432 17970 6488
rect 12525 6430 17970 6432
rect 12525 6427 12591 6430
rect 8109 6354 8175 6357
rect 17910 6354 17970 6430
rect 20161 6354 20227 6357
rect 8109 6352 17418 6354
rect 8109 6296 8114 6352
rect 8170 6296 17418 6352
rect 8109 6294 17418 6296
rect 17910 6352 20227 6354
rect 17910 6296 20166 6352
rect 20222 6296 20227 6352
rect 17910 6294 20227 6296
rect 8109 6291 8175 6294
rect 7833 6218 7899 6221
rect 12525 6218 12591 6221
rect 7833 6216 12591 6218
rect 7833 6160 7838 6216
rect 7894 6160 12530 6216
rect 12586 6160 12591 6216
rect 7833 6158 12591 6160
rect 7833 6155 7899 6158
rect 12525 6155 12591 6158
rect 12985 6218 13051 6221
rect 14825 6218 14891 6221
rect 12985 6216 14891 6218
rect 12985 6160 12990 6216
rect 13046 6160 14830 6216
rect 14886 6160 14891 6216
rect 12985 6158 14891 6160
rect 17358 6218 17418 6294
rect 20161 6291 20227 6294
rect 22200 6218 23000 6248
rect 17358 6158 23000 6218
rect 12985 6155 13051 6158
rect 14825 6155 14891 6158
rect 22200 6128 23000 6158
rect 9397 6082 9463 6085
rect 14549 6082 14615 6085
rect 9397 6080 14615 6082
rect 9397 6024 9402 6080
rect 9458 6024 14554 6080
rect 14610 6024 14615 6080
rect 9397 6022 14615 6024
rect 9397 6019 9463 6022
rect 14549 6019 14615 6022
rect 7874 6016 8194 6017
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8194 6016
rect 7874 5951 8194 5952
rect 14805 6016 15125 6017
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 5951 15125 5952
rect 10869 5946 10935 5949
rect 12893 5946 12959 5949
rect 10869 5944 12959 5946
rect 10869 5888 10874 5944
rect 10930 5888 12898 5944
rect 12954 5888 12959 5944
rect 10869 5886 12959 5888
rect 10869 5883 10935 5886
rect 12893 5883 12959 5886
rect 0 5810 800 5840
rect 1577 5810 1643 5813
rect 0 5808 1643 5810
rect 0 5752 1582 5808
rect 1638 5752 1643 5808
rect 0 5750 1643 5752
rect 0 5720 800 5750
rect 1577 5747 1643 5750
rect 6913 5810 6979 5813
rect 12249 5810 12315 5813
rect 15561 5810 15627 5813
rect 6913 5808 12315 5810
rect 6913 5752 6918 5808
rect 6974 5752 12254 5808
rect 12310 5752 12315 5808
rect 6913 5750 12315 5752
rect 6913 5747 6979 5750
rect 12249 5747 12315 5750
rect 12390 5808 15627 5810
rect 12390 5752 15566 5808
rect 15622 5752 15627 5808
rect 12390 5750 15627 5752
rect 7373 5674 7439 5677
rect 7557 5674 7623 5677
rect 10317 5674 10383 5677
rect 12390 5674 12450 5750
rect 15561 5747 15627 5750
rect 18689 5810 18755 5813
rect 22200 5810 23000 5840
rect 18689 5808 23000 5810
rect 18689 5752 18694 5808
rect 18750 5752 23000 5808
rect 18689 5750 23000 5752
rect 18689 5747 18755 5750
rect 22200 5720 23000 5750
rect 7373 5672 7482 5674
rect 7373 5616 7378 5672
rect 7434 5616 7482 5672
rect 7373 5611 7482 5616
rect 7557 5672 12450 5674
rect 7557 5616 7562 5672
rect 7618 5616 10322 5672
rect 10378 5616 12450 5672
rect 7557 5614 12450 5616
rect 18094 5614 18890 5674
rect 7557 5611 7623 5614
rect 10317 5611 10383 5614
rect 7422 5538 7482 5611
rect 9581 5538 9647 5541
rect 7422 5536 9647 5538
rect 7422 5480 9586 5536
rect 9642 5480 9647 5536
rect 7422 5478 9647 5480
rect 9581 5475 9647 5478
rect 12433 5538 12499 5541
rect 17309 5538 17375 5541
rect 12433 5536 17375 5538
rect 12433 5480 12438 5536
rect 12494 5480 17314 5536
rect 17370 5480 17375 5536
rect 12433 5478 17375 5480
rect 12433 5475 12499 5478
rect 17309 5475 17375 5478
rect 4409 5472 4729 5473
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 5407 4729 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 9857 5402 9923 5405
rect 10869 5402 10935 5405
rect 18094 5402 18154 5614
rect 18830 5538 18890 5614
rect 21081 5538 21147 5541
rect 18830 5536 21147 5538
rect 18830 5480 21086 5536
rect 21142 5480 21147 5536
rect 18830 5478 21147 5480
rect 21081 5475 21147 5478
rect 18270 5472 18590 5473
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18590 5472
rect 18270 5407 18590 5408
rect 9857 5400 10935 5402
rect 9857 5344 9862 5400
rect 9918 5344 10874 5400
rect 10930 5344 10935 5400
rect 9857 5342 10935 5344
rect 9857 5339 9923 5342
rect 10869 5339 10935 5342
rect 12390 5342 18154 5402
rect 10317 5266 10383 5269
rect 12390 5266 12450 5342
rect 10317 5264 12450 5266
rect 10317 5208 10322 5264
rect 10378 5208 12450 5264
rect 10317 5206 12450 5208
rect 18137 5266 18203 5269
rect 22200 5266 23000 5296
rect 18137 5264 23000 5266
rect 18137 5208 18142 5264
rect 18198 5208 23000 5264
rect 18137 5206 23000 5208
rect 10317 5203 10383 5206
rect 18137 5203 18203 5206
rect 22200 5176 23000 5206
rect 7649 5130 7715 5133
rect 20621 5130 20687 5133
rect 7649 5128 20687 5130
rect 7649 5072 7654 5128
rect 7710 5072 20626 5128
rect 20682 5072 20687 5128
rect 7649 5070 20687 5072
rect 7649 5067 7715 5070
rect 20621 5067 20687 5070
rect 9213 4994 9279 4997
rect 11881 4994 11947 4997
rect 9213 4992 11947 4994
rect 9213 4936 9218 4992
rect 9274 4936 11886 4992
rect 11942 4936 11947 4992
rect 9213 4934 11947 4936
rect 9213 4931 9279 4934
rect 11881 4931 11947 4934
rect 12065 4992 12131 4997
rect 12065 4936 12070 4992
rect 12126 4936 12131 4992
rect 12065 4931 12131 4936
rect 7874 4928 8194 4929
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8194 4928
rect 7874 4863 8194 4864
rect 9029 4858 9095 4861
rect 12068 4858 12128 4931
rect 14805 4928 15125 4929
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 14805 4863 15125 4864
rect 9029 4856 12128 4858
rect 9029 4800 9034 4856
rect 9090 4800 12128 4856
rect 9029 4798 12128 4800
rect 18597 4858 18663 4861
rect 22200 4858 23000 4888
rect 18597 4856 23000 4858
rect 18597 4800 18602 4856
rect 18658 4800 23000 4856
rect 18597 4798 23000 4800
rect 9029 4795 9095 4798
rect 18597 4795 18663 4798
rect 22200 4768 23000 4798
rect 8569 4722 8635 4725
rect 18505 4722 18571 4725
rect 19149 4724 19215 4725
rect 19149 4722 19196 4724
rect 8569 4720 18571 4722
rect 8569 4664 8574 4720
rect 8630 4664 18510 4720
rect 18566 4664 18571 4720
rect 8569 4662 18571 4664
rect 19104 4720 19196 4722
rect 19104 4664 19154 4720
rect 19104 4662 19196 4664
rect 8569 4659 8635 4662
rect 18505 4659 18571 4662
rect 19149 4660 19196 4662
rect 19260 4660 19266 4724
rect 19149 4659 19215 4660
rect 7281 4586 7347 4589
rect 12198 4586 12204 4588
rect 7281 4584 12204 4586
rect 7281 4528 7286 4584
rect 7342 4528 12204 4584
rect 7281 4526 12204 4528
rect 7281 4523 7347 4526
rect 12198 4524 12204 4526
rect 12268 4524 12274 4588
rect 14641 4586 14707 4589
rect 15929 4586 15995 4589
rect 14641 4584 15995 4586
rect 14641 4528 14646 4584
rect 14702 4528 15934 4584
rect 15990 4528 15995 4584
rect 14641 4526 15995 4528
rect 14641 4523 14707 4526
rect 15929 4523 15995 4526
rect 9305 4450 9371 4453
rect 10593 4450 10659 4453
rect 9305 4448 10659 4450
rect 9305 4392 9310 4448
rect 9366 4392 10598 4448
rect 10654 4392 10659 4448
rect 9305 4390 10659 4392
rect 9305 4387 9371 4390
rect 10593 4387 10659 4390
rect 18689 4450 18755 4453
rect 22200 4450 23000 4480
rect 18689 4448 23000 4450
rect 18689 4392 18694 4448
rect 18750 4392 23000 4448
rect 18689 4390 23000 4392
rect 18689 4387 18755 4390
rect 4409 4384 4729 4385
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 4319 4729 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 18270 4384 18590 4385
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18590 4384
rect 22200 4360 23000 4390
rect 18270 4319 18590 4320
rect 8017 4314 8083 4317
rect 8477 4314 8543 4317
rect 10133 4314 10199 4317
rect 8017 4312 10199 4314
rect 8017 4256 8022 4312
rect 8078 4256 8482 4312
rect 8538 4256 10138 4312
rect 10194 4256 10199 4312
rect 8017 4254 10199 4256
rect 8017 4251 8083 4254
rect 8477 4251 8543 4254
rect 10133 4251 10199 4254
rect 8937 4178 9003 4181
rect 9438 4178 9444 4180
rect 8937 4176 9444 4178
rect 8937 4120 8942 4176
rect 8998 4120 9444 4176
rect 8937 4118 9444 4120
rect 8937 4115 9003 4118
rect 9438 4116 9444 4118
rect 9508 4116 9514 4180
rect 9622 4116 9628 4180
rect 9692 4178 9698 4180
rect 9692 4118 12266 4178
rect 9692 4116 9698 4118
rect 8477 4042 8543 4045
rect 12065 4042 12131 4045
rect 8477 4040 12131 4042
rect 8477 3984 8482 4040
rect 8538 3984 12070 4040
rect 12126 3984 12131 4040
rect 8477 3982 12131 3984
rect 8477 3979 8543 3982
rect 12065 3979 12131 3982
rect 8293 3906 8359 3909
rect 12065 3906 12131 3909
rect 8293 3904 12131 3906
rect 8293 3848 8298 3904
rect 8354 3848 12070 3904
rect 12126 3848 12131 3904
rect 8293 3846 12131 3848
rect 12206 3906 12266 4118
rect 12801 4042 12867 4045
rect 12801 4040 19350 4042
rect 12801 3984 12806 4040
rect 12862 3984 19350 4040
rect 12801 3982 19350 3984
rect 12801 3979 12867 3982
rect 13813 3906 13879 3909
rect 12206 3904 13879 3906
rect 12206 3848 13818 3904
rect 13874 3848 13879 3904
rect 12206 3846 13879 3848
rect 19290 3906 19350 3982
rect 22200 3906 23000 3936
rect 19290 3846 23000 3906
rect 8293 3843 8359 3846
rect 12065 3843 12131 3846
rect 13813 3843 13879 3846
rect 7874 3840 8194 3841
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8194 3840
rect 7874 3775 8194 3776
rect 14805 3840 15125 3841
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 22200 3816 23000 3846
rect 14805 3775 15125 3776
rect 12157 3770 12223 3773
rect 8342 3768 12223 3770
rect 8342 3712 12162 3768
rect 12218 3712 12223 3768
rect 8342 3710 12223 3712
rect 7465 3634 7531 3637
rect 8342 3634 8402 3710
rect 12157 3707 12223 3710
rect 7465 3632 8402 3634
rect 7465 3576 7470 3632
rect 7526 3576 8402 3632
rect 7465 3574 8402 3576
rect 9305 3634 9371 3637
rect 12341 3634 12407 3637
rect 9305 3632 12407 3634
rect 9305 3576 9310 3632
rect 9366 3576 12346 3632
rect 12402 3576 12407 3632
rect 9305 3574 12407 3576
rect 7465 3571 7531 3574
rect 9305 3571 9371 3574
rect 12341 3571 12407 3574
rect 15469 3634 15535 3637
rect 19149 3634 19215 3637
rect 15469 3632 19215 3634
rect 15469 3576 15474 3632
rect 15530 3576 19154 3632
rect 19210 3576 19215 3632
rect 15469 3574 19215 3576
rect 15469 3571 15535 3574
rect 19149 3571 19215 3574
rect 7097 3498 7163 3501
rect 8845 3498 8911 3501
rect 7097 3496 8911 3498
rect 7097 3440 7102 3496
rect 7158 3440 8850 3496
rect 8906 3440 8911 3496
rect 7097 3438 8911 3440
rect 7097 3435 7163 3438
rect 8845 3435 8911 3438
rect 9489 3498 9555 3501
rect 18781 3498 18847 3501
rect 9489 3496 18847 3498
rect 9489 3440 9494 3496
rect 9550 3440 18786 3496
rect 18842 3440 18847 3496
rect 9489 3438 18847 3440
rect 9489 3435 9555 3438
rect 18781 3435 18847 3438
rect 20713 3498 20779 3501
rect 22200 3498 23000 3528
rect 20713 3496 23000 3498
rect 20713 3440 20718 3496
rect 20774 3440 23000 3496
rect 20713 3438 23000 3440
rect 20713 3435 20779 3438
rect 22200 3408 23000 3438
rect 7005 3362 7071 3365
rect 10685 3362 10751 3365
rect 7005 3360 10751 3362
rect 7005 3304 7010 3360
rect 7066 3304 10690 3360
rect 10746 3304 10751 3360
rect 7005 3302 10751 3304
rect 7005 3299 7071 3302
rect 10685 3299 10751 3302
rect 12065 3362 12131 3365
rect 15837 3362 15903 3365
rect 12065 3360 15903 3362
rect 12065 3304 12070 3360
rect 12126 3304 15842 3360
rect 15898 3304 15903 3360
rect 12065 3302 15903 3304
rect 12065 3299 12131 3302
rect 15837 3299 15903 3302
rect 4409 3296 4729 3297
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 3231 4729 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 18270 3296 18590 3297
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18590 3296
rect 18270 3231 18590 3232
rect 6913 3226 6979 3229
rect 10910 3226 10916 3228
rect 6913 3224 10916 3226
rect 6913 3168 6918 3224
rect 6974 3168 10916 3224
rect 6913 3166 10916 3168
rect 6913 3163 6979 3166
rect 10910 3164 10916 3166
rect 10980 3164 10986 3228
rect 11789 3226 11855 3229
rect 16297 3226 16363 3229
rect 11789 3224 16363 3226
rect 11789 3168 11794 3224
rect 11850 3168 16302 3224
rect 16358 3168 16363 3224
rect 11789 3166 16363 3168
rect 11789 3163 11855 3166
rect 16297 3163 16363 3166
rect 4429 3090 4495 3093
rect 12065 3090 12131 3093
rect 20345 3090 20411 3093
rect 4429 3088 12131 3090
rect 4429 3032 4434 3088
rect 4490 3032 12070 3088
rect 12126 3032 12131 3088
rect 4429 3030 12131 3032
rect 4429 3027 4495 3030
rect 12065 3027 12131 3030
rect 12390 3088 20411 3090
rect 12390 3032 20350 3088
rect 20406 3032 20411 3088
rect 12390 3030 20411 3032
rect 6913 2954 6979 2957
rect 7649 2954 7715 2957
rect 12390 2954 12450 3030
rect 20345 3027 20411 3030
rect 6913 2952 12450 2954
rect 6913 2896 6918 2952
rect 6974 2896 7654 2952
rect 7710 2896 12450 2952
rect 6913 2894 12450 2896
rect 12525 2954 12591 2957
rect 14089 2954 14155 2957
rect 12525 2952 14155 2954
rect 12525 2896 12530 2952
rect 12586 2896 14094 2952
rect 14150 2896 14155 2952
rect 12525 2894 14155 2896
rect 6913 2891 6979 2894
rect 7649 2891 7715 2894
rect 12525 2891 12591 2894
rect 14089 2891 14155 2894
rect 18873 2954 18939 2957
rect 19793 2954 19859 2957
rect 18873 2952 19859 2954
rect 18873 2896 18878 2952
rect 18934 2896 19798 2952
rect 19854 2896 19859 2952
rect 18873 2894 19859 2896
rect 18873 2891 18939 2894
rect 19793 2891 19859 2894
rect 21265 2954 21331 2957
rect 22200 2954 23000 2984
rect 21265 2952 23000 2954
rect 21265 2896 21270 2952
rect 21326 2896 23000 2952
rect 21265 2894 23000 2896
rect 21265 2891 21331 2894
rect 22200 2864 23000 2894
rect 8845 2818 8911 2821
rect 8845 2816 10794 2818
rect 8845 2760 8850 2816
rect 8906 2760 10794 2816
rect 8845 2758 10794 2760
rect 8845 2755 8911 2758
rect 7874 2752 8194 2753
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8194 2752
rect 7874 2687 8194 2688
rect 9489 2684 9555 2685
rect 9438 2620 9444 2684
rect 9508 2682 9555 2684
rect 9508 2680 9600 2682
rect 9550 2624 9600 2680
rect 9508 2622 9600 2624
rect 9508 2620 9555 2622
rect 9806 2620 9812 2684
rect 9876 2682 9882 2684
rect 9949 2682 10015 2685
rect 9876 2680 10015 2682
rect 9876 2624 9954 2680
rect 10010 2624 10015 2680
rect 9876 2622 10015 2624
rect 10734 2682 10794 2758
rect 10910 2756 10916 2820
rect 10980 2818 10986 2820
rect 18781 2818 18847 2821
rect 10980 2758 14658 2818
rect 10980 2756 10986 2758
rect 11789 2682 11855 2685
rect 10734 2680 11855 2682
rect 10734 2624 11794 2680
rect 11850 2624 11855 2680
rect 10734 2622 11855 2624
rect 9876 2620 9882 2622
rect 9489 2619 9555 2620
rect 9949 2619 10015 2622
rect 11789 2619 11855 2622
rect 7741 2546 7807 2549
rect 12433 2546 12499 2549
rect 7741 2544 12499 2546
rect 7741 2488 7746 2544
rect 7802 2488 12438 2544
rect 12494 2488 12499 2544
rect 7741 2486 12499 2488
rect 14598 2546 14658 2758
rect 15334 2816 18847 2818
rect 15334 2760 18786 2816
rect 18842 2760 18847 2816
rect 15334 2758 18847 2760
rect 14805 2752 15125 2753
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2687 15125 2688
rect 15334 2546 15394 2758
rect 18781 2755 18847 2758
rect 19057 2818 19123 2821
rect 19190 2818 19196 2820
rect 19057 2816 19196 2818
rect 19057 2760 19062 2816
rect 19118 2760 19196 2816
rect 19057 2758 19196 2760
rect 19057 2755 19123 2758
rect 19190 2756 19196 2758
rect 19260 2756 19266 2820
rect 14598 2486 15394 2546
rect 19517 2546 19583 2549
rect 22200 2546 23000 2576
rect 19517 2544 23000 2546
rect 19517 2488 19522 2544
rect 19578 2488 23000 2544
rect 19517 2486 23000 2488
rect 7741 2483 7807 2486
rect 12433 2483 12499 2486
rect 19517 2483 19583 2486
rect 22200 2456 23000 2486
rect 9581 2410 9647 2413
rect 15285 2410 15351 2413
rect 9581 2408 15351 2410
rect 9581 2352 9586 2408
rect 9642 2352 15290 2408
rect 15346 2352 15351 2408
rect 9581 2350 15351 2352
rect 9581 2347 9647 2350
rect 15285 2347 15351 2350
rect 4409 2208 4729 2209
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2143 4729 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 18270 2208 18590 2209
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18590 2208
rect 18270 2143 18590 2144
rect 20713 2002 20779 2005
rect 22200 2002 23000 2032
rect 20713 2000 23000 2002
rect 20713 1944 20718 2000
rect 20774 1944 23000 2000
rect 20713 1942 23000 1944
rect 20713 1939 20779 1942
rect 22200 1912 23000 1942
rect 20897 1594 20963 1597
rect 22200 1594 23000 1624
rect 20897 1592 23000 1594
rect 20897 1536 20902 1592
rect 20958 1536 23000 1592
rect 20897 1534 23000 1536
rect 20897 1531 20963 1534
rect 22200 1504 23000 1534
rect 22001 1050 22067 1053
rect 22200 1050 23000 1080
rect 22001 1048 23000 1050
rect 22001 992 22006 1048
rect 22062 992 23000 1048
rect 22001 990 23000 992
rect 22001 987 22067 990
rect 22200 960 23000 990
rect 21357 642 21423 645
rect 22200 642 23000 672
rect 21357 640 23000 642
rect 21357 584 21362 640
rect 21418 584 23000 640
rect 21357 582 23000 584
rect 21357 579 21423 582
rect 22200 552 23000 582
rect 21909 234 21975 237
rect 22200 234 23000 264
rect 21909 232 23000 234
rect 21909 176 21914 232
rect 21970 176 23000 232
rect 21909 174 23000 176
rect 21909 171 21975 174
rect 22200 144 23000 174
<< via3 >>
rect 4417 20700 4481 20704
rect 4417 20644 4421 20700
rect 4421 20644 4477 20700
rect 4477 20644 4481 20700
rect 4417 20640 4481 20644
rect 4497 20700 4561 20704
rect 4497 20644 4501 20700
rect 4501 20644 4557 20700
rect 4557 20644 4561 20700
rect 4497 20640 4561 20644
rect 4577 20700 4641 20704
rect 4577 20644 4581 20700
rect 4581 20644 4637 20700
rect 4637 20644 4641 20700
rect 4577 20640 4641 20644
rect 4657 20700 4721 20704
rect 4657 20644 4661 20700
rect 4661 20644 4717 20700
rect 4717 20644 4721 20700
rect 4657 20640 4721 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 18278 20700 18342 20704
rect 18278 20644 18282 20700
rect 18282 20644 18338 20700
rect 18338 20644 18342 20700
rect 18278 20640 18342 20644
rect 18358 20700 18422 20704
rect 18358 20644 18362 20700
rect 18362 20644 18418 20700
rect 18418 20644 18422 20700
rect 18358 20640 18422 20644
rect 18438 20700 18502 20704
rect 18438 20644 18442 20700
rect 18442 20644 18498 20700
rect 18498 20644 18502 20700
rect 18438 20640 18502 20644
rect 18518 20700 18582 20704
rect 18518 20644 18522 20700
rect 18522 20644 18578 20700
rect 18578 20644 18582 20700
rect 18518 20640 18582 20644
rect 7882 20156 7946 20160
rect 7882 20100 7886 20156
rect 7886 20100 7942 20156
rect 7942 20100 7946 20156
rect 7882 20096 7946 20100
rect 7962 20156 8026 20160
rect 7962 20100 7966 20156
rect 7966 20100 8022 20156
rect 8022 20100 8026 20156
rect 7962 20096 8026 20100
rect 8042 20156 8106 20160
rect 8042 20100 8046 20156
rect 8046 20100 8102 20156
rect 8102 20100 8106 20156
rect 8042 20096 8106 20100
rect 8122 20156 8186 20160
rect 8122 20100 8126 20156
rect 8126 20100 8182 20156
rect 8182 20100 8186 20156
rect 8122 20096 8186 20100
rect 14813 20156 14877 20160
rect 14813 20100 14817 20156
rect 14817 20100 14873 20156
rect 14873 20100 14877 20156
rect 14813 20096 14877 20100
rect 14893 20156 14957 20160
rect 14893 20100 14897 20156
rect 14897 20100 14953 20156
rect 14953 20100 14957 20156
rect 14893 20096 14957 20100
rect 14973 20156 15037 20160
rect 14973 20100 14977 20156
rect 14977 20100 15033 20156
rect 15033 20100 15037 20156
rect 14973 20096 15037 20100
rect 15053 20156 15117 20160
rect 15053 20100 15057 20156
rect 15057 20100 15113 20156
rect 15113 20100 15117 20156
rect 15053 20096 15117 20100
rect 4417 19612 4481 19616
rect 4417 19556 4421 19612
rect 4421 19556 4477 19612
rect 4477 19556 4481 19612
rect 4417 19552 4481 19556
rect 4497 19612 4561 19616
rect 4497 19556 4501 19612
rect 4501 19556 4557 19612
rect 4557 19556 4561 19612
rect 4497 19552 4561 19556
rect 4577 19612 4641 19616
rect 4577 19556 4581 19612
rect 4581 19556 4637 19612
rect 4637 19556 4641 19612
rect 4577 19552 4641 19556
rect 4657 19612 4721 19616
rect 4657 19556 4661 19612
rect 4661 19556 4717 19612
rect 4717 19556 4721 19612
rect 4657 19552 4721 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 18278 19612 18342 19616
rect 18278 19556 18282 19612
rect 18282 19556 18338 19612
rect 18338 19556 18342 19612
rect 18278 19552 18342 19556
rect 18358 19612 18422 19616
rect 18358 19556 18362 19612
rect 18362 19556 18418 19612
rect 18418 19556 18422 19612
rect 18358 19552 18422 19556
rect 18438 19612 18502 19616
rect 18438 19556 18442 19612
rect 18442 19556 18498 19612
rect 18498 19556 18502 19612
rect 18438 19552 18502 19556
rect 18518 19612 18582 19616
rect 18518 19556 18522 19612
rect 18522 19556 18578 19612
rect 18578 19556 18582 19612
rect 18518 19552 18582 19556
rect 7882 19068 7946 19072
rect 7882 19012 7886 19068
rect 7886 19012 7942 19068
rect 7942 19012 7946 19068
rect 7882 19008 7946 19012
rect 7962 19068 8026 19072
rect 7962 19012 7966 19068
rect 7966 19012 8022 19068
rect 8022 19012 8026 19068
rect 7962 19008 8026 19012
rect 8042 19068 8106 19072
rect 8042 19012 8046 19068
rect 8046 19012 8102 19068
rect 8102 19012 8106 19068
rect 8042 19008 8106 19012
rect 8122 19068 8186 19072
rect 8122 19012 8126 19068
rect 8126 19012 8182 19068
rect 8182 19012 8186 19068
rect 8122 19008 8186 19012
rect 14813 19068 14877 19072
rect 14813 19012 14817 19068
rect 14817 19012 14873 19068
rect 14873 19012 14877 19068
rect 14813 19008 14877 19012
rect 14893 19068 14957 19072
rect 14893 19012 14897 19068
rect 14897 19012 14953 19068
rect 14953 19012 14957 19068
rect 14893 19008 14957 19012
rect 14973 19068 15037 19072
rect 14973 19012 14977 19068
rect 14977 19012 15033 19068
rect 15033 19012 15037 19068
rect 14973 19008 15037 19012
rect 15053 19068 15117 19072
rect 15053 19012 15057 19068
rect 15057 19012 15113 19068
rect 15113 19012 15117 19068
rect 15053 19008 15117 19012
rect 4417 18524 4481 18528
rect 4417 18468 4421 18524
rect 4421 18468 4477 18524
rect 4477 18468 4481 18524
rect 4417 18464 4481 18468
rect 4497 18524 4561 18528
rect 4497 18468 4501 18524
rect 4501 18468 4557 18524
rect 4557 18468 4561 18524
rect 4497 18464 4561 18468
rect 4577 18524 4641 18528
rect 4577 18468 4581 18524
rect 4581 18468 4637 18524
rect 4637 18468 4641 18524
rect 4577 18464 4641 18468
rect 4657 18524 4721 18528
rect 4657 18468 4661 18524
rect 4661 18468 4717 18524
rect 4717 18468 4721 18524
rect 4657 18464 4721 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 18278 18524 18342 18528
rect 18278 18468 18282 18524
rect 18282 18468 18338 18524
rect 18338 18468 18342 18524
rect 18278 18464 18342 18468
rect 18358 18524 18422 18528
rect 18358 18468 18362 18524
rect 18362 18468 18418 18524
rect 18418 18468 18422 18524
rect 18358 18464 18422 18468
rect 18438 18524 18502 18528
rect 18438 18468 18442 18524
rect 18442 18468 18498 18524
rect 18498 18468 18502 18524
rect 18438 18464 18502 18468
rect 18518 18524 18582 18528
rect 18518 18468 18522 18524
rect 18522 18468 18578 18524
rect 18578 18468 18582 18524
rect 18518 18464 18582 18468
rect 9628 17988 9692 18052
rect 7882 17980 7946 17984
rect 7882 17924 7886 17980
rect 7886 17924 7942 17980
rect 7942 17924 7946 17980
rect 7882 17920 7946 17924
rect 7962 17980 8026 17984
rect 7962 17924 7966 17980
rect 7966 17924 8022 17980
rect 8022 17924 8026 17980
rect 7962 17920 8026 17924
rect 8042 17980 8106 17984
rect 8042 17924 8046 17980
rect 8046 17924 8102 17980
rect 8102 17924 8106 17980
rect 8042 17920 8106 17924
rect 8122 17980 8186 17984
rect 8122 17924 8126 17980
rect 8126 17924 8182 17980
rect 8182 17924 8186 17980
rect 8122 17920 8186 17924
rect 14813 17980 14877 17984
rect 14813 17924 14817 17980
rect 14817 17924 14873 17980
rect 14873 17924 14877 17980
rect 14813 17920 14877 17924
rect 14893 17980 14957 17984
rect 14893 17924 14897 17980
rect 14897 17924 14953 17980
rect 14953 17924 14957 17980
rect 14893 17920 14957 17924
rect 14973 17980 15037 17984
rect 14973 17924 14977 17980
rect 14977 17924 15033 17980
rect 15033 17924 15037 17980
rect 14973 17920 15037 17924
rect 15053 17980 15117 17984
rect 15053 17924 15057 17980
rect 15057 17924 15113 17980
rect 15113 17924 15117 17980
rect 15053 17920 15117 17924
rect 4417 17436 4481 17440
rect 4417 17380 4421 17436
rect 4421 17380 4477 17436
rect 4477 17380 4481 17436
rect 4417 17376 4481 17380
rect 4497 17436 4561 17440
rect 4497 17380 4501 17436
rect 4501 17380 4557 17436
rect 4557 17380 4561 17436
rect 4497 17376 4561 17380
rect 4577 17436 4641 17440
rect 4577 17380 4581 17436
rect 4581 17380 4637 17436
rect 4637 17380 4641 17436
rect 4577 17376 4641 17380
rect 4657 17436 4721 17440
rect 4657 17380 4661 17436
rect 4661 17380 4717 17436
rect 4717 17380 4721 17436
rect 4657 17376 4721 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 18278 17436 18342 17440
rect 18278 17380 18282 17436
rect 18282 17380 18338 17436
rect 18338 17380 18342 17436
rect 18278 17376 18342 17380
rect 18358 17436 18422 17440
rect 18358 17380 18362 17436
rect 18362 17380 18418 17436
rect 18418 17380 18422 17436
rect 18358 17376 18422 17380
rect 18438 17436 18502 17440
rect 18438 17380 18442 17436
rect 18442 17380 18498 17436
rect 18498 17380 18502 17436
rect 18438 17376 18502 17380
rect 18518 17436 18582 17440
rect 18518 17380 18522 17436
rect 18522 17380 18578 17436
rect 18578 17380 18582 17436
rect 18518 17376 18582 17380
rect 7882 16892 7946 16896
rect 7882 16836 7886 16892
rect 7886 16836 7942 16892
rect 7942 16836 7946 16892
rect 7882 16832 7946 16836
rect 7962 16892 8026 16896
rect 7962 16836 7966 16892
rect 7966 16836 8022 16892
rect 8022 16836 8026 16892
rect 7962 16832 8026 16836
rect 8042 16892 8106 16896
rect 8042 16836 8046 16892
rect 8046 16836 8102 16892
rect 8102 16836 8106 16892
rect 8042 16832 8106 16836
rect 8122 16892 8186 16896
rect 8122 16836 8126 16892
rect 8126 16836 8182 16892
rect 8182 16836 8186 16892
rect 8122 16832 8186 16836
rect 14813 16892 14877 16896
rect 14813 16836 14817 16892
rect 14817 16836 14873 16892
rect 14873 16836 14877 16892
rect 14813 16832 14877 16836
rect 14893 16892 14957 16896
rect 14893 16836 14897 16892
rect 14897 16836 14953 16892
rect 14953 16836 14957 16892
rect 14893 16832 14957 16836
rect 14973 16892 15037 16896
rect 14973 16836 14977 16892
rect 14977 16836 15033 16892
rect 15033 16836 15037 16892
rect 14973 16832 15037 16836
rect 15053 16892 15117 16896
rect 15053 16836 15057 16892
rect 15057 16836 15113 16892
rect 15113 16836 15117 16892
rect 15053 16832 15117 16836
rect 7604 16764 7668 16828
rect 4417 16348 4481 16352
rect 4417 16292 4421 16348
rect 4421 16292 4477 16348
rect 4477 16292 4481 16348
rect 4417 16288 4481 16292
rect 4497 16348 4561 16352
rect 4497 16292 4501 16348
rect 4501 16292 4557 16348
rect 4557 16292 4561 16348
rect 4497 16288 4561 16292
rect 4577 16348 4641 16352
rect 4577 16292 4581 16348
rect 4581 16292 4637 16348
rect 4637 16292 4641 16348
rect 4577 16288 4641 16292
rect 4657 16348 4721 16352
rect 4657 16292 4661 16348
rect 4661 16292 4717 16348
rect 4717 16292 4721 16348
rect 4657 16288 4721 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 18278 16348 18342 16352
rect 18278 16292 18282 16348
rect 18282 16292 18338 16348
rect 18338 16292 18342 16348
rect 18278 16288 18342 16292
rect 18358 16348 18422 16352
rect 18358 16292 18362 16348
rect 18362 16292 18418 16348
rect 18418 16292 18422 16348
rect 18358 16288 18422 16292
rect 18438 16348 18502 16352
rect 18438 16292 18442 16348
rect 18442 16292 18498 16348
rect 18498 16292 18502 16348
rect 18438 16288 18502 16292
rect 18518 16348 18582 16352
rect 18518 16292 18522 16348
rect 18522 16292 18578 16348
rect 18578 16292 18582 16348
rect 18518 16288 18582 16292
rect 7882 15804 7946 15808
rect 7882 15748 7886 15804
rect 7886 15748 7942 15804
rect 7942 15748 7946 15804
rect 7882 15744 7946 15748
rect 7962 15804 8026 15808
rect 7962 15748 7966 15804
rect 7966 15748 8022 15804
rect 8022 15748 8026 15804
rect 7962 15744 8026 15748
rect 8042 15804 8106 15808
rect 8042 15748 8046 15804
rect 8046 15748 8102 15804
rect 8102 15748 8106 15804
rect 8042 15744 8106 15748
rect 8122 15804 8186 15808
rect 8122 15748 8126 15804
rect 8126 15748 8182 15804
rect 8182 15748 8186 15804
rect 8122 15744 8186 15748
rect 14813 15804 14877 15808
rect 14813 15748 14817 15804
rect 14817 15748 14873 15804
rect 14873 15748 14877 15804
rect 14813 15744 14877 15748
rect 14893 15804 14957 15808
rect 14893 15748 14897 15804
rect 14897 15748 14953 15804
rect 14953 15748 14957 15804
rect 14893 15744 14957 15748
rect 14973 15804 15037 15808
rect 14973 15748 14977 15804
rect 14977 15748 15033 15804
rect 15033 15748 15037 15804
rect 14973 15744 15037 15748
rect 15053 15804 15117 15808
rect 15053 15748 15057 15804
rect 15057 15748 15113 15804
rect 15113 15748 15117 15804
rect 15053 15744 15117 15748
rect 9812 15404 9876 15468
rect 4417 15260 4481 15264
rect 4417 15204 4421 15260
rect 4421 15204 4477 15260
rect 4477 15204 4481 15260
rect 4417 15200 4481 15204
rect 4497 15260 4561 15264
rect 4497 15204 4501 15260
rect 4501 15204 4557 15260
rect 4557 15204 4561 15260
rect 4497 15200 4561 15204
rect 4577 15260 4641 15264
rect 4577 15204 4581 15260
rect 4581 15204 4637 15260
rect 4637 15204 4641 15260
rect 4577 15200 4641 15204
rect 4657 15260 4721 15264
rect 4657 15204 4661 15260
rect 4661 15204 4717 15260
rect 4717 15204 4721 15260
rect 4657 15200 4721 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 18278 15260 18342 15264
rect 18278 15204 18282 15260
rect 18282 15204 18338 15260
rect 18338 15204 18342 15260
rect 18278 15200 18342 15204
rect 18358 15260 18422 15264
rect 18358 15204 18362 15260
rect 18362 15204 18418 15260
rect 18418 15204 18422 15260
rect 18358 15200 18422 15204
rect 18438 15260 18502 15264
rect 18438 15204 18442 15260
rect 18442 15204 18498 15260
rect 18498 15204 18502 15260
rect 18438 15200 18502 15204
rect 18518 15260 18582 15264
rect 18518 15204 18522 15260
rect 18522 15204 18578 15260
rect 18578 15204 18582 15260
rect 18518 15200 18582 15204
rect 9996 15056 10060 15060
rect 9996 15000 10010 15056
rect 10010 15000 10060 15056
rect 9996 14996 10060 15000
rect 7882 14716 7946 14720
rect 7882 14660 7886 14716
rect 7886 14660 7942 14716
rect 7942 14660 7946 14716
rect 7882 14656 7946 14660
rect 7962 14716 8026 14720
rect 7962 14660 7966 14716
rect 7966 14660 8022 14716
rect 8022 14660 8026 14716
rect 7962 14656 8026 14660
rect 8042 14716 8106 14720
rect 8042 14660 8046 14716
rect 8046 14660 8102 14716
rect 8102 14660 8106 14716
rect 8042 14656 8106 14660
rect 8122 14716 8186 14720
rect 8122 14660 8126 14716
rect 8126 14660 8182 14716
rect 8182 14660 8186 14716
rect 8122 14656 8186 14660
rect 14813 14716 14877 14720
rect 14813 14660 14817 14716
rect 14817 14660 14873 14716
rect 14873 14660 14877 14716
rect 14813 14656 14877 14660
rect 14893 14716 14957 14720
rect 14893 14660 14897 14716
rect 14897 14660 14953 14716
rect 14953 14660 14957 14716
rect 14893 14656 14957 14660
rect 14973 14716 15037 14720
rect 14973 14660 14977 14716
rect 14977 14660 15033 14716
rect 15033 14660 15037 14716
rect 14973 14656 15037 14660
rect 15053 14716 15117 14720
rect 15053 14660 15057 14716
rect 15057 14660 15113 14716
rect 15113 14660 15117 14716
rect 15053 14656 15117 14660
rect 4417 14172 4481 14176
rect 4417 14116 4421 14172
rect 4421 14116 4477 14172
rect 4477 14116 4481 14172
rect 4417 14112 4481 14116
rect 4497 14172 4561 14176
rect 4497 14116 4501 14172
rect 4501 14116 4557 14172
rect 4557 14116 4561 14172
rect 4497 14112 4561 14116
rect 4577 14172 4641 14176
rect 4577 14116 4581 14172
rect 4581 14116 4637 14172
rect 4637 14116 4641 14172
rect 4577 14112 4641 14116
rect 4657 14172 4721 14176
rect 4657 14116 4661 14172
rect 4661 14116 4717 14172
rect 4717 14116 4721 14172
rect 4657 14112 4721 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 18278 14172 18342 14176
rect 18278 14116 18282 14172
rect 18282 14116 18338 14172
rect 18338 14116 18342 14172
rect 18278 14112 18342 14116
rect 18358 14172 18422 14176
rect 18358 14116 18362 14172
rect 18362 14116 18418 14172
rect 18418 14116 18422 14172
rect 18358 14112 18422 14116
rect 18438 14172 18502 14176
rect 18438 14116 18442 14172
rect 18442 14116 18498 14172
rect 18498 14116 18502 14172
rect 18438 14112 18502 14116
rect 18518 14172 18582 14176
rect 18518 14116 18522 14172
rect 18522 14116 18578 14172
rect 18578 14116 18582 14172
rect 18518 14112 18582 14116
rect 9628 14044 9692 14108
rect 9812 13772 9876 13836
rect 7882 13628 7946 13632
rect 7882 13572 7886 13628
rect 7886 13572 7942 13628
rect 7942 13572 7946 13628
rect 7882 13568 7946 13572
rect 7962 13628 8026 13632
rect 7962 13572 7966 13628
rect 7966 13572 8022 13628
rect 8022 13572 8026 13628
rect 7962 13568 8026 13572
rect 8042 13628 8106 13632
rect 8042 13572 8046 13628
rect 8046 13572 8102 13628
rect 8102 13572 8106 13628
rect 8042 13568 8106 13572
rect 8122 13628 8186 13632
rect 8122 13572 8126 13628
rect 8126 13572 8182 13628
rect 8182 13572 8186 13628
rect 8122 13568 8186 13572
rect 14813 13628 14877 13632
rect 14813 13572 14817 13628
rect 14817 13572 14873 13628
rect 14873 13572 14877 13628
rect 14813 13568 14877 13572
rect 14893 13628 14957 13632
rect 14893 13572 14897 13628
rect 14897 13572 14953 13628
rect 14953 13572 14957 13628
rect 14893 13568 14957 13572
rect 14973 13628 15037 13632
rect 14973 13572 14977 13628
rect 14977 13572 15033 13628
rect 15033 13572 15037 13628
rect 14973 13568 15037 13572
rect 15053 13628 15117 13632
rect 15053 13572 15057 13628
rect 15057 13572 15113 13628
rect 15113 13572 15117 13628
rect 15053 13568 15117 13572
rect 4417 13084 4481 13088
rect 4417 13028 4421 13084
rect 4421 13028 4477 13084
rect 4477 13028 4481 13084
rect 4417 13024 4481 13028
rect 4497 13084 4561 13088
rect 4497 13028 4501 13084
rect 4501 13028 4557 13084
rect 4557 13028 4561 13084
rect 4497 13024 4561 13028
rect 4577 13084 4641 13088
rect 4577 13028 4581 13084
rect 4581 13028 4637 13084
rect 4637 13028 4641 13084
rect 4577 13024 4641 13028
rect 4657 13084 4721 13088
rect 4657 13028 4661 13084
rect 4661 13028 4717 13084
rect 4717 13028 4721 13084
rect 4657 13024 4721 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 18278 13084 18342 13088
rect 18278 13028 18282 13084
rect 18282 13028 18338 13084
rect 18338 13028 18342 13084
rect 18278 13024 18342 13028
rect 18358 13084 18422 13088
rect 18358 13028 18362 13084
rect 18362 13028 18418 13084
rect 18418 13028 18422 13084
rect 18358 13024 18422 13028
rect 18438 13084 18502 13088
rect 18438 13028 18442 13084
rect 18442 13028 18498 13084
rect 18498 13028 18502 13084
rect 18438 13024 18502 13028
rect 18518 13084 18582 13088
rect 18518 13028 18522 13084
rect 18522 13028 18578 13084
rect 18578 13028 18582 13084
rect 18518 13024 18582 13028
rect 9996 13016 10060 13020
rect 9996 12960 10010 13016
rect 10010 12960 10060 13016
rect 9996 12956 10060 12960
rect 7882 12540 7946 12544
rect 7882 12484 7886 12540
rect 7886 12484 7942 12540
rect 7942 12484 7946 12540
rect 7882 12480 7946 12484
rect 7962 12540 8026 12544
rect 7962 12484 7966 12540
rect 7966 12484 8022 12540
rect 8022 12484 8026 12540
rect 7962 12480 8026 12484
rect 8042 12540 8106 12544
rect 8042 12484 8046 12540
rect 8046 12484 8102 12540
rect 8102 12484 8106 12540
rect 8042 12480 8106 12484
rect 8122 12540 8186 12544
rect 8122 12484 8126 12540
rect 8126 12484 8182 12540
rect 8182 12484 8186 12540
rect 8122 12480 8186 12484
rect 14813 12540 14877 12544
rect 14813 12484 14817 12540
rect 14817 12484 14873 12540
rect 14873 12484 14877 12540
rect 14813 12480 14877 12484
rect 14893 12540 14957 12544
rect 14893 12484 14897 12540
rect 14897 12484 14953 12540
rect 14953 12484 14957 12540
rect 14893 12480 14957 12484
rect 14973 12540 15037 12544
rect 14973 12484 14977 12540
rect 14977 12484 15033 12540
rect 15033 12484 15037 12540
rect 14973 12480 15037 12484
rect 15053 12540 15117 12544
rect 15053 12484 15057 12540
rect 15057 12484 15113 12540
rect 15113 12484 15117 12540
rect 15053 12480 15117 12484
rect 4417 11996 4481 12000
rect 4417 11940 4421 11996
rect 4421 11940 4477 11996
rect 4477 11940 4481 11996
rect 4417 11936 4481 11940
rect 4497 11996 4561 12000
rect 4497 11940 4501 11996
rect 4501 11940 4557 11996
rect 4557 11940 4561 11996
rect 4497 11936 4561 11940
rect 4577 11996 4641 12000
rect 4577 11940 4581 11996
rect 4581 11940 4637 11996
rect 4637 11940 4641 11996
rect 4577 11936 4641 11940
rect 4657 11996 4721 12000
rect 4657 11940 4661 11996
rect 4661 11940 4717 11996
rect 4717 11940 4721 11996
rect 4657 11936 4721 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 18278 11996 18342 12000
rect 18278 11940 18282 11996
rect 18282 11940 18338 11996
rect 18338 11940 18342 11996
rect 18278 11936 18342 11940
rect 18358 11996 18422 12000
rect 18358 11940 18362 11996
rect 18362 11940 18418 11996
rect 18418 11940 18422 11996
rect 18358 11936 18422 11940
rect 18438 11996 18502 12000
rect 18438 11940 18442 11996
rect 18442 11940 18498 11996
rect 18498 11940 18502 11996
rect 18438 11936 18502 11940
rect 18518 11996 18582 12000
rect 18518 11940 18522 11996
rect 18522 11940 18578 11996
rect 18578 11940 18582 11996
rect 18518 11936 18582 11940
rect 7882 11452 7946 11456
rect 7882 11396 7886 11452
rect 7886 11396 7942 11452
rect 7942 11396 7946 11452
rect 7882 11392 7946 11396
rect 7962 11452 8026 11456
rect 7962 11396 7966 11452
rect 7966 11396 8022 11452
rect 8022 11396 8026 11452
rect 7962 11392 8026 11396
rect 8042 11452 8106 11456
rect 8042 11396 8046 11452
rect 8046 11396 8102 11452
rect 8102 11396 8106 11452
rect 8042 11392 8106 11396
rect 8122 11452 8186 11456
rect 8122 11396 8126 11452
rect 8126 11396 8182 11452
rect 8182 11396 8186 11452
rect 8122 11392 8186 11396
rect 14813 11452 14877 11456
rect 14813 11396 14817 11452
rect 14817 11396 14873 11452
rect 14873 11396 14877 11452
rect 14813 11392 14877 11396
rect 14893 11452 14957 11456
rect 14893 11396 14897 11452
rect 14897 11396 14953 11452
rect 14953 11396 14957 11452
rect 14893 11392 14957 11396
rect 14973 11452 15037 11456
rect 14973 11396 14977 11452
rect 14977 11396 15033 11452
rect 15033 11396 15037 11452
rect 14973 11392 15037 11396
rect 15053 11452 15117 11456
rect 15053 11396 15057 11452
rect 15057 11396 15113 11452
rect 15113 11396 15117 11452
rect 15053 11392 15117 11396
rect 4417 10908 4481 10912
rect 4417 10852 4421 10908
rect 4421 10852 4477 10908
rect 4477 10852 4481 10908
rect 4417 10848 4481 10852
rect 4497 10908 4561 10912
rect 4497 10852 4501 10908
rect 4501 10852 4557 10908
rect 4557 10852 4561 10908
rect 4497 10848 4561 10852
rect 4577 10908 4641 10912
rect 4577 10852 4581 10908
rect 4581 10852 4637 10908
rect 4637 10852 4641 10908
rect 4577 10848 4641 10852
rect 4657 10908 4721 10912
rect 4657 10852 4661 10908
rect 4661 10852 4717 10908
rect 4717 10852 4721 10908
rect 4657 10848 4721 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 18278 10908 18342 10912
rect 18278 10852 18282 10908
rect 18282 10852 18338 10908
rect 18338 10852 18342 10908
rect 18278 10848 18342 10852
rect 18358 10908 18422 10912
rect 18358 10852 18362 10908
rect 18362 10852 18418 10908
rect 18418 10852 18422 10908
rect 18358 10848 18422 10852
rect 18438 10908 18502 10912
rect 18438 10852 18442 10908
rect 18442 10852 18498 10908
rect 18498 10852 18502 10908
rect 18438 10848 18502 10852
rect 18518 10908 18582 10912
rect 18518 10852 18522 10908
rect 18522 10852 18578 10908
rect 18578 10852 18582 10908
rect 18518 10848 18582 10852
rect 7882 10364 7946 10368
rect 7882 10308 7886 10364
rect 7886 10308 7942 10364
rect 7942 10308 7946 10364
rect 7882 10304 7946 10308
rect 7962 10364 8026 10368
rect 7962 10308 7966 10364
rect 7966 10308 8022 10364
rect 8022 10308 8026 10364
rect 7962 10304 8026 10308
rect 8042 10364 8106 10368
rect 8042 10308 8046 10364
rect 8046 10308 8102 10364
rect 8102 10308 8106 10364
rect 8042 10304 8106 10308
rect 8122 10364 8186 10368
rect 8122 10308 8126 10364
rect 8126 10308 8182 10364
rect 8182 10308 8186 10364
rect 8122 10304 8186 10308
rect 14813 10364 14877 10368
rect 14813 10308 14817 10364
rect 14817 10308 14873 10364
rect 14873 10308 14877 10364
rect 14813 10304 14877 10308
rect 14893 10364 14957 10368
rect 14893 10308 14897 10364
rect 14897 10308 14953 10364
rect 14953 10308 14957 10364
rect 14893 10304 14957 10308
rect 14973 10364 15037 10368
rect 14973 10308 14977 10364
rect 14977 10308 15033 10364
rect 15033 10308 15037 10364
rect 14973 10304 15037 10308
rect 15053 10364 15117 10368
rect 15053 10308 15057 10364
rect 15057 10308 15113 10364
rect 15113 10308 15117 10364
rect 15053 10304 15117 10308
rect 7604 10236 7668 10300
rect 4417 9820 4481 9824
rect 4417 9764 4421 9820
rect 4421 9764 4477 9820
rect 4477 9764 4481 9820
rect 4417 9760 4481 9764
rect 4497 9820 4561 9824
rect 4497 9764 4501 9820
rect 4501 9764 4557 9820
rect 4557 9764 4561 9820
rect 4497 9760 4561 9764
rect 4577 9820 4641 9824
rect 4577 9764 4581 9820
rect 4581 9764 4637 9820
rect 4637 9764 4641 9820
rect 4577 9760 4641 9764
rect 4657 9820 4721 9824
rect 4657 9764 4661 9820
rect 4661 9764 4717 9820
rect 4717 9764 4721 9820
rect 4657 9760 4721 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 18278 9820 18342 9824
rect 18278 9764 18282 9820
rect 18282 9764 18338 9820
rect 18338 9764 18342 9820
rect 18278 9760 18342 9764
rect 18358 9820 18422 9824
rect 18358 9764 18362 9820
rect 18362 9764 18418 9820
rect 18418 9764 18422 9820
rect 18358 9760 18422 9764
rect 18438 9820 18502 9824
rect 18438 9764 18442 9820
rect 18442 9764 18498 9820
rect 18498 9764 18502 9820
rect 18438 9760 18502 9764
rect 18518 9820 18582 9824
rect 18518 9764 18522 9820
rect 18522 9764 18578 9820
rect 18578 9764 18582 9820
rect 18518 9760 18582 9764
rect 7882 9276 7946 9280
rect 7882 9220 7886 9276
rect 7886 9220 7942 9276
rect 7942 9220 7946 9276
rect 7882 9216 7946 9220
rect 7962 9276 8026 9280
rect 7962 9220 7966 9276
rect 7966 9220 8022 9276
rect 8022 9220 8026 9276
rect 7962 9216 8026 9220
rect 8042 9276 8106 9280
rect 8042 9220 8046 9276
rect 8046 9220 8102 9276
rect 8102 9220 8106 9276
rect 8042 9216 8106 9220
rect 8122 9276 8186 9280
rect 8122 9220 8126 9276
rect 8126 9220 8182 9276
rect 8182 9220 8186 9276
rect 8122 9216 8186 9220
rect 14813 9276 14877 9280
rect 14813 9220 14817 9276
rect 14817 9220 14873 9276
rect 14873 9220 14877 9276
rect 14813 9216 14877 9220
rect 14893 9276 14957 9280
rect 14893 9220 14897 9276
rect 14897 9220 14953 9276
rect 14953 9220 14957 9276
rect 14893 9216 14957 9220
rect 14973 9276 15037 9280
rect 14973 9220 14977 9276
rect 14977 9220 15033 9276
rect 15033 9220 15037 9276
rect 14973 9216 15037 9220
rect 15053 9276 15117 9280
rect 15053 9220 15057 9276
rect 15057 9220 15113 9276
rect 15113 9220 15117 9276
rect 15053 9216 15117 9220
rect 9628 9012 9692 9076
rect 4417 8732 4481 8736
rect 4417 8676 4421 8732
rect 4421 8676 4477 8732
rect 4477 8676 4481 8732
rect 4417 8672 4481 8676
rect 4497 8732 4561 8736
rect 4497 8676 4501 8732
rect 4501 8676 4557 8732
rect 4557 8676 4561 8732
rect 4497 8672 4561 8676
rect 4577 8732 4641 8736
rect 4577 8676 4581 8732
rect 4581 8676 4637 8732
rect 4637 8676 4641 8732
rect 4577 8672 4641 8676
rect 4657 8732 4721 8736
rect 4657 8676 4661 8732
rect 4661 8676 4717 8732
rect 4717 8676 4721 8732
rect 4657 8672 4721 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 18278 8732 18342 8736
rect 18278 8676 18282 8732
rect 18282 8676 18338 8732
rect 18338 8676 18342 8732
rect 18278 8672 18342 8676
rect 18358 8732 18422 8736
rect 18358 8676 18362 8732
rect 18362 8676 18418 8732
rect 18418 8676 18422 8732
rect 18358 8672 18422 8676
rect 18438 8732 18502 8736
rect 18438 8676 18442 8732
rect 18442 8676 18498 8732
rect 18498 8676 18502 8732
rect 18438 8672 18502 8676
rect 18518 8732 18582 8736
rect 18518 8676 18522 8732
rect 18522 8676 18578 8732
rect 18578 8676 18582 8732
rect 18518 8672 18582 8676
rect 7882 8188 7946 8192
rect 7882 8132 7886 8188
rect 7886 8132 7942 8188
rect 7942 8132 7946 8188
rect 7882 8128 7946 8132
rect 7962 8188 8026 8192
rect 7962 8132 7966 8188
rect 7966 8132 8022 8188
rect 8022 8132 8026 8188
rect 7962 8128 8026 8132
rect 8042 8188 8106 8192
rect 8042 8132 8046 8188
rect 8046 8132 8102 8188
rect 8102 8132 8106 8188
rect 8042 8128 8106 8132
rect 8122 8188 8186 8192
rect 8122 8132 8126 8188
rect 8126 8132 8182 8188
rect 8182 8132 8186 8188
rect 8122 8128 8186 8132
rect 14813 8188 14877 8192
rect 14813 8132 14817 8188
rect 14817 8132 14873 8188
rect 14873 8132 14877 8188
rect 14813 8128 14877 8132
rect 14893 8188 14957 8192
rect 14893 8132 14897 8188
rect 14897 8132 14953 8188
rect 14953 8132 14957 8188
rect 14893 8128 14957 8132
rect 14973 8188 15037 8192
rect 14973 8132 14977 8188
rect 14977 8132 15033 8188
rect 15033 8132 15037 8188
rect 14973 8128 15037 8132
rect 15053 8188 15117 8192
rect 15053 8132 15057 8188
rect 15057 8132 15113 8188
rect 15113 8132 15117 8188
rect 15053 8128 15117 8132
rect 9812 7984 9876 7988
rect 9812 7928 9826 7984
rect 9826 7928 9876 7984
rect 9812 7924 9876 7928
rect 4417 7644 4481 7648
rect 4417 7588 4421 7644
rect 4421 7588 4477 7644
rect 4477 7588 4481 7644
rect 4417 7584 4481 7588
rect 4497 7644 4561 7648
rect 4497 7588 4501 7644
rect 4501 7588 4557 7644
rect 4557 7588 4561 7644
rect 4497 7584 4561 7588
rect 4577 7644 4641 7648
rect 4577 7588 4581 7644
rect 4581 7588 4637 7644
rect 4637 7588 4641 7644
rect 4577 7584 4641 7588
rect 4657 7644 4721 7648
rect 4657 7588 4661 7644
rect 4661 7588 4717 7644
rect 4717 7588 4721 7644
rect 4657 7584 4721 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 18278 7644 18342 7648
rect 18278 7588 18282 7644
rect 18282 7588 18338 7644
rect 18338 7588 18342 7644
rect 18278 7584 18342 7588
rect 18358 7644 18422 7648
rect 18358 7588 18362 7644
rect 18362 7588 18418 7644
rect 18418 7588 18422 7644
rect 18358 7584 18422 7588
rect 18438 7644 18502 7648
rect 18438 7588 18442 7644
rect 18442 7588 18498 7644
rect 18498 7588 18502 7644
rect 18438 7584 18502 7588
rect 18518 7644 18582 7648
rect 18518 7588 18522 7644
rect 18522 7588 18578 7644
rect 18578 7588 18582 7644
rect 18518 7584 18582 7588
rect 12204 7516 12268 7580
rect 7882 7100 7946 7104
rect 7882 7044 7886 7100
rect 7886 7044 7942 7100
rect 7942 7044 7946 7100
rect 7882 7040 7946 7044
rect 7962 7100 8026 7104
rect 7962 7044 7966 7100
rect 7966 7044 8022 7100
rect 8022 7044 8026 7100
rect 7962 7040 8026 7044
rect 8042 7100 8106 7104
rect 8042 7044 8046 7100
rect 8046 7044 8102 7100
rect 8102 7044 8106 7100
rect 8042 7040 8106 7044
rect 8122 7100 8186 7104
rect 8122 7044 8126 7100
rect 8126 7044 8182 7100
rect 8182 7044 8186 7100
rect 8122 7040 8186 7044
rect 14813 7100 14877 7104
rect 14813 7044 14817 7100
rect 14817 7044 14873 7100
rect 14873 7044 14877 7100
rect 14813 7040 14877 7044
rect 14893 7100 14957 7104
rect 14893 7044 14897 7100
rect 14897 7044 14953 7100
rect 14953 7044 14957 7100
rect 14893 7040 14957 7044
rect 14973 7100 15037 7104
rect 14973 7044 14977 7100
rect 14977 7044 15033 7100
rect 15033 7044 15037 7100
rect 14973 7040 15037 7044
rect 15053 7100 15117 7104
rect 15053 7044 15057 7100
rect 15057 7044 15113 7100
rect 15113 7044 15117 7100
rect 15053 7040 15117 7044
rect 4417 6556 4481 6560
rect 4417 6500 4421 6556
rect 4421 6500 4477 6556
rect 4477 6500 4481 6556
rect 4417 6496 4481 6500
rect 4497 6556 4561 6560
rect 4497 6500 4501 6556
rect 4501 6500 4557 6556
rect 4557 6500 4561 6556
rect 4497 6496 4561 6500
rect 4577 6556 4641 6560
rect 4577 6500 4581 6556
rect 4581 6500 4637 6556
rect 4637 6500 4641 6556
rect 4577 6496 4641 6500
rect 4657 6556 4721 6560
rect 4657 6500 4661 6556
rect 4661 6500 4717 6556
rect 4717 6500 4721 6556
rect 4657 6496 4721 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 18278 6556 18342 6560
rect 18278 6500 18282 6556
rect 18282 6500 18338 6556
rect 18338 6500 18342 6556
rect 18278 6496 18342 6500
rect 18358 6556 18422 6560
rect 18358 6500 18362 6556
rect 18362 6500 18418 6556
rect 18418 6500 18422 6556
rect 18358 6496 18422 6500
rect 18438 6556 18502 6560
rect 18438 6500 18442 6556
rect 18442 6500 18498 6556
rect 18498 6500 18502 6556
rect 18438 6496 18502 6500
rect 18518 6556 18582 6560
rect 18518 6500 18522 6556
rect 18522 6500 18578 6556
rect 18578 6500 18582 6556
rect 18518 6496 18582 6500
rect 7882 6012 7946 6016
rect 7882 5956 7886 6012
rect 7886 5956 7942 6012
rect 7942 5956 7946 6012
rect 7882 5952 7946 5956
rect 7962 6012 8026 6016
rect 7962 5956 7966 6012
rect 7966 5956 8022 6012
rect 8022 5956 8026 6012
rect 7962 5952 8026 5956
rect 8042 6012 8106 6016
rect 8042 5956 8046 6012
rect 8046 5956 8102 6012
rect 8102 5956 8106 6012
rect 8042 5952 8106 5956
rect 8122 6012 8186 6016
rect 8122 5956 8126 6012
rect 8126 5956 8182 6012
rect 8182 5956 8186 6012
rect 8122 5952 8186 5956
rect 14813 6012 14877 6016
rect 14813 5956 14817 6012
rect 14817 5956 14873 6012
rect 14873 5956 14877 6012
rect 14813 5952 14877 5956
rect 14893 6012 14957 6016
rect 14893 5956 14897 6012
rect 14897 5956 14953 6012
rect 14953 5956 14957 6012
rect 14893 5952 14957 5956
rect 14973 6012 15037 6016
rect 14973 5956 14977 6012
rect 14977 5956 15033 6012
rect 15033 5956 15037 6012
rect 14973 5952 15037 5956
rect 15053 6012 15117 6016
rect 15053 5956 15057 6012
rect 15057 5956 15113 6012
rect 15113 5956 15117 6012
rect 15053 5952 15117 5956
rect 4417 5468 4481 5472
rect 4417 5412 4421 5468
rect 4421 5412 4477 5468
rect 4477 5412 4481 5468
rect 4417 5408 4481 5412
rect 4497 5468 4561 5472
rect 4497 5412 4501 5468
rect 4501 5412 4557 5468
rect 4557 5412 4561 5468
rect 4497 5408 4561 5412
rect 4577 5468 4641 5472
rect 4577 5412 4581 5468
rect 4581 5412 4637 5468
rect 4637 5412 4641 5468
rect 4577 5408 4641 5412
rect 4657 5468 4721 5472
rect 4657 5412 4661 5468
rect 4661 5412 4717 5468
rect 4717 5412 4721 5468
rect 4657 5408 4721 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 18278 5468 18342 5472
rect 18278 5412 18282 5468
rect 18282 5412 18338 5468
rect 18338 5412 18342 5468
rect 18278 5408 18342 5412
rect 18358 5468 18422 5472
rect 18358 5412 18362 5468
rect 18362 5412 18418 5468
rect 18418 5412 18422 5468
rect 18358 5408 18422 5412
rect 18438 5468 18502 5472
rect 18438 5412 18442 5468
rect 18442 5412 18498 5468
rect 18498 5412 18502 5468
rect 18438 5408 18502 5412
rect 18518 5468 18582 5472
rect 18518 5412 18522 5468
rect 18522 5412 18578 5468
rect 18578 5412 18582 5468
rect 18518 5408 18582 5412
rect 7882 4924 7946 4928
rect 7882 4868 7886 4924
rect 7886 4868 7942 4924
rect 7942 4868 7946 4924
rect 7882 4864 7946 4868
rect 7962 4924 8026 4928
rect 7962 4868 7966 4924
rect 7966 4868 8022 4924
rect 8022 4868 8026 4924
rect 7962 4864 8026 4868
rect 8042 4924 8106 4928
rect 8042 4868 8046 4924
rect 8046 4868 8102 4924
rect 8102 4868 8106 4924
rect 8042 4864 8106 4868
rect 8122 4924 8186 4928
rect 8122 4868 8126 4924
rect 8126 4868 8182 4924
rect 8182 4868 8186 4924
rect 8122 4864 8186 4868
rect 14813 4924 14877 4928
rect 14813 4868 14817 4924
rect 14817 4868 14873 4924
rect 14873 4868 14877 4924
rect 14813 4864 14877 4868
rect 14893 4924 14957 4928
rect 14893 4868 14897 4924
rect 14897 4868 14953 4924
rect 14953 4868 14957 4924
rect 14893 4864 14957 4868
rect 14973 4924 15037 4928
rect 14973 4868 14977 4924
rect 14977 4868 15033 4924
rect 15033 4868 15037 4924
rect 14973 4864 15037 4868
rect 15053 4924 15117 4928
rect 15053 4868 15057 4924
rect 15057 4868 15113 4924
rect 15113 4868 15117 4924
rect 15053 4864 15117 4868
rect 19196 4720 19260 4724
rect 19196 4664 19210 4720
rect 19210 4664 19260 4720
rect 19196 4660 19260 4664
rect 12204 4524 12268 4588
rect 4417 4380 4481 4384
rect 4417 4324 4421 4380
rect 4421 4324 4477 4380
rect 4477 4324 4481 4380
rect 4417 4320 4481 4324
rect 4497 4380 4561 4384
rect 4497 4324 4501 4380
rect 4501 4324 4557 4380
rect 4557 4324 4561 4380
rect 4497 4320 4561 4324
rect 4577 4380 4641 4384
rect 4577 4324 4581 4380
rect 4581 4324 4637 4380
rect 4637 4324 4641 4380
rect 4577 4320 4641 4324
rect 4657 4380 4721 4384
rect 4657 4324 4661 4380
rect 4661 4324 4717 4380
rect 4717 4324 4721 4380
rect 4657 4320 4721 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 18278 4380 18342 4384
rect 18278 4324 18282 4380
rect 18282 4324 18338 4380
rect 18338 4324 18342 4380
rect 18278 4320 18342 4324
rect 18358 4380 18422 4384
rect 18358 4324 18362 4380
rect 18362 4324 18418 4380
rect 18418 4324 18422 4380
rect 18358 4320 18422 4324
rect 18438 4380 18502 4384
rect 18438 4324 18442 4380
rect 18442 4324 18498 4380
rect 18498 4324 18502 4380
rect 18438 4320 18502 4324
rect 18518 4380 18582 4384
rect 18518 4324 18522 4380
rect 18522 4324 18578 4380
rect 18578 4324 18582 4380
rect 18518 4320 18582 4324
rect 9444 4116 9508 4180
rect 9628 4116 9692 4180
rect 7882 3836 7946 3840
rect 7882 3780 7886 3836
rect 7886 3780 7942 3836
rect 7942 3780 7946 3836
rect 7882 3776 7946 3780
rect 7962 3836 8026 3840
rect 7962 3780 7966 3836
rect 7966 3780 8022 3836
rect 8022 3780 8026 3836
rect 7962 3776 8026 3780
rect 8042 3836 8106 3840
rect 8042 3780 8046 3836
rect 8046 3780 8102 3836
rect 8102 3780 8106 3836
rect 8042 3776 8106 3780
rect 8122 3836 8186 3840
rect 8122 3780 8126 3836
rect 8126 3780 8182 3836
rect 8182 3780 8186 3836
rect 8122 3776 8186 3780
rect 14813 3836 14877 3840
rect 14813 3780 14817 3836
rect 14817 3780 14873 3836
rect 14873 3780 14877 3836
rect 14813 3776 14877 3780
rect 14893 3836 14957 3840
rect 14893 3780 14897 3836
rect 14897 3780 14953 3836
rect 14953 3780 14957 3836
rect 14893 3776 14957 3780
rect 14973 3836 15037 3840
rect 14973 3780 14977 3836
rect 14977 3780 15033 3836
rect 15033 3780 15037 3836
rect 14973 3776 15037 3780
rect 15053 3836 15117 3840
rect 15053 3780 15057 3836
rect 15057 3780 15113 3836
rect 15113 3780 15117 3836
rect 15053 3776 15117 3780
rect 4417 3292 4481 3296
rect 4417 3236 4421 3292
rect 4421 3236 4477 3292
rect 4477 3236 4481 3292
rect 4417 3232 4481 3236
rect 4497 3292 4561 3296
rect 4497 3236 4501 3292
rect 4501 3236 4557 3292
rect 4557 3236 4561 3292
rect 4497 3232 4561 3236
rect 4577 3292 4641 3296
rect 4577 3236 4581 3292
rect 4581 3236 4637 3292
rect 4637 3236 4641 3292
rect 4577 3232 4641 3236
rect 4657 3292 4721 3296
rect 4657 3236 4661 3292
rect 4661 3236 4717 3292
rect 4717 3236 4721 3292
rect 4657 3232 4721 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 18278 3292 18342 3296
rect 18278 3236 18282 3292
rect 18282 3236 18338 3292
rect 18338 3236 18342 3292
rect 18278 3232 18342 3236
rect 18358 3292 18422 3296
rect 18358 3236 18362 3292
rect 18362 3236 18418 3292
rect 18418 3236 18422 3292
rect 18358 3232 18422 3236
rect 18438 3292 18502 3296
rect 18438 3236 18442 3292
rect 18442 3236 18498 3292
rect 18498 3236 18502 3292
rect 18438 3232 18502 3236
rect 18518 3292 18582 3296
rect 18518 3236 18522 3292
rect 18522 3236 18578 3292
rect 18578 3236 18582 3292
rect 18518 3232 18582 3236
rect 10916 3164 10980 3228
rect 7882 2748 7946 2752
rect 7882 2692 7886 2748
rect 7886 2692 7942 2748
rect 7942 2692 7946 2748
rect 7882 2688 7946 2692
rect 7962 2748 8026 2752
rect 7962 2692 7966 2748
rect 7966 2692 8022 2748
rect 8022 2692 8026 2748
rect 7962 2688 8026 2692
rect 8042 2748 8106 2752
rect 8042 2692 8046 2748
rect 8046 2692 8102 2748
rect 8102 2692 8106 2748
rect 8042 2688 8106 2692
rect 8122 2748 8186 2752
rect 8122 2692 8126 2748
rect 8126 2692 8182 2748
rect 8182 2692 8186 2748
rect 8122 2688 8186 2692
rect 9444 2680 9508 2684
rect 9444 2624 9494 2680
rect 9494 2624 9508 2680
rect 9444 2620 9508 2624
rect 9812 2620 9876 2684
rect 10916 2756 10980 2820
rect 14813 2748 14877 2752
rect 14813 2692 14817 2748
rect 14817 2692 14873 2748
rect 14873 2692 14877 2748
rect 14813 2688 14877 2692
rect 14893 2748 14957 2752
rect 14893 2692 14897 2748
rect 14897 2692 14953 2748
rect 14953 2692 14957 2748
rect 14893 2688 14957 2692
rect 14973 2748 15037 2752
rect 14973 2692 14977 2748
rect 14977 2692 15033 2748
rect 15033 2692 15037 2748
rect 14973 2688 15037 2692
rect 15053 2748 15117 2752
rect 15053 2692 15057 2748
rect 15057 2692 15113 2748
rect 15113 2692 15117 2748
rect 15053 2688 15117 2692
rect 19196 2756 19260 2820
rect 4417 2204 4481 2208
rect 4417 2148 4421 2204
rect 4421 2148 4477 2204
rect 4477 2148 4481 2204
rect 4417 2144 4481 2148
rect 4497 2204 4561 2208
rect 4497 2148 4501 2204
rect 4501 2148 4557 2204
rect 4557 2148 4561 2204
rect 4497 2144 4561 2148
rect 4577 2204 4641 2208
rect 4577 2148 4581 2204
rect 4581 2148 4637 2204
rect 4637 2148 4641 2204
rect 4577 2144 4641 2148
rect 4657 2204 4721 2208
rect 4657 2148 4661 2204
rect 4661 2148 4717 2204
rect 4717 2148 4721 2204
rect 4657 2144 4721 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 18278 2204 18342 2208
rect 18278 2148 18282 2204
rect 18282 2148 18338 2204
rect 18338 2148 18342 2204
rect 18278 2144 18342 2148
rect 18358 2204 18422 2208
rect 18358 2148 18362 2204
rect 18362 2148 18418 2204
rect 18418 2148 18422 2204
rect 18358 2144 18422 2148
rect 18438 2204 18502 2208
rect 18438 2148 18442 2204
rect 18442 2148 18498 2204
rect 18498 2148 18502 2204
rect 18438 2144 18502 2148
rect 18518 2204 18582 2208
rect 18518 2148 18522 2204
rect 18522 2148 18578 2204
rect 18578 2148 18582 2204
rect 18518 2144 18582 2148
<< metal4 >>
rect 4409 20704 4729 20720
rect 4409 20640 4417 20704
rect 4481 20640 4497 20704
rect 4561 20640 4577 20704
rect 4641 20640 4657 20704
rect 4721 20640 4729 20704
rect 4409 19616 4729 20640
rect 4409 19552 4417 19616
rect 4481 19552 4497 19616
rect 4561 19552 4577 19616
rect 4641 19552 4657 19616
rect 4721 19552 4729 19616
rect 4409 18528 4729 19552
rect 4409 18464 4417 18528
rect 4481 18464 4497 18528
rect 4561 18464 4577 18528
rect 4641 18464 4657 18528
rect 4721 18464 4729 18528
rect 4409 17440 4729 18464
rect 4409 17376 4417 17440
rect 4481 17376 4497 17440
rect 4561 17376 4577 17440
rect 4641 17376 4657 17440
rect 4721 17376 4729 17440
rect 4409 16352 4729 17376
rect 7874 20160 8195 20720
rect 7874 20096 7882 20160
rect 7946 20096 7962 20160
rect 8026 20096 8042 20160
rect 8106 20096 8122 20160
rect 8186 20096 8195 20160
rect 7874 19072 8195 20096
rect 7874 19008 7882 19072
rect 7946 19008 7962 19072
rect 8026 19008 8042 19072
rect 8106 19008 8122 19072
rect 8186 19008 8195 19072
rect 7874 17984 8195 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9627 18052 9693 18053
rect 9627 17988 9628 18052
rect 9692 17988 9693 18052
rect 9627 17987 9693 17988
rect 7874 17920 7882 17984
rect 7946 17920 7962 17984
rect 8026 17920 8042 17984
rect 8106 17920 8122 17984
rect 8186 17920 8195 17984
rect 7874 16896 8195 17920
rect 7874 16832 7882 16896
rect 7946 16832 7962 16896
rect 8026 16832 8042 16896
rect 8106 16832 8122 16896
rect 8186 16832 8195 16896
rect 7603 16828 7669 16829
rect 7603 16764 7604 16828
rect 7668 16764 7669 16828
rect 7603 16763 7669 16764
rect 4409 16288 4417 16352
rect 4481 16288 4497 16352
rect 4561 16288 4577 16352
rect 4641 16288 4657 16352
rect 4721 16288 4729 16352
rect 4409 15264 4729 16288
rect 4409 15200 4417 15264
rect 4481 15200 4497 15264
rect 4561 15200 4577 15264
rect 4641 15200 4657 15264
rect 4721 15200 4729 15264
rect 4409 14176 4729 15200
rect 4409 14112 4417 14176
rect 4481 14112 4497 14176
rect 4561 14112 4577 14176
rect 4641 14112 4657 14176
rect 4721 14112 4729 14176
rect 4409 13088 4729 14112
rect 4409 13024 4417 13088
rect 4481 13024 4497 13088
rect 4561 13024 4577 13088
rect 4641 13024 4657 13088
rect 4721 13024 4729 13088
rect 4409 12000 4729 13024
rect 4409 11936 4417 12000
rect 4481 11936 4497 12000
rect 4561 11936 4577 12000
rect 4641 11936 4657 12000
rect 4721 11936 4729 12000
rect 4409 10912 4729 11936
rect 4409 10848 4417 10912
rect 4481 10848 4497 10912
rect 4561 10848 4577 10912
rect 4641 10848 4657 10912
rect 4721 10848 4729 10912
rect 4409 9824 4729 10848
rect 7606 10301 7666 16763
rect 7874 15808 8195 16832
rect 7874 15744 7882 15808
rect 7946 15744 7962 15808
rect 8026 15744 8042 15808
rect 8106 15744 8122 15808
rect 8186 15744 8195 15808
rect 7874 14720 8195 15744
rect 7874 14656 7882 14720
rect 7946 14656 7962 14720
rect 8026 14656 8042 14720
rect 8106 14656 8122 14720
rect 8186 14656 8195 14720
rect 7874 13632 8195 14656
rect 9630 14109 9690 17987
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 9811 15468 9877 15469
rect 9811 15404 9812 15468
rect 9876 15404 9877 15468
rect 9811 15403 9877 15404
rect 9627 14108 9693 14109
rect 9627 14044 9628 14108
rect 9692 14044 9693 14108
rect 9627 14043 9693 14044
rect 9814 13837 9874 15403
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 9995 15060 10061 15061
rect 9995 14996 9996 15060
rect 10060 14996 10061 15060
rect 9995 14995 10061 14996
rect 9811 13836 9877 13837
rect 9811 13772 9812 13836
rect 9876 13772 9877 13836
rect 9811 13771 9877 13772
rect 7874 13568 7882 13632
rect 7946 13568 7962 13632
rect 8026 13568 8042 13632
rect 8106 13568 8122 13632
rect 8186 13568 8195 13632
rect 7874 12544 8195 13568
rect 9998 13021 10058 14995
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 9995 13020 10061 13021
rect 9995 12956 9996 13020
rect 10060 12956 10061 13020
rect 9995 12955 10061 12956
rect 7874 12480 7882 12544
rect 7946 12480 7962 12544
rect 8026 12480 8042 12544
rect 8106 12480 8122 12544
rect 8186 12480 8195 12544
rect 7874 11456 8195 12480
rect 7874 11392 7882 11456
rect 7946 11392 7962 11456
rect 8026 11392 8042 11456
rect 8106 11392 8122 11456
rect 8186 11392 8195 11456
rect 7874 10368 8195 11392
rect 7874 10304 7882 10368
rect 7946 10304 7962 10368
rect 8026 10304 8042 10368
rect 8106 10304 8122 10368
rect 8186 10304 8195 10368
rect 7603 10300 7669 10301
rect 7603 10236 7604 10300
rect 7668 10236 7669 10300
rect 7603 10235 7669 10236
rect 4409 9760 4417 9824
rect 4481 9760 4497 9824
rect 4561 9760 4577 9824
rect 4641 9760 4657 9824
rect 4721 9760 4729 9824
rect 4409 8736 4729 9760
rect 4409 8672 4417 8736
rect 4481 8672 4497 8736
rect 4561 8672 4577 8736
rect 4641 8672 4657 8736
rect 4721 8672 4729 8736
rect 4409 7648 4729 8672
rect 4409 7584 4417 7648
rect 4481 7584 4497 7648
rect 4561 7584 4577 7648
rect 4641 7584 4657 7648
rect 4721 7584 4729 7648
rect 4409 6560 4729 7584
rect 4409 6496 4417 6560
rect 4481 6496 4497 6560
rect 4561 6496 4577 6560
rect 4641 6496 4657 6560
rect 4721 6496 4729 6560
rect 4409 5472 4729 6496
rect 4409 5408 4417 5472
rect 4481 5408 4497 5472
rect 4561 5408 4577 5472
rect 4641 5408 4657 5472
rect 4721 5408 4729 5472
rect 4409 4384 4729 5408
rect 4409 4320 4417 4384
rect 4481 4320 4497 4384
rect 4561 4320 4577 4384
rect 4641 4320 4657 4384
rect 4721 4320 4729 4384
rect 4409 3296 4729 4320
rect 4409 3232 4417 3296
rect 4481 3232 4497 3296
rect 4561 3232 4577 3296
rect 4641 3232 4657 3296
rect 4721 3232 4729 3296
rect 4409 2208 4729 3232
rect 4409 2144 4417 2208
rect 4481 2144 4497 2208
rect 4561 2144 4577 2208
rect 4641 2144 4657 2208
rect 4721 2144 4729 2208
rect 4409 2128 4729 2144
rect 7874 9280 8195 10304
rect 7874 9216 7882 9280
rect 7946 9216 7962 9280
rect 8026 9216 8042 9280
rect 8106 9216 8122 9280
rect 8186 9216 8195 9280
rect 7874 8192 8195 9216
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 9627 9076 9693 9077
rect 9627 9012 9628 9076
rect 9692 9012 9693 9076
rect 9627 9011 9693 9012
rect 7874 8128 7882 8192
rect 7946 8128 7962 8192
rect 8026 8128 8042 8192
rect 8106 8128 8122 8192
rect 8186 8128 8195 8192
rect 7874 7104 8195 8128
rect 7874 7040 7882 7104
rect 7946 7040 7962 7104
rect 8026 7040 8042 7104
rect 8106 7040 8122 7104
rect 8186 7040 8195 7104
rect 7874 6016 8195 7040
rect 7874 5952 7882 6016
rect 7946 5952 7962 6016
rect 8026 5952 8042 6016
rect 8106 5952 8122 6016
rect 8186 5952 8195 6016
rect 7874 4928 8195 5952
rect 7874 4864 7882 4928
rect 7946 4864 7962 4928
rect 8026 4864 8042 4928
rect 8106 4864 8122 4928
rect 8186 4864 8195 4928
rect 7874 3840 8195 4864
rect 9630 4181 9690 9011
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 9811 7988 9877 7989
rect 9811 7924 9812 7988
rect 9876 7924 9877 7988
rect 9811 7923 9877 7924
rect 9443 4180 9509 4181
rect 9443 4116 9444 4180
rect 9508 4116 9509 4180
rect 9443 4115 9509 4116
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 7874 3776 7882 3840
rect 7946 3776 7962 3840
rect 8026 3776 8042 3840
rect 8106 3776 8122 3840
rect 8186 3776 8195 3840
rect 7874 2752 8195 3776
rect 7874 2688 7882 2752
rect 7946 2688 7962 2752
rect 8026 2688 8042 2752
rect 8106 2688 8122 2752
rect 8186 2688 8195 2752
rect 7874 2128 8195 2688
rect 9446 2685 9506 4115
rect 9814 2685 9874 7923
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 14805 20160 15125 20720
rect 14805 20096 14813 20160
rect 14877 20096 14893 20160
rect 14957 20096 14973 20160
rect 15037 20096 15053 20160
rect 15117 20096 15125 20160
rect 14805 19072 15125 20096
rect 14805 19008 14813 19072
rect 14877 19008 14893 19072
rect 14957 19008 14973 19072
rect 15037 19008 15053 19072
rect 15117 19008 15125 19072
rect 14805 17984 15125 19008
rect 14805 17920 14813 17984
rect 14877 17920 14893 17984
rect 14957 17920 14973 17984
rect 15037 17920 15053 17984
rect 15117 17920 15125 17984
rect 14805 16896 15125 17920
rect 14805 16832 14813 16896
rect 14877 16832 14893 16896
rect 14957 16832 14973 16896
rect 15037 16832 15053 16896
rect 15117 16832 15125 16896
rect 14805 15808 15125 16832
rect 14805 15744 14813 15808
rect 14877 15744 14893 15808
rect 14957 15744 14973 15808
rect 15037 15744 15053 15808
rect 15117 15744 15125 15808
rect 14805 14720 15125 15744
rect 14805 14656 14813 14720
rect 14877 14656 14893 14720
rect 14957 14656 14973 14720
rect 15037 14656 15053 14720
rect 15117 14656 15125 14720
rect 14805 13632 15125 14656
rect 14805 13568 14813 13632
rect 14877 13568 14893 13632
rect 14957 13568 14973 13632
rect 15037 13568 15053 13632
rect 15117 13568 15125 13632
rect 14805 12544 15125 13568
rect 14805 12480 14813 12544
rect 14877 12480 14893 12544
rect 14957 12480 14973 12544
rect 15037 12480 15053 12544
rect 15117 12480 15125 12544
rect 14805 11456 15125 12480
rect 14805 11392 14813 11456
rect 14877 11392 14893 11456
rect 14957 11392 14973 11456
rect 15037 11392 15053 11456
rect 15117 11392 15125 11456
rect 14805 10368 15125 11392
rect 14805 10304 14813 10368
rect 14877 10304 14893 10368
rect 14957 10304 14973 10368
rect 15037 10304 15053 10368
rect 15117 10304 15125 10368
rect 14805 9280 15125 10304
rect 14805 9216 14813 9280
rect 14877 9216 14893 9280
rect 14957 9216 14973 9280
rect 15037 9216 15053 9280
rect 15117 9216 15125 9280
rect 14805 8192 15125 9216
rect 14805 8128 14813 8192
rect 14877 8128 14893 8192
rect 14957 8128 14973 8192
rect 15037 8128 15053 8192
rect 15117 8128 15125 8192
rect 12203 7580 12269 7581
rect 12203 7516 12204 7580
rect 12268 7516 12269 7580
rect 12203 7515 12269 7516
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 12206 4589 12266 7515
rect 14805 7104 15125 8128
rect 14805 7040 14813 7104
rect 14877 7040 14893 7104
rect 14957 7040 14973 7104
rect 15037 7040 15053 7104
rect 15117 7040 15125 7104
rect 14805 6016 15125 7040
rect 14805 5952 14813 6016
rect 14877 5952 14893 6016
rect 14957 5952 14973 6016
rect 15037 5952 15053 6016
rect 15117 5952 15125 6016
rect 14805 4928 15125 5952
rect 14805 4864 14813 4928
rect 14877 4864 14893 4928
rect 14957 4864 14973 4928
rect 15037 4864 15053 4928
rect 15117 4864 15125 4928
rect 12203 4588 12269 4589
rect 12203 4524 12204 4588
rect 12268 4524 12269 4588
rect 12203 4523 12269 4524
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10915 3228 10981 3229
rect 10915 3164 10916 3228
rect 10980 3164 10981 3228
rect 10915 3163 10981 3164
rect 10918 2821 10978 3163
rect 10915 2820 10981 2821
rect 10915 2756 10916 2820
rect 10980 2756 10981 2820
rect 10915 2755 10981 2756
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 9811 2684 9877 2685
rect 9811 2620 9812 2684
rect 9876 2620 9877 2684
rect 9811 2619 9877 2620
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 14805 3840 15125 4864
rect 14805 3776 14813 3840
rect 14877 3776 14893 3840
rect 14957 3776 14973 3840
rect 15037 3776 15053 3840
rect 15117 3776 15125 3840
rect 14805 2752 15125 3776
rect 14805 2688 14813 2752
rect 14877 2688 14893 2752
rect 14957 2688 14973 2752
rect 15037 2688 15053 2752
rect 15117 2688 15125 2752
rect 14805 2128 15125 2688
rect 18270 20704 18591 20720
rect 18270 20640 18278 20704
rect 18342 20640 18358 20704
rect 18422 20640 18438 20704
rect 18502 20640 18518 20704
rect 18582 20640 18591 20704
rect 18270 19616 18591 20640
rect 18270 19552 18278 19616
rect 18342 19552 18358 19616
rect 18422 19552 18438 19616
rect 18502 19552 18518 19616
rect 18582 19552 18591 19616
rect 18270 18528 18591 19552
rect 18270 18464 18278 18528
rect 18342 18464 18358 18528
rect 18422 18464 18438 18528
rect 18502 18464 18518 18528
rect 18582 18464 18591 18528
rect 18270 17440 18591 18464
rect 18270 17376 18278 17440
rect 18342 17376 18358 17440
rect 18422 17376 18438 17440
rect 18502 17376 18518 17440
rect 18582 17376 18591 17440
rect 18270 16352 18591 17376
rect 18270 16288 18278 16352
rect 18342 16288 18358 16352
rect 18422 16288 18438 16352
rect 18502 16288 18518 16352
rect 18582 16288 18591 16352
rect 18270 15264 18591 16288
rect 18270 15200 18278 15264
rect 18342 15200 18358 15264
rect 18422 15200 18438 15264
rect 18502 15200 18518 15264
rect 18582 15200 18591 15264
rect 18270 14176 18591 15200
rect 18270 14112 18278 14176
rect 18342 14112 18358 14176
rect 18422 14112 18438 14176
rect 18502 14112 18518 14176
rect 18582 14112 18591 14176
rect 18270 13088 18591 14112
rect 18270 13024 18278 13088
rect 18342 13024 18358 13088
rect 18422 13024 18438 13088
rect 18502 13024 18518 13088
rect 18582 13024 18591 13088
rect 18270 12000 18591 13024
rect 18270 11936 18278 12000
rect 18342 11936 18358 12000
rect 18422 11936 18438 12000
rect 18502 11936 18518 12000
rect 18582 11936 18591 12000
rect 18270 10912 18591 11936
rect 18270 10848 18278 10912
rect 18342 10848 18358 10912
rect 18422 10848 18438 10912
rect 18502 10848 18518 10912
rect 18582 10848 18591 10912
rect 18270 9824 18591 10848
rect 18270 9760 18278 9824
rect 18342 9760 18358 9824
rect 18422 9760 18438 9824
rect 18502 9760 18518 9824
rect 18582 9760 18591 9824
rect 18270 8736 18591 9760
rect 18270 8672 18278 8736
rect 18342 8672 18358 8736
rect 18422 8672 18438 8736
rect 18502 8672 18518 8736
rect 18582 8672 18591 8736
rect 18270 7648 18591 8672
rect 18270 7584 18278 7648
rect 18342 7584 18358 7648
rect 18422 7584 18438 7648
rect 18502 7584 18518 7648
rect 18582 7584 18591 7648
rect 18270 6560 18591 7584
rect 18270 6496 18278 6560
rect 18342 6496 18358 6560
rect 18422 6496 18438 6560
rect 18502 6496 18518 6560
rect 18582 6496 18591 6560
rect 18270 5472 18591 6496
rect 18270 5408 18278 5472
rect 18342 5408 18358 5472
rect 18422 5408 18438 5472
rect 18502 5408 18518 5472
rect 18582 5408 18591 5472
rect 18270 4384 18591 5408
rect 19195 4724 19261 4725
rect 19195 4660 19196 4724
rect 19260 4660 19261 4724
rect 19195 4659 19261 4660
rect 18270 4320 18278 4384
rect 18342 4320 18358 4384
rect 18422 4320 18438 4384
rect 18502 4320 18518 4384
rect 18582 4320 18591 4384
rect 18270 3296 18591 4320
rect 18270 3232 18278 3296
rect 18342 3232 18358 3296
rect 18422 3232 18438 3296
rect 18502 3232 18518 3296
rect 18582 3232 18591 3296
rect 18270 2208 18591 3232
rect 19198 2821 19258 4659
rect 19195 2820 19261 2821
rect 19195 2756 19196 2820
rect 19260 2756 19261 2820
rect 19195 2755 19261 2756
rect 18270 2144 18278 2208
rect 18342 2144 18358 2208
rect 18422 2144 18438 2208
rect 18502 2144 18518 2208
rect 18582 2144 18591 2208
rect 18270 2128 18591 2144
use sky130_fd_sc_hd__buf_1  input23 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1380 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1624635492
transform 1 0 1380 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1624635492
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1656 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp 1624635492
transform 1 0 1656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1624635492
transform 1 0 1840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1624635492
transform 1 0 2116 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13
timestamp 1624635492
transform 1 0 2300 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1624635492
transform 1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_15
timestamp 1624635492
transform 1 0 2484 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp 1624635492
transform 1 0 2760 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1624635492
transform -1 0 2852 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1624635492
transform 1 0 2484 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1624635492
transform 1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3404 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1624635492
transform -1 0 3588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1624635492
transform -1 0 3220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1624635492
transform 1 0 3036 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_27
timestamp 1624635492
transform 1 0 3588 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30
timestamp 1624635492
transform 1 0 3864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1624635492
transform -1 0 4048 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_68 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_32
timestamp 1624635492
transform 1 0 4048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1624635492
transform 1 0 4048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_37
timestamp 1624635492
transform 1 0 4508 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36
timestamp 1624635492
transform 1 0 4416 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input40 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 4968 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1624635492
transform 1 0 4600 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_46
timestamp 1624635492
transform 1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_42
timestamp 1624635492
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42
timestamp 1624635492
transform 1 0 4968 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1624635492
transform -1 0 5336 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1624635492
transform 1 0 5244 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_50
timestamp 1624635492
transform 1 0 5704 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49
timestamp 1624635492
transform 1 0 5612 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1624635492
transform -1 0 5704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1624635492
transform -1 0 6164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_55
timestamp 1624635492
transform 1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55
timestamp 1624635492
transform 1 0 6164 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1624635492
transform -1 0 6164 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_61
timestamp 1624635492
transform 1 0 6716 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 6440 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59
timestamp 1624635492
transform 1 0 6532 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1624635492
transform -1 0 6716 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1624635492
transform 1 0 6716 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1624635492
transform 1 0 6348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_69
timestamp 1624635492
transform 1 0 6440 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_67
timestamp 1624635492
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1624635492
transform 1 0 7084 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1624635492
transform -1 0 7268 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1624635492
transform 1 0 7728 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1624635492
transform 1 0 7452 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1624635492
transform -1 0 7728 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1624635492
transform -1 0 7912 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_77
timestamp 1624635492
transform 1 0 8188 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74
timestamp 1624635492
transform 1 0 7912 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1624635492
transform 1 0 8096 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1624635492
transform -1 0 8188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_80
timestamp 1624635492
transform 1 0 8464 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1624635492
transform -1 0 8648 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_82
timestamp 1624635492
transform 1 0 8648 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8924 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_87
timestamp 1624635492
transform 1 0 9108 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 1624635492
transform 1 0 9200 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1624635492
transform 1 0 8924 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1624635492
transform 1 0 9108 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1624635492
transform -1 0 9108 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1624635492
transform 1 0 9568 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1624635492
transform 1 0 9384 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1624635492
transform -1 0 9568 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_97
timestamp 1624635492
transform 1 0 10028 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1624635492
transform 1 0 9752 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1624635492
transform 1 0 9936 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1624635492
transform -1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 1624635492
transform 1 0 10488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_100
timestamp 1624635492
transform 1 0 10304 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1624635492
transform 1 0 10488 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1624635492
transform -1 0 10488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1624635492
transform -1 0 10948 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_112
timestamp 1624635492
transform 1 0 11408 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_107
timestamp 1624635492
transform 1 0 10948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_112
timestamp 1624635492
transform 1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_106
timestamp 1624635492
transform 1 0 10856 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1624635492
transform -1 0 11408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1624635492
transform 1 0 11592 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1624635492
transform -1 0 11408 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_115
timestamp 1624635492
transform 1 0 11684 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1624635492
transform 1 0 12420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1624635492
transform 1 0 11868 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output93
timestamp 1624635492
transform -1 0 12420 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1624635492
transform 1 0 11776 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 11868 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13524 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1624635492
transform 1 0 14444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output98
timestamp 1624635492
transform 1 0 13892 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output99
timestamp 1624635492
transform 1 0 13340 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output103
timestamp 1624635492
transform 1 0 12788 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_131
timestamp 1624635492
transform 1 0 13156 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_137
timestamp 1624635492
transform 1 0 13708 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_143
timestamp 1624635492
transform 1 0 14260 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1624635492
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _040_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 14720 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 15180 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16560 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output95
timestamp 1624635492
transform 1 0 15180 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_146
timestamp 1624635492
transform 1 0 14536 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1624635492
transform 1 0 14996 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1624635492
transform 1 0 15548 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_151
timestamp 1624635492
transform 1 0 14996 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_172
timestamp 1624635492
transform 1 0 16928 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_169
timestamp 1624635492
transform 1 0 16652 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_177
timestamp 1624635492
transform 1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_172
timestamp 1624635492
transform 1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_168
timestamp 1624635492
transform 1 0 16560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1624635492
transform -1 0 17388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1624635492
transform -1 0 16928 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1624635492
transform 1 0 16836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1624635492
transform 1 0 17112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18400 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17112 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_1_190
timestamp 1624635492
transform 1 0 18584 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_194
timestamp 1624635492
transform 1 0 18952 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 1624635492
transform 1 0 18400 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output94
timestamp 1624635492
transform -1 0 18952 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1624635492
transform -1 0 19596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18768 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1624635492
transform 1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_201
timestamp 1624635492
transform 1 0 19596 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 1624635492
transform 1 0 19872 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1624635492
transform 1 0 19596 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output96
timestamp 1624635492
transform -1 0 20148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1624635492
transform 1 0 19780 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1624635492
transform 1 0 20056 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1624635492
transform 1 0 20332 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1624635492
transform -1 0 20884 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1624635492
transform -1 0 20884 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1624635492
transform 1 0 20884 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1624635492
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1624635492
transform -1 0 21436 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1624635492
transform -1 0 21436 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1624635492
transform 1 0 21436 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1624635492
transform 1 0 21436 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1624635492
transform -1 0 21896 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1624635492
transform -1 0 21896 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1624635492
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1624635492
transform -1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1624635492
transform -1 0 1932 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5
timestamp 1624635492
transform 1 0 1564 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 1932 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1624635492
transform 1 0 3772 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 3036 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_30
timestamp 1624635492
transform 1 0 3864 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_38
timestamp 1624635492
transform 1 0 4600 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1624635492
transform -1 0 5796 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1624635492
transform -1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1624635492
transform -1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1624635492
transform -1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 1624635492
transform 1 0 5060 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_47
timestamp 1624635492
transform 1 0 5428 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1624635492
transform 1 0 5796 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1624635492
transform 1 0 6348 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1624635492
transform 1 0 6716 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8372 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1624635492
transform -1 0 7452 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1624635492
transform -1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1624635492
transform -1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_65
timestamp 1624635492
transform 1 0 7084 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_69
timestamp 1624635492
transform 1 0 7452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_74
timestamp 1624635492
transform 1 0 7912 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_79
timestamp 1624635492
transform 1 0 8372 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_87
timestamp 1624635492
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_84
timestamp 1624635492
transform 1 0 8832 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1624635492
transform 1 0 9016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1624635492
transform -1 0 9568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1624635492
transform 1 0 9568 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1624635492
transform -1 0 10028 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_97
timestamp 1624635492
transform 1 0 10028 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_102
timestamp 1624635492
transform 1 0 10488 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1624635492
transform -1 0 10488 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1624635492
transform -1 0 10948 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1624635492
transform 1 0 12144 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11960 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output104
timestamp 1624635492
transform -1 0 12972 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_107
timestamp 1624635492
transform 1 0 10948 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_118
timestamp 1624635492
transform 1 0 11960 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_123
timestamp 1624635492
transform 1 0 12420 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1624635492
transform 1 0 14260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_129
timestamp 1624635492
transform 1 0 12972 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1624635492
transform 1 0 14076 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1624635492
transform 1 0 14352 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 14536 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16284 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_2_162
timestamp 1624635492
transform 1 0 16008 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17480 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_174
timestamp 1624635492
transform 1 0 17112 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1624635492
transform 1 0 19504 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output97
timestamp 1624635492
transform -1 0 20148 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1624635492
transform -1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1624635492
transform 1 0 18952 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_198
timestamp 1624635492
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_201
timestamp 1624635492
transform 1 0 19596 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_207
timestamp 1624635492
transform 1 0 20148 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1624635492
transform -1 0 21896 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1624635492
transform -1 0 21436 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1624635492
transform -1 0 20884 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 1624635492
transform 1 0 20884 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1624635492
transform 1 0 21436 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1624635492
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1624635492
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1624635492
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1624635492
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_39
timestamp 1624635492
transform 1 0 4692 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1624635492
transform 1 0 6348 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1624635492
transform -1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1624635492
transform -1 0 6624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1624635492
transform -1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1624635492
transform 1 0 5612 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 1624635492
transform 1 0 5428 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_51
timestamp 1624635492
transform 1 0 5796 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_55
timestamp 1624635492
transform 1 0 6164 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_60
timestamp 1624635492
transform 1 0 6624 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_64
timestamp 1624635492
transform 1 0 6992 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 7176 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1624635492
transform 1 0 7360 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1624635492
transform -1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1624635492
transform 1 0 7728 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1624635492
transform -1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_76
timestamp 1624635492
transform 1 0 8096 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_81
timestamp 1624635492
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1624635492
transform -1 0 8556 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9016 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1624635492
transform -1 0 10396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9936 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11408 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_86
timestamp 1624635492
transform 1 0 9016 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_91
timestamp 1624635492
transform 1 0 9476 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_96
timestamp 1624635492
transform 1 0 9936 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_101
timestamp 1624635492
transform 1 0 10396 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1624635492
transform 1 0 11868 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1624635492
transform 1 0 11592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_112
timestamp 1624635492
transform 1 0 11408 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_115
timestamp 1624635492
transform 1 0 11684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12880 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  mux_right_track_30.mux_l2_in_0_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 13984 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_126
timestamp 1624635492
transform 1 0 12696 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_137
timestamp 1624635492
transform 1 0 13708 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15732 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  output107
timestamp 1624635492
transform -1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_149
timestamp 1624635492
transform 1 0 14812 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_155
timestamp 1624635492
transform 1 0 15364 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18308 0 1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1624635492
transform 1 0 16836 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output110
timestamp 1624635492
transform -1 0 17480 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output111
timestamp 1624635492
transform -1 0 18032 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_168
timestamp 1624635492
transform 1 0 16560 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1624635492
transform 1 0 16928 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1624635492
transform 1 0 17480 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp 1624635492
transform 1 0 18032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20792 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1624635492
transform 1 0 19780 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1624635492
transform -1 0 21896 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1624635492
transform -1 0 21436 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp 1624635492
transform 1 0 20792 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1624635492
transform 1 0 21436 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1624635492
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1624635492
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1624635492
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1624635492
transform 1 0 3772 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_27
timestamp 1624635492
transform 1 0 3588 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_30
timestamp 1624635492
transform 1 0 3864 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1624635492
transform -1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1624635492
transform 1 0 6440 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6072 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_42
timestamp 1624635492
transform 1 0 4968 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_56
timestamp 1624635492
transform 1 0 6256 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1624635492
transform 1 0 6624 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_64
timestamp 1624635492
transform 1 0 6992 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1624635492
transform 1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1624635492
transform -1 0 7360 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1624635492
transform 1 0 7728 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_76
timestamp 1624635492
transform 1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1624635492
transform -1 0 8096 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1624635492
transform -1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_80
timestamp 1624635492
transform 1 0 8464 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1624635492
transform -1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9752 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1624635492
transform 1 0 9016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1624635492
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_84
timestamp 1624635492
transform 1 0 8832 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1624635492
transform 1 0 9108 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1624635492
transform 1 0 9568 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11408 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1624635492
transform 1 0 11224 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1624635492
transform 1 0 14260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output105
timestamp 1624635492
transform -1 0 13524 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output106
timestamp 1624635492
transform -1 0 14076 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1624635492
transform -1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_128
timestamp 1624635492
transform 1 0 12880 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_135
timestamp 1624635492
transform 1 0 13524 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_141
timestamp 1624635492
transform 1 0 14076 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_144
timestamp 1624635492
transform 1 0 14352 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 15916 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_2  output108
timestamp 1624635492
transform -1 0 15180 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output109
timestamp 1624635492
transform -1 0 15732 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_147
timestamp 1624635492
transform 1 0 14628 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_153
timestamp 1624635492
transform 1 0 15180 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_159
timestamp 1624635492
transform 1 0 15732 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output112
timestamp 1624635492
transform -1 0 17940 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_177
timestamp 1624635492
transform 1 0 17388 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_183
timestamp 1624635492
transform 1 0 17940 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_187
timestamp 1624635492
transform 1 0 18308 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 19780 0 -1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1624635492
transform 1 0 19504 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output101
timestamp 1624635492
transform 1 0 18952 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output102
timestamp 1624635492
transform 1 0 18400 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_192
timestamp 1624635492
transform 1 0 18768 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_198
timestamp 1624635492
transform 1 0 19320 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1624635492
transform 1 0 19596 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1624635492
transform -1 0 21896 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1624635492
transform 1 0 21252 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1624635492
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1624635492
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1624635492
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1624635492
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1624635492
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1624635492
transform 1 0 6348 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 1624635492
transform 1 0 5796 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_55
timestamp 1624635492
transform 1 0 6164 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_58
timestamp 1624635492
transform 1 0 6440 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_61
timestamp 1624635492
transform 1 0 6716 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_65
timestamp 1624635492
transform 1 0 7084 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6900 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_69
timestamp 1624635492
transform 1 0 7452 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7268 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1624635492
transform 1 0 7820 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7636 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1624635492
transform 1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1624635492
transform -1 0 8188 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_81
timestamp 1624635492
transform 1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1624635492
transform -1 0 8556 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 9016 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11408 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1624635492
transform 1 0 10120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1624635492
transform 1 0 9660 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1624635492
transform 1 0 9200 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_86
timestamp 1624635492
transform 1 0 9016 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 1624635492
transform 1 0 9476 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_96
timestamp 1624635492
transform 1 0 9936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_101
timestamp 1624635492
transform 1 0 10396 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1624635492
transform 1 0 11592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_112
timestamp 1624635492
transform 1 0 11408 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1624635492
transform 1 0 11684 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 13064 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_5_126
timestamp 1624635492
transform 1 0 12696 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1624635492
transform -1 0 16652 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14720 0 1 4896
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_5_146
timestamp 1624635492
transform 1 0 14536 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_164
timestamp 1624635492
transform 1 0 16192 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1624635492
transform 1 0 16836 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1624635492
transform -1 0 18308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_169
timestamp 1624635492
transform 1 0 16652 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1624635492
transform 1 0 16928 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_183
timestamp 1624635492
transform 1 0 17940 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_187
timestamp 1624635492
transform 1 0 18308 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1624635492
transform -1 0 18768 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1624635492
transform -1 0 19412 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1624635492
transform 1 0 19596 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_5_192
timestamp 1624635492
transform 1 0 18768 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_199
timestamp 1624635492
transform 1 0 19412 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1624635492
transform 1 0 20608 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1624635492
transform -1 0 21896 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1624635492
transform 1 0 20424 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1624635492
transform 1 0 21436 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1624635492
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1624635492
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1624635492
transform -1 0 1840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1624635492
transform -1 0 2208 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1624635492
transform 1 0 1380 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_8
timestamp 1624635492
transform 1 0 1840 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_12
timestamp 1624635492
transform 1 0 2208 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1624635492
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1624635492
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1624635492
transform 1 0 3772 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_24
timestamp 1624635492
transform 1 0 3312 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_28
timestamp 1624635492
transform 1 0 3680 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_30
timestamp 1624635492
transform 1 0 3864 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1624635492
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1624635492
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_51
timestamp 1624635492
transform 1 0 5796 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_50
timestamp 1624635492
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_42
timestamp 1624635492
transform 1 0 4968 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1624635492
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_61
timestamp 1624635492
transform 1 0 6716 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_58
timestamp 1624635492
transform 1 0 6440 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_55
timestamp 1624635492
transform 1 0 6164 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_57
timestamp 1624635492
transform 1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_53
timestamp 1624635492
transform 1 0 5980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 5980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1624635492
transform -1 0 6348 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1624635492
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 6532 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7636 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1624635492
transform 1 0 8556 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1624635492
transform -1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1624635492
transform 1 0 8004 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1624635492
transform 1 0 8372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1624635492
transform 1 0 7084 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_69
timestamp 1624635492
transform 1 0 7452 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_87
timestamp 1624635492
transform 1 0 9108 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1624635492
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_87
timestamp 1624635492
transform 1 0 9108 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_84
timestamp 1624635492
transform 1 0 8832 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1624635492
transform -1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1624635492
transform 1 0 9016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 9568 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 9292 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1624635492
transform 1 0 10120 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_101
timestamp 1624635492
transform 1 0 10396 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1624635492
transform 1 0 10304 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 12144 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1624635492
transform -1 0 12880 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1624635492
transform 1 0 11592 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1624635492
transform -1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11684 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1624635492
transform 1 0 12144 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1624635492
transform 1 0 12512 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_109
timestamp 1624635492
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_113
timestamp 1624635492
transform 1 0 11500 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_117
timestamp 1624635492
transform 1 0 11868 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1624635492
transform -1 0 12972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 14536 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13156 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1624635492
transform 1 0 14260 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_129
timestamp 1624635492
transform 1 0 12972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_140
timestamp 1624635492
transform 1 0 13984 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_144
timestamp 1624635492
transform 1 0 14352 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1624635492
transform 1 0 12880 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1624635492
transform 1 0 14996 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_146
timestamp 1624635492
transform 1 0 14536 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_149
timestamp 1624635492
transform 1 0 14812 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1624635492
transform -1 0 16008 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1624635492
transform -1 0 16008 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1624635492
transform -1 0 14812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1624635492
transform 1 0 14720 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_162
timestamp 1624635492
transform 1 0 16008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_162
timestamp 1624635492
transform 1 0 16008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1624635492
transform 1 0 16192 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1624635492
transform -1 0 16468 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 18768 0 -1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17296 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1624635492
transform 1 0 16836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1624635492
transform -1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_173
timestamp 1624635492
transform 1 0 17020 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_167
timestamp 1624635492
transform 1 0 16468 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_174
timestamp 1624635492
transform 1 0 17112 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1624635492
transform 1 0 18952 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 18952 0 1 5984
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20608 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1624635492
transform 1 0 19504 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_192
timestamp 1624635492
transform 1 0 18768 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 1624635492
transform 1 0 19228 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_201
timestamp 1624635492
transform 1 0 19596 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1624635492
transform 1 0 18768 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1624635492
transform 1 0 20608 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1624635492
transform -1 0 21896 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1624635492
transform -1 0 21896 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output100
timestamp 1624635492
transform -1 0 21344 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1624635492
transform 1 0 20608 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1624635492
transform 1 0 21344 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1624635492
transform 1 0 20424 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1624635492
transform 1 0 21436 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1624635492
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1624635492
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1624635492
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1624635492
transform 1 0 3772 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_27
timestamp 1624635492
transform 1 0 3588 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_30
timestamp 1624635492
transform 1 0 3864 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6532 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1624635492
transform 1 0 6164 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_42
timestamp 1624635492
transform 1 0 4968 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_54
timestamp 1624635492
transform 1 0 6072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1624635492
transform 1 0 6348 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1624635492
transform 1 0 6716 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1624635492
transform -1 0 8832 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1624635492
transform -1 0 8372 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1624635492
transform -1 0 7912 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1624635492
transform -1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1624635492
transform -1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1624635492
transform 1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_69
timestamp 1624635492
transform 1 0 7452 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_74
timestamp 1624635492
transform 1 0 7912 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_79
timestamp 1624635492
transform 1 0 8372 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 10488 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1624635492
transform -1 0 10120 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1624635492
transform 1 0 9016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_84
timestamp 1624635492
transform 1 0 8832 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1624635492
transform 1 0 9108 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_98
timestamp 1624635492
transform 1 0 10120 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 12972 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_8_111
timestamp 1624635492
transform 1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1624635492
transform 1 0 13248 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1624635492
transform 1 0 14260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_129
timestamp 1624635492
transform 1 0 12972 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1624635492
transform 1 0 14076 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1624635492
transform 1 0 14352 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1624635492
transform -1 0 15824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16008 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1624635492
transform 1 0 14536 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp 1624635492
transform 1 0 15364 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_160
timestamp 1624635492
transform 1 0 15824 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1624635492
transform 1 0 18032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1624635492
transform 1 0 17020 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_8_171
timestamp 1624635492
transform 1 0 16836 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1624635492
transform 1 0 17848 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_187
timestamp 1624635492
transform 1 0 18308 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 19780 0 -1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1624635492
transform -1 0 19320 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1624635492
transform 1 0 19504 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_198
timestamp 1624635492
transform 1 0 19320 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1624635492
transform 1 0 19596 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1624635492
transform -1 0 21896 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1624635492
transform 1 0 21252 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1624635492
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1624635492
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1624635492
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1624635492
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1624635492
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1624635492
transform 1 0 6348 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform 1 0 5796 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_58
timestamp 1624635492
transform 1 0 6440 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_62
timestamp 1624635492
transform 1 0 6808 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 8096 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7636 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1624635492
transform 1 0 7268 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6900 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1624635492
transform 1 0 7084 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_69
timestamp 1624635492
transform 1 0 7452 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1624635492
transform 1 0 7912 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9752 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_9_92
timestamp 1624635492
transform 1 0 9568 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12604 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1624635492
transform 1 0 11592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1624635492
transform 1 0 12144 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1624635492
transform -1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_110
timestamp 1624635492
transform 1 0 11224 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_115
timestamp 1624635492
transform 1 0 11684 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_118
timestamp 1624635492
transform 1 0 11960 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_123
timestamp 1624635492
transform 1 0 12420 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1624635492
transform 1 0 13616 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_134
timestamp 1624635492
transform 1 0 13432 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 1624635492
transform 1 0 14444 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 16560 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 14628 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_150
timestamp 1624635492
transform 1 0 14904 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18584 0 1 7072
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1624635492
transform 1 0 16836 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_168
timestamp 1624635492
transform 1 0 16560 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1624635492
transform 1 0 16928 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18768 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19872 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 1624635492
transform 1 0 18584 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp 1624635492
transform 1 0 19596 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1624635492
transform 1 0 20884 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1624635492
transform -1 0 21896 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp 1624635492
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_218
timestamp 1624635492
transform 1 0 21160 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1624635492
transform 1 0 21528 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1624635492
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1624635492
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1624635492
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1624635492
transform 1 0 3772 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_27
timestamp 1624635492
transform 1 0 3588 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_10_30
timestamp 1624635492
transform 1 0 3864 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_42
timestamp 1624635492
transform 1 0 4968 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_54
timestamp 1624635492
transform 1 0 6072 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_62
timestamp 1624635492
transform 1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1624635492
transform -1 0 8832 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1624635492
transform 1 0 8096 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1624635492
transform -1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1624635492
transform -1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6992 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_66
timestamp 1624635492
transform 1 0 7176 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1624635492
transform 1 0 7544 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_74
timestamp 1624635492
transform 1 0 7912 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1624635492
transform 1 0 8372 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9292 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11132 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1624635492
transform 1 0 9016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_84
timestamp 1624635492
transform 1 0 8832 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_87
timestamp 1624635492
transform 1 0 9108 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_98
timestamp 1624635492
transform 1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12512 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 12144 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_109
timestamp 1624635492
transform 1 0 11132 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_120
timestamp 1624635492
transform 1 0 12144 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1624635492
transform 1 0 14260 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1624635492
transform -1 0 14536 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_140
timestamp 1624635492
transform 1 0 13984 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 16376 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_10_146
timestamp 1624635492
transform 1 0 14536 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_166
timestamp 1624635492
transform 1 0 16376 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1624635492
transform 1 0 16836 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18216 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_170
timestamp 1624635492
transform 1 0 16744 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_174
timestamp 1624635492
transform 1 0 17112 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_186
timestamp 1624635492
transform 1 0 18216 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19780 0 -1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1624635492
transform -1 0 19228 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1624635492
transform 1 0 19504 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 1624635492
transform 1 0 19228 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_201
timestamp 1624635492
transform 1 0 19596 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1624635492
transform -1 0 21896 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_219
timestamp 1624635492
transform 1 0 21252 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1624635492
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1624635492
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1624635492
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1624635492
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1624635492
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1624635492
transform 1 0 6348 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_51
timestamp 1624635492
transform 1 0 5796 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_58
timestamp 1624635492
transform 1 0 6440 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_64
timestamp 1624635492
transform 1 0 6992 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1624635492
transform 1 0 7084 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_67
timestamp 1624635492
transform 1 0 7268 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1624635492
transform 1 0 7636 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_75
timestamp 1624635492
transform 1 0 8004 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8464 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1624635492
transform 1 0 8464 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1624635492
transform 1 0 8648 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11040 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9108 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1624635492
transform 1 0 8924 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_90
timestamp 1624635492
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 12144 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1624635492
transform 1 0 11592 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 11224 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 11684 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_108
timestamp 1624635492
transform 1 0 11040 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_112
timestamp 1624635492
transform 1 0 11408 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_117
timestamp 1624635492
transform 1 0 11868 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14260 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1624635492
transform -1 0 14076 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_136
timestamp 1624635492
transform 1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_141
timestamp 1624635492
transform 1 0 14076 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1624635492
transform -1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15824 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1624635492
transform 1 0 15088 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_157
timestamp 1624635492
transform 1 0 15548 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1624635492
transform -1 0 17388 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18400 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1624635492
transform 1 0 16836 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1624635492
transform 1 0 16652 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1624635492
transform 1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1624635492
transform 1 0 17388 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 21252 0 1 8160
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18768 0 1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_11_188
timestamp 1624635492
transform 1 0 18400 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_201
timestamp 1624635492
transform 1 0 19596 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1624635492
transform -1 0 21896 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1624635492
transform 1 0 21252 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1624635492
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1624635492
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1624635492
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1624635492
transform 1 0 3772 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_27
timestamp 1624635492
transform 1 0 3588 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_12_30
timestamp 1624635492
transform 1 0 3864 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_42
timestamp 1624635492
transform 1 0 4968 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_54
timestamp 1624635492
transform 1 0 6072 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8556 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 8188 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7820 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_66
timestamp 1624635492
transform 1 0 7176 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_72
timestamp 1624635492
transform 1 0 7728 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_75
timestamp 1624635492
transform 1 0 8004 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_79
timestamp 1624635492
transform 1 0 8372 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 9660 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1624635492
transform 1 0 9016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1624635492
transform -1 0 9292 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_84
timestamp 1624635492
transform 1 0 8832 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_89
timestamp 1624635492
transform 1 0 9292 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1624635492
transform 1 0 12328 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 12144 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_109
timestamp 1624635492
transform 1 0 11132 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1624635492
transform 1 0 12144 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_125
timestamp 1624635492
transform 1 0 12604 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13156 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1624635492
transform 1 0 14260 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 12788 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1624635492
transform 1 0 12972 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_140
timestamp 1624635492
transform 1 0 13984 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 1624635492
transform 1 0 14352 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 14536 0 -1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1624635492
transform 1 0 16192 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_162
timestamp 1624635492
transform 1 0 16008 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1624635492
transform -1 0 18032 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18216 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_12_173
timestamp 1624635492
transform 1 0 17020 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_184
timestamp 1624635492
transform 1 0 18032 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19964 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1624635492
transform 1 0 19504 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1624635492
transform -1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_195
timestamp 1624635492
transform 1 0 19044 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_199
timestamp 1624635492
transform 1 0 19412 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_203
timestamp 1624635492
transform 1 0 19780 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1624635492
transform 1 0 20976 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1624635492
transform -1 0 21896 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_214
timestamp 1624635492
transform 1 0 20792 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1624635492
transform 1 0 21252 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1624635492
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1624635492
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1624635492
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1624635492
transform 1 0 2484 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1624635492
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1624635492
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1624635492
transform 1 0 3772 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1624635492
transform 1 0 3588 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1624635492
transform 1 0 4692 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_27
timestamp 1624635492
transform 1 0 3588 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_30
timestamp 1624635492
transform 1 0 3864 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1624635492
transform 1 0 6348 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_51
timestamp 1624635492
transform 1 0 5796 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_58
timestamp 1624635492
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_42
timestamp 1624635492
transform 1 0 4968 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_54
timestamp 1624635492
transform 1 0 6072 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_70
timestamp 1624635492
transform 1 0 7544 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_80
timestamp 1624635492
transform 1 0 8464 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1624635492
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_77
timestamp 1624635492
transform 1 0 8188 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_74
timestamp 1624635492
transform 1 0 7912 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8004 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 8372 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 8280 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 8740 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1624635492
transform -1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_66
timestamp 1624635492
transform 1 0 7176 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_92
timestamp 1624635492
transform 1 0 9568 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_87
timestamp 1624635492
transform 1 0 9108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_84
timestamp 1624635492
transform 1 0 8832 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_89
timestamp 1624635492
transform 1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_85
timestamp 1624635492
transform 1 0 8924 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1624635492
transform -1 0 9292 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1624635492
transform -1 0 9568 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1624635492
transform -1 0 9752 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1624635492
transform 1 0 9016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_103
timestamp 1624635492
transform 1 0 10580 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1624635492
transform 1 0 10212 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_94
timestamp 1624635492
transform 1 0 9752 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1624635492
transform -1 0 10580 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 10212 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11224 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 10764 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12420 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1624635492
transform 1 0 11592 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_110
timestamp 1624635492
transform 1 0 11224 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1624635492
transform 1 0 11684 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1624635492
transform 1 0 12236 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13984 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13800 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1624635492
transform 1 0 14260 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_126
timestamp 1624635492
transform 1 0 12696 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_138
timestamp 1624635492
transform 1 0 13800 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_139
timestamp 1624635492
transform 1 0 13892 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1624635492
transform 1 0 14352 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_155
timestamp 1624635492
transform 1 0 15364 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_149
timestamp 1624635492
transform 1 0 14812 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14536 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1624635492
transform 1 0 14996 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_14_162
timestamp 1624635492
transform 1 0 16008 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_164
timestamp 1624635492
transform 1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1624635492
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1624635492
transform -1 0 16192 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 16008 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1624635492
transform -1 0 16652 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 16192 0 -1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 17112 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1624635492
transform 1 0 17848 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1624635492
transform 1 0 16836 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1624635492
transform 1 0 16652 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1624635492
transform 1 0 16928 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_180
timestamp 1624635492
transform 1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18768 0 1 9248
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 18860 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1624635492
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_190
timestamp 1624635492
transform 1 0 18584 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1624635492
transform 1 0 20240 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_191
timestamp 1624635492
transform 1 0 18676 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_196
timestamp 1624635492
transform 1 0 19136 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_201
timestamp 1624635492
transform 1 0 19596 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1624635492
transform -1 0 21068 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1624635492
transform 1 0 20424 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1624635492
transform -1 0 21896 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1624635492
transform -1 0 21896 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1624635492
transform -1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1624635492
transform 1 0 21252 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_212
timestamp 1624635492
transform 1 0 20608 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1624635492
transform 1 0 21068 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1624635492
transform 1 0 21436 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1624635492
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1624635492
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1624635492
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1624635492
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1624635492
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1624635492
transform 1 0 6348 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_51
timestamp 1624635492
transform 1 0 5796 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_58
timestamp 1624635492
transform 1 0 6440 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8740 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1624635492
transform -1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 7728 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7360 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_66
timestamp 1624635492
transform 1 0 7176 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1624635492
transform 1 0 7544 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1624635492
transform 1 0 7912 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1624635492
transform 1 0 8280 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_83
timestamp 1624635492
transform 1 0 8740 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9844 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1624635492
transform -1 0 9660 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 9200 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1624635492
transform 1 0 9200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_93
timestamp 1624635492
transform 1 0 9660 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1624635492
transform -1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1624635492
transform -1 0 13248 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1624635492
transform 1 0 11592 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_111
timestamp 1624635492
transform 1 0 11316 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_115
timestamp 1624635492
transform 1 0 11684 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_120
timestamp 1624635492
transform 1 0 12144 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1624635492
transform -1 0 14260 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_15_132
timestamp 1624635492
transform 1 0 13248 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_143
timestamp 1624635492
transform 1 0 14260 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1624635492
transform -1 0 16652 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 14720 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_15_147
timestamp 1624635492
transform 1 0 14628 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_157
timestamp 1624635492
transform 1 0 15548 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1624635492
transform -1 0 17940 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1624635492
transform 1 0 16836 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_169
timestamp 1624635492
transform 1 0 16652 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1624635492
transform 1 0 16928 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_183
timestamp 1624635492
transform 1 0 17940 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_187
timestamp 1624635492
transform 1 0 18308 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1624635492
transform -1 0 18676 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 20332 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1624635492
transform 1 0 18676 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20516 0 1 10336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1624635492
transform -1 0 21896 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_209
timestamp 1624635492
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_220
timestamp 1624635492
transform 1 0 21344 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1624635492
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1624635492
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1624635492
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1624635492
transform 1 0 3772 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1624635492
transform 1 0 3588 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1624635492
transform 1 0 3864 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1624635492
transform 1 0 4968 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_54
timestamp 1624635492
transform 1 0 6072 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1624635492
transform 1 0 6808 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1624635492
transform 1 0 8556 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1624635492
transform 1 0 8096 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1624635492
transform -1 0 7912 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 7360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6992 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_66
timestamp 1624635492
transform 1 0 7176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_70
timestamp 1624635492
transform 1 0 7544 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_74
timestamp 1624635492
transform 1 0 7912 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_79
timestamp 1624635492
transform 1 0 8372 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1624635492
transform 1 0 9016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_84
timestamp 1624635492
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1624635492
transform 1 0 9108 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1624635492
transform -1 0 11776 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11960 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1624635492
transform 1 0 10764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1624635492
transform 1 0 11776 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1624635492
transform -1 0 13800 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1624635492
transform 1 0 14260 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1624635492
transform 1 0 12788 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_138
timestamp 1624635492
transform 1 0 13800 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_142
timestamp 1624635492
transform 1 0 14168 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_144
timestamp 1624635492
transform 1 0 14352 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 16376 0 -1 11424
box -38 -48 1878 592
use sky130_fd_sc_hd__fill_2  FILLER_16_166
timestamp 1624635492
transform 1 0 16376 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 16560 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_16_184
timestamp 1624635492
transform 1 0 18032 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 19780 0 -1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1624635492
transform 1 0 18492 0 -1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1624635492
transform 1 0 19504 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_188
timestamp 1624635492
transform 1 0 18400 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1624635492
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_201
timestamp 1624635492
transform 1 0 19596 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1624635492
transform -1 0 21896 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1624635492
transform 1 0 21252 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1624635492
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1624635492
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1624635492
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1624635492
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1624635492
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1624635492
transform 1 0 6348 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_51
timestamp 1624635492
transform 1 0 5796 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_58
timestamp 1624635492
transform 1 0 6440 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 8372 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1624635492
transform -1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1624635492
transform -1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_70
timestamp 1624635492
transform 1 0 7544 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_73
timestamp 1624635492
transform 1 0 7820 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1624635492
transform 1 0 8188 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1624635492
transform 1 0 10028 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1624635492
transform 1 0 9844 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1624635492
transform 1 0 11040 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 11868 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1624635492
transform 1 0 11592 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1624635492
transform 1 0 10856 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_111
timestamp 1624635492
transform 1 0 11316 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_115
timestamp 1624635492
transform 1 0 11684 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1624635492
transform 1 0 13524 0 1 11424
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1624635492
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1624635492
transform 1 0 14352 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1624635492
transform 1 0 16376 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14720 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_17_164
timestamp 1624635492
transform 1 0 16192 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 19320 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 17388 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1624635492
transform 1 0 16836 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1624635492
transform 1 0 16652 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1624635492
transform 1 0 16928 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_177
timestamp 1624635492
transform 1 0 17388 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_181
timestamp 1624635492
transform 1 0 17756 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 21436 0 1 11424
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 19504 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_198
timestamp 1624635492
transform 1 0 19320 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1624635492
transform 1 0 19780 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1624635492
transform -1 0 21896 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1624635492
transform 1 0 21436 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1624635492
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1624635492
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1624635492
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1624635492
transform 1 0 3772 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_27
timestamp 1624635492
transform 1 0 3588 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_30
timestamp 1624635492
transform 1 0 3864 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_42
timestamp 1624635492
transform 1 0 4968 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_54
timestamp 1624635492
transform 1 0 6072 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_62
timestamp 1624635492
transform 1 0 6808 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8832 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1624635492
transform 1 0 8096 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1624635492
transform 1 0 7636 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1624635492
transform -1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6900 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_65
timestamp 1624635492
transform 1 0 7084 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_69
timestamp 1624635492
transform 1 0 7452 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_74
timestamp 1624635492
transform 1 0 7912 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_79
timestamp 1624635492
transform 1 0 8372 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10120 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 10764 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1624635492
transform 1 0 9016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_84
timestamp 1624635492
transform 1 0 8832 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1624635492
transform 1 0 9108 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_98
timestamp 1624635492
transform 1 0 10120 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1624635492
transform -1 0 12328 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12512 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1624635492
transform -1 0 11776 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_105
timestamp 1624635492
transform 1 0 10764 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_116
timestamp 1624635492
transform 1 0 11776 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1624635492
transform 1 0 12328 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1624635492
transform 1 0 14260 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_140
timestamp 1624635492
transform 1 0 13984 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_144
timestamp 1624635492
transform 1 0 14352 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 16008 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_18_162
timestamp 1624635492
transform 1 0 16008 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_166
timestamp 1624635492
transform 1 0 16376 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1624635492
transform 1 0 16468 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17480 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_18_176
timestamp 1624635492
transform 1 0 17296 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1624635492
transform 1 0 18308 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 21344 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1624635492
transform 1 0 18492 0 -1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1624635492
transform 1 0 19504 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_198
timestamp 1624635492
transform 1 0 19320 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_201
timestamp 1624635492
transform 1 0 19596 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1624635492
transform -1 0 21896 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1624635492
transform 1 0 21344 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1624635492
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1624635492
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1624635492
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1624635492
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1624635492
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1624635492
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1624635492
transform 1 0 3772 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1624635492
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1624635492
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_27
timestamp 1624635492
transform 1 0 3588 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_30
timestamp 1624635492
transform 1 0 3864 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1624635492
transform 1 0 6348 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6624 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_51
timestamp 1624635492
transform 1 0 5796 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_58
timestamp 1624635492
transform 1 0 6440 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 1624635492
transform 1 0 6808 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_42
timestamp 1624635492
transform 1 0 4968 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_54
timestamp 1624635492
transform 1 0 6072 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1624635492
transform 1 0 6808 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6900 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 6992 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1624635492
transform 1 0 7084 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_66
timestamp 1624635492
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7268 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7360 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_69
timestamp 1624635492
transform 1 0 7452 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1624635492
transform 1 0 7544 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 7912 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7728 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_79
timestamp 1624635492
transform 1 0 8372 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_74
timestamp 1624635492
transform 1 0 7912 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1624635492
transform 1 0 7912 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8096 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1624635492
transform 1 0 8556 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 9568 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_20_89
timestamp 1624635492
transform 1 0 9292 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_84
timestamp 1624635492
transform 1 0 8832 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_92
timestamp 1624635492
transform 1 0 9568 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1624635492
transform 1 0 9108 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1624635492
transform 1 0 9016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9476 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_98
timestamp 1624635492
transform 1 0 10120 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1624635492
transform 1 0 9752 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1624635492
transform 1 0 10396 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_96
timestamp 1624635492
transform 1 0 9936 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 9752 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 10120 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11408 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 11684 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1624635492
transform 1 0 11868 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1624635492
transform 1 0 11868 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 12420 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1624635492
transform 1 0 11592 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1624635492
transform 1 0 11408 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1624635492
transform 1 0 11684 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_120
timestamp 1624635492
transform 1 0 12144 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1624635492
transform 1 0 11684 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1624635492
transform 1 0 13064 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_126
timestamp 1624635492
transform 1 0 12696 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_132
timestamp 1624635492
transform 1 0 13248 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 12880 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13248 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 13432 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1624635492
transform 1 0 14352 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_141
timestamp 1624635492
transform 1 0 14076 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1624635492
transform 1 0 14260 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1624635492
transform 1 0 14260 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1624635492
transform -1 0 15272 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_153
timestamp 1624635492
transform 1 0 15180 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_148
timestamp 1624635492
transform 1 0 14720 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1624635492
transform 1 0 15272 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 14536 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 15180 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1624635492
transform 1 0 15364 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1624635492
transform 1 0 16192 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_158
timestamp 1624635492
transform 1 0 15640 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1624635492
transform 1 0 15732 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17848 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1624635492
transform -1 0 18216 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1624635492
transform 1 0 18032 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1624635492
transform 1 0 16836 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 16928 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_168
timestamp 1624635492
transform 1 0 16560 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_174
timestamp 1624635492
transform 1 0 17112 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_186
timestamp 1624635492
transform 1 0 18216 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1624635492
transform 1 0 17848 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_193
timestamp 1624635492
transform 1 0 18860 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1624635492
transform -1 0 19320 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_204
timestamp 1624635492
transform 1 0 19872 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_201
timestamp 1624635492
transform 1 0 19596 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_198
timestamp 1624635492
transform 1 0 19320 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_205
timestamp 1624635492
transform 1 0 19964 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 19688 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1624635492
transform 1 0 19504 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1624635492
transform 1 0 20056 0 -1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 19964 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1624635492
transform 1 0 20424 0 1 12512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1624635492
transform -1 0 21896 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1624635492
transform -1 0 21896 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output73
timestamp 1624635492
transform 1 0 21068 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_209
timestamp 1624635492
transform 1 0 20332 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1624635492
transform 1 0 21252 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_215
timestamp 1624635492
transform 1 0 20884 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1624635492
transform 1 0 21436 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1624635492
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1624635492
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1624635492
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1624635492
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1624635492
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1624635492
transform 1 0 6348 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6716 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_51
timestamp 1624635492
transform 1 0 5796 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_58
timestamp 1624635492
transform 1 0 6440 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_63
timestamp 1624635492
transform 1 0 6900 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 7084 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_67
timestamp 1624635492
transform 1 0 7268 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1624635492
transform 1 0 7452 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_71
timestamp 1624635492
transform 1 0 7636 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 7820 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 1624635492
transform 1 0 8004 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8464 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_80
timestamp 1624635492
transform 1 0 8464 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 8648 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11040 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9384 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_85
timestamp 1624635492
transform 1 0 8924 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1624635492
transform 1 0 9384 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12420 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12236 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1624635492
transform 1 0 11592 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1624635492
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_108
timestamp 1624635492
transform 1 0 11040 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_112
timestamp 1624635492
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_115
timestamp 1624635492
transform 1 0 11684 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1624635492
transform 1 0 12236 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1624635492
transform 1 0 14076 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1624635492
transform 1 0 13892 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1624635492
transform 1 0 15088 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1624635492
transform 1 0 15824 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_21_150
timestamp 1624635492
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_155
timestamp 1624635492
transform 1 0 15364 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_159
timestamp 1624635492
transform 1 0 15732 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 18584 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1624635492
transform 1 0 16836 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1624635492
transform 1 0 16652 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1624635492
transform 1 0 16928 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19872 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1624635492
transform 1 0 18860 0 1 13600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_21_190
timestamp 1624635492
transform 1 0 18584 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1624635492
transform 1 0 19688 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1624635492
transform -1 0 21896 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output84
timestamp 1624635492
transform 1 0 21068 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_213
timestamp 1624635492
transform 1 0 20700 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1624635492
transform 1 0 21436 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1624635492
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1624635492
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1624635492
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1624635492
transform 1 0 3772 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_27
timestamp 1624635492
transform 1 0 3588 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_30
timestamp 1624635492
transform 1 0 3864 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 6716 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 6348 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 5980 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5612 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_42
timestamp 1624635492
transform 1 0 4968 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_48
timestamp 1624635492
transform 1 0 5520 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1624635492
transform 1 0 5796 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1624635492
transform 1 0 6164 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_59
timestamp 1624635492
transform 1 0 6532 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1624635492
transform 1 0 7912 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform 1 0 7452 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7084 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_63
timestamp 1624635492
transform 1 0 6900 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_67
timestamp 1624635492
transform 1 0 7268 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1624635492
transform 1 0 7728 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_83
timestamp 1624635492
transform 1 0 8740 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9476 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1624635492
transform 1 0 9016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 9108 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1624635492
transform 1 0 9292 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13432 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12420 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11132 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1624635492
transform 1 0 10948 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 1624635492
transform 1 0 11960 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_123
timestamp 1624635492
transform 1 0 12420 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14076 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1624635492
transform 1 0 14260 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1624635492
transform 1 0 14352 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_134
timestamp 1624635492
transform 1 0 13432 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_141
timestamp 1624635492
transform 1 0 14076 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 14996 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1624635492
transform 1 0 15180 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_22_146
timestamp 1624635492
transform 1 0 14536 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1624635492
transform 1 0 14996 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_162
timestamp 1624635492
transform 1 0 16008 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_166
timestamp 1624635492
transform 1 0 16376 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1624635492
transform -1 0 18400 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 17940 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1624635492
transform 1 0 17940 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1624635492
transform -1 0 19320 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1624635492
transform -1 0 18860 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1624635492
transform 1 0 20056 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1624635492
transform 1 0 19504 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1624635492
transform -1 0 19780 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_188
timestamp 1624635492
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_193
timestamp 1624635492
transform 1 0 18860 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_198
timestamp 1624635492
transform 1 0 19320 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_203
timestamp 1624635492
transform 1 0 19780 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1624635492
transform -1 0 21896 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output85
timestamp 1624635492
transform 1 0 21068 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1624635492
transform 1 0 20884 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1624635492
transform 1 0 21436 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1624635492
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1624635492
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1624635492
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1624635492
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1624635492
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1624635492
transform 1 0 6348 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1624635492
transform -1 0 6716 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_51
timestamp 1624635492
transform 1 0 5796 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_58
timestamp 1624635492
transform 1 0 6440 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_61
timestamp 1624635492
transform 1 0 6716 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1624635492
transform 1 0 8096 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 7636 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 7268 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 6900 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1624635492
transform 1 0 7084 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_69
timestamp 1624635492
transform 1 0 7452 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1624635492
transform 1 0 7912 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1624635492
transform -1 0 11408 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1624635492
transform -1 0 10396 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9384 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 1624635492
transform 1 0 8924 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1624635492
transform 1 0 9384 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_101
timestamp 1624635492
transform 1 0 10396 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11868 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1624635492
transform 1 0 11592 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_112
timestamp 1624635492
transform 1 0 11408 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1624635492
transform 1 0 11684 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1624635492
transform 1 0 12880 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 13524 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_126
timestamp 1624635492
transform 1 0 12696 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_131
timestamp 1624635492
transform 1 0 13156 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15180 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_151
timestamp 1624635492
transform 1 0 14996 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1624635492
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1624635492
transform -1 0 18584 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1624635492
transform -1 0 18124 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1624635492
transform 1 0 16836 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_169
timestamp 1624635492
transform 1 0 16652 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_172
timestamp 1624635492
transform 1 0 16928 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1624635492
transform 1 0 17388 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1624635492
transform 1 0 17756 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1624635492
transform 1 0 18124 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1624635492
transform -1 0 19044 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 20700 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_23_190
timestamp 1624635492
transform 1 0 18584 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_195
timestamp 1624635492
transform 1 0 19044 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1624635492
transform -1 0 21896 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output86
timestamp 1624635492
transform 1 0 21068 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_213
timestamp 1624635492
transform 1 0 20700 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1624635492
transform 1 0 21436 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1624635492
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1624635492
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1624635492
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1624635492
transform 1 0 3772 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1624635492
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_30
timestamp 1624635492
transform 1 0 3864 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1624635492
transform -1 0 7176 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 5980 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1624635492
transform 1 0 5612 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_42
timestamp 1624635492
transform 1 0 4968 0 -1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_48
timestamp 1624635492
transform 1 0 5520 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_51
timestamp 1624635492
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_55
timestamp 1624635492
transform 1 0 6164 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 8832 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_66
timestamp 1624635492
transform 1 0 7176 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1624635492
transform 1 0 9292 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9936 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1624635492
transform 1 0 9016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_84
timestamp 1624635492
transform 1 0 8832 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1624635492
transform 1 0 9108 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_92
timestamp 1624635492
transform 1 0 9568 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 12052 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1624635492
transform 1 0 12236 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1624635492
transform 1 0 11408 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_119
timestamp 1624635492
transform 1 0 12052 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14076 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1624635492
transform 1 0 14260 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1624635492
transform 1 0 13064 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_141
timestamp 1624635492
transform 1 0 14076 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 1624635492
transform 1 0 14352 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1624635492
transform -1 0 15364 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1624635492
transform 1 0 15732 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_155
timestamp 1624635492
transform 1 0 15364 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1624635492
transform -1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 18768 0 -1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_24_168
timestamp 1624635492
transform 1 0 16560 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_173
timestamp 1624635492
transform 1 0 17020 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1624635492
transform 1 0 18952 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1624635492
transform 1 0 19504 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_192
timestamp 1624635492
transform 1 0 18768 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_197
timestamp 1624635492
transform 1 0 19228 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_201
timestamp 1624635492
transform 1 0 19596 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1624635492
transform -1 0 21896 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output87
timestamp 1624635492
transform 1 0 21068 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1624635492
transform 1 0 20608 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_216
timestamp 1624635492
transform 1 0 20976 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1624635492
transform 1 0 21436 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1624635492
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1624635492
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1624635492
transform 1 0 2484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1624635492
transform 1 0 4876 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1624635492
transform 1 0 3588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1624635492
transform 1 0 4692 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_43
timestamp 1624635492
transform 1 0 5060 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1624635492
transform -1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_47
timestamp 1624635492
transform 1 0 5428 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5612 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_51
timestamp 1624635492
transform 1 0 5796 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5980 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_55
timestamp 1624635492
transform 1 0 6164 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1624635492
transform 1 0 6348 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1624635492
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1624635492
transform 1 0 6716 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 8556 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1624635492
transform 1 0 8740 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_63
timestamp 1624635492
transform 1 0 6900 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1624635492
transform 1 0 8556 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10856 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 1624635492
transform 1 0 9568 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_96
timestamp 1624635492
transform 1 0 9936 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 11408 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1624635492
transform 1 0 11592 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_106
timestamp 1624635492
transform 1 0 10856 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1624635492
transform 1 0 11408 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_115
timestamp 1624635492
transform 1 0 11684 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 14536 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_25_126
timestamp 1624635492
transform 1 0 12696 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1624635492
transform -1 0 15548 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1624635492
transform 1 0 15732 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_25_146
timestamp 1624635492
transform 1 0 14536 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1624635492
transform 1 0 15548 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18308 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1624635492
transform 1 0 17296 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1624635492
transform 1 0 16836 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_168
timestamp 1624635492
transform 1 0 16560 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_174
timestamp 1624635492
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1624635492
transform 1 0 18124 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1624635492
transform 1 0 20056 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_25_203
timestamp 1624635492
transform 1 0 19780 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1624635492
transform -1 0 21896 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output88
timestamp 1624635492
transform 1 0 21068 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1624635492
transform 1 0 20884 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1624635492
transform 1 0 21436 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1624635492
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1624635492
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output72
timestamp 1624635492
transform -1 0 1932 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1624635492
transform -1 0 2300 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1624635492
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1624635492
transform 1 0 2484 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1624635492
transform 1 0 1380 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1624635492
transform 1 0 1932 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_13
timestamp 1624635492
transform 1 0 2300 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1624635492
transform 1 0 3772 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_27
timestamp 1624635492
transform 1 0 3588 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_30
timestamp 1624635492
transform 1 0 3864 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1624635492
transform 1 0 3404 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_37
timestamp 1624635492
transform 1 0 4508 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_51
timestamp 1624635492
transform 1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_47
timestamp 1624635492
transform 1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1624635492
transform 1 0 5888 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_48
timestamp 1624635492
transform 1 0 5520 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_42
timestamp 1624635492
transform 1 0 4968 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1624635492
transform -1 0 5428 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1624635492
transform 1 0 5336 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 5704 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 5796 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1624635492
transform 1 0 6716 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_58
timestamp 1624635492
transform 1 0 6440 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_55
timestamp 1624635492
transform 1 0 6164 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1624635492
transform 1 0 6348 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 5980 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1624635492
transform -1 0 6716 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 6348 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1624635492
transform 1 0 6348 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8004 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform -1 0 8372 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8832 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1624635492
transform -1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_75
timestamp 1624635492
transform 1 0 8004 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_79
timestamp 1624635492
transform 1 0 8372 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1624635492
transform 1 0 8372 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1624635492
transform 1 0 8740 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp 1624635492
transform 1 0 9108 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1624635492
transform 1 0 9292 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_84
timestamp 1624635492
transform 1 0 8832 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1624635492
transform 1 0 9108 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1624635492
transform 1 0 9016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 9108 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform 1 0 9476 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1624635492
transform -1 0 10120 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1624635492
transform 1 0 10120 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_99
timestamp 1624635492
transform 1 0 10212 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1624635492
transform 1 0 9752 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1624635492
transform 1 0 10304 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1624635492
transform -1 0 10212 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 11960 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1624635492
transform -1 0 12512 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 12144 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1624635492
transform 1 0 11592 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1624635492
transform -1 0 11868 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_118
timestamp 1624635492
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_109
timestamp 1624635492
transform 1 0 11132 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1624635492
transform 1 0 11500 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_117
timestamp 1624635492
transform 1 0 11868 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_124
timestamp 1624635492
transform 1 0 12512 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1624635492
transform 1 0 13800 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 12696 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1624635492
transform 1 0 14260 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1624635492
transform 1 0 14352 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_136
timestamp 1624635492
transform 1 0 13616 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1624635492
transform 1 0 14076 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_144
timestamp 1624635492
transform 1 0 14352 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_142
timestamp 1624635492
transform 1 0 14168 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_146
timestamp 1624635492
transform 1 0 14536 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_155
timestamp 1624635492
transform 1 0 15364 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1624635492
transform 1 0 14720 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1624635492
transform -1 0 15364 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_27_157
timestamp 1624635492
transform 1 0 15548 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1624635492
transform 1 0 16284 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_160
timestamp 1624635492
transform 1 0 15824 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1624635492
transform 1 0 15824 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1624635492
transform -1 0 16284 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1624635492
transform 1 0 15548 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1624635492
transform 1 0 16928 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_169
timestamp 1624635492
transform 1 0 16652 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1624635492
transform 1 0 17296 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1624635492
transform 1 0 16836 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1624635492
transform 1 0 17112 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1624635492
transform 1 0 16468 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_27_183
timestamp 1624635492
transform 1 0 17940 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_185
timestamp 1624635492
transform 1 0 18124 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_181
timestamp 1624635492
transform 1 0 17756 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17940 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1624635492
transform 1 0 18308 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1624635492
transform 1 0 17480 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 18124 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1624635492
transform 1 0 19780 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1624635492
transform -1 0 20608 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1624635492
transform 1 0 19504 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 20240 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_196
timestamp 1624635492
transform 1 0 19136 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_201
timestamp 1624635492
transform 1 0 19596 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1624635492
transform 1 0 20056 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1624635492
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1624635492
transform 1 0 20608 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1624635492
transform 1 0 20424 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1624635492
transform -1 0 20884 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1624635492
transform 1 0 20976 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1624635492
transform 1 0 20884 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output90
timestamp 1624635492
transform 1 0 21068 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output89
timestamp 1624635492
transform 1 0 21068 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1624635492
transform 1 0 21436 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1624635492
transform 1 0 21436 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1624635492
transform -1 0 21896 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1624635492
transform -1 0 21896 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1624635492
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1624635492
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1624635492
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1624635492
transform 1 0 3772 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_27
timestamp 1624635492
transform 1 0 3588 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_30
timestamp 1624635492
transform 1 0 3864 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1624635492
transform -1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1624635492
transform 1 0 6348 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1624635492
transform 1 0 5980 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_42
timestamp 1624635492
transform 1 0 4968 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_48
timestamp 1624635492
transform 1 0 5520 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1624635492
transform 1 0 5796 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_55
timestamp 1624635492
transform 1 0 6164 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_59
timestamp 1624635492
transform 1 0 6532 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1624635492
transform -1 0 8280 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_mem_bottom_track_1.prog_clk
timestamp 1624635492
transform -1 0 8832 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1624635492
transform -1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1624635492
transform 1 0 6900 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1624635492
transform 1 0 7268 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_78
timestamp 1624635492
transform 1 0 8280 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform -1 0 10764 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1624635492
transform 1 0 9016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_84
timestamp 1624635492
transform 1 0 8832 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_87
timestamp 1624635492
transform 1 0 9108 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1624635492
transform -1 0 11776 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1624635492
transform -1 0 11316 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11960 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_28_105
timestamp 1624635492
transform 1 0 10764 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1624635492
transform 1 0 11316 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1624635492
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13800 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1624635492
transform 1 0 14260 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1624635492
transform 1 0 12788 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_138
timestamp 1624635492
transform 1 0 13800 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_142
timestamp 1624635492
transform 1 0 14168 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_144
timestamp 1624635492
transform 1 0 14352 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform -1 0 17388 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1624635492
transform 1 0 14536 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1624635492
transform -1 0 15732 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_155
timestamp 1624635492
transform 1 0 15364 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_159
timestamp 1624635492
transform 1 0 15732 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 17572 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1624635492
transform 1 0 17388 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1624635492
transform 1 0 19780 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1624635492
transform 1 0 19504 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_195
timestamp 1624635492
transform 1 0 19044 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_199
timestamp 1624635492
transform 1 0 19412 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_201
timestamp 1624635492
transform 1 0 19596 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1624635492
transform -1 0 21896 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output91
timestamp 1624635492
transform 1 0 21068 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_212
timestamp 1624635492
transform 1 0 20608 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_216
timestamp 1624635492
transform 1 0 20976 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1624635492
transform 1 0 21436 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1624635492
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1624635492
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1624635492
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1624635492
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1624635492
transform 1 0 4692 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1624635492
transform 1 0 5060 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_47
timestamp 1624635492
transform 1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 5428 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1624635492
transform 1 0 5612 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_51
timestamp 1624635492
transform 1 0 5796 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1624635492
transform -1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_55
timestamp 1624635492
transform 1 0 6164 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_58
timestamp 1624635492
transform 1 0 6440 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1624635492
transform 1 0 6348 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_61
timestamp 1624635492
transform 1 0 6716 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1624635492
transform -1 0 6716 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 7636 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1624635492
transform -1 0 7452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1624635492
transform -1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1624635492
transform 1 0 7084 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_69
timestamp 1624635492
transform 1 0 7452 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1624635492
transform -1 0 10948 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1624635492
transform 1 0 9384 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_29_87
timestamp 1624635492
transform 1 0 9108 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_99
timestamp 1624635492
transform 1 0 10212 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_103
timestamp 1624635492
transform 1 0 10580 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1624635492
transform -1 0 11408 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1624635492
transform 1 0 11868 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1624635492
transform 1 0 11592 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_107
timestamp 1624635492
transform 1 0 10948 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_112
timestamp 1624635492
transform 1 0 11408 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_115
timestamp 1624635492
transform 1 0 11684 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1624635492
transform -1 0 14904 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1624635492
transform 1 0 13064 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1624635492
transform 1 0 12696 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1624635492
transform 1 0 13892 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 15180 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_29_150
timestamp 1624635492
transform 1 0 14904 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1624635492
transform -1 0 17664 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 17848 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1624635492
transform 1 0 16836 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1624635492
transform 1 0 17020 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_169
timestamp 1624635492
transform 1 0 16652 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_172
timestamp 1624635492
transform 1 0 16928 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1624635492
transform 1 0 17204 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_180
timestamp 1624635492
transform 1 0 17664 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1624635492
transform -1 0 20332 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_29_198
timestamp 1624635492
transform 1 0 19320 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1624635492
transform -1 0 21896 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output74
timestamp 1624635492
transform 1 0 21068 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output92
timestamp 1624635492
transform 1 0 20516 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1624635492
transform 1 0 20332 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1624635492
transform 1 0 20884 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1624635492
transform 1 0 21436 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1624635492
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1624635492
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1624635492
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1624635492
transform 1 0 3772 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1624635492
transform -1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1624635492
transform -1 0 4692 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1624635492
transform -1 0 4324 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_27
timestamp 1624635492
transform 1 0 3588 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_30
timestamp 1624635492
transform 1 0 3864 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1624635492
transform 1 0 4324 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_39
timestamp 1624635492
transform 1 0 4692 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1624635492
transform -1 0 6532 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1624635492
transform -1 0 6164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1624635492
transform -1 0 5796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1624635492
transform -1 0 5428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1624635492
transform 1 0 5060 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1624635492
transform 1 0 5428 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_51
timestamp 1624635492
transform 1 0 5796 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_55
timestamp 1624635492
transform 1 0 6164 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_59
timestamp 1624635492
transform 1 0 6532 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1624635492
transform -1 0 8832 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 8372 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 7912 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1624635492
transform -1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1624635492
transform -1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_65
timestamp 1624635492
transform 1 0 7084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_69
timestamp 1624635492
transform 1 0 7452 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_74
timestamp 1624635492
transform 1 0 7912 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_79
timestamp 1624635492
transform 1 0 8372 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 9292 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1624635492
transform 1 0 9016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_84
timestamp 1624635492
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_87
timestamp 1624635492
transform 1 0 9108 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1624635492
transform -1 0 11776 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1624635492
transform 1 0 11960 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_105
timestamp 1624635492
transform 1 0 10764 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_116
timestamp 1624635492
transform 1 0 11776 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1624635492
transform 1 0 12972 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1624635492
transform 1 0 13432 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1624635492
transform 1 0 14260 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1624635492
transform -1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_127
timestamp 1624635492
transform 1 0 12788 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_132
timestamp 1624635492
transform 1 0 13248 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_137
timestamp 1624635492
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_141
timestamp 1624635492
transform 1 0 14076 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1624635492
transform 1 0 14352 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 14536 0 -1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1624635492
transform 1 0 16192 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_30_162
timestamp 1624635492
transform 1 0 16008 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1624635492
transform -1 0 18400 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1624635492
transform 1 0 17664 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1624635492
transform 1 0 17204 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_173
timestamp 1624635492
transform 1 0 17020 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1624635492
transform 1 0 17480 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1624635492
transform 1 0 17940 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1624635492
transform -1 0 19320 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1624635492
transform -1 0 18860 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1624635492
transform 1 0 19504 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output123
timestamp 1624635492
transform 1 0 19964 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1624635492
transform -1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1624635492
transform 1 0 18400 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_193
timestamp 1624635492
transform 1 0 18860 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_198
timestamp 1624635492
transform 1 0 19320 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1624635492
transform 1 0 19780 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1624635492
transform -1 0 21896 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output75
timestamp 1624635492
transform 1 0 21068 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output120
timestamp 1624635492
transform 1 0 20516 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1624635492
transform 1 0 20332 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1624635492
transform 1 0 20884 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1624635492
transform 1 0 21436 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1624635492
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1624635492
transform -1 0 2116 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1624635492
transform -1 0 2576 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1624635492
transform -1 0 1564 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_5
timestamp 1624635492
transform 1 0 1564 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_31_11
timestamp 1624635492
transform 1 0 2116 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_16
timestamp 1624635492
transform 1 0 2576 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1624635492
transform -1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1624635492
transform -1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_28
timestamp 1624635492
transform 1 0 3680 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_36
timestamp 1624635492
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_40
timestamp 1624635492
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_44
timestamp 1624635492
transform 1 0 5152 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1624635492
transform -1 0 5152 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_51
timestamp 1624635492
transform 1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_48
timestamp 1624635492
transform 1 0 5520 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1624635492
transform -1 0 5796 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_55
timestamp 1624635492
transform 1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1624635492
transform -1 0 6164 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_61
timestamp 1624635492
transform 1 0 6716 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_58
timestamp 1624635492
transform 1 0 6440 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1624635492
transform -1 0 6716 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1624635492
transform 1 0 6348 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1624635492
transform -1 0 8832 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1624635492
transform -1 0 8372 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1624635492
transform -1 0 7912 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 7452 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_65
timestamp 1624635492
transform 1 0 7084 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_69
timestamp 1624635492
transform 1 0 7452 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1624635492
transform 1 0 7912 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_79
timestamp 1624635492
transform 1 0 8372 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1624635492
transform -1 0 9752 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1624635492
transform -1 0 9292 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 9936 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_84
timestamp 1624635492
transform 1 0 8832 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_89
timestamp 1624635492
transform 1 0 9292 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_94
timestamp 1624635492
transform 1 0 9752 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1624635492
transform 1 0 11868 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1624635492
transform 1 0 11592 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_112
timestamp 1624635492
transform 1 0 11408 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_115
timestamp 1624635492
transform 1 0 11684 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1624635492
transform 1 0 13524 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_31_133
timestamp 1624635492
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1624635492
transform 1 0 16192 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1624635492
transform -1 0 16008 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_31_151
timestamp 1624635492
transform 1 0 14996 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_162
timestamp 1624635492
transform 1 0 16008 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1624635492
transform -1 0 18216 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1624635492
transform -1 0 17756 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1624635492
transform 1 0 16836 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1624635492
transform -1 0 17112 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_167
timestamp 1624635492
transform 1 0 16468 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_174
timestamp 1624635492
transform 1 0 17112 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_181
timestamp 1624635492
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_186
timestamp 1624635492
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1624635492
transform -1 0 19596 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1624635492
transform -1 0 19136 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1624635492
transform -1 0 18676 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1624635492
transform -1 0 20884 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1624635492
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1624635492
transform 1 0 19136 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 1624635492
transform 1 0 19596 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1624635492
transform -1 0 21896 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output76
timestamp 1624635492
transform 1 0 21068 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1624635492
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1624635492
transform 1 0 21436 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1624635492
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1624635492
transform 1 0 2116 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1624635492
transform 1 0 2576 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1624635492
transform 1 0 1564 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1624635492
transform 1 0 1380 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_9
timestamp 1624635492
transform 1 0 1932 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_14
timestamp 1624635492
transform 1 0 2392 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_19
timestamp 1624635492
transform 1 0 2852 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_23
timestamp 1624635492
transform 1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1624635492
transform -1 0 3220 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_27
timestamp 1624635492
transform 1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1624635492
transform -1 0 3588 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_32
timestamp 1624635492
transform 1 0 4048 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1624635492
transform -1 0 4048 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1624635492
transform 1 0 3772 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1624635492
transform -1 0 4508 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_37
timestamp 1624635492
transform 1 0 4508 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1624635492
transform -1 0 4968 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1624635492
transform -1 0 6808 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1624635492
transform -1 0 6348 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1624635492
transform -1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1624635492
transform -1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1624635492
transform 1 0 4968 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_48
timestamp 1624635492
transform 1 0 5520 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_52
timestamp 1624635492
transform 1 0 5888 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_57
timestamp 1624635492
transform 1 0 6348 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_62
timestamp 1624635492
transform 1 0 6808 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1624635492
transform -1 0 8832 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1624635492
transform -1 0 8372 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1624635492
transform -1 0 7912 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1624635492
transform -1 0 7268 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_67
timestamp 1624635492
transform 1 0 7268 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_74
timestamp 1624635492
transform 1 0 7912 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_79
timestamp 1624635492
transform 1 0 8372 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1624635492
transform -1 0 9660 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1624635492
transform -1 0 10672 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1624635492
transform 1 0 9016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_84
timestamp 1624635492
transform 1 0 8832 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_87
timestamp 1624635492
transform 1 0 9108 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1624635492
transform 1 0 9660 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_104
timestamp 1624635492
transform 1 0 10672 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1624635492
transform 1 0 10948 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1624635492
transform 1 0 12420 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1624635492
transform 1 0 13800 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1624635492
transform -1 0 13616 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1624635492
transform 1 0 14260 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1624635492
transform 1 0 13616 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1624635492
transform 1 0 14076 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1624635492
transform 1 0 14352 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  output127
timestamp 1624635492
transform -1 0 14904 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output128
timestamp 1624635492
transform -1 0 15456 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output129
timestamp 1624635492
transform -1 0 16008 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output130
timestamp 1624635492
transform -1 0 16560 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_150
timestamp 1624635492
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_156
timestamp 1624635492
transform 1 0 15456 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1624635492
transform 1 0 16008 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1624635492
transform -1 0 18216 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output131
timestamp 1624635492
transform -1 0 17112 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output132
timestamp 1624635492
transform -1 0 17664 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1624635492
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_174
timestamp 1624635492
transform 1 0 17112 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_180
timestamp 1624635492
transform 1 0 17664 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1624635492
transform 1 0 18216 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1624635492
transform 1 0 19504 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output117
timestamp 1624635492
transform -1 0 20148 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output121
timestamp 1624635492
transform 1 0 18952 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output122
timestamp 1624635492
transform 1 0 18400 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_192
timestamp 1624635492
transform 1 0 18768 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_198
timestamp 1624635492
transform 1 0 19320 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1624635492
transform 1 0 19596 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_207
timestamp 1624635492
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1624635492
transform -1 0 21896 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output77
timestamp 1624635492
transform 1 0 21068 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output118
timestamp 1624635492
transform -1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_213
timestamp 1624635492
transform 1 0 20700 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1624635492
transform 1 0 21436 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1624635492
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1624635492
transform 1 0 2484 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1624635492
transform 1 0 1932 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1624635492
transform 1 0 1564 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1624635492
transform 1 0 1380 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1624635492
transform 1 0 1748 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1624635492
transform 1 0 2300 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_18
timestamp 1624635492
transform 1 0 2760 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1624635492
transform 1 0 3772 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1624635492
transform 1 0 3036 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1624635492
transform 1 0 4048 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1624635492
transform 1 0 4600 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_25
timestamp 1624635492
transform 1 0 3404 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_30
timestamp 1624635492
transform 1 0 3864 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_36
timestamp 1624635492
transform 1 0 4416 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1624635492
transform 1 0 6440 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1624635492
transform 1 0 6716 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1624635492
transform 1 0 5244 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1624635492
transform -1 0 6164 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_42
timestamp 1624635492
transform 1 0 4968 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1624635492
transform 1 0 5612 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_55
timestamp 1624635492
transform 1 0 6164 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1624635492
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1624635492
transform -1 0 8924 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1624635492
transform 1 0 7544 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1624635492
transform 1 0 8096 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_65
timestamp 1624635492
transform 1 0 7084 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_69
timestamp 1624635492
transform 1 0 7452 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1624635492
transform 1 0 7912 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_80
timestamp 1624635492
transform 1 0 8464 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1624635492
transform 1 0 9108 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1624635492
transform -1 0 9752 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1624635492
transform 1 0 9936 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1624635492
transform -1 0 10856 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1624635492
transform 1 0 8924 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_88
timestamp 1624635492
transform 1 0 9200 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_94
timestamp 1624635492
transform 1 0 9752 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_100
timestamp 1624635492
transform 1 0 10304 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1624635492
transform 1 0 11776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1624635492
transform -1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output113
timestamp 1624635492
transform -1 0 12420 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output124
timestamp 1624635492
transform -1 0 12972 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_106
timestamp 1624635492
transform 1 0 10856 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_112
timestamp 1624635492
transform 1 0 11408 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1624635492
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1624635492
transform 1 0 12420 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1624635492
transform 1 0 14444 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output125
timestamp 1624635492
transform -1 0 13524 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output126
timestamp 1624635492
transform -1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_129
timestamp 1624635492
transform 1 0 12972 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_135
timestamp 1624635492
transform 1 0 13524 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1624635492
transform 1 0 14076 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output115
timestamp 1624635492
transform 1 0 16008 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output116
timestamp 1624635492
transform 1 0 15456 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output119
timestamp 1624635492
transform 1 0 14904 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1624635492
transform -1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_148
timestamp 1624635492
transform 1 0 14720 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1624635492
transform 1 0 15272 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1624635492
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1624635492
transform 1 0 16376 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1624635492
transform 1 0 17112 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output82
timestamp 1624635492
transform 1 0 18124 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output83
timestamp 1624635492
transform 1 0 17572 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output114
timestamp 1624635492
transform 1 0 16560 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1624635492
transform -1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_172
timestamp 1624635492
transform 1 0 16928 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1624635492
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_183
timestamp 1624635492
transform 1 0 17940 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1624635492
transform -1 0 20332 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1624635492
transform 1 0 19780 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output80
timestamp 1624635492
transform 1 0 19228 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output81
timestamp 1624635492
transform 1 0 18676 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1624635492
transform 1 0 18492 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_195
timestamp 1624635492
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1624635492
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_204
timestamp 1624635492
transform 1 0 19872 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1624635492
transform -1 0 21896 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output78
timestamp 1624635492
transform 1 0 21068 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output79
timestamp 1624635492
transform 1 0 20516 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1624635492
transform 1 0 20332 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1624635492
transform 1 0 20884 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1624635492
transform 1 0 21436 0 1 20128
box -38 -48 222 592
<< labels >>
rlabel metal2 s 294 0 350 800 6 bottom_left_grid_pin_1_
port 0 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 1 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 2 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 3 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 4 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 5 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 6 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 7 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 8 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 9 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 10 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 11 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 12 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 13 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 14 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 15 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 16 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 17 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 18 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 19 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 20 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 21 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 22 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 23 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 24 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 25 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 26 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 27 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 28 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 29 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 30 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 31 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 32 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 33 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 34 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 35 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 36 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 37 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 38 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 39 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 40 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 41 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 42 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 chany_bottom_in[0]
port 43 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[10]
port 44 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[11]
port 45 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[12]
port 46 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[13]
port 47 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[14]
port 48 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[15]
port 49 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[16]
port 50 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[17]
port 51 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[18]
port 52 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[19]
port 53 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_in[1]
port 54 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 chany_bottom_in[2]
port 55 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_in[3]
port 56 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_in[4]
port 57 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_in[5]
port 58 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[6]
port 59 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[7]
port 60 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[8]
port 61 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[9]
port 62 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_out[0]
port 63 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[10]
port 64 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[11]
port 65 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[12]
port 66 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[13]
port 67 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 68 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[15]
port 69 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[16]
port 70 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[17]
port 71 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[18]
port 72 nsew signal tristate
rlabel metal2 s 22650 0 22706 800 6 chany_bottom_out[19]
port 73 nsew signal tristate
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_out[1]
port 74 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[2]
port 75 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[3]
port 76 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 77 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 78 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[6]
port 79 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 80 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[8]
port 81 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[9]
port 82 nsew signal tristate
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 83 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 84 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 85 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 86 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 87 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 88 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 89 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 90 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 91 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 92 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 93 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 94 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 95 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 96 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 97 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 98 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 99 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 100 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 101 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 102 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 103 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 104 nsew signal tristate
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 105 nsew signal tristate
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 106 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 107 nsew signal tristate
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 108 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 109 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 110 nsew signal tristate
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 111 nsew signal tristate
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 112 nsew signal tristate
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 113 nsew signal tristate
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 114 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 115 nsew signal tristate
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 116 nsew signal tristate
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 117 nsew signal tristate
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 118 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 119 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 120 nsew signal tristate
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 121 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 122 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 123 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 124 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 125 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 126 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 127 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 128 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 129 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 130 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 131 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 132 nsew signal input
rlabel metal4 s 18271 2128 18591 20720 6 VPWR
port 133 nsew power bidirectional
rlabel metal4 s 11340 2128 11660 20720 6 VPWR
port 134 nsew power bidirectional
rlabel metal4 s 4409 2128 4729 20720 6 VPWR
port 135 nsew power bidirectional
rlabel metal4 s 14805 2128 15125 20720 6 VGND
port 136 nsew ground bidirectional
rlabel metal4 s 7875 2128 8195 20720 6 VGND
port 137 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
