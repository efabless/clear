magic
tech sky130A
magscale 1 2
timestamp 1679319512
<< viali >>
rect 45201 54281 45235 54315
rect 3249 54213 3283 54247
rect 5825 54213 5859 54247
rect 8401 54213 8435 54247
rect 10977 54213 11011 54247
rect 13553 54213 13587 54247
rect 16129 54213 16163 54247
rect 18705 54213 18739 54247
rect 21005 54213 21039 54247
rect 28733 54213 28767 54247
rect 32965 54213 32999 54247
rect 33701 54213 33735 54247
rect 37565 54213 37599 54247
rect 42717 54213 42751 54247
rect 2237 54145 2271 54179
rect 4169 54145 4203 54179
rect 4813 54145 4847 54179
rect 7389 54145 7423 54179
rect 9781 54145 9815 54179
rect 12541 54145 12575 54179
rect 15117 54145 15151 54179
rect 17693 54145 17727 54179
rect 20269 54145 20303 54179
rect 22753 54145 22787 54179
rect 24777 54145 24811 54179
rect 25513 54145 25547 54179
rect 26433 54145 26467 54179
rect 27169 54145 27203 54179
rect 27905 54145 27939 54179
rect 29929 54145 29963 54179
rect 30665 54145 30699 54179
rect 31401 54145 31435 54179
rect 34897 54145 34931 54179
rect 35817 54145 35851 54179
rect 36553 54145 36587 54179
rect 38761 54145 38795 54179
rect 40049 54145 40083 54179
rect 40785 54145 40819 54179
rect 41705 54145 41739 54179
rect 43729 54145 43763 54179
rect 44373 54145 44407 54179
rect 45385 54145 45419 54179
rect 46581 54145 46615 54179
rect 47225 54145 47259 54179
rect 47961 54145 47995 54179
rect 23029 54077 23063 54111
rect 48421 54077 48455 54111
rect 28917 54009 28951 54043
rect 33149 54009 33183 54043
rect 33885 54009 33919 54043
rect 42993 54009 43027 54043
rect 3985 53941 4019 53975
rect 24961 53941 24995 53975
rect 25697 53941 25731 53975
rect 26249 53941 26283 53975
rect 27353 53941 27387 53975
rect 28089 53941 28123 53975
rect 30113 53941 30147 53975
rect 30849 53941 30883 53975
rect 31585 53941 31619 53975
rect 35081 53941 35115 53975
rect 36001 53941 36035 53975
rect 36737 53941 36771 53975
rect 37657 53941 37691 53975
rect 38945 53941 38979 53975
rect 40233 53941 40267 53975
rect 40969 53941 41003 53975
rect 41521 53941 41555 53975
rect 43545 53941 43579 53975
rect 44189 53941 44223 53975
rect 46397 53941 46431 53975
rect 47041 53941 47075 53975
rect 23673 53669 23707 53703
rect 2421 53601 2455 53635
rect 5733 53601 5767 53635
rect 7573 53601 7607 53635
rect 10885 53601 10919 53635
rect 12725 53601 12759 53635
rect 16129 53601 16163 53635
rect 18337 53601 18371 53635
rect 20453 53601 20487 53635
rect 22293 53601 22327 53635
rect 47317 53601 47351 53635
rect 2145 53533 2179 53567
rect 5457 53533 5491 53567
rect 7297 53533 7331 53567
rect 10425 53533 10459 53567
rect 12357 53533 12391 53567
rect 15853 53533 15887 53567
rect 17693 53533 17727 53567
rect 20177 53533 20211 53567
rect 22017 53533 22051 53567
rect 23857 53533 23891 53567
rect 24685 53533 24719 53567
rect 29929 53533 29963 53567
rect 32321 53533 32355 53567
rect 35265 53533 35299 53567
rect 38209 53533 38243 53567
rect 41889 53533 41923 53567
rect 46857 53533 46891 53567
rect 49249 53533 49283 53567
rect 24869 53465 24903 53499
rect 29745 53397 29779 53431
rect 32137 53397 32171 53431
rect 35081 53397 35115 53431
rect 38025 53397 38059 53431
rect 41705 53397 41739 53431
rect 49065 53397 49099 53431
rect 46121 53193 46155 53227
rect 46857 53193 46891 53227
rect 49157 53125 49191 53159
rect 1685 53057 1719 53091
rect 2881 53057 2915 53091
rect 4813 53057 4847 53091
rect 8033 53057 8067 53091
rect 9781 53057 9815 53091
rect 13185 53057 13219 53091
rect 15025 53057 15059 53091
rect 17601 53057 17635 53091
rect 19625 53057 19659 53091
rect 46305 53057 46339 53091
rect 47041 53057 47075 53091
rect 48145 53057 48179 53091
rect 3157 52989 3191 53023
rect 5089 52989 5123 53023
rect 8309 52989 8343 53023
rect 10241 52989 10275 53023
rect 13461 52989 13495 53023
rect 15393 52989 15427 53023
rect 17877 52989 17911 53023
rect 20085 52989 20119 53023
rect 1777 52853 1811 52887
rect 2053 52513 2087 52547
rect 4629 52513 4663 52547
rect 9781 52513 9815 52547
rect 14933 52513 14967 52547
rect 1777 52445 1811 52479
rect 4353 52445 4387 52479
rect 9505 52445 9539 52479
rect 14657 52445 14691 52479
rect 49341 52445 49375 52479
rect 49157 52309 49191 52343
rect 23581 52105 23615 52139
rect 2789 52037 2823 52071
rect 1593 51969 1627 52003
rect 23765 51969 23799 52003
rect 49065 51969 49099 52003
rect 49249 51765 49283 51799
rect 13093 51561 13127 51595
rect 14473 51561 14507 51595
rect 24685 51561 24719 51595
rect 24869 51357 24903 51391
rect 49065 51357 49099 51391
rect 13001 51289 13035 51323
rect 14381 51289 14415 51323
rect 49249 51221 49283 51255
rect 22201 51017 22235 51051
rect 23305 50949 23339 50983
rect 1685 50881 1719 50915
rect 22109 50881 22143 50915
rect 23121 50881 23155 50915
rect 48973 50881 49007 50915
rect 1869 50745 1903 50779
rect 49065 50677 49099 50711
rect 20269 50473 20303 50507
rect 49065 50269 49099 50303
rect 20177 50201 20211 50235
rect 49249 50133 49283 50167
rect 12357 49929 12391 49963
rect 14749 49929 14783 49963
rect 49249 49929 49283 49963
rect 12265 49861 12299 49895
rect 14657 49793 14691 49827
rect 49065 49793 49099 49827
rect 18061 49385 18095 49419
rect 20361 49385 20395 49419
rect 17969 49181 18003 49215
rect 49065 49181 49099 49215
rect 20269 49113 20303 49147
rect 49249 49045 49283 49079
rect 49065 48705 49099 48739
rect 49249 48501 49283 48535
rect 47961 48229 47995 48263
rect 48881 48229 48915 48263
rect 10149 48161 10183 48195
rect 48145 48093 48179 48127
rect 48697 48093 48731 48127
rect 1685 48025 1719 48059
rect 1869 48025 1903 48059
rect 10425 48025 10459 48059
rect 12173 48025 12207 48059
rect 24685 47753 24719 47787
rect 24869 47617 24903 47651
rect 49065 47617 49099 47651
rect 49249 47413 49283 47447
rect 48237 47209 48271 47243
rect 48789 47209 48823 47243
rect 48973 47005 49007 47039
rect 48145 46937 48179 46971
rect 49341 46529 49375 46563
rect 49157 46325 49191 46359
rect 18429 46121 18463 46155
rect 26709 46121 26743 46155
rect 18613 45917 18647 45951
rect 19717 45917 19751 45951
rect 26893 45917 26927 45951
rect 48145 45917 48179 45951
rect 1685 45849 1719 45883
rect 49157 45849 49191 45883
rect 1777 45781 1811 45815
rect 19533 45781 19567 45815
rect 48605 45577 48639 45611
rect 15117 45509 15151 45543
rect 33885 45509 33919 45543
rect 33977 45509 34011 45543
rect 14933 45441 14967 45475
rect 32689 45441 32723 45475
rect 32781 45441 32815 45475
rect 48145 45441 48179 45475
rect 48789 45441 48823 45475
rect 32873 45373 32907 45407
rect 34161 45373 34195 45407
rect 47961 45305 47995 45339
rect 32321 45237 32355 45271
rect 33517 45237 33551 45271
rect 22937 45033 22971 45067
rect 25053 45033 25087 45067
rect 35357 44897 35391 44931
rect 35541 44897 35575 44931
rect 48789 44897 48823 44931
rect 23121 44829 23155 44863
rect 25237 44829 25271 44863
rect 48513 44829 48547 44863
rect 35265 44761 35299 44795
rect 34897 44693 34931 44727
rect 14381 44489 14415 44523
rect 36553 44489 36587 44523
rect 36645 44489 36679 44523
rect 39221 44489 39255 44523
rect 14289 44353 14323 44387
rect 39129 44353 39163 44387
rect 49341 44353 49375 44387
rect 36829 44285 36863 44319
rect 39313 44285 39347 44319
rect 36185 44149 36219 44183
rect 38761 44149 38795 44183
rect 49157 44149 49191 44183
rect 13553 43945 13587 43979
rect 16221 43945 16255 43979
rect 16957 43945 16991 43979
rect 20453 43945 20487 43979
rect 21281 43945 21315 43979
rect 22293 43945 22327 43979
rect 28457 43945 28491 43979
rect 12449 43877 12483 43911
rect 22937 43877 22971 43911
rect 28917 43809 28951 43843
rect 29009 43809 29043 43843
rect 30389 43809 30423 43843
rect 34069 43809 34103 43843
rect 37933 43809 37967 43843
rect 1777 43741 1811 43775
rect 12265 43741 12299 43775
rect 22477 43741 22511 43775
rect 30113 43741 30147 43775
rect 32321 43741 32355 43775
rect 37749 43741 37783 43775
rect 48513 43741 48547 43775
rect 48789 43741 48823 43775
rect 13461 43673 13495 43707
rect 16129 43673 16163 43707
rect 16865 43673 16899 43707
rect 20361 43673 20395 43707
rect 21189 43673 21223 43707
rect 22201 43673 22235 43707
rect 22753 43673 22787 43707
rect 28825 43673 28859 43707
rect 32597 43673 32631 43707
rect 37657 43673 37691 43707
rect 1593 43605 1627 43639
rect 31861 43605 31895 43639
rect 37289 43605 37323 43639
rect 2053 43401 2087 43435
rect 12173 43401 12207 43435
rect 16865 43401 16899 43435
rect 19165 43401 19199 43435
rect 20361 43401 20395 43435
rect 20913 43401 20947 43435
rect 25881 43401 25915 43435
rect 40325 43401 40359 43435
rect 34805 43333 34839 43367
rect 2237 43265 2271 43299
rect 12081 43265 12115 43299
rect 17049 43265 17083 43299
rect 19073 43265 19107 43299
rect 20269 43265 20303 43299
rect 21097 43265 21131 43299
rect 26249 43265 26283 43299
rect 32321 43265 32355 43299
rect 34529 43265 34563 43299
rect 40233 43265 40267 43299
rect 48789 43265 48823 43299
rect 26341 43197 26375 43231
rect 26525 43197 26559 43231
rect 28825 43197 28859 43231
rect 29101 43197 29135 43231
rect 32597 43197 32631 43231
rect 40509 43197 40543 43231
rect 48513 43197 48547 43231
rect 30573 43061 30607 43095
rect 34069 43061 34103 43095
rect 36277 43061 36311 43095
rect 39865 43061 39899 43095
rect 27353 42857 27387 42891
rect 35909 42721 35943 42755
rect 40601 42721 40635 42755
rect 25605 42653 25639 42687
rect 35633 42653 35667 42687
rect 40509 42653 40543 42687
rect 48513 42653 48547 42687
rect 48789 42653 48823 42687
rect 25881 42585 25915 42619
rect 37381 42517 37415 42551
rect 40049 42517 40083 42551
rect 40417 42517 40451 42551
rect 7297 42313 7331 42347
rect 9229 42313 9263 42347
rect 17325 42313 17359 42347
rect 20637 42313 20671 42347
rect 22201 42313 22235 42347
rect 25881 42313 25915 42347
rect 40049 42313 40083 42347
rect 41613 42313 41647 42347
rect 8125 42245 8159 42279
rect 24409 42245 24443 42279
rect 27997 42245 28031 42279
rect 30297 42245 30331 42279
rect 7205 42177 7239 42211
rect 7941 42177 7975 42211
rect 9137 42177 9171 42211
rect 17233 42177 17267 42211
rect 20821 42177 20855 42211
rect 22385 42177 22419 42211
rect 33885 42177 33919 42211
rect 41521 42177 41555 42211
rect 48789 42177 48823 42211
rect 24133 42109 24167 42143
rect 27721 42109 27755 42143
rect 30021 42109 30055 42143
rect 34161 42109 34195 42143
rect 38301 42109 38335 42143
rect 38577 42109 38611 42143
rect 41797 42109 41831 42143
rect 48513 42109 48547 42143
rect 29469 41973 29503 42007
rect 31769 41973 31803 42007
rect 35633 41973 35667 42007
rect 41153 41973 41187 42007
rect 21281 41769 21315 41803
rect 22004 41769 22038 41803
rect 26985 41769 27019 41803
rect 36645 41769 36679 41803
rect 38853 41769 38887 41803
rect 48605 41769 48639 41803
rect 21741 41633 21775 41667
rect 27537 41633 27571 41667
rect 34897 41633 34931 41667
rect 37105 41633 37139 41667
rect 23765 41565 23799 41599
rect 31401 41565 31435 41599
rect 48789 41565 48823 41599
rect 1685 41497 1719 41531
rect 27445 41497 27479 41531
rect 31677 41497 31711 41531
rect 35173 41497 35207 41531
rect 37381 41497 37415 41531
rect 1777 41429 1811 41463
rect 27353 41429 27387 41463
rect 33149 41429 33183 41463
rect 5825 41225 5859 41259
rect 9873 41225 9907 41259
rect 10793 41225 10827 41259
rect 22017 41225 22051 41259
rect 29469 41225 29503 41259
rect 29837 41157 29871 41191
rect 33425 41157 33459 41191
rect 5733 41089 5767 41123
rect 9781 41089 9815 41123
rect 10701 41089 10735 41123
rect 21281 41089 21315 41123
rect 22385 41089 22419 41123
rect 24777 41089 24811 41123
rect 27261 41089 27295 41123
rect 29929 41089 29963 41123
rect 38209 41089 38243 41123
rect 48789 41089 48823 41123
rect 22477 41021 22511 41055
rect 22661 41021 22695 41055
rect 25053 41021 25087 41055
rect 26525 41021 26559 41055
rect 27537 41021 27571 41055
rect 30021 41021 30055 41055
rect 33149 41021 33183 41055
rect 48513 41021 48547 41055
rect 23213 40885 23247 40919
rect 29009 40885 29043 40919
rect 34897 40885 34931 40919
rect 38472 40885 38506 40919
rect 39957 40885 39991 40919
rect 23305 40681 23339 40715
rect 35265 40681 35299 40715
rect 38761 40681 38795 40715
rect 25513 40613 25547 40647
rect 23949 40545 23983 40579
rect 25973 40545 26007 40579
rect 26157 40545 26191 40579
rect 27261 40545 27295 40579
rect 30021 40545 30055 40579
rect 32689 40545 32723 40579
rect 32781 40545 32815 40579
rect 34069 40545 34103 40579
rect 34161 40545 34195 40579
rect 35817 40545 35851 40579
rect 39221 40545 39255 40579
rect 39405 40545 39439 40579
rect 48789 40545 48823 40579
rect 27077 40477 27111 40511
rect 29745 40477 29779 40511
rect 32597 40477 32631 40511
rect 35725 40477 35759 40511
rect 48513 40477 48547 40511
rect 25881 40409 25915 40443
rect 33977 40409 34011 40443
rect 35633 40409 35667 40443
rect 23673 40341 23707 40375
rect 23765 40341 23799 40375
rect 26709 40341 26743 40375
rect 27169 40341 27203 40375
rect 31493 40341 31527 40375
rect 32229 40341 32263 40375
rect 33609 40341 33643 40375
rect 39129 40341 39163 40375
rect 25053 40137 25087 40171
rect 36461 40137 36495 40171
rect 40325 40137 40359 40171
rect 40785 40137 40819 40171
rect 41153 40069 41187 40103
rect 32321 40001 32355 40035
rect 34713 40001 34747 40035
rect 38577 40001 38611 40035
rect 41245 40001 41279 40035
rect 23305 39933 23339 39967
rect 23581 39933 23615 39967
rect 28181 39933 28215 39967
rect 28457 39933 28491 39967
rect 32597 39933 32631 39967
rect 34069 39933 34103 39967
rect 34989 39933 35023 39967
rect 38853 39933 38887 39967
rect 41429 39933 41463 39967
rect 48513 39933 48547 39967
rect 48789 39933 48823 39967
rect 29929 39797 29963 39831
rect 22017 39593 22051 39627
rect 30462 39593 30496 39627
rect 32597 39593 32631 39627
rect 42625 39593 42659 39627
rect 22477 39457 22511 39491
rect 22569 39457 22603 39491
rect 24593 39457 24627 39491
rect 24869 39457 24903 39491
rect 31953 39457 31987 39491
rect 33149 39457 33183 39491
rect 36277 39457 36311 39491
rect 41153 39457 41187 39491
rect 48789 39457 48823 39491
rect 30205 39389 30239 39423
rect 36001 39389 36035 39423
rect 38485 39389 38519 39423
rect 40877 39389 40911 39423
rect 48513 39389 48547 39423
rect 32965 39321 32999 39355
rect 21465 39253 21499 39287
rect 22385 39253 22419 39287
rect 26341 39253 26375 39287
rect 33057 39253 33091 39287
rect 37749 39253 37783 39287
rect 24501 39049 24535 39083
rect 25881 39049 25915 39083
rect 26341 39049 26375 39083
rect 27353 39049 27387 39083
rect 28917 39049 28951 39083
rect 32413 39049 32447 39083
rect 33609 39049 33643 39083
rect 33977 39049 34011 39083
rect 34805 39049 34839 39083
rect 35449 39049 35483 39083
rect 36645 39049 36679 39083
rect 37933 39049 37967 39083
rect 38853 39049 38887 39083
rect 39313 39049 39347 39083
rect 23305 38981 23339 39015
rect 24869 38981 24903 39015
rect 24961 38981 24995 39015
rect 27813 38981 27847 39015
rect 31585 38981 31619 39015
rect 32781 38981 32815 39015
rect 1777 38913 1811 38947
rect 22385 38913 22419 38947
rect 23213 38913 23247 38947
rect 26249 38913 26283 38947
rect 27721 38913 27755 38947
rect 35357 38913 35391 38947
rect 36553 38913 36587 38947
rect 37841 38913 37875 38947
rect 39681 38913 39715 38947
rect 40325 38913 40359 38947
rect 23489 38845 23523 38879
rect 25053 38845 25087 38879
rect 26525 38845 26559 38879
rect 27905 38845 27939 38879
rect 29009 38845 29043 38879
rect 29101 38845 29135 38879
rect 31033 38845 31067 38879
rect 32873 38845 32907 38879
rect 32965 38845 32999 38879
rect 34069 38845 34103 38879
rect 34253 38845 34287 38879
rect 35541 38845 35575 38879
rect 36737 38845 36771 38879
rect 38025 38845 38059 38879
rect 38945 38845 38979 38879
rect 39129 38845 39163 38879
rect 39773 38845 39807 38879
rect 39865 38845 39899 38879
rect 40601 38845 40635 38879
rect 1593 38709 1627 38743
rect 22845 38709 22879 38743
rect 28549 38709 28583 38743
rect 34989 38709 35023 38743
rect 36185 38709 36219 38743
rect 37473 38709 37507 38743
rect 38485 38709 38519 38743
rect 42073 38709 42107 38743
rect 23305 38505 23339 38539
rect 27077 38505 27111 38539
rect 32873 38505 32907 38539
rect 36645 38505 36679 38539
rect 40049 38505 40083 38539
rect 43269 38505 43303 38539
rect 22845 38437 22879 38471
rect 28457 38437 28491 38471
rect 21097 38369 21131 38403
rect 23857 38369 23891 38403
rect 27629 38369 27663 38403
rect 28917 38369 28951 38403
rect 29009 38369 29043 38403
rect 29745 38369 29779 38403
rect 33333 38369 33367 38403
rect 33425 38369 33459 38403
rect 34897 38369 34931 38403
rect 39221 38369 39255 38403
rect 40601 38369 40635 38403
rect 31861 38301 31895 38335
rect 40509 38301 40543 38335
rect 41245 38301 41279 38335
rect 41521 38301 41555 38335
rect 49341 38301 49375 38335
rect 21373 38233 21407 38267
rect 26617 38233 26651 38267
rect 27445 38233 27479 38267
rect 30021 38233 30055 38267
rect 31769 38233 31803 38267
rect 32597 38233 32631 38267
rect 35173 38233 35207 38267
rect 37105 38233 37139 38267
rect 37933 38233 37967 38267
rect 41797 38233 41831 38267
rect 23673 38165 23707 38199
rect 23765 38165 23799 38199
rect 27537 38165 27571 38199
rect 28825 38165 28859 38199
rect 33241 38165 33275 38199
rect 40417 38165 40451 38199
rect 49157 38165 49191 38199
rect 33977 37961 34011 37995
rect 37473 37961 37507 37995
rect 41245 37961 41279 37995
rect 43085 37961 43119 37995
rect 31309 37893 31343 37927
rect 36001 37893 36035 37927
rect 41337 37893 41371 37927
rect 23121 37825 23155 37859
rect 27169 37825 27203 37859
rect 30481 37825 30515 37859
rect 32689 37825 32723 37859
rect 33885 37825 33919 37859
rect 36737 37825 36771 37859
rect 37841 37825 37875 37859
rect 42993 37825 43027 37859
rect 49341 37825 49375 37859
rect 23397 37757 23431 37791
rect 27445 37757 27479 37791
rect 29193 37757 29227 37791
rect 32781 37757 32815 37791
rect 32965 37757 32999 37791
rect 34069 37757 34103 37791
rect 37933 37757 37967 37791
rect 38117 37757 38151 37791
rect 38669 37757 38703 37791
rect 38945 37757 38979 37791
rect 41429 37757 41463 37791
rect 43177 37757 43211 37791
rect 40877 37689 40911 37723
rect 49157 37689 49191 37723
rect 22661 37621 22695 37655
rect 24869 37621 24903 37655
rect 30021 37621 30055 37655
rect 32321 37621 32355 37655
rect 33517 37621 33551 37655
rect 40417 37621 40451 37655
rect 42625 37621 42659 37655
rect 22109 37417 22143 37451
rect 25513 37417 25547 37451
rect 28549 37417 28583 37451
rect 29745 37349 29779 37383
rect 22753 37281 22787 37315
rect 23765 37281 23799 37315
rect 23857 37281 23891 37315
rect 26065 37281 26099 37315
rect 26801 37281 26835 37315
rect 30297 37281 30331 37315
rect 31493 37281 31527 37315
rect 32689 37281 32723 37315
rect 33977 37281 34011 37315
rect 39221 37281 39255 37315
rect 40601 37281 40635 37315
rect 41429 37281 41463 37315
rect 42165 37281 42199 37315
rect 48053 37281 48087 37315
rect 48513 37281 48547 37315
rect 22477 37213 22511 37247
rect 22569 37213 22603 37247
rect 23673 37213 23707 37247
rect 24777 37213 24811 37247
rect 29193 37213 29227 37247
rect 30113 37213 30147 37247
rect 31309 37213 31343 37247
rect 32597 37213 32631 37247
rect 38945 37213 38979 37247
rect 40509 37213 40543 37247
rect 48789 37213 48823 37247
rect 27077 37145 27111 37179
rect 31401 37145 31435 37179
rect 33885 37145 33919 37179
rect 40417 37145 40451 37179
rect 42441 37145 42475 37179
rect 23305 37077 23339 37111
rect 25881 37077 25915 37111
rect 25973 37077 26007 37111
rect 30205 37077 30239 37111
rect 30941 37077 30975 37111
rect 32137 37077 32171 37111
rect 32505 37077 32539 37111
rect 33425 37077 33459 37111
rect 33793 37077 33827 37111
rect 38577 37077 38611 37111
rect 39037 37077 39071 37111
rect 40049 37077 40083 37111
rect 43913 37077 43947 37111
rect 19441 36873 19475 36907
rect 27629 36873 27663 36907
rect 32321 36873 32355 36907
rect 32781 36873 32815 36907
rect 37841 36873 37875 36907
rect 41429 36873 41463 36907
rect 43085 36873 43119 36907
rect 26341 36805 26375 36839
rect 30389 36805 30423 36839
rect 1777 36737 1811 36771
rect 19809 36737 19843 36771
rect 19901 36737 19935 36771
rect 26249 36737 26283 36771
rect 27537 36737 27571 36771
rect 30297 36737 30331 36771
rect 31769 36737 31803 36771
rect 32689 36737 32723 36771
rect 42993 36737 43027 36771
rect 49341 36737 49375 36771
rect 20085 36669 20119 36703
rect 23397 36669 23431 36703
rect 23673 36669 23707 36703
rect 25421 36669 25455 36703
rect 26433 36669 26467 36703
rect 27721 36669 27755 36703
rect 30573 36669 30607 36703
rect 32965 36669 32999 36703
rect 34345 36669 34379 36703
rect 34621 36669 34655 36703
rect 37933 36669 37967 36703
rect 38117 36669 38151 36703
rect 39681 36669 39715 36703
rect 39957 36669 39991 36703
rect 43269 36669 43303 36703
rect 37473 36601 37507 36635
rect 1593 36533 1627 36567
rect 22937 36533 22971 36567
rect 25881 36533 25915 36567
rect 27169 36533 27203 36567
rect 29929 36533 29963 36567
rect 36093 36533 36127 36567
rect 42625 36533 42659 36567
rect 49157 36533 49191 36567
rect 21925 36329 21959 36363
rect 22477 36329 22511 36363
rect 27353 36329 27387 36363
rect 32045 36329 32079 36363
rect 37473 36329 37507 36363
rect 40141 36329 40175 36363
rect 36277 36261 36311 36295
rect 23029 36193 23063 36227
rect 28457 36193 28491 36227
rect 32689 36193 32723 36227
rect 35541 36193 35575 36227
rect 35633 36193 35667 36227
rect 36737 36193 36771 36227
rect 36829 36193 36863 36227
rect 38025 36193 38059 36227
rect 40785 36193 40819 36227
rect 41797 36193 41831 36227
rect 41889 36193 41923 36227
rect 43177 36193 43211 36227
rect 22845 36125 22879 36159
rect 28181 36125 28215 36159
rect 28273 36125 28307 36159
rect 32413 36125 32447 36159
rect 42993 36125 43027 36159
rect 35449 36057 35483 36091
rect 36645 36057 36679 36091
rect 37841 36057 37875 36091
rect 40509 36057 40543 36091
rect 41705 36057 41739 36091
rect 22937 35989 22971 36023
rect 27813 35989 27847 36023
rect 32505 35989 32539 36023
rect 35081 35989 35115 36023
rect 37933 35989 37967 36023
rect 40601 35989 40635 36023
rect 41337 35989 41371 36023
rect 42533 35989 42567 36023
rect 42901 35989 42935 36023
rect 21281 35785 21315 35819
rect 23765 35785 23799 35819
rect 30849 35785 30883 35819
rect 32321 35785 32355 35819
rect 35633 35785 35667 35819
rect 36093 35785 36127 35819
rect 39957 35785 39991 35819
rect 24961 35717 24995 35751
rect 40785 35717 40819 35751
rect 42901 35717 42935 35751
rect 19533 35649 19567 35683
rect 24685 35649 24719 35683
rect 29101 35649 29135 35683
rect 31769 35649 31803 35683
rect 32689 35649 32723 35683
rect 34805 35649 34839 35683
rect 34897 35649 34931 35683
rect 36001 35649 36035 35683
rect 38209 35649 38243 35683
rect 40877 35649 40911 35683
rect 42625 35649 42659 35683
rect 49341 35649 49375 35683
rect 19809 35581 19843 35615
rect 22017 35581 22051 35615
rect 22293 35581 22327 35615
rect 26433 35581 26467 35615
rect 29377 35581 29411 35615
rect 32781 35581 32815 35615
rect 32873 35581 32907 35615
rect 35081 35581 35115 35615
rect 36185 35581 36219 35615
rect 40969 35581 41003 35615
rect 33517 35513 33551 35547
rect 34437 35513 34471 35547
rect 49157 35513 49191 35547
rect 27353 35445 27387 35479
rect 38466 35445 38500 35479
rect 40417 35445 40451 35479
rect 44373 35445 44407 35479
rect 24593 35241 24627 35275
rect 26065 35241 26099 35275
rect 29009 35241 29043 35275
rect 33977 35241 34011 35275
rect 23489 35173 23523 35207
rect 21741 35105 21775 35139
rect 25145 35105 25179 35139
rect 26709 35105 26743 35139
rect 27261 35105 27295 35139
rect 27537 35105 27571 35139
rect 31493 35105 31527 35139
rect 31677 35105 31711 35139
rect 32229 35105 32263 35139
rect 32505 35105 32539 35139
rect 36645 35105 36679 35139
rect 37841 35105 37875 35139
rect 37933 35105 37967 35139
rect 39221 35105 39255 35139
rect 42073 35105 42107 35139
rect 42717 35105 42751 35139
rect 42993 35105 43027 35139
rect 44465 35105 44499 35139
rect 25053 35037 25087 35071
rect 26433 35037 26467 35071
rect 36461 35037 36495 35071
rect 37749 35037 37783 35071
rect 49341 35037 49375 35071
rect 22017 34969 22051 35003
rect 24961 34969 24995 35003
rect 30573 34969 30607 35003
rect 31401 34969 31435 35003
rect 38945 34969 38979 35003
rect 41889 34969 41923 35003
rect 26525 34901 26559 34935
rect 31033 34901 31067 34935
rect 36001 34901 36035 34935
rect 36369 34901 36403 34935
rect 37381 34901 37415 34935
rect 38577 34901 38611 34935
rect 39037 34901 39071 34935
rect 41429 34901 41463 34935
rect 41797 34901 41831 34935
rect 49157 34901 49191 34935
rect 1593 34697 1627 34731
rect 25421 34697 25455 34731
rect 30113 34697 30147 34731
rect 30481 34697 30515 34731
rect 31401 34697 31435 34731
rect 32321 34697 32355 34731
rect 35817 34697 35851 34731
rect 39037 34697 39071 34731
rect 39497 34697 39531 34731
rect 43361 34697 43395 34731
rect 31493 34629 31527 34663
rect 43453 34629 43487 34663
rect 1777 34561 1811 34595
rect 25789 34561 25823 34595
rect 28273 34561 28307 34595
rect 32689 34561 32723 34595
rect 32781 34561 32815 34595
rect 33517 34561 33551 34595
rect 39405 34561 39439 34595
rect 40601 34561 40635 34595
rect 40693 34561 40727 34595
rect 41981 34561 42015 34595
rect 49341 34561 49375 34595
rect 23121 34493 23155 34527
rect 23397 34493 23431 34527
rect 24869 34493 24903 34527
rect 25881 34493 25915 34527
rect 26065 34493 26099 34527
rect 28549 34493 28583 34527
rect 30021 34493 30055 34527
rect 30573 34493 30607 34527
rect 30665 34493 30699 34527
rect 31585 34493 31619 34527
rect 32965 34493 32999 34527
rect 34069 34493 34103 34527
rect 39681 34493 39715 34527
rect 40785 34493 40819 34527
rect 43545 34493 43579 34527
rect 31033 34425 31067 34459
rect 42993 34425 43027 34459
rect 49157 34425 49191 34459
rect 34332 34357 34366 34391
rect 40233 34357 40267 34391
rect 23305 34153 23339 34187
rect 32505 34153 32539 34187
rect 36829 34153 36863 34187
rect 22845 34085 22879 34119
rect 24593 34085 24627 34119
rect 30757 34085 30791 34119
rect 38301 34085 38335 34119
rect 21097 34017 21131 34051
rect 23949 34017 23983 34051
rect 25237 34017 25271 34051
rect 26249 34017 26283 34051
rect 31401 34017 31435 34051
rect 36185 34017 36219 34051
rect 37749 34017 37783 34051
rect 38761 34017 38795 34051
rect 38945 34017 38979 34051
rect 42349 34017 42383 34051
rect 29929 33949 29963 33983
rect 42165 33949 42199 33983
rect 49341 33949 49375 33983
rect 21373 33881 21407 33915
rect 24961 33881 24995 33915
rect 26525 33881 26559 33915
rect 36461 33881 36495 33915
rect 23673 33813 23707 33847
rect 23765 33813 23799 33847
rect 25053 33813 25087 33847
rect 27997 33813 28031 33847
rect 31125 33813 31159 33847
rect 31217 33813 31251 33847
rect 35541 33813 35575 33847
rect 36369 33813 36403 33847
rect 38669 33813 38703 33847
rect 41797 33813 41831 33847
rect 42257 33813 42291 33847
rect 49157 33813 49191 33847
rect 23673 33609 23707 33643
rect 28733 33609 28767 33643
rect 29101 33609 29135 33643
rect 37473 33609 37507 33643
rect 34253 33541 34287 33575
rect 37933 33541 37967 33575
rect 39221 33541 39255 33575
rect 24041 33473 24075 33507
rect 24133 33473 24167 33507
rect 30297 33473 30331 33507
rect 31309 33473 31343 33507
rect 33977 33473 34011 33507
rect 37841 33473 37875 33507
rect 38761 33473 38795 33507
rect 24225 33405 24259 33439
rect 29193 33405 29227 33439
rect 29377 33405 29411 33439
rect 30389 33405 30423 33439
rect 30481 33405 30515 33439
rect 38117 33405 38151 33439
rect 39313 33405 39347 33439
rect 39405 33405 39439 33439
rect 40325 33405 40359 33439
rect 40601 33405 40635 33439
rect 36185 33337 36219 33371
rect 29929 33269 29963 33303
rect 35725 33269 35759 33303
rect 38853 33269 38887 33303
rect 42073 33269 42107 33303
rect 28457 33065 28491 33099
rect 37657 33065 37691 33099
rect 29745 32997 29779 33031
rect 34897 32997 34931 33031
rect 38393 32997 38427 33031
rect 22569 32929 22603 32963
rect 24041 32929 24075 32963
rect 27077 32929 27111 32963
rect 27261 32929 27295 32963
rect 29009 32929 29043 32963
rect 30205 32929 30239 32963
rect 30297 32929 30331 32963
rect 31401 32929 31435 32963
rect 31493 32929 31527 32963
rect 35541 32929 35575 32963
rect 38853 32929 38887 32963
rect 38945 32929 38979 32963
rect 40969 32929 41003 32963
rect 42073 32929 42107 32963
rect 42257 32929 42291 32963
rect 22293 32861 22327 32895
rect 28825 32861 28859 32895
rect 34529 32861 34563 32895
rect 35265 32861 35299 32895
rect 35909 32861 35943 32895
rect 40785 32861 40819 32895
rect 41981 32861 42015 32895
rect 43821 32861 43855 32895
rect 49341 32861 49375 32895
rect 26065 32793 26099 32827
rect 26985 32793 27019 32827
rect 28917 32793 28951 32827
rect 36185 32793 36219 32827
rect 26617 32725 26651 32759
rect 30113 32725 30147 32759
rect 30941 32725 30975 32759
rect 31309 32725 31343 32759
rect 35357 32725 35391 32759
rect 38761 32725 38795 32759
rect 40417 32725 40451 32759
rect 40877 32725 40911 32759
rect 41613 32725 41647 32759
rect 43637 32725 43671 32759
rect 49157 32725 49191 32759
rect 17233 32521 17267 32555
rect 25697 32521 25731 32555
rect 27261 32521 27295 32555
rect 35081 32521 35115 32555
rect 27721 32453 27755 32487
rect 28457 32453 28491 32487
rect 35173 32453 35207 32487
rect 1777 32385 1811 32419
rect 17601 32385 17635 32419
rect 18797 32385 18831 32419
rect 27629 32385 27663 32419
rect 44833 32385 44867 32419
rect 48789 32385 48823 32419
rect 17693 32317 17727 32351
rect 17877 32317 17911 32351
rect 23949 32317 23983 32351
rect 24225 32317 24259 32351
rect 27905 32317 27939 32351
rect 28825 32317 28859 32351
rect 32505 32317 32539 32351
rect 32781 32317 32815 32351
rect 35265 32317 35299 32351
rect 39497 32317 39531 32351
rect 39773 32317 39807 32351
rect 48513 32317 48547 32351
rect 34253 32249 34287 32283
rect 1593 32181 1627 32215
rect 18521 32181 18555 32215
rect 34713 32181 34747 32215
rect 41245 32181 41279 32215
rect 42809 32181 42843 32215
rect 44649 32181 44683 32215
rect 24041 31977 24075 32011
rect 28457 31977 28491 32011
rect 39313 31977 39347 32011
rect 43637 31977 43671 32011
rect 32321 31909 32355 31943
rect 35357 31909 35391 31943
rect 37933 31909 37967 31943
rect 22293 31841 22327 31875
rect 22569 31841 22603 31875
rect 25789 31841 25823 31875
rect 26065 31841 26099 31875
rect 27813 31841 27847 31875
rect 29009 31841 29043 31875
rect 32781 31841 32815 31875
rect 32965 31841 32999 31875
rect 35817 31841 35851 31875
rect 36001 31841 36035 31875
rect 38485 31841 38519 31875
rect 41889 31841 41923 31875
rect 42165 31841 42199 31875
rect 48789 31841 48823 31875
rect 21833 31773 21867 31807
rect 24777 31773 24811 31807
rect 28917 31773 28951 31807
rect 38301 31773 38335 31807
rect 38393 31773 38427 31807
rect 39497 31773 39531 31807
rect 48053 31773 48087 31807
rect 48513 31773 48547 31807
rect 35725 31705 35759 31739
rect 28825 31637 28859 31671
rect 31861 31637 31895 31671
rect 32689 31637 32723 31671
rect 23489 31433 23523 31467
rect 23857 31433 23891 31467
rect 26617 31433 26651 31467
rect 36185 31433 36219 31467
rect 38577 31433 38611 31467
rect 42993 31433 43027 31467
rect 43085 31365 43119 31399
rect 21465 31297 21499 31331
rect 22385 31297 22419 31331
rect 24869 31297 24903 31331
rect 33333 31297 33367 31331
rect 33425 31297 33459 31331
rect 37749 31297 37783 31331
rect 40785 31297 40819 31331
rect 45569 31297 45603 31331
rect 48789 31297 48823 31331
rect 22477 31229 22511 31263
rect 22661 31229 22695 31263
rect 23949 31229 23983 31263
rect 24133 31229 24167 31263
rect 25145 31229 25179 31263
rect 33517 31229 33551 31263
rect 34437 31229 34471 31263
rect 34713 31229 34747 31263
rect 38669 31229 38703 31263
rect 38761 31229 38795 31263
rect 43177 31229 43211 31263
rect 48513 31229 48547 31263
rect 37565 31161 37599 31195
rect 40601 31161 40635 31195
rect 22017 31093 22051 31127
rect 32965 31093 32999 31127
rect 38209 31093 38243 31127
rect 42625 31093 42659 31127
rect 45385 31093 45419 31127
rect 21465 30889 21499 30923
rect 23213 30889 23247 30923
rect 29745 30889 29779 30923
rect 36185 30889 36219 30923
rect 37381 30889 37415 30923
rect 26617 30821 26651 30855
rect 33057 30821 33091 30855
rect 22109 30753 22143 30787
rect 23857 30753 23891 30787
rect 27077 30753 27111 30787
rect 30297 30753 30331 30787
rect 35633 30753 35667 30787
rect 36737 30753 36771 30787
rect 37841 30753 37875 30787
rect 37933 30753 37967 30787
rect 39221 30753 39255 30787
rect 40509 30753 40543 30787
rect 40601 30753 40635 30787
rect 21833 30685 21867 30719
rect 24869 30685 24903 30719
rect 31309 30685 31343 30719
rect 35357 30685 35391 30719
rect 39129 30685 39163 30719
rect 40417 30685 40451 30719
rect 41521 30685 41555 30719
rect 42165 30685 42199 30719
rect 43177 30685 43211 30719
rect 20913 30617 20947 30651
rect 21925 30617 21959 30651
rect 23673 30617 23707 30651
rect 25145 30617 25179 30651
rect 27353 30617 27387 30651
rect 30113 30617 30147 30651
rect 31585 30617 31619 30651
rect 36645 30617 36679 30651
rect 39037 30617 39071 30651
rect 23581 30549 23615 30583
rect 28825 30549 28859 30583
rect 30205 30549 30239 30583
rect 34989 30549 35023 30583
rect 35449 30549 35483 30583
rect 36553 30549 36587 30583
rect 37749 30549 37783 30583
rect 38669 30549 38703 30583
rect 40049 30549 40083 30583
rect 41337 30549 41371 30583
rect 41981 30549 42015 30583
rect 42993 30549 43027 30583
rect 23857 30345 23891 30379
rect 24869 30345 24903 30379
rect 28733 30345 28767 30379
rect 24777 30277 24811 30311
rect 25605 30277 25639 30311
rect 30757 30277 30791 30311
rect 34161 30277 34195 30311
rect 35909 30277 35943 30311
rect 36001 30277 36035 30311
rect 37841 30277 37875 30311
rect 37933 30277 37967 30311
rect 41337 30277 41371 30311
rect 7389 30209 7423 30243
rect 24225 30209 24259 30243
rect 34069 30209 34103 30243
rect 41245 30209 41279 30243
rect 49341 30209 49375 30243
rect 7573 30141 7607 30175
rect 9137 30141 9171 30175
rect 25053 30141 25087 30175
rect 28825 30141 28859 30175
rect 28917 30141 28951 30175
rect 30849 30141 30883 30175
rect 31033 30141 31067 30175
rect 34345 30141 34379 30175
rect 36093 30141 36127 30175
rect 38025 30141 38059 30175
rect 38669 30141 38703 30175
rect 38945 30141 38979 30175
rect 41429 30141 41463 30175
rect 24409 30073 24443 30107
rect 27813 30073 27847 30107
rect 33701 30073 33735 30107
rect 40877 30073 40911 30107
rect 49157 30073 49191 30107
rect 28365 30005 28399 30039
rect 30389 30005 30423 30039
rect 35541 30005 35575 30039
rect 37473 30005 37507 30039
rect 40417 30005 40451 30039
rect 42717 29801 42751 29835
rect 29745 29733 29779 29767
rect 2053 29665 2087 29699
rect 23213 29665 23247 29699
rect 25789 29665 25823 29699
rect 25973 29665 26007 29699
rect 30205 29665 30239 29699
rect 30297 29665 30331 29699
rect 32505 29665 32539 29699
rect 36369 29665 36403 29699
rect 41245 29665 41279 29699
rect 48789 29665 48823 29699
rect 1777 29597 1811 29631
rect 25697 29597 25731 29631
rect 26709 29597 26743 29631
rect 32321 29597 32355 29631
rect 40969 29597 41003 29631
rect 48513 29597 48547 29631
rect 22477 29529 22511 29563
rect 30113 29529 30147 29563
rect 36645 29529 36679 29563
rect 25329 29461 25363 29495
rect 31953 29461 31987 29495
rect 32413 29461 32447 29495
rect 38117 29461 38151 29495
rect 21189 29257 21223 29291
rect 22017 29257 22051 29291
rect 35725 29257 35759 29291
rect 39313 29257 39347 29291
rect 39681 29257 39715 29291
rect 39773 29257 39807 29291
rect 41245 29257 41279 29291
rect 49157 29257 49191 29291
rect 22477 29189 22511 29223
rect 27997 29189 28031 29223
rect 22385 29121 22419 29155
rect 23305 29121 23339 29155
rect 27721 29121 27755 29155
rect 30297 29121 30331 29155
rect 41153 29121 41187 29155
rect 49341 29121 49375 29155
rect 22661 29053 22695 29087
rect 29469 29053 29503 29087
rect 30389 29053 30423 29087
rect 30481 29053 30515 29087
rect 33977 29053 34011 29087
rect 39865 29053 39899 29087
rect 41429 29053 41463 29087
rect 29929 28985 29963 29019
rect 40785 28985 40819 29019
rect 34240 28917 34274 28951
rect 36369 28917 36403 28951
rect 38669 28917 38703 28951
rect 22937 28713 22971 28747
rect 38669 28713 38703 28747
rect 28365 28645 28399 28679
rect 23489 28577 23523 28611
rect 31217 28577 31251 28611
rect 34069 28577 34103 28611
rect 34161 28577 34195 28611
rect 35541 28577 35575 28611
rect 36645 28577 36679 28611
rect 37381 28577 37415 28611
rect 37565 28577 37599 28611
rect 39313 28577 39347 28611
rect 40509 28577 40543 28611
rect 40693 28577 40727 28611
rect 21005 28509 21039 28543
rect 29929 28509 29963 28543
rect 31033 28509 31067 28543
rect 33977 28509 34011 28543
rect 36461 28509 36495 28543
rect 39037 28509 39071 28543
rect 40417 28509 40451 28543
rect 49341 28509 49375 28543
rect 21741 28441 21775 28475
rect 27077 28441 27111 28475
rect 38117 28441 38151 28475
rect 39129 28441 39163 28475
rect 22385 28373 22419 28407
rect 23305 28373 23339 28407
rect 23397 28373 23431 28407
rect 30665 28373 30699 28407
rect 31125 28373 31159 28407
rect 33609 28373 33643 28407
rect 34897 28373 34931 28407
rect 35265 28373 35299 28407
rect 35357 28373 35391 28407
rect 36093 28373 36127 28407
rect 36553 28373 36587 28407
rect 36921 28373 36955 28407
rect 37289 28373 37323 28407
rect 40049 28373 40083 28407
rect 49157 28373 49191 28407
rect 4905 28169 4939 28203
rect 26341 28169 26375 28203
rect 31309 28169 31343 28203
rect 34069 28169 34103 28203
rect 36369 28169 36403 28203
rect 36461 28169 36495 28203
rect 39037 28169 39071 28203
rect 39497 28169 39531 28203
rect 22661 28101 22695 28135
rect 28181 28101 28215 28135
rect 38393 28101 38427 28135
rect 5089 28033 5123 28067
rect 7573 28033 7607 28067
rect 22385 28033 22419 28067
rect 31217 28033 31251 28067
rect 32321 28033 32355 28067
rect 37657 28033 37691 28067
rect 39405 28033 39439 28067
rect 48145 28033 48179 28067
rect 7757 27965 7791 27999
rect 9413 27965 9447 27999
rect 24593 27965 24627 27999
rect 24869 27965 24903 27999
rect 27905 27965 27939 27999
rect 31493 27965 31527 27999
rect 32597 27965 32631 27999
rect 36645 27965 36679 27999
rect 39681 27965 39715 27999
rect 24133 27829 24167 27863
rect 29653 27829 29687 27863
rect 30849 27829 30883 27863
rect 36001 27829 36035 27863
rect 48237 27829 48271 27863
rect 7803 27557 7837 27591
rect 27721 27557 27755 27591
rect 38669 27557 38703 27591
rect 41797 27557 41831 27591
rect 2053 27489 2087 27523
rect 28365 27489 28399 27523
rect 30757 27489 30791 27523
rect 32229 27489 32263 27523
rect 35357 27489 35391 27523
rect 35449 27489 35483 27523
rect 40049 27489 40083 27523
rect 1777 27421 1811 27455
rect 7700 27421 7734 27455
rect 23397 27421 23431 27455
rect 24869 27421 24903 27455
rect 28089 27421 28123 27455
rect 30665 27421 30699 27455
rect 32873 27421 32907 27455
rect 33701 27421 33735 27455
rect 36921 27421 36955 27455
rect 44005 27421 44039 27455
rect 47225 27421 47259 27455
rect 48513 27421 48547 27455
rect 48789 27421 48823 27455
rect 25145 27353 25179 27387
rect 32045 27353 32079 27387
rect 35265 27353 35299 27387
rect 37197 27353 37231 27387
rect 40325 27353 40359 27387
rect 47409 27353 47443 27387
rect 26617 27285 26651 27319
rect 28181 27285 28215 27319
rect 30205 27285 30239 27319
rect 30573 27285 30607 27319
rect 31677 27285 31711 27319
rect 32137 27285 32171 27319
rect 34897 27285 34931 27319
rect 43821 27285 43855 27319
rect 23121 27081 23155 27115
rect 23213 27081 23247 27115
rect 30297 27081 30331 27115
rect 35909 27081 35943 27115
rect 42073 27081 42107 27115
rect 27905 27013 27939 27047
rect 31125 27013 31159 27047
rect 33333 27013 33367 27047
rect 40601 27013 40635 27047
rect 47869 27013 47903 27047
rect 7849 26945 7883 26979
rect 24133 26945 24167 26979
rect 27169 26945 27203 26979
rect 28549 26945 28583 26979
rect 33425 26945 33459 26979
rect 36921 26945 36955 26979
rect 37473 26945 37507 26979
rect 40325 26945 40359 26979
rect 47041 26945 47075 26979
rect 8033 26877 8067 26911
rect 8953 26877 8987 26911
rect 23397 26877 23431 26911
rect 28825 26877 28859 26911
rect 31217 26877 31251 26911
rect 31309 26877 31343 26911
rect 33609 26877 33643 26911
rect 34161 26877 34195 26911
rect 34437 26877 34471 26911
rect 38301 26877 38335 26911
rect 48513 26877 48547 26911
rect 48789 26877 48823 26911
rect 22753 26741 22787 26775
rect 24225 26741 24259 26775
rect 30757 26741 30791 26775
rect 32965 26741 32999 26775
rect 36737 26741 36771 26775
rect 46857 26741 46891 26775
rect 47961 26741 47995 26775
rect 7895 26537 7929 26571
rect 9689 26537 9723 26571
rect 22372 26537 22406 26571
rect 33885 26537 33919 26571
rect 37381 26537 37415 26571
rect 23857 26469 23891 26503
rect 24593 26469 24627 26503
rect 9137 26401 9171 26435
rect 22109 26401 22143 26435
rect 25053 26401 25087 26435
rect 25145 26401 25179 26435
rect 26525 26401 26559 26435
rect 26709 26401 26743 26435
rect 31125 26401 31159 26435
rect 31217 26401 31251 26435
rect 37933 26401 37967 26435
rect 40049 26401 40083 26435
rect 41797 26401 41831 26435
rect 48789 26401 48823 26435
rect 7792 26333 7826 26367
rect 9321 26333 9355 26367
rect 24961 26333 24995 26367
rect 27261 26333 27295 26367
rect 32137 26333 32171 26367
rect 34897 26333 34931 26367
rect 37841 26333 37875 26367
rect 47409 26333 47443 26367
rect 48053 26333 48087 26367
rect 48513 26333 48547 26367
rect 28089 26265 28123 26299
rect 31033 26265 31067 26299
rect 32413 26265 32447 26299
rect 35633 26265 35667 26299
rect 40325 26265 40359 26299
rect 26065 26197 26099 26231
rect 26433 26197 26467 26231
rect 30665 26197 30699 26231
rect 37749 26197 37783 26231
rect 47225 26197 47259 26231
rect 27537 25993 27571 26027
rect 31309 25993 31343 26027
rect 31401 25993 31435 26027
rect 32321 25993 32355 26027
rect 32689 25993 32723 26027
rect 39037 25993 39071 26027
rect 39405 25993 39439 26027
rect 42073 25993 42107 26027
rect 32781 25925 32815 25959
rect 40601 25925 40635 25959
rect 46765 25925 46799 25959
rect 7665 25857 7699 25891
rect 24133 25857 24167 25891
rect 25145 25857 25179 25891
rect 26617 25857 26651 25891
rect 27629 25857 27663 25891
rect 35265 25857 35299 25891
rect 36277 25857 36311 25891
rect 38209 25857 38243 25891
rect 39497 25857 39531 25891
rect 40325 25857 40359 25891
rect 46029 25857 46063 25891
rect 49341 25857 49375 25891
rect 7849 25789 7883 25823
rect 9505 25789 9539 25823
rect 24225 25789 24259 25823
rect 24317 25789 24351 25823
rect 27721 25789 27755 25823
rect 28365 25789 28399 25823
rect 28641 25789 28675 25823
rect 31585 25789 31619 25823
rect 32873 25789 32907 25823
rect 35357 25789 35391 25823
rect 35541 25789 35575 25823
rect 38301 25789 38335 25823
rect 38393 25789 38427 25823
rect 39589 25789 39623 25823
rect 23765 25721 23799 25755
rect 36093 25721 36127 25755
rect 46213 25721 46247 25755
rect 46949 25721 46983 25755
rect 22845 25653 22879 25687
rect 25973 25653 26007 25687
rect 27169 25653 27203 25687
rect 30113 25653 30147 25687
rect 30941 25653 30975 25687
rect 34897 25653 34931 25687
rect 36921 25653 36955 25687
rect 37841 25653 37875 25687
rect 49157 25653 49191 25687
rect 4905 25449 4939 25483
rect 10793 25449 10827 25483
rect 11069 25449 11103 25483
rect 27721 25449 27755 25483
rect 39497 25449 39531 25483
rect 14289 25381 14323 25415
rect 30757 25381 30791 25415
rect 2053 25313 2087 25347
rect 22937 25313 22971 25347
rect 25237 25313 25271 25347
rect 25973 25313 26007 25347
rect 28917 25313 28951 25347
rect 31309 25313 31343 25347
rect 32505 25313 32539 25347
rect 33977 25313 34011 25347
rect 34069 25313 34103 25347
rect 35725 25313 35759 25347
rect 37013 25313 37047 25347
rect 37197 25313 37231 25347
rect 38025 25313 38059 25347
rect 40509 25313 40543 25347
rect 40693 25313 40727 25347
rect 1777 25245 1811 25279
rect 5089 25245 5123 25279
rect 10609 25245 10643 25279
rect 14473 25245 14507 25279
rect 22661 25245 22695 25279
rect 24041 25245 24075 25279
rect 24961 25245 24995 25279
rect 28733 25245 28767 25279
rect 28825 25245 28859 25279
rect 29929 25245 29963 25279
rect 31217 25245 31251 25279
rect 32413 25245 32447 25279
rect 33885 25245 33919 25279
rect 37749 25245 37783 25279
rect 45293 25245 45327 25279
rect 46029 25245 46063 25279
rect 22753 25177 22787 25211
rect 26249 25177 26283 25211
rect 32321 25177 32355 25211
rect 35633 25177 35667 25211
rect 36921 25177 36955 25211
rect 44373 25177 44407 25211
rect 45477 25177 45511 25211
rect 46213 25177 46247 25211
rect 22293 25109 22327 25143
rect 24593 25109 24627 25143
rect 25053 25109 25087 25143
rect 28365 25109 28399 25143
rect 31125 25109 31159 25143
rect 31953 25109 31987 25143
rect 33517 25109 33551 25143
rect 35173 25109 35207 25143
rect 35541 25109 35575 25143
rect 36553 25109 36587 25143
rect 40049 25109 40083 25143
rect 40417 25109 40451 25143
rect 44465 25109 44499 25143
rect 25789 24905 25823 24939
rect 28917 24905 28951 24939
rect 32781 24905 32815 24939
rect 37841 24905 37875 24939
rect 29653 24837 29687 24871
rect 34253 24837 34287 24871
rect 8452 24769 8486 24803
rect 27169 24769 27203 24803
rect 32873 24769 32907 24803
rect 33977 24769 34011 24803
rect 37933 24769 37967 24803
rect 40233 24769 40267 24803
rect 47961 24769 47995 24803
rect 8539 24701 8573 24735
rect 19717 24701 19751 24735
rect 19993 24701 20027 24735
rect 25881 24701 25915 24735
rect 26065 24701 26099 24735
rect 27445 24701 27479 24735
rect 29377 24701 29411 24735
rect 31125 24701 31159 24735
rect 32965 24701 32999 24735
rect 36001 24701 36035 24735
rect 38117 24701 38151 24735
rect 49157 24701 49191 24735
rect 21465 24565 21499 24599
rect 25421 24565 25455 24599
rect 32413 24565 32447 24599
rect 37473 24565 37507 24599
rect 10885 24361 10919 24395
rect 16405 24361 16439 24395
rect 27629 24361 27663 24395
rect 29745 24293 29779 24327
rect 14657 24225 14691 24259
rect 20821 24225 20855 24259
rect 25605 24225 25639 24259
rect 26893 24225 26927 24259
rect 27077 24225 27111 24259
rect 28273 24225 28307 24259
rect 30205 24225 30239 24259
rect 30297 24225 30331 24259
rect 34069 24225 34103 24259
rect 34253 24225 34287 24259
rect 37749 24225 37783 24259
rect 40509 24225 40543 24259
rect 40693 24225 40727 24259
rect 10609 24157 10643 24191
rect 25513 24157 25547 24191
rect 26249 24157 26283 24191
rect 27997 24157 28031 24191
rect 33977 24157 34011 24191
rect 34989 24157 35023 24191
rect 37657 24157 37691 24191
rect 40417 24157 40451 24191
rect 47961 24157 47995 24191
rect 14933 24089 14967 24123
rect 21097 24089 21131 24123
rect 35265 24089 35299 24123
rect 49157 24089 49191 24123
rect 11069 24021 11103 24055
rect 22569 24021 22603 24055
rect 25053 24021 25087 24055
rect 25421 24021 25455 24055
rect 26433 24021 26467 24055
rect 26801 24021 26835 24055
rect 28089 24021 28123 24055
rect 30113 24021 30147 24055
rect 33609 24021 33643 24055
rect 36737 24021 36771 24055
rect 37197 24021 37231 24055
rect 37565 24021 37599 24055
rect 40049 24021 40083 24055
rect 9413 23817 9447 23851
rect 19349 23817 19383 23851
rect 19717 23817 19751 23851
rect 20729 23817 20763 23851
rect 21097 23817 21131 23851
rect 26249 23817 26283 23851
rect 22293 23749 22327 23783
rect 34989 23749 35023 23783
rect 39037 23749 39071 23783
rect 8769 23681 8803 23715
rect 12909 23681 12943 23715
rect 22017 23681 22051 23715
rect 25421 23681 25455 23715
rect 28641 23681 28675 23715
rect 28733 23681 28767 23715
rect 34897 23681 34931 23715
rect 38761 23681 38795 23715
rect 47961 23681 47995 23715
rect 8953 23613 8987 23647
rect 13185 23613 13219 23647
rect 14657 23613 14691 23647
rect 19809 23613 19843 23647
rect 19993 23613 20027 23647
rect 21189 23613 21223 23647
rect 21281 23613 21315 23647
rect 24041 23613 24075 23647
rect 26341 23613 26375 23647
rect 26525 23613 26559 23647
rect 28825 23613 28859 23647
rect 32321 23613 32355 23647
rect 35173 23613 35207 23647
rect 49157 23613 49191 23647
rect 34069 23545 34103 23579
rect 24777 23477 24811 23511
rect 25881 23477 25915 23511
rect 28273 23477 28307 23511
rect 32584 23477 32618 23511
rect 34529 23477 34563 23511
rect 40509 23477 40543 23511
rect 5181 23273 5215 23307
rect 22569 23273 22603 23307
rect 28917 23273 28951 23307
rect 31861 23273 31895 23307
rect 34069 23273 34103 23307
rect 36645 23273 36679 23307
rect 37473 23273 37507 23307
rect 2053 23137 2087 23171
rect 9275 23137 9309 23171
rect 17141 23137 17175 23171
rect 19441 23137 19475 23171
rect 23489 23137 23523 23171
rect 23673 23137 23707 23171
rect 25237 23137 25271 23171
rect 27169 23137 27203 23171
rect 30113 23137 30147 23171
rect 30389 23137 30423 23171
rect 32321 23137 32355 23171
rect 34897 23137 34931 23171
rect 38761 23137 38795 23171
rect 1777 23069 1811 23103
rect 4169 23069 4203 23103
rect 9188 23069 9222 23103
rect 23397 23069 23431 23103
rect 24961 23069 24995 23103
rect 37657 23069 37691 23103
rect 38577 23069 38611 23103
rect 40233 23069 40267 23103
rect 44189 23069 44223 23103
rect 47961 23069 47995 23103
rect 5089 23001 5123 23035
rect 17417 23001 17451 23035
rect 19717 23001 19751 23035
rect 27445 23001 27479 23035
rect 32597 23001 32631 23035
rect 35173 23001 35207 23035
rect 38669 23001 38703 23035
rect 44373 23001 44407 23035
rect 49157 23001 49191 23035
rect 4261 22933 4295 22967
rect 18889 22933 18923 22967
rect 21189 22933 21223 22967
rect 23029 22933 23063 22967
rect 24593 22933 24627 22967
rect 25053 22933 25087 22967
rect 38209 22933 38243 22967
rect 17785 22729 17819 22763
rect 19349 22729 19383 22763
rect 19717 22729 19751 22763
rect 23673 22729 23707 22763
rect 30021 22729 30055 22763
rect 30113 22729 30147 22763
rect 31033 22729 31067 22763
rect 34069 22729 34103 22763
rect 21189 22661 21223 22695
rect 23765 22661 23799 22695
rect 27445 22661 27479 22695
rect 31493 22661 31527 22695
rect 34161 22661 34195 22695
rect 37933 22661 37967 22695
rect 21097 22593 21131 22627
rect 24961 22593 24995 22627
rect 25973 22593 26007 22627
rect 31401 22593 31435 22627
rect 32505 22593 32539 22627
rect 37657 22593 37691 22627
rect 17877 22525 17911 22559
rect 17969 22525 18003 22559
rect 19809 22525 19843 22559
rect 19901 22525 19935 22559
rect 21281 22525 21315 22559
rect 23949 22525 23983 22559
rect 25053 22525 25087 22559
rect 25145 22525 25179 22559
rect 27169 22525 27203 22559
rect 28917 22525 28951 22559
rect 30205 22525 30239 22559
rect 31677 22525 31711 22559
rect 34253 22525 34287 22559
rect 39681 22525 39715 22559
rect 20729 22457 20763 22491
rect 29653 22457 29687 22491
rect 17417 22389 17451 22423
rect 23305 22389 23339 22423
rect 24593 22389 24627 22423
rect 33701 22389 33735 22423
rect 12817 22185 12851 22219
rect 15006 22185 15040 22219
rect 16497 22185 16531 22219
rect 19704 22185 19738 22219
rect 23305 22185 23339 22219
rect 35614 22185 35648 22219
rect 5549 22117 5583 22151
rect 14749 22049 14783 22083
rect 19441 22049 19475 22083
rect 21189 22049 21223 22083
rect 22661 22049 22695 22083
rect 23949 22049 23983 22083
rect 25145 22049 25179 22083
rect 26249 22049 26283 22083
rect 28917 22049 28951 22083
rect 29009 22049 29043 22083
rect 37105 22049 37139 22083
rect 12541 21981 12575 22015
rect 13645 21981 13679 22015
rect 25973 21981 26007 22015
rect 26065 21981 26099 22015
rect 29929 21981 29963 22015
rect 35357 21981 35391 22015
rect 37841 21981 37875 22015
rect 47961 21981 47995 22015
rect 49157 21981 49191 22015
rect 5365 21913 5399 21947
rect 23673 21913 23707 21947
rect 13001 21845 13035 21879
rect 13461 21845 13495 21879
rect 22109 21845 22143 21879
rect 22477 21845 22511 21879
rect 22569 21845 22603 21879
rect 23765 21845 23799 21879
rect 25605 21845 25639 21879
rect 28457 21845 28491 21879
rect 28825 21845 28859 21879
rect 37657 21845 37691 21879
rect 10241 21641 10275 21675
rect 19441 21641 19475 21675
rect 20729 21641 20763 21675
rect 25145 21641 25179 21675
rect 25513 21641 25547 21675
rect 29009 21641 29043 21675
rect 34253 21641 34287 21675
rect 40233 21641 40267 21675
rect 22753 21573 22787 21607
rect 38761 21573 38795 21607
rect 43821 21573 43855 21607
rect 9597 21505 9631 21539
rect 14473 21505 14507 21539
rect 19809 21505 19843 21539
rect 21097 21505 21131 21539
rect 21189 21505 21223 21539
rect 28181 21505 28215 21539
rect 29101 21505 29135 21539
rect 29837 21505 29871 21539
rect 32505 21505 32539 21539
rect 35357 21505 35391 21539
rect 36001 21505 36035 21539
rect 38485 21505 38519 21539
rect 47961 21505 47995 21539
rect 9781 21437 9815 21471
rect 19901 21437 19935 21471
rect 20085 21437 20119 21471
rect 21373 21437 21407 21471
rect 22477 21437 22511 21471
rect 25605 21437 25639 21471
rect 25697 21437 25731 21471
rect 29285 21437 29319 21471
rect 30113 21437 30147 21471
rect 31585 21437 31619 21471
rect 32781 21437 32815 21471
rect 49157 21437 49191 21471
rect 14289 21369 14323 21403
rect 27997 21369 28031 21403
rect 35173 21369 35207 21403
rect 44005 21369 44039 21403
rect 24225 21301 24259 21335
rect 28641 21301 28675 21335
rect 35817 21301 35851 21335
rect 9689 21097 9723 21131
rect 36645 21029 36679 21063
rect 9137 20961 9171 20995
rect 30941 20961 30975 20995
rect 38393 20961 38427 20995
rect 4169 20893 4203 20927
rect 9321 20893 9355 20927
rect 30665 20893 30699 20927
rect 31677 20893 31711 20927
rect 32321 20893 32355 20927
rect 36829 20893 36863 20927
rect 38209 20893 38243 20927
rect 47961 20893 47995 20927
rect 49157 20825 49191 20859
rect 4261 20757 4295 20791
rect 30297 20757 30331 20791
rect 30757 20757 30791 20791
rect 32137 20757 32171 20791
rect 37841 20757 37875 20791
rect 38301 20757 38335 20791
rect 21189 20553 21223 20587
rect 26249 20553 26283 20587
rect 30021 20553 30055 20587
rect 30481 20553 30515 20587
rect 32873 20553 32907 20587
rect 30389 20485 30423 20519
rect 32781 20485 32815 20519
rect 1777 20417 1811 20451
rect 21097 20417 21131 20451
rect 23029 20417 23063 20451
rect 26157 20417 26191 20451
rect 36921 20417 36955 20451
rect 47961 20417 47995 20451
rect 2053 20349 2087 20383
rect 21373 20349 21407 20383
rect 23305 20349 23339 20383
rect 26433 20349 26467 20383
rect 30665 20349 30699 20383
rect 33057 20349 33091 20383
rect 49157 20349 49191 20383
rect 20729 20213 20763 20247
rect 24777 20213 24811 20247
rect 25789 20213 25823 20247
rect 32413 20213 32447 20247
rect 36737 20213 36771 20247
rect 14289 20009 14323 20043
rect 19888 20009 19922 20043
rect 25237 20009 25271 20043
rect 26709 20009 26743 20043
rect 18153 19941 18187 19975
rect 21373 19941 21407 19975
rect 35633 19941 35667 19975
rect 18797 19873 18831 19907
rect 19625 19873 19659 19907
rect 21833 19873 21867 19907
rect 22109 19873 22143 19907
rect 23581 19873 23615 19907
rect 25789 19873 25823 19907
rect 27353 19873 27387 19907
rect 14473 19805 14507 19839
rect 32321 19805 32355 19839
rect 33149 19805 33183 19839
rect 33885 19805 33919 19839
rect 34989 19805 35023 19839
rect 35817 19805 35851 19839
rect 44097 19805 44131 19839
rect 27077 19737 27111 19771
rect 34069 19737 34103 19771
rect 44281 19737 44315 19771
rect 18521 19669 18555 19703
rect 18613 19669 18647 19703
rect 25605 19669 25639 19703
rect 25697 19669 25731 19703
rect 27169 19669 27203 19703
rect 32413 19669 32447 19703
rect 33241 19669 33275 19703
rect 35081 19669 35115 19703
rect 19901 19465 19935 19499
rect 23397 19465 23431 19499
rect 23765 19465 23799 19499
rect 39221 19465 39255 19499
rect 20361 19397 20395 19431
rect 26617 19397 26651 19431
rect 27537 19397 27571 19431
rect 20269 19329 20303 19363
rect 23857 19329 23891 19363
rect 24593 19329 24627 19363
rect 28733 19329 28767 19363
rect 33701 19329 33735 19363
rect 37473 19329 37507 19363
rect 47961 19329 47995 19363
rect 49157 19329 49191 19363
rect 20545 19261 20579 19295
rect 23949 19261 23983 19295
rect 24869 19261 24903 19295
rect 27629 19261 27663 19295
rect 27813 19261 27847 19295
rect 28825 19261 28859 19295
rect 28917 19261 28951 19295
rect 33977 19261 34011 19295
rect 37749 19261 37783 19295
rect 27169 19193 27203 19227
rect 28365 19193 28399 19227
rect 22845 19125 22879 19159
rect 35449 19125 35483 19159
rect 18153 18921 18187 18955
rect 20269 18921 20303 18955
rect 22477 18921 22511 18955
rect 24593 18921 24627 18955
rect 38669 18921 38703 18955
rect 18337 18853 18371 18887
rect 23305 18853 23339 18887
rect 30941 18853 30975 18887
rect 20913 18785 20947 18819
rect 23121 18785 23155 18819
rect 23857 18785 23891 18819
rect 25145 18785 25179 18819
rect 26617 18785 26651 18819
rect 29009 18785 29043 18819
rect 31401 18785 31435 18819
rect 31585 18785 31619 18819
rect 36921 18785 36955 18819
rect 4629 18717 4663 18751
rect 17877 18717 17911 18751
rect 22937 18717 22971 18751
rect 23673 18717 23707 18751
rect 26433 18717 26467 18751
rect 31309 18717 31343 18751
rect 44189 18717 44223 18751
rect 47961 18717 47995 18751
rect 20729 18649 20763 18683
rect 21465 18649 21499 18683
rect 22293 18649 22327 18683
rect 28273 18649 28307 18683
rect 36277 18649 36311 18683
rect 36461 18649 36495 18683
rect 37197 18649 37231 18683
rect 44373 18649 44407 18683
rect 49157 18649 49191 18683
rect 4721 18581 4755 18615
rect 20637 18581 20671 18615
rect 22845 18581 22879 18615
rect 23765 18581 23799 18615
rect 24961 18581 24995 18615
rect 25053 18581 25087 18615
rect 25973 18581 26007 18615
rect 26341 18581 26375 18615
rect 19809 18377 19843 18411
rect 27261 18377 27295 18411
rect 27629 18377 27663 18411
rect 34069 18377 34103 18411
rect 37933 18377 37967 18411
rect 20545 18309 20579 18343
rect 23305 18309 23339 18343
rect 28457 18309 28491 18343
rect 32597 18309 32631 18343
rect 1777 18241 1811 18275
rect 19717 18241 19751 18275
rect 23029 18241 23063 18275
rect 25053 18241 25087 18275
rect 27721 18241 27755 18275
rect 30205 18241 30239 18275
rect 30297 18241 30331 18275
rect 37841 18241 37875 18275
rect 47961 18241 47995 18275
rect 2053 18173 2087 18207
rect 19993 18173 20027 18207
rect 21281 18173 21315 18207
rect 27813 18173 27847 18207
rect 29285 18173 29319 18207
rect 30389 18173 30423 18207
rect 32321 18173 32355 18207
rect 34529 18173 34563 18207
rect 34805 18173 34839 18207
rect 38117 18173 38151 18207
rect 49157 18173 49191 18207
rect 19349 18037 19383 18071
rect 29837 18037 29871 18071
rect 36277 18037 36311 18071
rect 37473 18037 37507 18071
rect 19441 17833 19475 17867
rect 27353 17833 27387 17867
rect 32413 17833 32447 17867
rect 37289 17833 37323 17867
rect 18153 17765 18187 17799
rect 43177 17765 43211 17799
rect 18797 17697 18831 17731
rect 20085 17697 20119 17731
rect 21281 17697 21315 17731
rect 23029 17697 23063 17731
rect 27905 17697 27939 17731
rect 30665 17697 30699 17731
rect 33701 17697 33735 17731
rect 33885 17697 33919 17731
rect 35541 17697 35575 17731
rect 37749 17697 37783 17731
rect 38025 17697 38059 17731
rect 44649 17697 44683 17731
rect 21005 17629 21039 17663
rect 23673 17629 23707 17663
rect 27721 17629 27755 17663
rect 33609 17629 33643 17663
rect 43913 17629 43947 17663
rect 47961 17629 47995 17663
rect 18613 17561 18647 17595
rect 30021 17561 30055 17595
rect 30941 17561 30975 17595
rect 35817 17561 35851 17595
rect 42993 17561 43027 17595
rect 43729 17561 43763 17595
rect 44465 17561 44499 17595
rect 49157 17561 49191 17595
rect 18521 17493 18555 17527
rect 19809 17493 19843 17527
rect 19901 17493 19935 17527
rect 27813 17493 27847 17527
rect 30113 17493 30147 17527
rect 33241 17493 33275 17527
rect 39497 17493 39531 17527
rect 21465 17289 21499 17323
rect 22937 17289 22971 17323
rect 23305 17289 23339 17323
rect 23397 17289 23431 17323
rect 27261 17289 27295 17323
rect 27721 17289 27755 17323
rect 28825 17289 28859 17323
rect 35173 17289 35207 17323
rect 25053 17221 25087 17255
rect 27629 17221 27663 17255
rect 33977 17221 34011 17255
rect 43729 17221 43763 17255
rect 32505 17153 32539 17187
rect 33885 17153 33919 17187
rect 35081 17153 35115 17187
rect 36093 17153 36127 17187
rect 19717 17085 19751 17119
rect 19993 17085 20027 17119
rect 23581 17085 23615 17119
rect 24777 17085 24811 17119
rect 27813 17085 27847 17119
rect 28917 17085 28951 17119
rect 29101 17085 29135 17119
rect 30021 17085 30055 17119
rect 30297 17085 30331 17119
rect 31769 17085 31803 17119
rect 34161 17085 34195 17119
rect 35265 17085 35299 17119
rect 33517 17017 33551 17051
rect 34713 17017 34747 17051
rect 43913 17017 43947 17051
rect 26525 16949 26559 16983
rect 28457 16949 28491 16983
rect 32321 16949 32355 16983
rect 38117 16949 38151 16983
rect 19698 16745 19732 16779
rect 26249 16745 26283 16779
rect 23397 16677 23431 16711
rect 19441 16609 19475 16643
rect 21649 16609 21683 16643
rect 25053 16609 25087 16643
rect 25145 16609 25179 16643
rect 27721 16609 27755 16643
rect 34069 16609 34103 16643
rect 34253 16609 34287 16643
rect 34897 16609 34931 16643
rect 35173 16609 35207 16643
rect 38025 16609 38059 16643
rect 24961 16541 24995 16575
rect 26157 16541 26191 16575
rect 27537 16541 27571 16575
rect 33977 16541 34011 16575
rect 37933 16541 37967 16575
rect 47961 16541 47995 16575
rect 5549 16473 5583 16507
rect 21925 16473 21959 16507
rect 49157 16473 49191 16507
rect 5641 16405 5675 16439
rect 21189 16405 21223 16439
rect 24593 16405 24627 16439
rect 27169 16405 27203 16439
rect 27629 16405 27663 16439
rect 33609 16405 33643 16439
rect 36645 16405 36679 16439
rect 37473 16405 37507 16439
rect 37841 16405 37875 16439
rect 25697 16201 25731 16235
rect 25789 16201 25823 16235
rect 27169 16201 27203 16235
rect 27537 16201 27571 16235
rect 32965 16201 32999 16235
rect 23029 16133 23063 16167
rect 24777 16133 24811 16167
rect 1777 16065 1811 16099
rect 22753 16065 22787 16099
rect 27629 16065 27663 16099
rect 28825 16065 28859 16099
rect 33333 16065 33367 16099
rect 34345 16065 34379 16099
rect 36277 16065 36311 16099
rect 38853 16065 38887 16099
rect 47961 16065 47995 16099
rect 2053 15997 2087 16031
rect 25973 15997 26007 16031
rect 27721 15997 27755 16031
rect 29101 15997 29135 16031
rect 33425 15997 33459 16031
rect 33609 15997 33643 16031
rect 49157 15997 49191 16031
rect 25329 15861 25363 15895
rect 30573 15861 30607 15895
rect 34989 15861 35023 15895
rect 36093 15861 36127 15895
rect 37657 15861 37691 15895
rect 38669 15861 38703 15895
rect 26433 15657 26467 15691
rect 33057 15657 33091 15691
rect 29193 15589 29227 15623
rect 26985 15521 27019 15555
rect 28089 15521 28123 15555
rect 28273 15521 28307 15555
rect 29745 15521 29779 15555
rect 33609 15521 33643 15555
rect 35909 15521 35943 15555
rect 36185 15521 36219 15555
rect 27997 15453 28031 15487
rect 29009 15453 29043 15487
rect 32597 15453 32631 15487
rect 33425 15453 33459 15487
rect 33517 15453 33551 15487
rect 47961 15453 47995 15487
rect 24685 15385 24719 15419
rect 26801 15385 26835 15419
rect 30021 15385 30055 15419
rect 49157 15385 49191 15419
rect 24777 15317 24811 15351
rect 26893 15317 26927 15351
rect 27629 15317 27663 15351
rect 31493 15317 31527 15351
rect 32413 15317 32447 15351
rect 37657 15317 37691 15351
rect 20913 15113 20947 15147
rect 25881 15113 25915 15147
rect 29377 15113 29411 15147
rect 32781 15113 32815 15147
rect 37841 15113 37875 15147
rect 26249 15045 26283 15079
rect 29929 15045 29963 15079
rect 31585 15045 31619 15079
rect 37933 15045 37967 15079
rect 20821 14977 20855 15011
rect 22477 14977 22511 15011
rect 27629 14977 27663 15011
rect 32689 14977 32723 15011
rect 41797 14977 41831 15011
rect 47961 14977 47995 15011
rect 21097 14909 21131 14943
rect 22753 14909 22787 14943
rect 24225 14909 24259 14943
rect 26341 14909 26375 14943
rect 26525 14909 26559 14943
rect 27905 14909 27939 14943
rect 30113 14909 30147 14943
rect 32873 14909 32907 14943
rect 38025 14909 38059 14943
rect 49157 14909 49191 14943
rect 31769 14841 31803 14875
rect 32321 14841 32355 14875
rect 20453 14773 20487 14807
rect 30757 14773 30791 14807
rect 37473 14773 37507 14807
rect 41613 14773 41647 14807
rect 27629 14569 27663 14603
rect 32229 14569 32263 14603
rect 32689 14501 32723 14535
rect 37197 14501 37231 14535
rect 25881 14433 25915 14467
rect 30389 14433 30423 14467
rect 33149 14433 33183 14467
rect 33333 14433 33367 14467
rect 37657 14433 37691 14467
rect 37749 14433 37783 14467
rect 30205 14365 30239 14399
rect 33057 14365 33091 14399
rect 34989 14365 35023 14399
rect 37565 14365 37599 14399
rect 38577 14365 38611 14399
rect 40233 14365 40267 14399
rect 26157 14297 26191 14331
rect 35173 14297 35207 14331
rect 29837 14229 29871 14263
rect 30297 14229 30331 14263
rect 40049 14229 40083 14263
rect 36737 14025 36771 14059
rect 37565 13957 37599 13991
rect 37749 13957 37783 13991
rect 38301 13957 38335 13991
rect 1777 13889 1811 13923
rect 29009 13889 29043 13923
rect 30665 13889 30699 13923
rect 33885 13889 33919 13923
rect 36921 13889 36955 13923
rect 39129 13889 39163 13923
rect 41797 13889 41831 13923
rect 47961 13889 47995 13923
rect 2789 13821 2823 13855
rect 29193 13821 29227 13855
rect 35633 13821 35667 13855
rect 38485 13821 38519 13855
rect 49157 13821 49191 13855
rect 30481 13753 30515 13787
rect 38945 13753 38979 13787
rect 41613 13753 41647 13787
rect 34148 13685 34182 13719
rect 28273 13481 28307 13515
rect 36645 13481 36679 13515
rect 28825 13345 28859 13379
rect 34897 13345 34931 13379
rect 35173 13345 35207 13379
rect 25697 13277 25731 13311
rect 28733 13277 28767 13311
rect 34161 13277 34195 13311
rect 37197 13277 37231 13311
rect 38025 13277 38059 13311
rect 38669 13277 38703 13311
rect 40601 13277 40635 13311
rect 47961 13277 47995 13311
rect 28641 13209 28675 13243
rect 37381 13209 37415 13243
rect 49157 13209 49191 13243
rect 25789 13141 25823 13175
rect 34253 13141 34287 13175
rect 38485 13141 38519 13175
rect 40693 13141 40727 13175
rect 28825 12937 28859 12971
rect 29285 12937 29319 12971
rect 30481 12937 30515 12971
rect 35449 12937 35483 12971
rect 36277 12937 36311 12971
rect 27261 12869 27295 12903
rect 27997 12869 28031 12903
rect 29193 12869 29227 12903
rect 33977 12869 34011 12903
rect 43729 12869 43763 12903
rect 30389 12801 30423 12835
rect 33701 12801 33735 12835
rect 47961 12801 47995 12835
rect 29469 12733 29503 12767
rect 30573 12733 30607 12767
rect 36369 12733 36403 12767
rect 36461 12733 36495 12767
rect 49157 12733 49191 12767
rect 28181 12665 28215 12699
rect 30021 12665 30055 12699
rect 43913 12665 43947 12699
rect 27353 12597 27387 12631
rect 35909 12597 35943 12631
rect 28825 12189 28859 12223
rect 38945 12189 38979 12223
rect 41245 12189 41279 12223
rect 44465 12189 44499 12223
rect 47961 12189 47995 12223
rect 29009 12121 29043 12155
rect 39129 12121 39163 12155
rect 49157 12121 49191 12155
rect 41061 12053 41095 12087
rect 44281 12053 44315 12087
rect 46305 11781 46339 11815
rect 41613 11713 41647 11747
rect 44833 11713 44867 11747
rect 45569 11713 45603 11747
rect 45017 11577 45051 11611
rect 45753 11577 45787 11611
rect 41429 11509 41463 11543
rect 46397 11509 46431 11543
rect 13001 11305 13035 11339
rect 13645 11169 13679 11203
rect 13369 11101 13403 11135
rect 14473 11101 14507 11135
rect 47961 11101 47995 11135
rect 49157 11101 49191 11135
rect 12449 11033 12483 11067
rect 13461 11033 13495 11067
rect 46305 11033 46339 11067
rect 46489 11033 46523 11067
rect 24501 10693 24535 10727
rect 40785 10625 40819 10659
rect 47961 10625 47995 10659
rect 49157 10557 49191 10591
rect 24685 10489 24719 10523
rect 40601 10421 40635 10455
rect 28733 10013 28767 10047
rect 31861 10013 31895 10047
rect 47961 10013 47995 10047
rect 28917 9945 28951 9979
rect 49157 9945 49191 9979
rect 31953 9877 31987 9911
rect 32413 9605 32447 9639
rect 35909 9605 35943 9639
rect 46305 9537 46339 9571
rect 47961 9537 47995 9571
rect 49157 9469 49191 9503
rect 32597 9401 32631 9435
rect 36093 9401 36127 9435
rect 46121 9333 46155 9367
rect 46029 8925 46063 8959
rect 48881 8925 48915 8959
rect 46213 8857 46247 8891
rect 47961 8857 47995 8891
rect 48697 8857 48731 8891
rect 48053 8789 48087 8823
rect 36553 8517 36587 8551
rect 37841 8517 37875 8551
rect 45753 8517 45787 8551
rect 9137 8449 9171 8483
rect 47961 8449 47995 8483
rect 9413 8381 9447 8415
rect 11161 8381 11195 8415
rect 36737 8381 36771 8415
rect 49157 8381 49191 8415
rect 38025 8313 38059 8347
rect 45937 8313 45971 8347
rect 47961 7837 47995 7871
rect 49157 7769 49191 7803
rect 35725 7429 35759 7463
rect 37565 7361 37599 7395
rect 47961 7361 47995 7395
rect 35909 7293 35943 7327
rect 49157 7293 49191 7327
rect 37749 7225 37783 7259
rect 37749 6749 37783 6783
rect 47961 6749 47995 6783
rect 37565 6681 37599 6715
rect 38301 6681 38335 6715
rect 38485 6681 38519 6715
rect 49157 6681 49191 6715
rect 47961 5661 47995 5695
rect 49157 5661 49191 5695
rect 30113 5185 30147 5219
rect 29469 4981 29503 5015
rect 30205 4981 30239 5015
rect 49341 4981 49375 5015
rect 47961 4573 47995 4607
rect 49157 4505 49191 4539
rect 33977 4097 34011 4131
rect 39129 4097 39163 4131
rect 43545 4097 43579 4131
rect 46029 4097 46063 4131
rect 48697 4097 48731 4131
rect 34437 4029 34471 4063
rect 39589 4029 39623 4063
rect 44005 4029 44039 4063
rect 48881 3961 48915 3995
rect 45845 3893 45879 3927
rect 1593 3689 1627 3723
rect 25053 3553 25087 3587
rect 30205 3553 30239 3587
rect 32045 3553 32079 3587
rect 35357 3553 35391 3587
rect 37197 3553 37231 3587
rect 40509 3553 40543 3587
rect 42349 3553 42383 3587
rect 45661 3553 45695 3587
rect 1777 3485 1811 3519
rect 24777 3485 24811 3519
rect 29745 3485 29779 3519
rect 31585 3485 31619 3519
rect 34897 3485 34931 3519
rect 36737 3485 36771 3519
rect 40049 3485 40083 3519
rect 41889 3485 41923 3519
rect 45201 3485 45235 3519
rect 47961 3485 47995 3519
rect 49157 3417 49191 3451
rect 2329 3145 2363 3179
rect 10609 3145 10643 3179
rect 47133 3145 47167 3179
rect 12909 3077 12943 3111
rect 1593 3009 1627 3043
rect 2513 3009 2547 3043
rect 3893 3009 3927 3043
rect 5365 3009 5399 3043
rect 5733 3009 5767 3043
rect 6837 3009 6871 3043
rect 7021 3009 7055 3043
rect 10425 3009 10459 3043
rect 12725 3009 12759 3043
rect 14105 3009 14139 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 20913 3009 20947 3043
rect 22293 3009 22327 3043
rect 23397 3009 23431 3043
rect 25145 3009 25179 3043
rect 27537 3009 27571 3043
rect 29193 3009 29227 3043
rect 32321 3009 32355 3043
rect 34161 3009 34195 3043
rect 37657 3009 37691 3043
rect 39313 3009 39347 3043
rect 42625 3009 42659 3043
rect 44465 3009 44499 3043
rect 46949 3009 46983 3043
rect 47961 3009 47995 3043
rect 19257 2941 19291 2975
rect 19533 2941 19567 2975
rect 20637 2941 20671 2975
rect 22017 2941 22051 2975
rect 23765 2941 23799 2975
rect 25605 2941 25639 2975
rect 27813 2941 27847 2975
rect 29653 2941 29687 2975
rect 32781 2941 32815 2975
rect 34621 2941 34655 2975
rect 37933 2941 37967 2975
rect 39773 2941 39807 2975
rect 43085 2941 43119 2975
rect 44925 2941 44959 2975
rect 48421 2941 48455 2975
rect 1777 2873 1811 2907
rect 4077 2873 4111 2907
rect 14289 2873 14323 2907
rect 10057 2601 10091 2635
rect 11069 2601 11103 2635
rect 13645 2601 13679 2635
rect 14565 2601 14599 2635
rect 20085 2601 20119 2635
rect 46765 2601 46799 2635
rect 12265 2533 12299 2567
rect 9505 2465 9539 2499
rect 18061 2465 18095 2499
rect 20637 2465 20671 2499
rect 23121 2465 23155 2499
rect 25789 2465 25823 2499
rect 27629 2465 27663 2499
rect 30205 2465 30239 2499
rect 32781 2465 32815 2499
rect 37933 2465 37967 2499
rect 40509 2465 40543 2499
rect 43085 2465 43119 2499
rect 48329 2465 48363 2499
rect 2145 2397 2179 2431
rect 7297 2397 7331 2431
rect 10241 2397 10275 2431
rect 14381 2397 14415 2431
rect 18337 2397 18371 2431
rect 19809 2397 19843 2431
rect 20913 2397 20947 2431
rect 22661 2397 22695 2431
rect 25237 2397 25271 2431
rect 27169 2397 27203 2431
rect 29929 2397 29963 2431
rect 32321 2397 32355 2431
rect 34897 2397 34931 2431
rect 37473 2397 37507 2431
rect 40049 2397 40083 2431
rect 42625 2397 42659 2431
rect 47777 2397 47811 2431
rect 3065 2329 3099 2363
rect 4629 2329 4663 2363
rect 4997 2329 5031 2363
rect 5641 2329 5675 2363
rect 6009 2329 6043 2363
rect 8217 2329 8251 2363
rect 9229 2329 9263 2363
rect 10793 2329 10827 2363
rect 11989 2329 12023 2363
rect 13369 2329 13403 2363
rect 15209 2329 15243 2363
rect 15945 2329 15979 2363
rect 16313 2329 16347 2363
rect 17141 2329 17175 2363
rect 35817 2329 35851 2363
rect 45477 2329 45511 2363
rect 2421 2261 2455 2295
rect 3341 2261 3375 2295
rect 7573 2261 7607 2295
rect 8493 2261 8527 2295
rect 15301 2261 15335 2295
rect 17417 2261 17451 2295
<< metal1 >>
rect 382 55700 388 55752
rect 440 55740 446 55752
rect 2866 55740 2872 55752
rect 440 55712 2872 55740
rect 440 55700 446 55712
rect 2866 55700 2872 55712
rect 2924 55700 2930 55752
rect 46842 55700 46848 55752
rect 46900 55740 46906 55752
rect 50430 55740 50436 55752
rect 46900 55712 50436 55740
rect 46900 55700 46906 55712
rect 50430 55700 50436 55712
rect 50488 55700 50494 55752
rect 1104 54426 49864 54448
rect 1104 54374 7950 54426
rect 8002 54374 8014 54426
rect 8066 54374 8078 54426
rect 8130 54374 8142 54426
rect 8194 54374 8206 54426
rect 8258 54374 17950 54426
rect 18002 54374 18014 54426
rect 18066 54374 18078 54426
rect 18130 54374 18142 54426
rect 18194 54374 18206 54426
rect 18258 54374 27950 54426
rect 28002 54374 28014 54426
rect 28066 54374 28078 54426
rect 28130 54374 28142 54426
rect 28194 54374 28206 54426
rect 28258 54374 37950 54426
rect 38002 54374 38014 54426
rect 38066 54374 38078 54426
rect 38130 54374 38142 54426
rect 38194 54374 38206 54426
rect 38258 54374 47950 54426
rect 48002 54374 48014 54426
rect 48066 54374 48078 54426
rect 48130 54374 48142 54426
rect 48194 54374 48206 54426
rect 48258 54374 49864 54426
rect 1104 54352 49864 54374
rect 10042 54312 10048 54324
rect 4816 54284 10048 54312
rect 3237 54247 3295 54253
rect 3237 54213 3249 54247
rect 3283 54244 3295 54247
rect 3326 54244 3332 54256
rect 3283 54216 3332 54244
rect 3283 54213 3295 54216
rect 3237 54207 3295 54213
rect 3326 54204 3332 54216
rect 3384 54204 3390 54256
rect 2225 54179 2283 54185
rect 2225 54145 2237 54179
rect 2271 54145 2283 54179
rect 2225 54139 2283 54145
rect 2240 54108 2268 54139
rect 2774 54136 2780 54188
rect 2832 54176 2838 54188
rect 4816 54185 4844 54284
rect 10042 54272 10048 54284
rect 10100 54272 10106 54324
rect 41690 54272 41696 54324
rect 41748 54312 41754 54324
rect 45189 54315 45247 54321
rect 45189 54312 45201 54315
rect 41748 54284 45201 54312
rect 41748 54272 41754 54284
rect 45189 54281 45201 54284
rect 45235 54281 45247 54315
rect 45189 54275 45247 54281
rect 5813 54247 5871 54253
rect 5813 54213 5825 54247
rect 5859 54244 5871 54247
rect 6270 54244 6276 54256
rect 5859 54216 6276 54244
rect 5859 54213 5871 54216
rect 5813 54207 5871 54213
rect 6270 54204 6276 54216
rect 6328 54204 6334 54256
rect 8389 54247 8447 54253
rect 8389 54213 8401 54247
rect 8435 54244 8447 54247
rect 8478 54244 8484 54256
rect 8435 54216 8484 54244
rect 8435 54213 8447 54216
rect 8389 54207 8447 54213
rect 8478 54204 8484 54216
rect 8536 54204 8542 54256
rect 10965 54247 11023 54253
rect 9416 54216 9904 54244
rect 4157 54179 4215 54185
rect 4157 54176 4169 54179
rect 2832 54148 4169 54176
rect 2832 54136 2838 54148
rect 4157 54145 4169 54148
rect 4203 54145 4215 54179
rect 4157 54139 4215 54145
rect 4801 54179 4859 54185
rect 4801 54145 4813 54179
rect 4847 54145 4859 54179
rect 4801 54139 4859 54145
rect 7377 54179 7435 54185
rect 7377 54145 7389 54179
rect 7423 54176 7435 54179
rect 9416 54176 9444 54216
rect 7423 54148 9444 54176
rect 9769 54179 9827 54185
rect 7423 54145 7435 54148
rect 7377 54139 7435 54145
rect 9769 54145 9781 54179
rect 9815 54145 9827 54179
rect 9876 54176 9904 54216
rect 10965 54213 10977 54247
rect 11011 54244 11023 54247
rect 11422 54244 11428 54256
rect 11011 54216 11428 54244
rect 11011 54213 11023 54216
rect 10965 54207 11023 54213
rect 11422 54204 11428 54216
rect 11480 54204 11486 54256
rect 13541 54247 13599 54253
rect 13541 54213 13553 54247
rect 13587 54244 13599 54247
rect 13630 54244 13636 54256
rect 13587 54216 13636 54244
rect 13587 54213 13599 54216
rect 13541 54207 13599 54213
rect 13630 54204 13636 54216
rect 13688 54204 13694 54256
rect 16117 54247 16175 54253
rect 16117 54213 16129 54247
rect 16163 54244 16175 54247
rect 16574 54244 16580 54256
rect 16163 54216 16580 54244
rect 16163 54213 16175 54216
rect 16117 54207 16175 54213
rect 16574 54204 16580 54216
rect 16632 54204 16638 54256
rect 18693 54247 18751 54253
rect 18693 54213 18705 54247
rect 18739 54244 18751 54247
rect 18782 54244 18788 54256
rect 18739 54216 18788 54244
rect 18739 54213 18751 54216
rect 18693 54207 18751 54213
rect 18782 54204 18788 54216
rect 18840 54204 18846 54256
rect 20990 54204 20996 54256
rect 21048 54204 21054 54256
rect 28350 54204 28356 54256
rect 28408 54244 28414 54256
rect 28721 54247 28779 54253
rect 28721 54244 28733 54247
rect 28408 54216 28733 54244
rect 28408 54204 28414 54216
rect 28721 54213 28733 54216
rect 28767 54213 28779 54247
rect 28721 54207 28779 54213
rect 32766 54204 32772 54256
rect 32824 54244 32830 54256
rect 32953 54247 33011 54253
rect 32953 54244 32965 54247
rect 32824 54216 32965 54244
rect 32824 54204 32830 54216
rect 32953 54213 32965 54216
rect 32999 54213 33011 54247
rect 32953 54207 33011 54213
rect 33502 54204 33508 54256
rect 33560 54244 33566 54256
rect 33689 54247 33747 54253
rect 33689 54244 33701 54247
rect 33560 54216 33701 54244
rect 33560 54204 33566 54216
rect 33689 54213 33701 54216
rect 33735 54213 33747 54247
rect 33689 54207 33747 54213
rect 37182 54204 37188 54256
rect 37240 54244 37246 54256
rect 37553 54247 37611 54253
rect 37553 54244 37565 54247
rect 37240 54216 37565 54244
rect 37240 54204 37246 54216
rect 37553 54213 37565 54216
rect 37599 54213 37611 54247
rect 37553 54207 37611 54213
rect 42334 54204 42340 54256
rect 42392 54244 42398 54256
rect 42705 54247 42763 54253
rect 42705 54244 42717 54247
rect 42392 54216 42717 54244
rect 42392 54204 42398 54216
rect 42705 54213 42717 54216
rect 42751 54213 42763 54247
rect 42705 54207 42763 54213
rect 11698 54176 11704 54188
rect 9876 54148 11704 54176
rect 9769 54139 9827 54145
rect 2240 54080 6914 54108
rect 3970 53932 3976 53984
rect 4028 53932 4034 53984
rect 6886 53972 6914 54080
rect 9784 54040 9812 54139
rect 11698 54136 11704 54148
rect 11756 54136 11762 54188
rect 12529 54179 12587 54185
rect 12529 54145 12541 54179
rect 12575 54176 12587 54179
rect 14550 54176 14556 54188
rect 12575 54148 14556 54176
rect 12575 54145 12587 54148
rect 12529 54139 12587 54145
rect 14550 54136 14556 54148
rect 14608 54136 14614 54188
rect 15105 54179 15163 54185
rect 15105 54145 15117 54179
rect 15151 54145 15163 54179
rect 15105 54139 15163 54145
rect 15120 54108 15148 54139
rect 17678 54136 17684 54188
rect 17736 54136 17742 54188
rect 20257 54179 20315 54185
rect 20257 54145 20269 54179
rect 20303 54176 20315 54179
rect 20346 54176 20352 54188
rect 20303 54148 20352 54176
rect 20303 54145 20315 54148
rect 20257 54139 20315 54145
rect 20346 54136 20352 54148
rect 20404 54136 20410 54188
rect 22738 54136 22744 54188
rect 22796 54136 22802 54188
rect 24670 54136 24676 54188
rect 24728 54176 24734 54188
rect 24765 54179 24823 54185
rect 24765 54176 24777 54179
rect 24728 54148 24777 54176
rect 24728 54136 24734 54148
rect 24765 54145 24777 54148
rect 24811 54145 24823 54179
rect 24765 54139 24823 54145
rect 25406 54136 25412 54188
rect 25464 54176 25470 54188
rect 25501 54179 25559 54185
rect 25501 54176 25513 54179
rect 25464 54148 25513 54176
rect 25464 54136 25470 54148
rect 25501 54145 25513 54148
rect 25547 54145 25559 54179
rect 25501 54139 25559 54145
rect 26234 54136 26240 54188
rect 26292 54176 26298 54188
rect 26421 54179 26479 54185
rect 26421 54176 26433 54179
rect 26292 54148 26433 54176
rect 26292 54136 26298 54148
rect 26421 54145 26433 54148
rect 26467 54145 26479 54179
rect 26421 54139 26479 54145
rect 26878 54136 26884 54188
rect 26936 54176 26942 54188
rect 27157 54179 27215 54185
rect 27157 54176 27169 54179
rect 26936 54148 27169 54176
rect 26936 54136 26942 54148
rect 27157 54145 27169 54148
rect 27203 54145 27215 54179
rect 27157 54139 27215 54145
rect 27614 54136 27620 54188
rect 27672 54176 27678 54188
rect 27893 54179 27951 54185
rect 27893 54176 27905 54179
rect 27672 54148 27905 54176
rect 27672 54136 27678 54148
rect 27893 54145 27905 54148
rect 27939 54145 27951 54179
rect 27893 54139 27951 54145
rect 29822 54136 29828 54188
rect 29880 54176 29886 54188
rect 29917 54179 29975 54185
rect 29917 54176 29929 54179
rect 29880 54148 29929 54176
rect 29880 54136 29886 54148
rect 29917 54145 29929 54148
rect 29963 54145 29975 54179
rect 29917 54139 29975 54145
rect 30558 54136 30564 54188
rect 30616 54176 30622 54188
rect 30653 54179 30711 54185
rect 30653 54176 30665 54179
rect 30616 54148 30665 54176
rect 30616 54136 30622 54148
rect 30653 54145 30665 54148
rect 30699 54145 30711 54179
rect 30653 54139 30711 54145
rect 31294 54136 31300 54188
rect 31352 54176 31358 54188
rect 31389 54179 31447 54185
rect 31389 54176 31401 54179
rect 31352 54148 31401 54176
rect 31352 54136 31358 54148
rect 31389 54145 31401 54148
rect 31435 54145 31447 54179
rect 31389 54139 31447 54145
rect 34238 54136 34244 54188
rect 34296 54176 34302 54188
rect 34885 54179 34943 54185
rect 34885 54176 34897 54179
rect 34296 54148 34897 54176
rect 34296 54136 34302 54148
rect 34885 54145 34897 54148
rect 34931 54145 34943 54179
rect 34885 54139 34943 54145
rect 35710 54136 35716 54188
rect 35768 54176 35774 54188
rect 35805 54179 35863 54185
rect 35805 54176 35817 54179
rect 35768 54148 35817 54176
rect 35768 54136 35774 54148
rect 35805 54145 35817 54148
rect 35851 54145 35863 54179
rect 35805 54139 35863 54145
rect 36446 54136 36452 54188
rect 36504 54176 36510 54188
rect 36541 54179 36599 54185
rect 36541 54176 36553 54179
rect 36504 54148 36553 54176
rect 36504 54136 36510 54148
rect 36541 54145 36553 54148
rect 36587 54145 36599 54179
rect 36541 54139 36599 54145
rect 38654 54136 38660 54188
rect 38712 54176 38718 54188
rect 38749 54179 38807 54185
rect 38749 54176 38761 54179
rect 38712 54148 38761 54176
rect 38712 54136 38718 54148
rect 38749 54145 38761 54148
rect 38795 54145 38807 54179
rect 38749 54139 38807 54145
rect 39390 54136 39396 54188
rect 39448 54176 39454 54188
rect 40037 54179 40095 54185
rect 40037 54176 40049 54179
rect 39448 54148 40049 54176
rect 39448 54136 39454 54148
rect 40037 54145 40049 54148
rect 40083 54145 40095 54179
rect 40037 54139 40095 54145
rect 40126 54136 40132 54188
rect 40184 54176 40190 54188
rect 40773 54179 40831 54185
rect 40773 54176 40785 54179
rect 40184 54148 40785 54176
rect 40184 54136 40190 54148
rect 40773 54145 40785 54148
rect 40819 54145 40831 54179
rect 40773 54139 40831 54145
rect 40862 54136 40868 54188
rect 40920 54176 40926 54188
rect 41693 54179 41751 54185
rect 41693 54176 41705 54179
rect 40920 54148 41705 54176
rect 40920 54136 40926 54148
rect 41693 54145 41705 54148
rect 41739 54145 41751 54179
rect 41693 54139 41751 54145
rect 43070 54136 43076 54188
rect 43128 54176 43134 54188
rect 43717 54179 43775 54185
rect 43717 54176 43729 54179
rect 43128 54148 43729 54176
rect 43128 54136 43134 54148
rect 43717 54145 43729 54148
rect 43763 54145 43775 54179
rect 43717 54139 43775 54145
rect 44082 54136 44088 54188
rect 44140 54176 44146 54188
rect 44361 54179 44419 54185
rect 44361 54176 44373 54179
rect 44140 54148 44373 54176
rect 44140 54136 44146 54148
rect 44361 54145 44373 54148
rect 44407 54145 44419 54179
rect 44361 54139 44419 54145
rect 44542 54136 44548 54188
rect 44600 54176 44606 54188
rect 45373 54179 45431 54185
rect 45373 54176 45385 54179
rect 44600 54148 45385 54176
rect 44600 54136 44606 54148
rect 45373 54145 45385 54148
rect 45419 54145 45431 54179
rect 45373 54139 45431 54145
rect 46569 54179 46627 54185
rect 46569 54145 46581 54179
rect 46615 54176 46627 54179
rect 46842 54176 46848 54188
rect 46615 54148 46848 54176
rect 46615 54145 46627 54148
rect 46569 54139 46627 54145
rect 46842 54136 46848 54148
rect 46900 54136 46906 54188
rect 47213 54179 47271 54185
rect 47213 54145 47225 54179
rect 47259 54176 47271 54179
rect 47486 54176 47492 54188
rect 47259 54148 47492 54176
rect 47259 54145 47271 54148
rect 47213 54139 47271 54145
rect 47486 54136 47492 54148
rect 47544 54136 47550 54188
rect 47854 54136 47860 54188
rect 47912 54176 47918 54188
rect 47949 54179 48007 54185
rect 47949 54176 47961 54179
rect 47912 54148 47961 54176
rect 47912 54136 47918 54148
rect 47949 54145 47961 54148
rect 47995 54145 48007 54179
rect 47949 54139 48007 54145
rect 20162 54108 20168 54120
rect 15120 54080 20168 54108
rect 20162 54068 20168 54080
rect 20220 54068 20226 54120
rect 22462 54068 22468 54120
rect 22520 54108 22526 54120
rect 23017 54111 23075 54117
rect 23017 54108 23029 54111
rect 22520 54080 23029 54108
rect 22520 54068 22526 54080
rect 23017 54077 23029 54080
rect 23063 54077 23075 54111
rect 23017 54071 23075 54077
rect 48222 54068 48228 54120
rect 48280 54108 48286 54120
rect 48409 54111 48467 54117
rect 48409 54108 48421 54111
rect 48280 54080 48421 54108
rect 48280 54068 48286 54080
rect 48409 54077 48421 54080
rect 48455 54077 48467 54111
rect 48409 54071 48467 54077
rect 14642 54040 14648 54052
rect 9784 54012 14648 54040
rect 14642 54000 14648 54012
rect 14700 54000 14706 54052
rect 28905 54043 28963 54049
rect 28905 54009 28917 54043
rect 28951 54040 28963 54043
rect 29638 54040 29644 54052
rect 28951 54012 29644 54040
rect 28951 54009 28963 54012
rect 28905 54003 28963 54009
rect 29638 54000 29644 54012
rect 29696 54000 29702 54052
rect 33137 54043 33195 54049
rect 33137 54009 33149 54043
rect 33183 54040 33195 54043
rect 33318 54040 33324 54052
rect 33183 54012 33324 54040
rect 33183 54009 33195 54012
rect 33137 54003 33195 54009
rect 33318 54000 33324 54012
rect 33376 54000 33382 54052
rect 33873 54043 33931 54049
rect 33873 54009 33885 54043
rect 33919 54040 33931 54043
rect 33962 54040 33968 54052
rect 33919 54012 33968 54040
rect 33919 54009 33931 54012
rect 33873 54003 33931 54009
rect 33962 54000 33968 54012
rect 34020 54000 34026 54052
rect 40310 54000 40316 54052
rect 40368 54040 40374 54052
rect 42981 54043 43039 54049
rect 40368 54012 41644 54040
rect 40368 54000 40374 54012
rect 12342 53972 12348 53984
rect 6886 53944 12348 53972
rect 12342 53932 12348 53944
rect 12400 53932 12406 53984
rect 24946 53932 24952 53984
rect 25004 53932 25010 53984
rect 25682 53932 25688 53984
rect 25740 53932 25746 53984
rect 26234 53932 26240 53984
rect 26292 53932 26298 53984
rect 27341 53975 27399 53981
rect 27341 53941 27353 53975
rect 27387 53972 27399 53975
rect 27430 53972 27436 53984
rect 27387 53944 27436 53972
rect 27387 53941 27399 53944
rect 27341 53935 27399 53941
rect 27430 53932 27436 53944
rect 27488 53932 27494 53984
rect 28077 53975 28135 53981
rect 28077 53941 28089 53975
rect 28123 53972 28135 53975
rect 28534 53972 28540 53984
rect 28123 53944 28540 53972
rect 28123 53941 28135 53944
rect 28077 53935 28135 53941
rect 28534 53932 28540 53944
rect 28592 53932 28598 53984
rect 30006 53932 30012 53984
rect 30064 53972 30070 53984
rect 30101 53975 30159 53981
rect 30101 53972 30113 53975
rect 30064 53944 30113 53972
rect 30064 53932 30070 53944
rect 30101 53941 30113 53944
rect 30147 53941 30159 53975
rect 30101 53935 30159 53941
rect 30742 53932 30748 53984
rect 30800 53972 30806 53984
rect 30837 53975 30895 53981
rect 30837 53972 30849 53975
rect 30800 53944 30849 53972
rect 30800 53932 30806 53944
rect 30837 53941 30849 53944
rect 30883 53941 30895 53975
rect 30837 53935 30895 53941
rect 31386 53932 31392 53984
rect 31444 53972 31450 53984
rect 31573 53975 31631 53981
rect 31573 53972 31585 53975
rect 31444 53944 31585 53972
rect 31444 53932 31450 53944
rect 31573 53941 31585 53944
rect 31619 53941 31631 53975
rect 31573 53935 31631 53941
rect 35066 53932 35072 53984
rect 35124 53932 35130 53984
rect 35989 53975 36047 53981
rect 35989 53941 36001 53975
rect 36035 53972 36047 53975
rect 36538 53972 36544 53984
rect 36035 53944 36544 53972
rect 36035 53941 36047 53944
rect 35989 53935 36047 53941
rect 36538 53932 36544 53944
rect 36596 53932 36602 53984
rect 36722 53932 36728 53984
rect 36780 53932 36786 53984
rect 37642 53932 37648 53984
rect 37700 53932 37706 53984
rect 38930 53932 38936 53984
rect 38988 53932 38994 53984
rect 40221 53975 40279 53981
rect 40221 53941 40233 53975
rect 40267 53972 40279 53975
rect 40402 53972 40408 53984
rect 40267 53944 40408 53972
rect 40267 53941 40279 53944
rect 40221 53935 40279 53941
rect 40402 53932 40408 53944
rect 40460 53932 40466 53984
rect 40957 53975 41015 53981
rect 40957 53941 40969 53975
rect 41003 53972 41015 53975
rect 41322 53972 41328 53984
rect 41003 53944 41328 53972
rect 41003 53941 41015 53944
rect 40957 53935 41015 53941
rect 41322 53932 41328 53944
rect 41380 53932 41386 53984
rect 41506 53932 41512 53984
rect 41564 53932 41570 53984
rect 41616 53972 41644 54012
rect 42981 54009 42993 54043
rect 43027 54040 43039 54043
rect 43622 54040 43628 54052
rect 43027 54012 43628 54040
rect 43027 54009 43039 54012
rect 42981 54003 43039 54009
rect 43622 54000 43628 54012
rect 43680 54000 43686 54052
rect 43533 53975 43591 53981
rect 43533 53972 43545 53975
rect 41616 53944 43545 53972
rect 43533 53941 43545 53944
rect 43579 53941 43591 53975
rect 43533 53935 43591 53941
rect 44174 53932 44180 53984
rect 44232 53932 44238 53984
rect 46382 53932 46388 53984
rect 46440 53932 46446 53984
rect 47026 53932 47032 53984
rect 47084 53932 47090 53984
rect 1104 53882 49864 53904
rect 1104 53830 2950 53882
rect 3002 53830 3014 53882
rect 3066 53830 3078 53882
rect 3130 53830 3142 53882
rect 3194 53830 3206 53882
rect 3258 53830 12950 53882
rect 13002 53830 13014 53882
rect 13066 53830 13078 53882
rect 13130 53830 13142 53882
rect 13194 53830 13206 53882
rect 13258 53830 22950 53882
rect 23002 53830 23014 53882
rect 23066 53830 23078 53882
rect 23130 53830 23142 53882
rect 23194 53830 23206 53882
rect 23258 53830 32950 53882
rect 33002 53830 33014 53882
rect 33066 53830 33078 53882
rect 33130 53830 33142 53882
rect 33194 53830 33206 53882
rect 33258 53830 42950 53882
rect 43002 53830 43014 53882
rect 43066 53830 43078 53882
rect 43130 53830 43142 53882
rect 43194 53830 43206 53882
rect 43258 53830 49864 53882
rect 1104 53808 49864 53830
rect 15838 53660 15844 53712
rect 15896 53660 15902 53712
rect 23661 53703 23719 53709
rect 23661 53669 23673 53703
rect 23707 53700 23719 53703
rect 27062 53700 27068 53712
rect 23707 53672 27068 53700
rect 23707 53669 23719 53672
rect 23661 53663 23719 53669
rect 27062 53660 27068 53672
rect 27120 53660 27126 53712
rect 1854 53592 1860 53644
rect 1912 53632 1918 53644
rect 2409 53635 2467 53641
rect 2409 53632 2421 53635
rect 1912 53604 2421 53632
rect 1912 53592 1918 53604
rect 2409 53601 2421 53604
rect 2455 53601 2467 53635
rect 2409 53595 2467 53601
rect 5534 53592 5540 53644
rect 5592 53632 5598 53644
rect 5721 53635 5779 53641
rect 5721 53632 5733 53635
rect 5592 53604 5733 53632
rect 5592 53592 5598 53604
rect 5721 53601 5733 53604
rect 5767 53601 5779 53635
rect 5721 53595 5779 53601
rect 7006 53592 7012 53644
rect 7064 53632 7070 53644
rect 7561 53635 7619 53641
rect 7561 53632 7573 53635
rect 7064 53604 7573 53632
rect 7064 53592 7070 53604
rect 7561 53601 7573 53604
rect 7607 53601 7619 53635
rect 7561 53595 7619 53601
rect 10686 53592 10692 53644
rect 10744 53632 10750 53644
rect 10873 53635 10931 53641
rect 10873 53632 10885 53635
rect 10744 53604 10885 53632
rect 10744 53592 10750 53604
rect 10873 53601 10885 53604
rect 10919 53601 10931 53635
rect 10873 53595 10931 53601
rect 12158 53592 12164 53644
rect 12216 53632 12222 53644
rect 12713 53635 12771 53641
rect 12713 53632 12725 53635
rect 12216 53604 12725 53632
rect 12216 53592 12222 53604
rect 12713 53601 12725 53604
rect 12759 53601 12771 53635
rect 15856 53632 15884 53660
rect 16117 53635 16175 53641
rect 16117 53632 16129 53635
rect 15856 53604 16129 53632
rect 12713 53595 12771 53601
rect 16117 53601 16129 53604
rect 16163 53601 16175 53635
rect 16117 53595 16175 53601
rect 18322 53592 18328 53644
rect 18380 53592 18386 53644
rect 20254 53592 20260 53644
rect 20312 53632 20318 53644
rect 20441 53635 20499 53641
rect 20441 53632 20453 53635
rect 20312 53604 20453 53632
rect 20312 53592 20318 53604
rect 20441 53601 20453 53604
rect 20487 53601 20499 53635
rect 20441 53595 20499 53601
rect 21726 53592 21732 53644
rect 21784 53632 21790 53644
rect 22281 53635 22339 53641
rect 22281 53632 22293 53635
rect 21784 53604 22293 53632
rect 21784 53592 21790 53604
rect 22281 53601 22293 53604
rect 22327 53601 22339 53635
rect 22281 53595 22339 53601
rect 46750 53592 46756 53644
rect 46808 53632 46814 53644
rect 47305 53635 47363 53641
rect 47305 53632 47317 53635
rect 46808 53604 47317 53632
rect 46808 53592 46814 53604
rect 47305 53601 47317 53604
rect 47351 53601 47363 53635
rect 47305 53595 47363 53601
rect 2133 53567 2191 53573
rect 2133 53533 2145 53567
rect 2179 53533 2191 53567
rect 2133 53527 2191 53533
rect 5445 53567 5503 53573
rect 5445 53533 5457 53567
rect 5491 53564 5503 53567
rect 7285 53567 7343 53573
rect 5491 53536 6914 53564
rect 5491 53533 5503 53536
rect 5445 53527 5503 53533
rect 2148 53496 2176 53527
rect 6362 53496 6368 53508
rect 2148 53468 6368 53496
rect 6362 53456 6368 53468
rect 6420 53456 6426 53508
rect 6886 53496 6914 53536
rect 7285 53533 7297 53567
rect 7331 53564 7343 53567
rect 8938 53564 8944 53576
rect 7331 53536 8944 53564
rect 7331 53533 7343 53536
rect 7285 53527 7343 53533
rect 8938 53524 8944 53536
rect 8996 53524 9002 53576
rect 10410 53524 10416 53576
rect 10468 53524 10474 53576
rect 12345 53567 12403 53573
rect 12345 53533 12357 53567
rect 12391 53564 12403 53567
rect 14734 53564 14740 53576
rect 12391 53536 14740 53564
rect 12391 53533 12403 53536
rect 12345 53527 12403 53533
rect 14734 53524 14740 53536
rect 14792 53524 14798 53576
rect 15841 53567 15899 53573
rect 15841 53533 15853 53567
rect 15887 53533 15899 53567
rect 15841 53527 15899 53533
rect 17681 53567 17739 53573
rect 17681 53533 17693 53567
rect 17727 53564 17739 53567
rect 18414 53564 18420 53576
rect 17727 53536 18420 53564
rect 17727 53533 17739 53536
rect 17681 53527 17739 53533
rect 10778 53496 10784 53508
rect 6886 53468 10784 53496
rect 10778 53456 10784 53468
rect 10836 53456 10842 53508
rect 15856 53428 15884 53527
rect 18414 53524 18420 53536
rect 18472 53524 18478 53576
rect 20165 53567 20223 53573
rect 20165 53533 20177 53567
rect 20211 53533 20223 53567
rect 20165 53527 20223 53533
rect 22005 53567 22063 53573
rect 22005 53533 22017 53567
rect 22051 53564 22063 53567
rect 22830 53564 22836 53576
rect 22051 53536 22836 53564
rect 22051 53533 22063 53536
rect 22005 53527 22063 53533
rect 20180 53496 20208 53527
rect 22830 53524 22836 53536
rect 22888 53524 22894 53576
rect 23290 53524 23296 53576
rect 23348 53564 23354 53576
rect 23845 53567 23903 53573
rect 23845 53564 23857 53567
rect 23348 53536 23857 53564
rect 23348 53524 23354 53536
rect 23845 53533 23857 53536
rect 23891 53533 23903 53567
rect 23845 53527 23903 53533
rect 23934 53524 23940 53576
rect 23992 53564 23998 53576
rect 24673 53567 24731 53573
rect 24673 53564 24685 53567
rect 23992 53536 24685 53564
rect 23992 53524 23998 53536
rect 24673 53533 24685 53536
rect 24719 53533 24731 53567
rect 24673 53527 24731 53533
rect 29086 53524 29092 53576
rect 29144 53564 29150 53576
rect 29917 53567 29975 53573
rect 29917 53564 29929 53567
rect 29144 53536 29929 53564
rect 29144 53524 29150 53536
rect 29917 53533 29929 53536
rect 29963 53533 29975 53567
rect 29917 53527 29975 53533
rect 32030 53524 32036 53576
rect 32088 53564 32094 53576
rect 32309 53567 32367 53573
rect 32309 53564 32321 53567
rect 32088 53536 32321 53564
rect 32088 53524 32094 53536
rect 32309 53533 32321 53536
rect 32355 53533 32367 53567
rect 32309 53527 32367 53533
rect 34974 53524 34980 53576
rect 35032 53564 35038 53576
rect 35253 53567 35311 53573
rect 35253 53564 35265 53567
rect 35032 53536 35265 53564
rect 35032 53524 35038 53536
rect 35253 53533 35265 53536
rect 35299 53533 35311 53567
rect 35253 53527 35311 53533
rect 37826 53524 37832 53576
rect 37884 53564 37890 53576
rect 38197 53567 38255 53573
rect 38197 53564 38209 53567
rect 37884 53536 38209 53564
rect 37884 53524 37890 53536
rect 38197 53533 38209 53536
rect 38243 53533 38255 53567
rect 38197 53527 38255 53533
rect 41598 53524 41604 53576
rect 41656 53564 41662 53576
rect 41877 53567 41935 53573
rect 41877 53564 41889 53567
rect 41656 53536 41889 53564
rect 41656 53524 41662 53536
rect 41877 53533 41889 53536
rect 41923 53533 41935 53567
rect 41877 53527 41935 53533
rect 46106 53524 46112 53576
rect 46164 53564 46170 53576
rect 46845 53567 46903 53573
rect 46845 53564 46857 53567
rect 46164 53536 46857 53564
rect 46164 53524 46170 53536
rect 46845 53533 46857 53536
rect 46891 53533 46903 53567
rect 46845 53527 46903 53533
rect 48958 53524 48964 53576
rect 49016 53564 49022 53576
rect 49237 53567 49295 53573
rect 49237 53564 49249 53567
rect 49016 53536 49249 53564
rect 49016 53524 49022 53536
rect 49237 53533 49249 53536
rect 49283 53533 49295 53567
rect 49237 53527 49295 53533
rect 22186 53496 22192 53508
rect 20180 53468 22192 53496
rect 22186 53456 22192 53468
rect 22244 53456 22250 53508
rect 24857 53499 24915 53505
rect 24857 53465 24869 53499
rect 24903 53496 24915 53499
rect 24946 53496 24952 53508
rect 24903 53468 24952 53496
rect 24903 53465 24915 53468
rect 24857 53459 24915 53465
rect 24946 53456 24952 53468
rect 25004 53456 25010 53508
rect 20438 53428 20444 53440
rect 15856 53400 20444 53428
rect 20438 53388 20444 53400
rect 20496 53388 20502 53440
rect 29730 53388 29736 53440
rect 29788 53388 29794 53440
rect 32122 53388 32128 53440
rect 32180 53388 32186 53440
rect 35069 53431 35127 53437
rect 35069 53397 35081 53431
rect 35115 53428 35127 53431
rect 35342 53428 35348 53440
rect 35115 53400 35348 53428
rect 35115 53397 35127 53400
rect 35069 53391 35127 53397
rect 35342 53388 35348 53400
rect 35400 53388 35406 53440
rect 36630 53388 36636 53440
rect 36688 53428 36694 53440
rect 38013 53431 38071 53437
rect 38013 53428 38025 53431
rect 36688 53400 38025 53428
rect 36688 53388 36694 53400
rect 38013 53397 38025 53400
rect 38059 53397 38071 53431
rect 38013 53391 38071 53397
rect 40678 53388 40684 53440
rect 40736 53428 40742 53440
rect 41693 53431 41751 53437
rect 41693 53428 41705 53431
rect 40736 53400 41705 53428
rect 40736 53388 40742 53400
rect 41693 53397 41705 53400
rect 41739 53397 41751 53431
rect 41693 53391 41751 53397
rect 48774 53388 48780 53440
rect 48832 53428 48838 53440
rect 49053 53431 49111 53437
rect 49053 53428 49065 53431
rect 48832 53400 49065 53428
rect 48832 53388 48838 53400
rect 49053 53397 49065 53400
rect 49099 53397 49111 53431
rect 49053 53391 49111 53397
rect 1104 53338 49864 53360
rect 1104 53286 7950 53338
rect 8002 53286 8014 53338
rect 8066 53286 8078 53338
rect 8130 53286 8142 53338
rect 8194 53286 8206 53338
rect 8258 53286 17950 53338
rect 18002 53286 18014 53338
rect 18066 53286 18078 53338
rect 18130 53286 18142 53338
rect 18194 53286 18206 53338
rect 18258 53286 27950 53338
rect 28002 53286 28014 53338
rect 28066 53286 28078 53338
rect 28130 53286 28142 53338
rect 28194 53286 28206 53338
rect 28258 53286 37950 53338
rect 38002 53286 38014 53338
rect 38066 53286 38078 53338
rect 38130 53286 38142 53338
rect 38194 53286 38206 53338
rect 38258 53286 47950 53338
rect 48002 53286 48014 53338
rect 48066 53286 48078 53338
rect 48130 53286 48142 53338
rect 48194 53286 48206 53338
rect 48258 53286 49864 53338
rect 1104 53264 49864 53286
rect 46106 53184 46112 53236
rect 46164 53184 46170 53236
rect 46845 53227 46903 53233
rect 46845 53193 46857 53227
rect 46891 53224 46903 53227
rect 47026 53224 47032 53236
rect 46891 53196 47032 53224
rect 46891 53193 46903 53196
rect 46845 53187 46903 53193
rect 47026 53184 47032 53196
rect 47084 53184 47090 53236
rect 6270 53156 6276 53168
rect 2884 53128 6276 53156
rect 934 53048 940 53100
rect 992 53088 998 53100
rect 2884 53097 2912 53128
rect 6270 53116 6276 53128
rect 6328 53116 6334 53168
rect 9858 53156 9864 53168
rect 6886 53128 9864 53156
rect 1673 53091 1731 53097
rect 1673 53088 1685 53091
rect 992 53060 1685 53088
rect 992 53048 998 53060
rect 1673 53057 1685 53060
rect 1719 53057 1731 53091
rect 1673 53051 1731 53057
rect 2869 53091 2927 53097
rect 2869 53057 2881 53091
rect 2915 53057 2927 53091
rect 2869 53051 2927 53057
rect 4801 53091 4859 53097
rect 4801 53057 4813 53091
rect 4847 53088 4859 53091
rect 6886 53088 6914 53128
rect 9858 53116 9864 53128
rect 9916 53116 9922 53168
rect 16942 53156 16948 53168
rect 13188 53128 16948 53156
rect 4847 53060 6914 53088
rect 8021 53091 8079 53097
rect 4847 53057 4859 53060
rect 4801 53051 4859 53057
rect 8021 53057 8033 53091
rect 8067 53088 8079 53091
rect 8067 53060 9720 53088
rect 8067 53057 8079 53060
rect 8021 53051 8079 53057
rect 2590 52980 2596 53032
rect 2648 53020 2654 53032
rect 3145 53023 3203 53029
rect 3145 53020 3157 53023
rect 2648 52992 3157 53020
rect 2648 52980 2654 52992
rect 3145 52989 3157 52992
rect 3191 52989 3203 53023
rect 3145 52983 3203 52989
rect 4890 52980 4896 53032
rect 4948 53020 4954 53032
rect 5077 53023 5135 53029
rect 5077 53020 5089 53023
rect 4948 52992 5089 53020
rect 4948 52980 4954 52992
rect 5077 52989 5089 52992
rect 5123 52989 5135 53023
rect 5077 52983 5135 52989
rect 7742 52980 7748 53032
rect 7800 53020 7806 53032
rect 8297 53023 8355 53029
rect 8297 53020 8309 53023
rect 7800 52992 8309 53020
rect 7800 52980 7806 52992
rect 8297 52989 8309 52992
rect 8343 52989 8355 53023
rect 8297 52983 8355 52989
rect 9692 52952 9720 53060
rect 9766 53048 9772 53100
rect 9824 53048 9830 53100
rect 13188 53097 13216 53128
rect 16942 53116 16948 53128
rect 17000 53116 17006 53168
rect 21266 53156 21272 53168
rect 17604 53128 21272 53156
rect 13173 53091 13231 53097
rect 13173 53057 13185 53091
rect 13219 53057 13231 53091
rect 13173 53051 13231 53057
rect 15013 53091 15071 53097
rect 15013 53057 15025 53091
rect 15059 53088 15071 53091
rect 15194 53088 15200 53100
rect 15059 53060 15200 53088
rect 15059 53057 15071 53060
rect 15013 53051 15071 53057
rect 15194 53048 15200 53060
rect 15252 53048 15258 53100
rect 17604 53097 17632 53128
rect 21266 53116 21272 53128
rect 21324 53116 21330 53168
rect 49145 53159 49203 53165
rect 49145 53125 49157 53159
rect 49191 53156 49203 53159
rect 49694 53156 49700 53168
rect 49191 53128 49700 53156
rect 49191 53125 49203 53128
rect 49145 53119 49203 53125
rect 49694 53116 49700 53128
rect 49752 53116 49758 53168
rect 17589 53091 17647 53097
rect 17589 53057 17601 53091
rect 17635 53057 17647 53091
rect 17589 53051 17647 53057
rect 19610 53048 19616 53100
rect 19668 53048 19674 53100
rect 46293 53091 46351 53097
rect 46293 53057 46305 53091
rect 46339 53088 46351 53091
rect 46934 53088 46940 53100
rect 46339 53060 46940 53088
rect 46339 53057 46351 53060
rect 46293 53051 46351 53057
rect 46934 53048 46940 53060
rect 46992 53088 46998 53100
rect 47029 53091 47087 53097
rect 47029 53088 47041 53091
rect 46992 53060 47041 53088
rect 46992 53048 46998 53060
rect 47029 53057 47041 53060
rect 47075 53057 47087 53091
rect 47029 53051 47087 53057
rect 48133 53091 48191 53097
rect 48133 53057 48145 53091
rect 48179 53088 48191 53091
rect 48314 53088 48320 53100
rect 48179 53060 48320 53088
rect 48179 53057 48191 53060
rect 48133 53051 48191 53057
rect 48314 53048 48320 53060
rect 48372 53048 48378 53100
rect 9950 52980 9956 53032
rect 10008 53020 10014 53032
rect 10229 53023 10287 53029
rect 10229 53020 10241 53023
rect 10008 52992 10241 53020
rect 10008 52980 10014 52992
rect 10229 52989 10241 52992
rect 10275 52989 10287 53023
rect 10229 52983 10287 52989
rect 12802 52980 12808 53032
rect 12860 53020 12866 53032
rect 13449 53023 13507 53029
rect 13449 53020 13461 53023
rect 12860 52992 13461 53020
rect 12860 52980 12866 52992
rect 13449 52989 13461 52992
rect 13495 52989 13507 53023
rect 13449 52983 13507 52989
rect 15102 52980 15108 53032
rect 15160 53020 15166 53032
rect 15381 53023 15439 53029
rect 15381 53020 15393 53023
rect 15160 52992 15393 53020
rect 15160 52980 15166 52992
rect 15381 52989 15393 52992
rect 15427 52989 15439 53023
rect 15381 52983 15439 52989
rect 17310 52980 17316 53032
rect 17368 53020 17374 53032
rect 17865 53023 17923 53029
rect 17865 53020 17877 53023
rect 17368 52992 17877 53020
rect 17368 52980 17374 52992
rect 17865 52989 17877 52992
rect 17911 52989 17923 53023
rect 17865 52983 17923 52989
rect 19518 52980 19524 53032
rect 19576 53020 19582 53032
rect 20073 53023 20131 53029
rect 20073 53020 20085 53023
rect 19576 52992 20085 53020
rect 19576 52980 19582 52992
rect 20073 52989 20085 52992
rect 20119 52989 20131 53023
rect 20073 52983 20131 52989
rect 12434 52952 12440 52964
rect 9692 52924 12440 52952
rect 12434 52912 12440 52924
rect 12492 52912 12498 52964
rect 1670 52844 1676 52896
rect 1728 52884 1734 52896
rect 1765 52887 1823 52893
rect 1765 52884 1777 52887
rect 1728 52856 1777 52884
rect 1728 52844 1734 52856
rect 1765 52853 1777 52856
rect 1811 52853 1823 52887
rect 1765 52847 1823 52853
rect 1104 52794 49864 52816
rect 1104 52742 2950 52794
rect 3002 52742 3014 52794
rect 3066 52742 3078 52794
rect 3130 52742 3142 52794
rect 3194 52742 3206 52794
rect 3258 52742 12950 52794
rect 13002 52742 13014 52794
rect 13066 52742 13078 52794
rect 13130 52742 13142 52794
rect 13194 52742 13206 52794
rect 13258 52742 22950 52794
rect 23002 52742 23014 52794
rect 23066 52742 23078 52794
rect 23130 52742 23142 52794
rect 23194 52742 23206 52794
rect 23258 52742 32950 52794
rect 33002 52742 33014 52794
rect 33066 52742 33078 52794
rect 33130 52742 33142 52794
rect 33194 52742 33206 52794
rect 33258 52742 42950 52794
rect 43002 52742 43014 52794
rect 43066 52742 43078 52794
rect 43130 52742 43142 52794
rect 43194 52742 43206 52794
rect 43258 52742 49864 52794
rect 1104 52720 49864 52742
rect 5810 52612 5816 52624
rect 3712 52584 5816 52612
rect 1118 52504 1124 52556
rect 1176 52544 1182 52556
rect 2041 52547 2099 52553
rect 2041 52544 2053 52547
rect 1176 52516 2053 52544
rect 1176 52504 1182 52516
rect 2041 52513 2053 52516
rect 2087 52513 2099 52547
rect 2041 52507 2099 52513
rect 1765 52479 1823 52485
rect 1765 52445 1777 52479
rect 1811 52476 1823 52479
rect 3712 52476 3740 52584
rect 5810 52572 5816 52584
rect 5868 52572 5874 52624
rect 9214 52572 9220 52624
rect 9272 52572 9278 52624
rect 4062 52504 4068 52556
rect 4120 52544 4126 52556
rect 4617 52547 4675 52553
rect 4617 52544 4629 52547
rect 4120 52516 4629 52544
rect 4120 52504 4126 52516
rect 4617 52513 4629 52516
rect 4663 52513 4675 52547
rect 9232 52544 9260 52572
rect 9769 52547 9827 52553
rect 9769 52544 9781 52547
rect 9232 52516 9781 52544
rect 4617 52507 4675 52513
rect 9769 52513 9781 52516
rect 9815 52513 9827 52547
rect 9769 52507 9827 52513
rect 14366 52504 14372 52556
rect 14424 52544 14430 52556
rect 14921 52547 14979 52553
rect 14921 52544 14933 52547
rect 14424 52516 14933 52544
rect 14424 52504 14430 52516
rect 14921 52513 14933 52516
rect 14967 52513 14979 52547
rect 14921 52507 14979 52513
rect 1811 52448 3740 52476
rect 4341 52479 4399 52485
rect 1811 52445 1823 52448
rect 1765 52439 1823 52445
rect 4341 52445 4353 52479
rect 4387 52476 4399 52479
rect 9214 52476 9220 52488
rect 4387 52448 9220 52476
rect 4387 52445 4399 52448
rect 4341 52439 4399 52445
rect 9214 52436 9220 52448
rect 9272 52436 9278 52488
rect 9493 52479 9551 52485
rect 9493 52445 9505 52479
rect 9539 52476 9551 52479
rect 14458 52476 14464 52488
rect 9539 52448 14464 52476
rect 9539 52445 9551 52448
rect 9493 52439 9551 52445
rect 14458 52436 14464 52448
rect 14516 52436 14522 52488
rect 14645 52479 14703 52485
rect 14645 52445 14657 52479
rect 14691 52476 14703 52479
rect 19150 52476 19156 52488
rect 14691 52448 19156 52476
rect 14691 52445 14703 52448
rect 14645 52439 14703 52445
rect 19150 52436 19156 52448
rect 19208 52436 19214 52488
rect 49326 52436 49332 52488
rect 49384 52436 49390 52488
rect 49142 52300 49148 52352
rect 49200 52300 49206 52352
rect 1104 52250 49864 52272
rect 1104 52198 7950 52250
rect 8002 52198 8014 52250
rect 8066 52198 8078 52250
rect 8130 52198 8142 52250
rect 8194 52198 8206 52250
rect 8258 52198 17950 52250
rect 18002 52198 18014 52250
rect 18066 52198 18078 52250
rect 18130 52198 18142 52250
rect 18194 52198 18206 52250
rect 18258 52198 27950 52250
rect 28002 52198 28014 52250
rect 28066 52198 28078 52250
rect 28130 52198 28142 52250
rect 28194 52198 28206 52250
rect 28258 52198 37950 52250
rect 38002 52198 38014 52250
rect 38066 52198 38078 52250
rect 38130 52198 38142 52250
rect 38194 52198 38206 52250
rect 38258 52198 47950 52250
rect 48002 52198 48014 52250
rect 48066 52198 48078 52250
rect 48130 52198 48142 52250
rect 48194 52198 48206 52250
rect 48258 52198 49864 52250
rect 1104 52176 49864 52198
rect 22738 52096 22744 52148
rect 22796 52136 22802 52148
rect 23569 52139 23627 52145
rect 23569 52136 23581 52139
rect 22796 52108 23581 52136
rect 22796 52096 22802 52108
rect 23569 52105 23581 52108
rect 23615 52105 23627 52139
rect 23569 52099 23627 52105
rect 2777 52071 2835 52077
rect 2777 52037 2789 52071
rect 2823 52068 2835 52071
rect 2866 52068 2872 52080
rect 2823 52040 2872 52068
rect 2823 52037 2835 52040
rect 2777 52031 2835 52037
rect 2866 52028 2872 52040
rect 2924 52028 2930 52080
rect 1578 51960 1584 52012
rect 1636 51960 1642 52012
rect 23750 51960 23756 52012
rect 23808 51960 23814 52012
rect 49050 51960 49056 52012
rect 49108 51960 49114 52012
rect 38378 51756 38384 51808
rect 38436 51796 38442 51808
rect 49237 51799 49295 51805
rect 49237 51796 49249 51799
rect 38436 51768 49249 51796
rect 38436 51756 38442 51768
rect 49237 51765 49249 51768
rect 49283 51765 49295 51799
rect 49237 51759 49295 51765
rect 1104 51706 49864 51728
rect 1104 51654 2950 51706
rect 3002 51654 3014 51706
rect 3066 51654 3078 51706
rect 3130 51654 3142 51706
rect 3194 51654 3206 51706
rect 3258 51654 12950 51706
rect 13002 51654 13014 51706
rect 13066 51654 13078 51706
rect 13130 51654 13142 51706
rect 13194 51654 13206 51706
rect 13258 51654 22950 51706
rect 23002 51654 23014 51706
rect 23066 51654 23078 51706
rect 23130 51654 23142 51706
rect 23194 51654 23206 51706
rect 23258 51654 32950 51706
rect 33002 51654 33014 51706
rect 33066 51654 33078 51706
rect 33130 51654 33142 51706
rect 33194 51654 33206 51706
rect 33258 51654 42950 51706
rect 43002 51654 43014 51706
rect 43066 51654 43078 51706
rect 43130 51654 43142 51706
rect 43194 51654 43206 51706
rect 43258 51654 49864 51706
rect 1104 51632 49864 51654
rect 10042 51552 10048 51604
rect 10100 51592 10106 51604
rect 13081 51595 13139 51601
rect 13081 51592 13093 51595
rect 10100 51564 13093 51592
rect 10100 51552 10106 51564
rect 13081 51561 13093 51564
rect 13127 51561 13139 51595
rect 13081 51555 13139 51561
rect 14458 51552 14464 51604
rect 14516 51552 14522 51604
rect 22830 51552 22836 51604
rect 22888 51592 22894 51604
rect 24673 51595 24731 51601
rect 24673 51592 24685 51595
rect 22888 51564 24685 51592
rect 22888 51552 22894 51564
rect 24673 51561 24685 51564
rect 24719 51561 24731 51595
rect 24673 51555 24731 51561
rect 24857 51391 24915 51397
rect 24857 51357 24869 51391
rect 24903 51388 24915 51391
rect 26694 51388 26700 51400
rect 24903 51360 26700 51388
rect 24903 51357 24915 51360
rect 24857 51351 24915 51357
rect 26694 51348 26700 51360
rect 26752 51348 26758 51400
rect 49050 51348 49056 51400
rect 49108 51348 49114 51400
rect 12989 51323 13047 51329
rect 12989 51289 13001 51323
rect 13035 51320 13047 51323
rect 14274 51320 14280 51332
rect 13035 51292 14280 51320
rect 13035 51289 13047 51292
rect 12989 51283 13047 51289
rect 14274 51280 14280 51292
rect 14332 51280 14338 51332
rect 14369 51323 14427 51329
rect 14369 51289 14381 51323
rect 14415 51320 14427 51323
rect 15930 51320 15936 51332
rect 14415 51292 15936 51320
rect 14415 51289 14427 51292
rect 14369 51283 14427 51289
rect 15930 51280 15936 51292
rect 15988 51280 15994 51332
rect 49237 51255 49295 51261
rect 49237 51221 49249 51255
rect 49283 51252 49295 51255
rect 49326 51252 49332 51264
rect 49283 51224 49332 51252
rect 49283 51221 49295 51224
rect 49237 51215 49295 51221
rect 49326 51212 49332 51224
rect 49384 51212 49390 51264
rect 1104 51162 49864 51184
rect 1104 51110 7950 51162
rect 8002 51110 8014 51162
rect 8066 51110 8078 51162
rect 8130 51110 8142 51162
rect 8194 51110 8206 51162
rect 8258 51110 17950 51162
rect 18002 51110 18014 51162
rect 18066 51110 18078 51162
rect 18130 51110 18142 51162
rect 18194 51110 18206 51162
rect 18258 51110 27950 51162
rect 28002 51110 28014 51162
rect 28066 51110 28078 51162
rect 28130 51110 28142 51162
rect 28194 51110 28206 51162
rect 28258 51110 37950 51162
rect 38002 51110 38014 51162
rect 38066 51110 38078 51162
rect 38130 51110 38142 51162
rect 38194 51110 38206 51162
rect 38258 51110 47950 51162
rect 48002 51110 48014 51162
rect 48066 51110 48078 51162
rect 48130 51110 48142 51162
rect 48194 51110 48206 51162
rect 48258 51110 49864 51162
rect 1104 51088 49864 51110
rect 22186 51008 22192 51060
rect 22244 51008 22250 51060
rect 20346 50940 20352 50992
rect 20404 50980 20410 50992
rect 23293 50983 23351 50989
rect 23293 50980 23305 50983
rect 20404 50952 23305 50980
rect 20404 50940 20410 50952
rect 23293 50949 23305 50952
rect 23339 50949 23351 50983
rect 23293 50943 23351 50949
rect 934 50872 940 50924
rect 992 50912 998 50924
rect 1673 50915 1731 50921
rect 1673 50912 1685 50915
rect 992 50884 1685 50912
rect 992 50872 998 50884
rect 1673 50881 1685 50884
rect 1719 50881 1731 50915
rect 1673 50875 1731 50881
rect 22097 50915 22155 50921
rect 22097 50881 22109 50915
rect 22143 50912 22155 50915
rect 22738 50912 22744 50924
rect 22143 50884 22744 50912
rect 22143 50881 22155 50884
rect 22097 50875 22155 50881
rect 22738 50872 22744 50884
rect 22796 50872 22802 50924
rect 23109 50915 23167 50921
rect 23109 50881 23121 50915
rect 23155 50912 23167 50915
rect 24118 50912 24124 50924
rect 23155 50884 24124 50912
rect 23155 50881 23167 50884
rect 23109 50875 23167 50881
rect 24118 50872 24124 50884
rect 24176 50872 24182 50924
rect 48958 50872 48964 50924
rect 49016 50872 49022 50924
rect 1857 50779 1915 50785
rect 1857 50745 1869 50779
rect 1903 50776 1915 50779
rect 1946 50776 1952 50788
rect 1903 50748 1952 50776
rect 1903 50745 1915 50748
rect 1857 50739 1915 50745
rect 1946 50736 1952 50748
rect 2004 50736 2010 50788
rect 38838 50668 38844 50720
rect 38896 50708 38902 50720
rect 49053 50711 49111 50717
rect 49053 50708 49065 50711
rect 38896 50680 49065 50708
rect 38896 50668 38902 50680
rect 49053 50677 49065 50680
rect 49099 50677 49111 50711
rect 49053 50671 49111 50677
rect 1104 50618 49864 50640
rect 1104 50566 2950 50618
rect 3002 50566 3014 50618
rect 3066 50566 3078 50618
rect 3130 50566 3142 50618
rect 3194 50566 3206 50618
rect 3258 50566 12950 50618
rect 13002 50566 13014 50618
rect 13066 50566 13078 50618
rect 13130 50566 13142 50618
rect 13194 50566 13206 50618
rect 13258 50566 22950 50618
rect 23002 50566 23014 50618
rect 23066 50566 23078 50618
rect 23130 50566 23142 50618
rect 23194 50566 23206 50618
rect 23258 50566 32950 50618
rect 33002 50566 33014 50618
rect 33066 50566 33078 50618
rect 33130 50566 33142 50618
rect 33194 50566 33206 50618
rect 33258 50566 42950 50618
rect 43002 50566 43014 50618
rect 43066 50566 43078 50618
rect 43130 50566 43142 50618
rect 43194 50566 43206 50618
rect 43258 50566 49864 50618
rect 1104 50544 49864 50566
rect 17678 50464 17684 50516
rect 17736 50504 17742 50516
rect 20257 50507 20315 50513
rect 20257 50504 20269 50507
rect 17736 50476 20269 50504
rect 17736 50464 17742 50476
rect 20257 50473 20269 50476
rect 20303 50473 20315 50507
rect 20257 50467 20315 50473
rect 49050 50260 49056 50312
rect 49108 50260 49114 50312
rect 20165 50235 20223 50241
rect 20165 50201 20177 50235
rect 20211 50232 20223 50235
rect 22278 50232 22284 50244
rect 20211 50204 22284 50232
rect 20211 50201 20223 50204
rect 20165 50195 20223 50201
rect 22278 50192 22284 50204
rect 22336 50192 22342 50244
rect 48866 50124 48872 50176
rect 48924 50164 48930 50176
rect 49237 50167 49295 50173
rect 49237 50164 49249 50167
rect 48924 50136 49249 50164
rect 48924 50124 48930 50136
rect 49237 50133 49249 50136
rect 49283 50133 49295 50167
rect 49237 50127 49295 50133
rect 1104 50074 49864 50096
rect 1104 50022 7950 50074
rect 8002 50022 8014 50074
rect 8066 50022 8078 50074
rect 8130 50022 8142 50074
rect 8194 50022 8206 50074
rect 8258 50022 17950 50074
rect 18002 50022 18014 50074
rect 18066 50022 18078 50074
rect 18130 50022 18142 50074
rect 18194 50022 18206 50074
rect 18258 50022 27950 50074
rect 28002 50022 28014 50074
rect 28066 50022 28078 50074
rect 28130 50022 28142 50074
rect 28194 50022 28206 50074
rect 28258 50022 37950 50074
rect 38002 50022 38014 50074
rect 38066 50022 38078 50074
rect 38130 50022 38142 50074
rect 38194 50022 38206 50074
rect 38258 50022 47950 50074
rect 48002 50022 48014 50074
rect 48066 50022 48078 50074
rect 48130 50022 48142 50074
rect 48194 50022 48206 50074
rect 48258 50022 49864 50074
rect 1104 50000 49864 50022
rect 12342 49920 12348 49972
rect 12400 49920 12406 49972
rect 14734 49920 14740 49972
rect 14792 49920 14798 49972
rect 46198 49920 46204 49972
rect 46256 49960 46262 49972
rect 49237 49963 49295 49969
rect 49237 49960 49249 49963
rect 46256 49932 49249 49960
rect 46256 49920 46262 49932
rect 49237 49929 49249 49932
rect 49283 49929 49295 49963
rect 49237 49923 49295 49929
rect 12253 49895 12311 49901
rect 12253 49861 12265 49895
rect 12299 49892 12311 49895
rect 20898 49892 20904 49904
rect 12299 49864 20904 49892
rect 12299 49861 12311 49864
rect 12253 49855 12311 49861
rect 20898 49852 20904 49864
rect 20956 49852 20962 49904
rect 14645 49827 14703 49833
rect 14645 49793 14657 49827
rect 14691 49824 14703 49827
rect 16850 49824 16856 49836
rect 14691 49796 16856 49824
rect 14691 49793 14703 49796
rect 14645 49787 14703 49793
rect 16850 49784 16856 49796
rect 16908 49784 16914 49836
rect 49053 49827 49111 49833
rect 49053 49793 49065 49827
rect 49099 49824 49111 49827
rect 49142 49824 49148 49836
rect 49099 49796 49148 49824
rect 49099 49793 49111 49796
rect 49053 49787 49111 49793
rect 49142 49784 49148 49796
rect 49200 49784 49206 49836
rect 1104 49530 49864 49552
rect 1104 49478 2950 49530
rect 3002 49478 3014 49530
rect 3066 49478 3078 49530
rect 3130 49478 3142 49530
rect 3194 49478 3206 49530
rect 3258 49478 12950 49530
rect 13002 49478 13014 49530
rect 13066 49478 13078 49530
rect 13130 49478 13142 49530
rect 13194 49478 13206 49530
rect 13258 49478 22950 49530
rect 23002 49478 23014 49530
rect 23066 49478 23078 49530
rect 23130 49478 23142 49530
rect 23194 49478 23206 49530
rect 23258 49478 32950 49530
rect 33002 49478 33014 49530
rect 33066 49478 33078 49530
rect 33130 49478 33142 49530
rect 33194 49478 33206 49530
rect 33258 49478 42950 49530
rect 43002 49478 43014 49530
rect 43066 49478 43078 49530
rect 43130 49478 43142 49530
rect 43194 49478 43206 49530
rect 43258 49478 49864 49530
rect 1104 49456 49864 49478
rect 15194 49376 15200 49428
rect 15252 49416 15258 49428
rect 18049 49419 18107 49425
rect 18049 49416 18061 49419
rect 15252 49388 18061 49416
rect 15252 49376 15258 49388
rect 18049 49385 18061 49388
rect 18095 49385 18107 49419
rect 18049 49379 18107 49385
rect 18414 49376 18420 49428
rect 18472 49416 18478 49428
rect 20349 49419 20407 49425
rect 20349 49416 20361 49419
rect 18472 49388 20361 49416
rect 18472 49376 18478 49388
rect 20349 49385 20361 49388
rect 20395 49385 20407 49419
rect 20349 49379 20407 49385
rect 17957 49215 18015 49221
rect 17957 49181 17969 49215
rect 18003 49212 18015 49215
rect 20622 49212 20628 49224
rect 18003 49184 20628 49212
rect 18003 49181 18015 49184
rect 17957 49175 18015 49181
rect 20622 49172 20628 49184
rect 20680 49172 20686 49224
rect 49053 49215 49111 49221
rect 49053 49181 49065 49215
rect 49099 49212 49111 49215
rect 49234 49212 49240 49224
rect 49099 49184 49240 49212
rect 49099 49181 49111 49184
rect 49053 49175 49111 49181
rect 49234 49172 49240 49184
rect 49292 49172 49298 49224
rect 20257 49147 20315 49153
rect 20257 49113 20269 49147
rect 20303 49144 20315 49147
rect 22186 49144 22192 49156
rect 20303 49116 22192 49144
rect 20303 49113 20315 49116
rect 20257 49107 20315 49113
rect 22186 49104 22192 49116
rect 22244 49104 22250 49156
rect 38654 49036 38660 49088
rect 38712 49076 38718 49088
rect 49237 49079 49295 49085
rect 49237 49076 49249 49079
rect 38712 49048 49249 49076
rect 38712 49036 38718 49048
rect 49237 49045 49249 49048
rect 49283 49045 49295 49079
rect 49237 49039 49295 49045
rect 1104 48986 49864 49008
rect 1104 48934 7950 48986
rect 8002 48934 8014 48986
rect 8066 48934 8078 48986
rect 8130 48934 8142 48986
rect 8194 48934 8206 48986
rect 8258 48934 17950 48986
rect 18002 48934 18014 48986
rect 18066 48934 18078 48986
rect 18130 48934 18142 48986
rect 18194 48934 18206 48986
rect 18258 48934 27950 48986
rect 28002 48934 28014 48986
rect 28066 48934 28078 48986
rect 28130 48934 28142 48986
rect 28194 48934 28206 48986
rect 28258 48934 37950 48986
rect 38002 48934 38014 48986
rect 38066 48934 38078 48986
rect 38130 48934 38142 48986
rect 38194 48934 38206 48986
rect 38258 48934 47950 48986
rect 48002 48934 48014 48986
rect 48066 48934 48078 48986
rect 48130 48934 48142 48986
rect 48194 48934 48206 48986
rect 48258 48934 49864 48986
rect 1104 48912 49864 48934
rect 49050 48696 49056 48748
rect 49108 48696 49114 48748
rect 40770 48492 40776 48544
rect 40828 48532 40834 48544
rect 49237 48535 49295 48541
rect 49237 48532 49249 48535
rect 40828 48504 49249 48532
rect 40828 48492 40834 48504
rect 49237 48501 49249 48504
rect 49283 48501 49295 48535
rect 49237 48495 49295 48501
rect 1104 48442 49864 48464
rect 1104 48390 2950 48442
rect 3002 48390 3014 48442
rect 3066 48390 3078 48442
rect 3130 48390 3142 48442
rect 3194 48390 3206 48442
rect 3258 48390 12950 48442
rect 13002 48390 13014 48442
rect 13066 48390 13078 48442
rect 13130 48390 13142 48442
rect 13194 48390 13206 48442
rect 13258 48390 22950 48442
rect 23002 48390 23014 48442
rect 23066 48390 23078 48442
rect 23130 48390 23142 48442
rect 23194 48390 23206 48442
rect 23258 48390 32950 48442
rect 33002 48390 33014 48442
rect 33066 48390 33078 48442
rect 33130 48390 33142 48442
rect 33194 48390 33206 48442
rect 33258 48390 42950 48442
rect 43002 48390 43014 48442
rect 43066 48390 43078 48442
rect 43130 48390 43142 48442
rect 43194 48390 43206 48442
rect 43258 48390 49864 48442
rect 1104 48368 49864 48390
rect 46382 48220 46388 48272
rect 46440 48260 46446 48272
rect 47949 48263 48007 48269
rect 47949 48260 47961 48263
rect 46440 48232 47961 48260
rect 46440 48220 46446 48232
rect 47949 48229 47961 48232
rect 47995 48229 48007 48263
rect 47949 48223 48007 48229
rect 48314 48220 48320 48272
rect 48372 48260 48378 48272
rect 48869 48263 48927 48269
rect 48869 48260 48881 48263
rect 48372 48232 48881 48260
rect 48372 48220 48378 48232
rect 48869 48229 48881 48232
rect 48915 48229 48927 48263
rect 48869 48223 48927 48229
rect 10137 48195 10195 48201
rect 10137 48161 10149 48195
rect 10183 48192 10195 48195
rect 21082 48192 21088 48204
rect 10183 48164 21088 48192
rect 10183 48161 10195 48164
rect 10137 48155 10195 48161
rect 21082 48152 21088 48164
rect 21140 48152 21146 48204
rect 47762 48084 47768 48136
rect 47820 48124 47826 48136
rect 48133 48127 48191 48133
rect 48133 48124 48145 48127
rect 47820 48096 48145 48124
rect 47820 48084 47826 48096
rect 48133 48093 48145 48096
rect 48179 48124 48191 48127
rect 48685 48127 48743 48133
rect 48685 48124 48697 48127
rect 48179 48096 48697 48124
rect 48179 48093 48191 48096
rect 48133 48087 48191 48093
rect 48685 48093 48697 48096
rect 48731 48093 48743 48127
rect 48685 48087 48743 48093
rect 934 48016 940 48068
rect 992 48056 998 48068
rect 1673 48059 1731 48065
rect 1673 48056 1685 48059
rect 992 48028 1685 48056
rect 992 48016 998 48028
rect 1673 48025 1685 48028
rect 1719 48025 1731 48059
rect 1673 48019 1731 48025
rect 1854 48016 1860 48068
rect 1912 48016 1918 48068
rect 3970 48016 3976 48068
rect 4028 48056 4034 48068
rect 10413 48059 10471 48065
rect 10413 48056 10425 48059
rect 4028 48028 10425 48056
rect 4028 48016 4034 48028
rect 10413 48025 10425 48028
rect 10459 48025 10471 48059
rect 11974 48056 11980 48068
rect 11638 48028 11980 48056
rect 10413 48019 10471 48025
rect 11974 48016 11980 48028
rect 12032 48016 12038 48068
rect 12161 48059 12219 48065
rect 12161 48025 12173 48059
rect 12207 48056 12219 48059
rect 22094 48056 22100 48068
rect 12207 48028 22100 48056
rect 12207 48025 12219 48028
rect 12161 48019 12219 48025
rect 22094 48016 22100 48028
rect 22152 48016 22158 48068
rect 1104 47898 49864 47920
rect 1104 47846 7950 47898
rect 8002 47846 8014 47898
rect 8066 47846 8078 47898
rect 8130 47846 8142 47898
rect 8194 47846 8206 47898
rect 8258 47846 17950 47898
rect 18002 47846 18014 47898
rect 18066 47846 18078 47898
rect 18130 47846 18142 47898
rect 18194 47846 18206 47898
rect 18258 47846 27950 47898
rect 28002 47846 28014 47898
rect 28066 47846 28078 47898
rect 28130 47846 28142 47898
rect 28194 47846 28206 47898
rect 28258 47846 37950 47898
rect 38002 47846 38014 47898
rect 38066 47846 38078 47898
rect 38130 47846 38142 47898
rect 38194 47846 38206 47898
rect 38258 47846 47950 47898
rect 48002 47846 48014 47898
rect 48066 47846 48078 47898
rect 48130 47846 48142 47898
rect 48194 47846 48206 47898
rect 48258 47846 49864 47898
rect 1104 47824 49864 47846
rect 23750 47744 23756 47796
rect 23808 47784 23814 47796
rect 24673 47787 24731 47793
rect 24673 47784 24685 47787
rect 23808 47756 24685 47784
rect 23808 47744 23814 47756
rect 24673 47753 24685 47756
rect 24719 47753 24731 47787
rect 24673 47747 24731 47753
rect 24854 47608 24860 47660
rect 24912 47608 24918 47660
rect 49050 47608 49056 47660
rect 49108 47608 49114 47660
rect 41046 47404 41052 47456
rect 41104 47444 41110 47456
rect 49237 47447 49295 47453
rect 49237 47444 49249 47447
rect 41104 47416 49249 47444
rect 41104 47404 41110 47416
rect 49237 47413 49249 47416
rect 49283 47413 49295 47447
rect 49237 47407 49295 47413
rect 1104 47354 49864 47376
rect 1104 47302 2950 47354
rect 3002 47302 3014 47354
rect 3066 47302 3078 47354
rect 3130 47302 3142 47354
rect 3194 47302 3206 47354
rect 3258 47302 12950 47354
rect 13002 47302 13014 47354
rect 13066 47302 13078 47354
rect 13130 47302 13142 47354
rect 13194 47302 13206 47354
rect 13258 47302 22950 47354
rect 23002 47302 23014 47354
rect 23066 47302 23078 47354
rect 23130 47302 23142 47354
rect 23194 47302 23206 47354
rect 23258 47302 32950 47354
rect 33002 47302 33014 47354
rect 33066 47302 33078 47354
rect 33130 47302 33142 47354
rect 33194 47302 33206 47354
rect 33258 47302 42950 47354
rect 43002 47302 43014 47354
rect 43066 47302 43078 47354
rect 43130 47302 43142 47354
rect 43194 47302 43206 47354
rect 43258 47302 49864 47354
rect 1104 47280 49864 47302
rect 47854 47200 47860 47252
rect 47912 47240 47918 47252
rect 48225 47243 48283 47249
rect 48225 47240 48237 47243
rect 47912 47212 48237 47240
rect 47912 47200 47918 47212
rect 48225 47209 48237 47212
rect 48271 47209 48283 47243
rect 48225 47203 48283 47209
rect 48774 47200 48780 47252
rect 48832 47200 48838 47252
rect 48961 47039 49019 47045
rect 48961 47036 48973 47039
rect 48424 47008 48973 47036
rect 48424 46980 48452 47008
rect 48961 47005 48973 47008
rect 49007 47005 49019 47039
rect 48961 46999 49019 47005
rect 48133 46971 48191 46977
rect 48133 46937 48145 46971
rect 48179 46968 48191 46971
rect 48406 46968 48412 46980
rect 48179 46940 48412 46968
rect 48179 46937 48191 46940
rect 48133 46931 48191 46937
rect 48406 46928 48412 46940
rect 48464 46928 48470 46980
rect 1104 46810 49864 46832
rect 1104 46758 7950 46810
rect 8002 46758 8014 46810
rect 8066 46758 8078 46810
rect 8130 46758 8142 46810
rect 8194 46758 8206 46810
rect 8258 46758 17950 46810
rect 18002 46758 18014 46810
rect 18066 46758 18078 46810
rect 18130 46758 18142 46810
rect 18194 46758 18206 46810
rect 18258 46758 27950 46810
rect 28002 46758 28014 46810
rect 28066 46758 28078 46810
rect 28130 46758 28142 46810
rect 28194 46758 28206 46810
rect 28258 46758 37950 46810
rect 38002 46758 38014 46810
rect 38066 46758 38078 46810
rect 38130 46758 38142 46810
rect 38194 46758 38206 46810
rect 38258 46758 47950 46810
rect 48002 46758 48014 46810
rect 48066 46758 48078 46810
rect 48130 46758 48142 46810
rect 48194 46758 48206 46810
rect 48258 46758 49864 46810
rect 1104 46736 49864 46758
rect 49326 46520 49332 46572
rect 49384 46520 49390 46572
rect 48682 46316 48688 46368
rect 48740 46356 48746 46368
rect 49145 46359 49203 46365
rect 49145 46356 49157 46359
rect 48740 46328 49157 46356
rect 48740 46316 48746 46328
rect 49145 46325 49157 46328
rect 49191 46325 49203 46359
rect 49145 46319 49203 46325
rect 1104 46266 49864 46288
rect 1104 46214 2950 46266
rect 3002 46214 3014 46266
rect 3066 46214 3078 46266
rect 3130 46214 3142 46266
rect 3194 46214 3206 46266
rect 3258 46214 12950 46266
rect 13002 46214 13014 46266
rect 13066 46214 13078 46266
rect 13130 46214 13142 46266
rect 13194 46214 13206 46266
rect 13258 46214 22950 46266
rect 23002 46214 23014 46266
rect 23066 46214 23078 46266
rect 23130 46214 23142 46266
rect 23194 46214 23206 46266
rect 23258 46214 32950 46266
rect 33002 46214 33014 46266
rect 33066 46214 33078 46266
rect 33130 46214 33142 46266
rect 33194 46214 33206 46266
rect 33258 46214 42950 46266
rect 43002 46214 43014 46266
rect 43066 46214 43078 46266
rect 43130 46214 43142 46266
rect 43194 46214 43206 46266
rect 43258 46214 49864 46266
rect 1104 46192 49864 46214
rect 15930 46112 15936 46164
rect 15988 46152 15994 46164
rect 18417 46155 18475 46161
rect 18417 46152 18429 46155
rect 15988 46124 18429 46152
rect 15988 46112 15994 46124
rect 18417 46121 18429 46124
rect 18463 46121 18475 46155
rect 18417 46115 18475 46121
rect 26694 46112 26700 46164
rect 26752 46112 26758 46164
rect 18601 45951 18659 45957
rect 18601 45917 18613 45951
rect 18647 45948 18659 45951
rect 19705 45951 19763 45957
rect 18647 45920 19656 45948
rect 18647 45917 18659 45920
rect 18601 45911 18659 45917
rect 934 45840 940 45892
rect 992 45880 998 45892
rect 1673 45883 1731 45889
rect 1673 45880 1685 45883
rect 992 45852 1685 45880
rect 992 45840 998 45852
rect 1673 45849 1685 45852
rect 1719 45849 1731 45883
rect 1673 45843 1731 45849
rect 14274 45840 14280 45892
rect 14332 45880 14338 45892
rect 19628 45880 19656 45920
rect 19705 45917 19717 45951
rect 19751 45948 19763 45951
rect 22002 45948 22008 45960
rect 19751 45920 22008 45948
rect 19751 45917 19763 45920
rect 19705 45911 19763 45917
rect 22002 45908 22008 45920
rect 22060 45908 22066 45960
rect 26881 45951 26939 45957
rect 26881 45917 26893 45951
rect 26927 45948 26939 45951
rect 27706 45948 27712 45960
rect 26927 45920 27712 45948
rect 26927 45917 26939 45920
rect 26881 45911 26939 45917
rect 27706 45908 27712 45920
rect 27764 45908 27770 45960
rect 48133 45951 48191 45957
rect 48133 45917 48145 45951
rect 48179 45948 48191 45951
rect 48590 45948 48596 45960
rect 48179 45920 48596 45948
rect 48179 45917 48191 45920
rect 48133 45911 48191 45917
rect 48590 45908 48596 45920
rect 48648 45908 48654 45960
rect 20530 45880 20536 45892
rect 14332 45852 19564 45880
rect 19628 45852 20536 45880
rect 14332 45840 14338 45852
rect 1762 45772 1768 45824
rect 1820 45772 1826 45824
rect 19536 45821 19564 45852
rect 20530 45840 20536 45852
rect 20588 45840 20594 45892
rect 49142 45840 49148 45892
rect 49200 45840 49206 45892
rect 19521 45815 19579 45821
rect 19521 45781 19533 45815
rect 19567 45781 19579 45815
rect 19521 45775 19579 45781
rect 1104 45722 49864 45744
rect 1104 45670 7950 45722
rect 8002 45670 8014 45722
rect 8066 45670 8078 45722
rect 8130 45670 8142 45722
rect 8194 45670 8206 45722
rect 8258 45670 17950 45722
rect 18002 45670 18014 45722
rect 18066 45670 18078 45722
rect 18130 45670 18142 45722
rect 18194 45670 18206 45722
rect 18258 45670 27950 45722
rect 28002 45670 28014 45722
rect 28066 45670 28078 45722
rect 28130 45670 28142 45722
rect 28194 45670 28206 45722
rect 28258 45670 37950 45722
rect 38002 45670 38014 45722
rect 38066 45670 38078 45722
rect 38130 45670 38142 45722
rect 38194 45670 38206 45722
rect 38258 45670 47950 45722
rect 48002 45670 48014 45722
rect 48066 45670 48078 45722
rect 48130 45670 48142 45722
rect 48194 45670 48206 45722
rect 48258 45670 49864 45722
rect 1104 45648 49864 45670
rect 1762 45568 1768 45620
rect 1820 45608 1826 45620
rect 22462 45608 22468 45620
rect 1820 45580 22468 45608
rect 1820 45568 1826 45580
rect 22462 45568 22468 45580
rect 22520 45568 22526 45620
rect 48590 45568 48596 45620
rect 48648 45568 48654 45620
rect 10410 45500 10416 45552
rect 10468 45540 10474 45552
rect 15105 45543 15163 45549
rect 15105 45540 15117 45543
rect 10468 45512 15117 45540
rect 10468 45500 10474 45512
rect 15105 45509 15117 45512
rect 15151 45509 15163 45543
rect 15105 45503 15163 45509
rect 32122 45500 32128 45552
rect 32180 45540 32186 45552
rect 33873 45543 33931 45549
rect 33873 45540 33885 45543
rect 32180 45512 33885 45540
rect 32180 45500 32186 45512
rect 33873 45509 33885 45512
rect 33919 45509 33931 45543
rect 33873 45503 33931 45509
rect 33962 45500 33968 45552
rect 34020 45500 34026 45552
rect 46934 45500 46940 45552
rect 46992 45540 46998 45552
rect 46992 45512 48820 45540
rect 46992 45500 46998 45512
rect 14918 45432 14924 45484
rect 14976 45432 14982 45484
rect 29730 45432 29736 45484
rect 29788 45472 29794 45484
rect 32677 45475 32735 45481
rect 32677 45472 32689 45475
rect 29788 45444 32689 45472
rect 29788 45432 29794 45444
rect 32677 45441 32689 45444
rect 32723 45441 32735 45475
rect 32677 45435 32735 45441
rect 32769 45475 32827 45481
rect 32769 45441 32781 45475
rect 32815 45472 32827 45475
rect 33318 45472 33324 45484
rect 32815 45444 33324 45472
rect 32815 45441 32827 45444
rect 32769 45435 32827 45441
rect 33318 45432 33324 45444
rect 33376 45432 33382 45484
rect 47854 45432 47860 45484
rect 47912 45472 47918 45484
rect 48792 45481 48820 45512
rect 48133 45475 48191 45481
rect 48133 45472 48145 45475
rect 47912 45444 48145 45472
rect 47912 45432 47918 45444
rect 48133 45441 48145 45444
rect 48179 45441 48191 45475
rect 48133 45435 48191 45441
rect 48777 45475 48835 45481
rect 48777 45441 48789 45475
rect 48823 45441 48835 45475
rect 48777 45435 48835 45441
rect 32858 45364 32864 45416
rect 32916 45364 32922 45416
rect 34146 45364 34152 45416
rect 34204 45364 34210 45416
rect 47949 45339 48007 45345
rect 47949 45305 47961 45339
rect 47995 45336 48007 45339
rect 49050 45336 49056 45348
rect 47995 45308 49056 45336
rect 47995 45305 48007 45308
rect 47949 45299 48007 45305
rect 49050 45296 49056 45308
rect 49108 45296 49114 45348
rect 32309 45271 32367 45277
rect 32309 45237 32321 45271
rect 32355 45268 32367 45271
rect 32674 45268 32680 45280
rect 32355 45240 32680 45268
rect 32355 45237 32367 45240
rect 32309 45231 32367 45237
rect 32674 45228 32680 45240
rect 32732 45228 32738 45280
rect 33502 45228 33508 45280
rect 33560 45228 33566 45280
rect 1104 45178 49864 45200
rect 1104 45126 2950 45178
rect 3002 45126 3014 45178
rect 3066 45126 3078 45178
rect 3130 45126 3142 45178
rect 3194 45126 3206 45178
rect 3258 45126 12950 45178
rect 13002 45126 13014 45178
rect 13066 45126 13078 45178
rect 13130 45126 13142 45178
rect 13194 45126 13206 45178
rect 13258 45126 22950 45178
rect 23002 45126 23014 45178
rect 23066 45126 23078 45178
rect 23130 45126 23142 45178
rect 23194 45126 23206 45178
rect 23258 45126 32950 45178
rect 33002 45126 33014 45178
rect 33066 45126 33078 45178
rect 33130 45126 33142 45178
rect 33194 45126 33206 45178
rect 33258 45126 42950 45178
rect 43002 45126 43014 45178
rect 43066 45126 43078 45178
rect 43130 45126 43142 45178
rect 43194 45126 43206 45178
rect 43258 45126 49864 45178
rect 1104 45104 49864 45126
rect 22738 45024 22744 45076
rect 22796 45064 22802 45076
rect 22925 45067 22983 45073
rect 22925 45064 22937 45067
rect 22796 45036 22937 45064
rect 22796 45024 22802 45036
rect 22925 45033 22937 45036
rect 22971 45033 22983 45067
rect 22925 45027 22983 45033
rect 24118 45024 24124 45076
rect 24176 45064 24182 45076
rect 25041 45067 25099 45073
rect 25041 45064 25053 45067
rect 24176 45036 25053 45064
rect 24176 45024 24182 45036
rect 25041 45033 25053 45036
rect 25087 45033 25099 45067
rect 25041 45027 25099 45033
rect 35342 44888 35348 44940
rect 35400 44888 35406 44940
rect 35526 44888 35532 44940
rect 35584 44888 35590 44940
rect 48777 44931 48835 44937
rect 48777 44928 48789 44931
rect 45526 44900 48789 44928
rect 23109 44863 23167 44869
rect 23109 44829 23121 44863
rect 23155 44860 23167 44863
rect 24486 44860 24492 44872
rect 23155 44832 24492 44860
rect 23155 44829 23167 44832
rect 23109 44823 23167 44829
rect 24486 44820 24492 44832
rect 24544 44820 24550 44872
rect 25225 44863 25283 44869
rect 25225 44829 25237 44863
rect 25271 44860 25283 44863
rect 27154 44860 27160 44872
rect 25271 44832 27160 44860
rect 25271 44829 25283 44832
rect 25225 44823 25283 44829
rect 27154 44820 27160 44832
rect 27212 44820 27218 44872
rect 38562 44820 38568 44872
rect 38620 44860 38626 44872
rect 45526 44860 45554 44900
rect 48777 44897 48789 44900
rect 48823 44897 48835 44931
rect 48777 44891 48835 44897
rect 38620 44832 45554 44860
rect 38620 44820 38626 44832
rect 48498 44820 48504 44872
rect 48556 44820 48562 44872
rect 32398 44752 32404 44804
rect 32456 44792 32462 44804
rect 35066 44792 35072 44804
rect 32456 44764 35072 44792
rect 32456 44752 32462 44764
rect 35066 44752 35072 44764
rect 35124 44792 35130 44804
rect 35253 44795 35311 44801
rect 35253 44792 35265 44795
rect 35124 44764 35265 44792
rect 35124 44752 35130 44764
rect 35253 44761 35265 44764
rect 35299 44761 35311 44795
rect 35253 44755 35311 44761
rect 34882 44684 34888 44736
rect 34940 44684 34946 44736
rect 1104 44634 49864 44656
rect 1104 44582 7950 44634
rect 8002 44582 8014 44634
rect 8066 44582 8078 44634
rect 8130 44582 8142 44634
rect 8194 44582 8206 44634
rect 8258 44582 17950 44634
rect 18002 44582 18014 44634
rect 18066 44582 18078 44634
rect 18130 44582 18142 44634
rect 18194 44582 18206 44634
rect 18258 44582 27950 44634
rect 28002 44582 28014 44634
rect 28066 44582 28078 44634
rect 28130 44582 28142 44634
rect 28194 44582 28206 44634
rect 28258 44582 37950 44634
rect 38002 44582 38014 44634
rect 38066 44582 38078 44634
rect 38130 44582 38142 44634
rect 38194 44582 38206 44634
rect 38258 44582 47950 44634
rect 48002 44582 48014 44634
rect 48066 44582 48078 44634
rect 48130 44582 48142 44634
rect 48194 44582 48206 44634
rect 48258 44582 49864 44634
rect 1104 44560 49864 44582
rect 9766 44480 9772 44532
rect 9824 44520 9830 44532
rect 14369 44523 14427 44529
rect 14369 44520 14381 44523
rect 9824 44492 14381 44520
rect 9824 44480 9830 44492
rect 14369 44489 14381 44492
rect 14415 44489 14427 44523
rect 14369 44483 14427 44489
rect 35434 44480 35440 44532
rect 35492 44520 35498 44532
rect 36538 44520 36544 44532
rect 35492 44492 36544 44520
rect 35492 44480 35498 44492
rect 36538 44480 36544 44492
rect 36596 44480 36602 44532
rect 36630 44480 36636 44532
rect 36688 44480 36694 44532
rect 39209 44523 39267 44529
rect 39209 44489 39221 44523
rect 39255 44520 39267 44523
rect 40678 44520 40684 44532
rect 39255 44492 40684 44520
rect 39255 44489 39267 44492
rect 39209 44483 39267 44489
rect 40678 44480 40684 44492
rect 40736 44480 40742 44532
rect 14277 44387 14335 44393
rect 14277 44353 14289 44387
rect 14323 44384 14335 44387
rect 14458 44384 14464 44396
rect 14323 44356 14464 44384
rect 14323 44353 14335 44356
rect 14277 44347 14335 44353
rect 14458 44344 14464 44356
rect 14516 44344 14522 44396
rect 37642 44344 37648 44396
rect 37700 44384 37706 44396
rect 39117 44387 39175 44393
rect 39117 44384 39129 44387
rect 37700 44356 39129 44384
rect 37700 44344 37706 44356
rect 39117 44353 39129 44356
rect 39163 44353 39175 44387
rect 39117 44347 39175 44353
rect 49326 44344 49332 44396
rect 49384 44344 49390 44396
rect 36817 44319 36875 44325
rect 36817 44285 36829 44319
rect 36863 44316 36875 44319
rect 36906 44316 36912 44328
rect 36863 44288 36912 44316
rect 36863 44285 36875 44288
rect 36817 44279 36875 44285
rect 36906 44276 36912 44288
rect 36964 44276 36970 44328
rect 39298 44276 39304 44328
rect 39356 44276 39362 44328
rect 36170 44140 36176 44192
rect 36228 44140 36234 44192
rect 36538 44140 36544 44192
rect 36596 44180 36602 44192
rect 37642 44180 37648 44192
rect 36596 44152 37648 44180
rect 36596 44140 36602 44152
rect 37642 44140 37648 44152
rect 37700 44140 37706 44192
rect 38746 44140 38752 44192
rect 38804 44140 38810 44192
rect 43438 44140 43444 44192
rect 43496 44180 43502 44192
rect 49145 44183 49203 44189
rect 49145 44180 49157 44183
rect 43496 44152 49157 44180
rect 43496 44140 43502 44152
rect 49145 44149 49157 44152
rect 49191 44149 49203 44183
rect 49145 44143 49203 44149
rect 1104 44090 49864 44112
rect 1104 44038 2950 44090
rect 3002 44038 3014 44090
rect 3066 44038 3078 44090
rect 3130 44038 3142 44090
rect 3194 44038 3206 44090
rect 3258 44038 12950 44090
rect 13002 44038 13014 44090
rect 13066 44038 13078 44090
rect 13130 44038 13142 44090
rect 13194 44038 13206 44090
rect 13258 44038 22950 44090
rect 23002 44038 23014 44090
rect 23066 44038 23078 44090
rect 23130 44038 23142 44090
rect 23194 44038 23206 44090
rect 23258 44038 32950 44090
rect 33002 44038 33014 44090
rect 33066 44038 33078 44090
rect 33130 44038 33142 44090
rect 33194 44038 33206 44090
rect 33258 44038 42950 44090
rect 43002 44038 43014 44090
rect 43066 44038 43078 44090
rect 43130 44038 43142 44090
rect 43194 44038 43206 44090
rect 43258 44038 49864 44090
rect 1104 44016 49864 44038
rect 11698 43936 11704 43988
rect 11756 43976 11762 43988
rect 13541 43979 13599 43985
rect 13541 43976 13553 43979
rect 11756 43948 13553 43976
rect 11756 43936 11762 43948
rect 13541 43945 13553 43948
rect 13587 43945 13599 43979
rect 13541 43939 13599 43945
rect 14642 43936 14648 43988
rect 14700 43976 14706 43988
rect 16209 43979 16267 43985
rect 16209 43976 16221 43979
rect 14700 43948 16221 43976
rect 14700 43936 14706 43948
rect 16209 43945 16221 43948
rect 16255 43945 16267 43979
rect 16209 43939 16267 43945
rect 16942 43936 16948 43988
rect 17000 43936 17006 43988
rect 20438 43936 20444 43988
rect 20496 43936 20502 43988
rect 21266 43936 21272 43988
rect 21324 43936 21330 43988
rect 22278 43936 22284 43988
rect 22336 43936 22342 43988
rect 28445 43979 28503 43985
rect 28445 43945 28457 43979
rect 28491 43976 28503 43979
rect 32030 43976 32036 43988
rect 28491 43948 32036 43976
rect 28491 43945 28503 43948
rect 28445 43939 28503 43945
rect 32030 43936 32036 43948
rect 32088 43936 32094 43988
rect 12434 43868 12440 43920
rect 12492 43868 12498 43920
rect 19610 43868 19616 43920
rect 19668 43908 19674 43920
rect 22925 43911 22983 43917
rect 22925 43908 22937 43911
rect 19668 43880 22937 43908
rect 19668 43868 19674 43880
rect 22925 43877 22937 43880
rect 22971 43877 22983 43911
rect 22925 43871 22983 43877
rect 28810 43868 28816 43920
rect 28868 43908 28874 43920
rect 28868 43880 28948 43908
rect 28868 43868 28874 43880
rect 28920 43849 28948 43880
rect 28905 43843 28963 43849
rect 28905 43809 28917 43843
rect 28951 43809 28963 43843
rect 28905 43803 28963 43809
rect 28994 43800 29000 43852
rect 29052 43800 29058 43852
rect 30377 43843 30435 43849
rect 30377 43809 30389 43843
rect 30423 43840 30435 43843
rect 32950 43840 32956 43852
rect 30423 43812 32956 43840
rect 30423 43809 30435 43812
rect 30377 43803 30435 43809
rect 32950 43800 32956 43812
rect 33008 43840 33014 43852
rect 34057 43843 34115 43849
rect 34057 43840 34069 43843
rect 33008 43812 34069 43840
rect 33008 43800 33014 43812
rect 34057 43809 34069 43812
rect 34103 43809 34115 43843
rect 34057 43803 34115 43809
rect 37921 43843 37979 43849
rect 37921 43809 37933 43843
rect 37967 43840 37979 43843
rect 38286 43840 38292 43852
rect 37967 43812 38292 43840
rect 37967 43809 37979 43812
rect 37921 43803 37979 43809
rect 38286 43800 38292 43812
rect 38344 43800 38350 43852
rect 934 43732 940 43784
rect 992 43772 998 43784
rect 1765 43775 1823 43781
rect 1765 43772 1777 43775
rect 992 43744 1777 43772
rect 992 43732 998 43744
rect 1765 43741 1777 43744
rect 1811 43741 1823 43775
rect 1765 43735 1823 43741
rect 12253 43775 12311 43781
rect 12253 43741 12265 43775
rect 12299 43772 12311 43775
rect 21910 43772 21916 43784
rect 12299 43744 21916 43772
rect 12299 43741 12311 43744
rect 12253 43735 12311 43741
rect 21910 43732 21916 43744
rect 21968 43732 21974 43784
rect 22465 43775 22523 43781
rect 22465 43741 22477 43775
rect 22511 43772 22523 43775
rect 23290 43772 23296 43784
rect 22511 43744 23296 43772
rect 22511 43741 22523 43744
rect 22465 43735 22523 43741
rect 23290 43732 23296 43744
rect 23348 43732 23354 43784
rect 26234 43732 26240 43784
rect 26292 43772 26298 43784
rect 26292 43744 27568 43772
rect 26292 43732 26298 43744
rect 13446 43664 13452 43716
rect 13504 43664 13510 43716
rect 16117 43707 16175 43713
rect 16117 43673 16129 43707
rect 16163 43704 16175 43707
rect 16853 43707 16911 43713
rect 16163 43676 16574 43704
rect 16163 43673 16175 43676
rect 16117 43667 16175 43673
rect 1581 43639 1639 43645
rect 1581 43605 1593 43639
rect 1627 43636 1639 43639
rect 2038 43636 2044 43648
rect 1627 43608 2044 43636
rect 1627 43605 1639 43608
rect 1581 43599 1639 43605
rect 2038 43596 2044 43608
rect 2096 43596 2102 43648
rect 16546 43636 16574 43676
rect 16853 43673 16865 43707
rect 16899 43704 16911 43707
rect 19978 43704 19984 43716
rect 16899 43676 19984 43704
rect 16899 43673 16911 43676
rect 16853 43667 16911 43673
rect 19978 43664 19984 43676
rect 20036 43664 20042 43716
rect 20349 43707 20407 43713
rect 20349 43673 20361 43707
rect 20395 43704 20407 43707
rect 20438 43704 20444 43716
rect 20395 43676 20444 43704
rect 20395 43673 20407 43676
rect 20349 43667 20407 43673
rect 20438 43664 20444 43676
rect 20496 43664 20502 43716
rect 21177 43707 21235 43713
rect 21177 43673 21189 43707
rect 21223 43673 21235 43707
rect 21177 43667 21235 43673
rect 22189 43707 22247 43713
rect 22189 43673 22201 43707
rect 22235 43704 22247 43707
rect 22741 43707 22799 43713
rect 22741 43704 22753 43707
rect 22235 43676 22753 43704
rect 22235 43673 22247 43676
rect 22189 43667 22247 43673
rect 22741 43673 22753 43676
rect 22787 43704 22799 43707
rect 27540 43704 27568 43744
rect 28626 43732 28632 43784
rect 28684 43772 28690 43784
rect 30101 43775 30159 43781
rect 30101 43772 30113 43775
rect 28684 43744 30113 43772
rect 28684 43732 28690 43744
rect 30101 43741 30113 43744
rect 30147 43741 30159 43775
rect 30101 43735 30159 43741
rect 32306 43732 32312 43784
rect 32364 43732 32370 43784
rect 37737 43775 37795 43781
rect 37737 43741 37749 43775
rect 37783 43772 37795 43775
rect 41506 43772 41512 43784
rect 37783 43744 41512 43772
rect 37783 43741 37795 43744
rect 37737 43735 37795 43741
rect 41506 43732 41512 43744
rect 41564 43732 41570 43784
rect 48498 43732 48504 43784
rect 48556 43732 48562 43784
rect 48777 43775 48835 43781
rect 48777 43741 48789 43775
rect 48823 43741 48835 43775
rect 48777 43735 48835 43741
rect 28813 43707 28871 43713
rect 28813 43704 28825 43707
rect 22787 43676 26234 43704
rect 27540 43676 28825 43704
rect 22787 43673 22799 43676
rect 22741 43667 22799 43673
rect 20990 43636 20996 43648
rect 16546 43608 20996 43636
rect 20990 43596 20996 43608
rect 21048 43596 21054 43648
rect 21192 43636 21220 43667
rect 24210 43636 24216 43648
rect 21192 43608 24216 43636
rect 24210 43596 24216 43608
rect 24268 43596 24274 43648
rect 26206 43636 26234 43676
rect 28813 43673 28825 43676
rect 28859 43673 28871 43707
rect 31662 43704 31668 43716
rect 31602 43676 31668 43704
rect 28813 43667 28871 43673
rect 31662 43664 31668 43676
rect 31720 43664 31726 43716
rect 32585 43707 32643 43713
rect 32585 43673 32597 43707
rect 32631 43673 32643 43707
rect 32585 43667 32643 43673
rect 30650 43636 30656 43648
rect 26206 43608 30656 43636
rect 30650 43596 30656 43608
rect 30708 43596 30714 43648
rect 31754 43596 31760 43648
rect 31812 43636 31818 43648
rect 31849 43639 31907 43645
rect 31849 43636 31861 43639
rect 31812 43608 31861 43636
rect 31812 43596 31818 43608
rect 31849 43605 31861 43608
rect 31895 43605 31907 43639
rect 32600 43636 32628 43667
rect 33594 43664 33600 43716
rect 33652 43664 33658 43716
rect 36722 43704 36728 43716
rect 35866 43676 36728 43704
rect 33318 43636 33324 43648
rect 32600 43608 33324 43636
rect 31849 43599 31907 43605
rect 33318 43596 33324 43608
rect 33376 43596 33382 43648
rect 33410 43596 33416 43648
rect 33468 43636 33474 43648
rect 35866 43636 35894 43676
rect 36722 43664 36728 43676
rect 36780 43704 36786 43716
rect 37645 43707 37703 43713
rect 37645 43704 37657 43707
rect 36780 43676 37657 43704
rect 36780 43664 36786 43676
rect 37645 43673 37657 43676
rect 37691 43673 37703 43707
rect 37645 43667 37703 43673
rect 40954 43664 40960 43716
rect 41012 43704 41018 43716
rect 48792 43704 48820 43735
rect 41012 43676 48820 43704
rect 41012 43664 41018 43676
rect 33468 43608 35894 43636
rect 33468 43596 33474 43608
rect 37274 43596 37280 43648
rect 37332 43596 37338 43648
rect 1104 43546 49864 43568
rect 1104 43494 7950 43546
rect 8002 43494 8014 43546
rect 8066 43494 8078 43546
rect 8130 43494 8142 43546
rect 8194 43494 8206 43546
rect 8258 43494 17950 43546
rect 18002 43494 18014 43546
rect 18066 43494 18078 43546
rect 18130 43494 18142 43546
rect 18194 43494 18206 43546
rect 18258 43494 27950 43546
rect 28002 43494 28014 43546
rect 28066 43494 28078 43546
rect 28130 43494 28142 43546
rect 28194 43494 28206 43546
rect 28258 43494 37950 43546
rect 38002 43494 38014 43546
rect 38066 43494 38078 43546
rect 38130 43494 38142 43546
rect 38194 43494 38206 43546
rect 38258 43494 47950 43546
rect 48002 43494 48014 43546
rect 48066 43494 48078 43546
rect 48130 43494 48142 43546
rect 48194 43494 48206 43546
rect 48258 43494 49864 43546
rect 1104 43472 49864 43494
rect 2038 43392 2044 43444
rect 2096 43392 2102 43444
rect 8938 43392 8944 43444
rect 8996 43432 9002 43444
rect 12161 43435 12219 43441
rect 12161 43432 12173 43435
rect 8996 43404 12173 43432
rect 8996 43392 9002 43404
rect 12161 43401 12173 43404
rect 12207 43401 12219 43435
rect 12161 43395 12219 43401
rect 16850 43392 16856 43444
rect 16908 43392 16914 43444
rect 19150 43392 19156 43444
rect 19208 43392 19214 43444
rect 20346 43392 20352 43444
rect 20404 43392 20410 43444
rect 20898 43392 20904 43444
rect 20956 43392 20962 43444
rect 20990 43392 20996 43444
rect 21048 43432 21054 43444
rect 24394 43432 24400 43444
rect 21048 43404 24400 43432
rect 21048 43392 21054 43404
rect 24394 43392 24400 43404
rect 24452 43392 24458 43444
rect 24854 43392 24860 43444
rect 24912 43432 24918 43444
rect 25869 43435 25927 43441
rect 25869 43432 25881 43435
rect 24912 43404 25881 43432
rect 24912 43392 24918 43404
rect 25869 43401 25881 43404
rect 25915 43401 25927 43435
rect 25869 43395 25927 43401
rect 28810 43392 28816 43444
rect 28868 43432 28874 43444
rect 31386 43432 31392 43444
rect 28868 43404 31392 43432
rect 28868 43392 28874 43404
rect 31386 43392 31392 43404
rect 31444 43392 31450 43444
rect 32306 43392 32312 43444
rect 32364 43432 32370 43444
rect 32364 43404 34560 43432
rect 32364 43392 32370 43404
rect 31662 43364 31668 43376
rect 30314 43336 31668 43364
rect 31662 43324 31668 43336
rect 31720 43324 31726 43376
rect 34532 43308 34560 43404
rect 40310 43392 40316 43444
rect 40368 43392 40374 43444
rect 34790 43324 34796 43376
rect 34848 43324 34854 43376
rect 2225 43299 2283 43305
rect 2225 43265 2237 43299
rect 2271 43296 2283 43299
rect 11974 43296 11980 43308
rect 2271 43268 11980 43296
rect 2271 43265 2283 43268
rect 2225 43259 2283 43265
rect 11974 43256 11980 43268
rect 12032 43256 12038 43308
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 17037 43299 17095 43305
rect 17037 43265 17049 43299
rect 17083 43265 17095 43299
rect 17037 43259 17095 43265
rect 17052 43228 17080 43259
rect 19058 43256 19064 43308
rect 19116 43256 19122 43308
rect 20254 43256 20260 43308
rect 20312 43256 20318 43308
rect 21085 43299 21143 43305
rect 21085 43265 21097 43299
rect 21131 43296 21143 43299
rect 21726 43296 21732 43308
rect 21131 43268 21732 43296
rect 21131 43265 21143 43268
rect 21085 43259 21143 43265
rect 21726 43256 21732 43268
rect 21784 43256 21790 43308
rect 25958 43256 25964 43308
rect 26016 43296 26022 43308
rect 26237 43299 26295 43305
rect 26237 43296 26249 43299
rect 26016 43268 26249 43296
rect 26016 43256 26022 43268
rect 26237 43265 26249 43268
rect 26283 43265 26295 43299
rect 26237 43259 26295 43265
rect 32306 43256 32312 43308
rect 32364 43256 32370 43308
rect 33594 43256 33600 43308
rect 33652 43296 33658 43308
rect 33652 43282 33718 43296
rect 33652 43268 33732 43282
rect 33652 43256 33658 43268
rect 19426 43228 19432 43240
rect 17052 43200 19432 43228
rect 19426 43188 19432 43200
rect 19484 43188 19490 43240
rect 26326 43188 26332 43240
rect 26384 43188 26390 43240
rect 26513 43231 26571 43237
rect 26513 43197 26525 43231
rect 26559 43228 26571 43231
rect 27338 43228 27344 43240
rect 26559 43200 27344 43228
rect 26559 43197 26571 43200
rect 26513 43191 26571 43197
rect 27338 43188 27344 43200
rect 27396 43188 27402 43240
rect 28626 43188 28632 43240
rect 28684 43228 28690 43240
rect 28813 43231 28871 43237
rect 28813 43228 28825 43231
rect 28684 43200 28825 43228
rect 28684 43188 28690 43200
rect 28813 43197 28825 43200
rect 28859 43197 28871 43231
rect 28813 43191 28871 43197
rect 29089 43231 29147 43237
rect 29089 43197 29101 43231
rect 29135 43228 29147 43231
rect 31846 43228 31852 43240
rect 29135 43200 31852 43228
rect 29135 43197 29147 43200
rect 29089 43191 29147 43197
rect 31846 43188 31852 43200
rect 31904 43188 31910 43240
rect 32585 43231 32643 43237
rect 32585 43197 32597 43231
rect 32631 43228 32643 43231
rect 33704 43228 33732 43268
rect 34514 43256 34520 43308
rect 34572 43256 34578 43308
rect 35912 43228 35940 43282
rect 38930 43256 38936 43308
rect 38988 43296 38994 43308
rect 39850 43296 39856 43308
rect 38988 43268 39856 43296
rect 38988 43256 38994 43268
rect 39850 43256 39856 43268
rect 39908 43296 39914 43308
rect 40221 43299 40279 43305
rect 40221 43296 40233 43299
rect 39908 43268 40233 43296
rect 39908 43256 39914 43268
rect 40221 43265 40233 43268
rect 40267 43265 40279 43299
rect 48777 43299 48835 43305
rect 48777 43296 48789 43299
rect 40221 43259 40279 43265
rect 45526 43268 48789 43296
rect 35986 43228 35992 43240
rect 32631 43200 33640 43228
rect 33704 43200 35992 43228
rect 32631 43197 32643 43200
rect 32585 43191 32643 43197
rect 13446 43120 13452 43172
rect 13504 43160 13510 43172
rect 24026 43160 24032 43172
rect 13504 43132 24032 43160
rect 13504 43120 13510 43132
rect 24026 43120 24032 43132
rect 24084 43120 24090 43172
rect 33612 43160 33640 43200
rect 35986 43188 35992 43200
rect 36044 43188 36050 43240
rect 40497 43231 40555 43237
rect 40497 43197 40509 43231
rect 40543 43228 40555 43231
rect 40586 43228 40592 43240
rect 40543 43200 40592 43228
rect 40543 43197 40555 43200
rect 40497 43191 40555 43197
rect 40586 43188 40592 43200
rect 40644 43188 40650 43240
rect 42058 43188 42064 43240
rect 42116 43228 42122 43240
rect 45526 43228 45554 43268
rect 48777 43265 48789 43268
rect 48823 43265 48835 43299
rect 48777 43259 48835 43265
rect 42116 43200 45554 43228
rect 42116 43188 42122 43200
rect 48498 43188 48504 43240
rect 48556 43188 48562 43240
rect 34146 43160 34152 43172
rect 33612 43132 34152 43160
rect 34146 43120 34152 43132
rect 34204 43120 34210 43172
rect 28902 43052 28908 43104
rect 28960 43092 28966 43104
rect 30561 43095 30619 43101
rect 30561 43092 30573 43095
rect 28960 43064 30573 43092
rect 28960 43052 28966 43064
rect 30561 43061 30573 43064
rect 30607 43061 30619 43095
rect 30561 43055 30619 43061
rect 34054 43052 34060 43104
rect 34112 43052 34118 43104
rect 34164 43092 34192 43120
rect 36265 43095 36323 43101
rect 36265 43092 36277 43095
rect 34164 43064 36277 43092
rect 36265 43061 36277 43064
rect 36311 43061 36323 43095
rect 36265 43055 36323 43061
rect 39853 43095 39911 43101
rect 39853 43061 39865 43095
rect 39899 43092 39911 43095
rect 41230 43092 41236 43104
rect 39899 43064 41236 43092
rect 39899 43061 39911 43064
rect 39853 43055 39911 43061
rect 41230 43052 41236 43064
rect 41288 43052 41294 43104
rect 1104 43002 49864 43024
rect 1104 42950 2950 43002
rect 3002 42950 3014 43002
rect 3066 42950 3078 43002
rect 3130 42950 3142 43002
rect 3194 42950 3206 43002
rect 3258 42950 12950 43002
rect 13002 42950 13014 43002
rect 13066 42950 13078 43002
rect 13130 42950 13142 43002
rect 13194 42950 13206 43002
rect 13258 42950 22950 43002
rect 23002 42950 23014 43002
rect 23066 42950 23078 43002
rect 23130 42950 23142 43002
rect 23194 42950 23206 43002
rect 23258 42950 32950 43002
rect 33002 42950 33014 43002
rect 33066 42950 33078 43002
rect 33130 42950 33142 43002
rect 33194 42950 33206 43002
rect 33258 42950 42950 43002
rect 43002 42950 43014 43002
rect 43066 42950 43078 43002
rect 43130 42950 43142 43002
rect 43194 42950 43206 43002
rect 43258 42950 49864 43002
rect 1104 42928 49864 42950
rect 12066 42848 12072 42900
rect 12124 42888 12130 42900
rect 21542 42888 21548 42900
rect 12124 42860 21548 42888
rect 12124 42848 12130 42860
rect 21542 42848 21548 42860
rect 21600 42848 21606 42900
rect 27338 42848 27344 42900
rect 27396 42848 27402 42900
rect 40034 42780 40040 42832
rect 40092 42820 40098 42832
rect 40092 42792 40632 42820
rect 40092 42780 40098 42792
rect 35897 42755 35955 42761
rect 35897 42721 35909 42755
rect 35943 42752 35955 42755
rect 36906 42752 36912 42764
rect 35943 42724 36912 42752
rect 35943 42721 35955 42724
rect 35897 42715 35955 42721
rect 36906 42712 36912 42724
rect 36964 42712 36970 42764
rect 40604 42761 40632 42792
rect 40589 42755 40647 42761
rect 40589 42721 40601 42755
rect 40635 42721 40647 42755
rect 40589 42715 40647 42721
rect 24118 42644 24124 42696
rect 24176 42684 24182 42696
rect 25593 42687 25651 42693
rect 25593 42684 25605 42687
rect 24176 42656 25605 42684
rect 24176 42644 24182 42656
rect 25593 42653 25605 42656
rect 25639 42653 25651 42687
rect 25593 42647 25651 42653
rect 25608 42548 25636 42647
rect 34514 42644 34520 42696
rect 34572 42684 34578 42696
rect 35621 42687 35679 42693
rect 35621 42684 35633 42687
rect 34572 42656 35633 42684
rect 34572 42644 34578 42656
rect 35621 42653 35633 42656
rect 35667 42653 35679 42687
rect 35621 42647 35679 42653
rect 36998 42644 37004 42696
rect 37056 42644 37062 42696
rect 40497 42687 40555 42693
rect 40497 42653 40509 42687
rect 40543 42684 40555 42687
rect 44174 42684 44180 42696
rect 40543 42656 44180 42684
rect 40543 42653 40555 42656
rect 40497 42647 40555 42653
rect 44174 42644 44180 42656
rect 44232 42644 44238 42696
rect 48498 42644 48504 42696
rect 48556 42644 48562 42696
rect 48777 42687 48835 42693
rect 48777 42653 48789 42687
rect 48823 42653 48835 42687
rect 48777 42647 48835 42653
rect 25866 42576 25872 42628
rect 25924 42576 25930 42628
rect 26142 42576 26148 42628
rect 26200 42616 26206 42628
rect 48792 42616 48820 42647
rect 26200 42588 26358 42616
rect 40512 42588 48820 42616
rect 26200 42576 26206 42588
rect 40512 42560 40540 42588
rect 27246 42548 27252 42560
rect 25608 42520 27252 42548
rect 27246 42508 27252 42520
rect 27304 42508 27310 42560
rect 36814 42508 36820 42560
rect 36872 42548 36878 42560
rect 37369 42551 37427 42557
rect 37369 42548 37381 42551
rect 36872 42520 37381 42548
rect 36872 42508 36878 42520
rect 37369 42517 37381 42520
rect 37415 42517 37427 42551
rect 37369 42511 37427 42517
rect 40037 42551 40095 42557
rect 40037 42517 40049 42551
rect 40083 42548 40095 42551
rect 40218 42548 40224 42560
rect 40083 42520 40224 42548
rect 40083 42517 40095 42520
rect 40037 42511 40095 42517
rect 40218 42508 40224 42520
rect 40276 42508 40282 42560
rect 40402 42508 40408 42560
rect 40460 42508 40466 42560
rect 40494 42508 40500 42560
rect 40552 42508 40558 42560
rect 1104 42458 49864 42480
rect 1104 42406 7950 42458
rect 8002 42406 8014 42458
rect 8066 42406 8078 42458
rect 8130 42406 8142 42458
rect 8194 42406 8206 42458
rect 8258 42406 17950 42458
rect 18002 42406 18014 42458
rect 18066 42406 18078 42458
rect 18130 42406 18142 42458
rect 18194 42406 18206 42458
rect 18258 42406 27950 42458
rect 28002 42406 28014 42458
rect 28066 42406 28078 42458
rect 28130 42406 28142 42458
rect 28194 42406 28206 42458
rect 28258 42406 37950 42458
rect 38002 42406 38014 42458
rect 38066 42406 38078 42458
rect 38130 42406 38142 42458
rect 38194 42406 38206 42458
rect 38258 42406 47950 42458
rect 48002 42406 48014 42458
rect 48066 42406 48078 42458
rect 48130 42406 48142 42458
rect 48194 42406 48206 42458
rect 48258 42406 49864 42458
rect 1104 42384 49864 42406
rect 6362 42304 6368 42356
rect 6420 42344 6426 42356
rect 7285 42347 7343 42353
rect 7285 42344 7297 42347
rect 6420 42316 7297 42344
rect 6420 42304 6426 42316
rect 7285 42313 7297 42316
rect 7331 42313 7343 42347
rect 7285 42307 7343 42313
rect 9214 42304 9220 42356
rect 9272 42304 9278 42356
rect 14550 42304 14556 42356
rect 14608 42344 14614 42356
rect 17313 42347 17371 42353
rect 17313 42344 17325 42347
rect 14608 42316 17325 42344
rect 14608 42304 14614 42316
rect 17313 42313 17325 42316
rect 17359 42313 17371 42347
rect 17313 42307 17371 42313
rect 20622 42304 20628 42356
rect 20680 42304 20686 42356
rect 22186 42304 22192 42356
rect 22244 42304 22250 42356
rect 25866 42304 25872 42356
rect 25924 42304 25930 42356
rect 31754 42344 31760 42356
rect 27264 42316 31760 42344
rect 6270 42236 6276 42288
rect 6328 42276 6334 42288
rect 8113 42279 8171 42285
rect 8113 42276 8125 42279
rect 6328 42248 8125 42276
rect 6328 42236 6334 42248
rect 8113 42245 8125 42248
rect 8159 42245 8171 42279
rect 8113 42239 8171 42245
rect 24302 42236 24308 42288
rect 24360 42276 24366 42288
rect 24397 42279 24455 42285
rect 24397 42276 24409 42279
rect 24360 42248 24409 42276
rect 24360 42236 24366 42248
rect 24397 42245 24409 42248
rect 24443 42245 24455 42279
rect 24397 42239 24455 42245
rect 24854 42236 24860 42288
rect 24912 42236 24918 42288
rect 7190 42168 7196 42220
rect 7248 42168 7254 42220
rect 7929 42211 7987 42217
rect 7929 42177 7941 42211
rect 7975 42177 7987 42211
rect 7929 42171 7987 42177
rect 7944 42140 7972 42171
rect 9122 42168 9128 42220
rect 9180 42168 9186 42220
rect 17221 42211 17279 42217
rect 17221 42177 17233 42211
rect 17267 42208 17279 42211
rect 17402 42208 17408 42220
rect 17267 42180 17408 42208
rect 17267 42177 17279 42180
rect 17221 42171 17279 42177
rect 17402 42168 17408 42180
rect 17460 42168 17466 42220
rect 20806 42168 20812 42220
rect 20864 42168 20870 42220
rect 22370 42168 22376 42220
rect 22428 42168 22434 42220
rect 27264 42208 27292 42316
rect 27338 42236 27344 42288
rect 27396 42276 27402 42288
rect 30300 42285 30328 42316
rect 31754 42304 31760 42316
rect 31812 42344 31818 42356
rect 32766 42344 32772 42356
rect 31812 42316 32772 42344
rect 31812 42304 31818 42316
rect 32766 42304 32772 42316
rect 32824 42304 32830 42356
rect 34514 42304 34520 42356
rect 34572 42304 34578 42356
rect 38286 42304 38292 42356
rect 38344 42344 38350 42356
rect 40037 42347 40095 42353
rect 40037 42344 40049 42347
rect 38344 42316 40049 42344
rect 38344 42304 38350 42316
rect 40037 42313 40049 42316
rect 40083 42313 40095 42347
rect 40037 42307 40095 42313
rect 41598 42304 41604 42356
rect 41656 42304 41662 42356
rect 27985 42279 28043 42285
rect 27985 42276 27997 42279
rect 27396 42248 27997 42276
rect 27396 42236 27402 42248
rect 27985 42245 27997 42248
rect 28031 42245 28043 42279
rect 27985 42239 28043 42245
rect 30285 42279 30343 42285
rect 30285 42245 30297 42279
rect 30331 42245 30343 42279
rect 31662 42276 31668 42288
rect 31510 42248 31668 42276
rect 30285 42239 30343 42245
rect 31662 42236 31668 42248
rect 31720 42236 31726 42288
rect 34532 42276 34560 42304
rect 35986 42276 35992 42288
rect 33888 42248 34560 42276
rect 35374 42248 35992 42276
rect 33888 42217 33916 42248
rect 35986 42236 35992 42248
rect 36044 42276 36050 42288
rect 36998 42276 37004 42288
rect 36044 42248 37004 42276
rect 36044 42236 36050 42248
rect 36998 42236 37004 42248
rect 37056 42236 37062 42288
rect 33873 42211 33931 42217
rect 27264 42180 27384 42208
rect 27356 42152 27384 42180
rect 17310 42140 17316 42152
rect 7944 42112 17316 42140
rect 17310 42100 17316 42112
rect 17368 42100 17374 42152
rect 24118 42100 24124 42152
rect 24176 42100 24182 42152
rect 27338 42100 27344 42152
rect 27396 42100 27402 42152
rect 27709 42143 27767 42149
rect 27709 42109 27721 42143
rect 27755 42109 27767 42143
rect 27709 42103 27767 42109
rect 1578 42032 1584 42084
rect 1636 42072 1642 42084
rect 23750 42072 23756 42084
rect 1636 42044 23756 42072
rect 1636 42032 1642 42044
rect 23750 42032 23756 42044
rect 23808 42032 23814 42084
rect 25866 41964 25872 42016
rect 25924 42004 25930 42016
rect 26510 42004 26516 42016
rect 25924 41976 26516 42004
rect 25924 41964 25930 41976
rect 26510 41964 26516 41976
rect 26568 41964 26574 42016
rect 27246 41964 27252 42016
rect 27304 42004 27310 42016
rect 27724 42004 27752 42103
rect 29104 42084 29132 42194
rect 33873 42177 33885 42211
rect 33919 42177 33931 42211
rect 33873 42171 33931 42177
rect 39666 42168 39672 42220
rect 39724 42168 39730 42220
rect 41322 42168 41328 42220
rect 41380 42208 41386 42220
rect 41509 42211 41567 42217
rect 41509 42208 41521 42211
rect 41380 42180 41521 42208
rect 41380 42168 41386 42180
rect 41509 42177 41521 42180
rect 41555 42177 41567 42211
rect 41509 42171 41567 42177
rect 46290 42168 46296 42220
rect 46348 42208 46354 42220
rect 48777 42211 48835 42217
rect 48777 42208 48789 42211
rect 46348 42180 48789 42208
rect 46348 42168 46354 42180
rect 48777 42177 48789 42180
rect 48823 42177 48835 42211
rect 48777 42171 48835 42177
rect 29178 42100 29184 42152
rect 29236 42140 29242 42152
rect 30009 42143 30067 42149
rect 30009 42140 30021 42143
rect 29236 42112 30021 42140
rect 29236 42100 29242 42112
rect 30009 42109 30021 42112
rect 30055 42140 30067 42143
rect 31294 42140 31300 42152
rect 30055 42112 31300 42140
rect 30055 42109 30067 42112
rect 30009 42103 30067 42109
rect 31294 42100 31300 42112
rect 31352 42100 31358 42152
rect 34149 42143 34207 42149
rect 34149 42109 34161 42143
rect 34195 42140 34207 42143
rect 35526 42140 35532 42152
rect 34195 42112 35532 42140
rect 34195 42109 34207 42112
rect 34149 42103 34207 42109
rect 35526 42100 35532 42112
rect 35584 42100 35590 42152
rect 37826 42100 37832 42152
rect 37884 42140 37890 42152
rect 38289 42143 38347 42149
rect 38289 42140 38301 42143
rect 37884 42112 38301 42140
rect 37884 42100 37890 42112
rect 38289 42109 38301 42112
rect 38335 42109 38347 42143
rect 38289 42103 38347 42109
rect 38565 42143 38623 42149
rect 38565 42109 38577 42143
rect 38611 42140 38623 42143
rect 40310 42140 40316 42152
rect 38611 42112 40316 42140
rect 38611 42109 38623 42112
rect 38565 42103 38623 42109
rect 40310 42100 40316 42112
rect 40368 42100 40374 42152
rect 41785 42143 41843 42149
rect 41785 42109 41797 42143
rect 41831 42140 41843 42143
rect 43898 42140 43904 42152
rect 41831 42112 43904 42140
rect 41831 42109 41843 42112
rect 41785 42103 41843 42109
rect 43898 42100 43904 42112
rect 43956 42100 43962 42152
rect 48498 42100 48504 42152
rect 48556 42100 48562 42152
rect 29086 42032 29092 42084
rect 29144 42072 29150 42084
rect 29144 42044 29960 42072
rect 29144 42032 29150 42044
rect 28626 42004 28632 42016
rect 27304 41976 28632 42004
rect 27304 41964 27310 41976
rect 28626 41964 28632 41976
rect 28684 42004 28690 42016
rect 29178 42004 29184 42016
rect 28684 41976 29184 42004
rect 28684 41964 28690 41976
rect 29178 41964 29184 41976
rect 29236 41964 29242 42016
rect 29457 42007 29515 42013
rect 29457 41973 29469 42007
rect 29503 42004 29515 42007
rect 29822 42004 29828 42016
rect 29503 41976 29828 42004
rect 29503 41973 29515 41976
rect 29457 41967 29515 41973
rect 29822 41964 29828 41976
rect 29880 41964 29886 42016
rect 29932 42004 29960 42044
rect 31386 42032 31392 42084
rect 31444 42072 31450 42084
rect 32490 42072 32496 42084
rect 31444 42044 32496 42072
rect 31444 42032 31450 42044
rect 32490 42032 32496 42044
rect 32548 42032 32554 42084
rect 31662 42004 31668 42016
rect 29932 41976 31668 42004
rect 31662 41964 31668 41976
rect 31720 41964 31726 42016
rect 31757 42007 31815 42013
rect 31757 41973 31769 42007
rect 31803 42004 31815 42007
rect 31846 42004 31852 42016
rect 31803 41976 31852 42004
rect 31803 41973 31815 41976
rect 31757 41967 31815 41973
rect 31846 41964 31852 41976
rect 31904 41964 31910 42016
rect 35618 41964 35624 42016
rect 35676 41964 35682 42016
rect 41141 42007 41199 42013
rect 41141 41973 41153 42007
rect 41187 42004 41199 42007
rect 43530 42004 43536 42016
rect 41187 41976 43536 42004
rect 41187 41973 41199 41976
rect 41141 41967 41199 41973
rect 43530 41964 43536 41976
rect 43588 41964 43594 42016
rect 1104 41914 49864 41936
rect 1104 41862 2950 41914
rect 3002 41862 3014 41914
rect 3066 41862 3078 41914
rect 3130 41862 3142 41914
rect 3194 41862 3206 41914
rect 3258 41862 12950 41914
rect 13002 41862 13014 41914
rect 13066 41862 13078 41914
rect 13130 41862 13142 41914
rect 13194 41862 13206 41914
rect 13258 41862 22950 41914
rect 23002 41862 23014 41914
rect 23066 41862 23078 41914
rect 23130 41862 23142 41914
rect 23194 41862 23206 41914
rect 23258 41862 32950 41914
rect 33002 41862 33014 41914
rect 33066 41862 33078 41914
rect 33130 41862 33142 41914
rect 33194 41862 33206 41914
rect 33258 41862 42950 41914
rect 43002 41862 43014 41914
rect 43066 41862 43078 41914
rect 43130 41862 43142 41914
rect 43194 41862 43206 41914
rect 43258 41862 49864 41914
rect 1104 41840 49864 41862
rect 21269 41803 21327 41809
rect 21269 41769 21281 41803
rect 21315 41800 21327 41803
rect 21992 41803 22050 41809
rect 21992 41800 22004 41803
rect 21315 41772 22004 41800
rect 21315 41769 21327 41772
rect 21269 41763 21327 41769
rect 21992 41769 22004 41772
rect 22038 41800 22050 41803
rect 22038 41772 26234 41800
rect 22038 41769 22050 41772
rect 21992 41763 22050 41769
rect 26206 41732 26234 41772
rect 26326 41760 26332 41812
rect 26384 41800 26390 41812
rect 26973 41803 27031 41809
rect 26973 41800 26985 41803
rect 26384 41772 26985 41800
rect 26384 41760 26390 41772
rect 26973 41769 26985 41772
rect 27019 41769 27031 41803
rect 26973 41763 27031 41769
rect 31662 41760 31668 41812
rect 31720 41800 31726 41812
rect 33042 41800 33048 41812
rect 31720 41772 33048 41800
rect 31720 41760 31726 41772
rect 33042 41760 33048 41772
rect 33100 41760 33106 41812
rect 35526 41760 35532 41812
rect 35584 41800 35590 41812
rect 36633 41803 36691 41809
rect 36633 41800 36645 41803
rect 35584 41772 36645 41800
rect 35584 41760 35590 41772
rect 36633 41769 36645 41772
rect 36679 41769 36691 41803
rect 36633 41763 36691 41769
rect 36906 41760 36912 41812
rect 36964 41800 36970 41812
rect 38841 41803 38899 41809
rect 38841 41800 38853 41803
rect 36964 41772 38853 41800
rect 36964 41760 36970 41772
rect 38841 41769 38853 41772
rect 38887 41769 38899 41803
rect 38841 41763 38899 41769
rect 48593 41803 48651 41809
rect 48593 41769 48605 41803
rect 48639 41800 48651 41803
rect 48682 41800 48688 41812
rect 48639 41772 48688 41800
rect 48639 41769 48651 41772
rect 48593 41763 48651 41769
rect 48682 41760 48688 41772
rect 48740 41760 48746 41812
rect 31386 41732 31392 41744
rect 26206 41704 31392 41732
rect 31386 41692 31392 41704
rect 31444 41692 31450 41744
rect 21729 41667 21787 41673
rect 21729 41633 21741 41667
rect 21775 41664 21787 41667
rect 24118 41664 24124 41676
rect 21775 41636 24124 41664
rect 21775 41633 21787 41636
rect 21729 41627 21787 41633
rect 24118 41624 24124 41636
rect 24176 41624 24182 41676
rect 26510 41624 26516 41676
rect 26568 41664 26574 41676
rect 27525 41667 27583 41673
rect 27525 41664 27537 41667
rect 26568 41636 27537 41664
rect 26568 41624 26574 41636
rect 27525 41633 27537 41636
rect 27571 41633 27583 41667
rect 34146 41664 34152 41676
rect 27525 41627 27583 41633
rect 31220 41636 34152 41664
rect 23750 41556 23756 41608
rect 23808 41596 23814 41608
rect 26418 41596 26424 41608
rect 23808 41568 26424 41596
rect 23808 41556 23814 41568
rect 26418 41556 26424 41568
rect 26476 41556 26482 41608
rect 31220 41540 31248 41636
rect 34146 41624 34152 41636
rect 34204 41624 34210 41676
rect 34514 41624 34520 41676
rect 34572 41664 34578 41676
rect 34698 41664 34704 41676
rect 34572 41636 34704 41664
rect 34572 41624 34578 41636
rect 34698 41624 34704 41636
rect 34756 41664 34762 41676
rect 34885 41667 34943 41673
rect 34885 41664 34897 41667
rect 34756 41636 34897 41664
rect 34756 41624 34762 41636
rect 34885 41633 34897 41636
rect 34931 41664 34943 41667
rect 37093 41667 37151 41673
rect 37093 41664 37105 41667
rect 34931 41636 37105 41664
rect 34931 41633 34943 41636
rect 34885 41627 34943 41633
rect 37093 41633 37105 41636
rect 37139 41664 37151 41667
rect 37826 41664 37832 41676
rect 37139 41636 37832 41664
rect 37139 41633 37151 41636
rect 37093 41627 37151 41633
rect 37826 41624 37832 41636
rect 37884 41624 37890 41676
rect 31294 41556 31300 41608
rect 31352 41596 31358 41608
rect 31389 41599 31447 41605
rect 31389 41596 31401 41599
rect 31352 41568 31401 41596
rect 31352 41556 31358 41568
rect 31389 41565 31401 41568
rect 31435 41565 31447 41599
rect 33042 41596 33048 41608
rect 32798 41568 33048 41596
rect 31389 41559 31447 41565
rect 33042 41556 33048 41568
rect 33100 41556 33106 41608
rect 48406 41556 48412 41608
rect 48464 41596 48470 41608
rect 48777 41599 48835 41605
rect 48777 41596 48789 41599
rect 48464 41568 48789 41596
rect 48464 41556 48470 41568
rect 48777 41565 48789 41568
rect 48823 41565 48835 41599
rect 48777 41559 48835 41565
rect 1670 41488 1676 41540
rect 1728 41488 1734 41540
rect 11974 41488 11980 41540
rect 12032 41528 12038 41540
rect 22462 41528 22468 41540
rect 12032 41500 22468 41528
rect 12032 41488 12038 41500
rect 22462 41488 22468 41500
rect 22520 41488 22526 41540
rect 27433 41531 27491 41537
rect 27433 41528 27445 41531
rect 26206 41500 27445 41528
rect 1765 41463 1823 41469
rect 1765 41429 1777 41463
rect 1811 41460 1823 41463
rect 10594 41460 10600 41472
rect 1811 41432 10600 41460
rect 1811 41429 1823 41432
rect 1765 41423 1823 41429
rect 10594 41420 10600 41432
rect 10652 41420 10658 41472
rect 22094 41420 22100 41472
rect 22152 41460 22158 41472
rect 26206 41460 26234 41500
rect 27433 41497 27445 41500
rect 27479 41497 27491 41531
rect 27433 41491 27491 41497
rect 31202 41488 31208 41540
rect 31260 41528 31266 41540
rect 31665 41531 31723 41537
rect 31665 41528 31677 41531
rect 31260 41500 31677 41528
rect 31260 41488 31266 41500
rect 31665 41497 31677 41500
rect 31711 41497 31723 41531
rect 35066 41528 35072 41540
rect 31665 41491 31723 41497
rect 32968 41500 35072 41528
rect 22152 41432 26234 41460
rect 27341 41463 27399 41469
rect 22152 41420 22158 41432
rect 27341 41429 27353 41463
rect 27387 41460 27399 41463
rect 32968 41460 32996 41500
rect 35066 41488 35072 41500
rect 35124 41488 35130 41540
rect 35161 41531 35219 41537
rect 35161 41497 35173 41531
rect 35207 41497 35219 41531
rect 36386 41500 36584 41528
rect 35161 41491 35219 41497
rect 27387 41432 32996 41460
rect 33137 41463 33195 41469
rect 27387 41429 27399 41432
rect 27341 41423 27399 41429
rect 33137 41429 33149 41463
rect 33183 41460 33195 41463
rect 33318 41460 33324 41472
rect 33183 41432 33324 41460
rect 33183 41429 33195 41432
rect 33137 41423 33195 41429
rect 33318 41420 33324 41432
rect 33376 41460 33382 41472
rect 34054 41460 34060 41472
rect 33376 41432 34060 41460
rect 33376 41420 33382 41432
rect 34054 41420 34060 41432
rect 34112 41420 34118 41472
rect 35176 41460 35204 41491
rect 35802 41460 35808 41472
rect 35176 41432 35808 41460
rect 35802 41420 35808 41432
rect 35860 41420 35866 41472
rect 36556 41460 36584 41500
rect 36630 41488 36636 41540
rect 36688 41528 36694 41540
rect 37369 41531 37427 41537
rect 37369 41528 37381 41531
rect 36688 41500 37381 41528
rect 36688 41488 36694 41500
rect 37369 41497 37381 41500
rect 37415 41497 37427 41531
rect 39666 41528 39672 41540
rect 38594 41500 39672 41528
rect 37369 41491 37427 41497
rect 36998 41460 37004 41472
rect 36556 41432 37004 41460
rect 36998 41420 37004 41432
rect 37056 41460 37062 41472
rect 38672 41460 38700 41500
rect 39666 41488 39672 41500
rect 39724 41488 39730 41540
rect 37056 41432 38700 41460
rect 37056 41420 37062 41432
rect 1104 41370 49864 41392
rect 1104 41318 7950 41370
rect 8002 41318 8014 41370
rect 8066 41318 8078 41370
rect 8130 41318 8142 41370
rect 8194 41318 8206 41370
rect 8258 41318 17950 41370
rect 18002 41318 18014 41370
rect 18066 41318 18078 41370
rect 18130 41318 18142 41370
rect 18194 41318 18206 41370
rect 18258 41318 27950 41370
rect 28002 41318 28014 41370
rect 28066 41318 28078 41370
rect 28130 41318 28142 41370
rect 28194 41318 28206 41370
rect 28258 41318 37950 41370
rect 38002 41318 38014 41370
rect 38066 41318 38078 41370
rect 38130 41318 38142 41370
rect 38194 41318 38206 41370
rect 38258 41318 47950 41370
rect 48002 41318 48014 41370
rect 48066 41318 48078 41370
rect 48130 41318 48142 41370
rect 48194 41318 48206 41370
rect 48258 41318 49864 41370
rect 1104 41296 49864 41318
rect 5810 41216 5816 41268
rect 5868 41216 5874 41268
rect 9858 41216 9864 41268
rect 9916 41216 9922 41268
rect 10778 41216 10784 41268
rect 10836 41216 10842 41268
rect 22005 41259 22063 41265
rect 22005 41225 22017 41259
rect 22051 41256 22063 41259
rect 22094 41256 22100 41268
rect 22051 41228 22100 41256
rect 22051 41225 22063 41228
rect 22005 41219 22063 41225
rect 22094 41216 22100 41228
rect 22152 41216 22158 41268
rect 22462 41216 22468 41268
rect 22520 41256 22526 41268
rect 24854 41256 24860 41268
rect 22520 41228 24860 41256
rect 22520 41216 22526 41228
rect 24854 41216 24860 41228
rect 24912 41216 24918 41268
rect 26050 41256 26056 41268
rect 25424 41228 26056 41256
rect 22186 41148 22192 41200
rect 22244 41188 22250 41200
rect 24872 41188 24900 41216
rect 25424 41188 25452 41228
rect 26050 41216 26056 41228
rect 26108 41256 26114 41268
rect 26108 41228 26372 41256
rect 26108 41216 26114 41228
rect 26344 41188 26372 41228
rect 27706 41216 27712 41268
rect 27764 41256 27770 41268
rect 29457 41259 29515 41265
rect 29457 41256 29469 41259
rect 27764 41228 29469 41256
rect 27764 41216 27770 41228
rect 29457 41225 29469 41228
rect 29503 41225 29515 41259
rect 29457 41219 29515 41225
rect 29546 41216 29552 41268
rect 29604 41256 29610 41268
rect 31938 41256 31944 41268
rect 29604 41228 31944 41256
rect 29604 41216 29610 41228
rect 31938 41216 31944 41228
rect 31996 41216 32002 41268
rect 27982 41188 27988 41200
rect 22244 41160 22692 41188
rect 24872 41160 25530 41188
rect 26344 41160 27988 41188
rect 22244 41148 22250 41160
rect 5718 41080 5724 41132
rect 5776 41080 5782 41132
rect 9766 41080 9772 41132
rect 9824 41080 9830 41132
rect 10686 41080 10692 41132
rect 10744 41080 10750 41132
rect 21269 41123 21327 41129
rect 21269 41120 21281 41123
rect 19306 41092 21281 41120
rect 1762 41012 1768 41064
rect 1820 41052 1826 41064
rect 19306 41052 19334 41092
rect 21269 41089 21281 41092
rect 21315 41120 21327 41123
rect 22370 41120 22376 41132
rect 21315 41092 22376 41120
rect 21315 41089 21327 41092
rect 21269 41083 21327 41089
rect 22370 41080 22376 41092
rect 22428 41080 22434 41132
rect 22664 41061 22692 41160
rect 27982 41148 27988 41160
rect 28040 41148 28046 41200
rect 29825 41191 29883 41197
rect 29825 41157 29837 41191
rect 29871 41188 29883 41191
rect 30834 41188 30840 41200
rect 29871 41160 30840 41188
rect 29871 41157 29883 41160
rect 29825 41151 29883 41157
rect 30834 41148 30840 41160
rect 30892 41148 30898 41200
rect 32858 41148 32864 41200
rect 32916 41188 32922 41200
rect 33413 41191 33471 41197
rect 33413 41188 33425 41191
rect 32916 41160 33425 41188
rect 32916 41148 32922 41160
rect 33413 41157 33425 41160
rect 33459 41157 33471 41191
rect 36998 41188 37004 41200
rect 34638 41174 37004 41188
rect 33413 41151 33471 41157
rect 34624 41160 37004 41174
rect 24118 41080 24124 41132
rect 24176 41120 24182 41132
rect 24578 41120 24584 41132
rect 24176 41092 24584 41120
rect 24176 41080 24182 41092
rect 24578 41080 24584 41092
rect 24636 41120 24642 41132
rect 24765 41123 24823 41129
rect 24765 41120 24777 41123
rect 24636 41092 24777 41120
rect 24636 41080 24642 41092
rect 24765 41089 24777 41092
rect 24811 41089 24823 41123
rect 24765 41083 24823 41089
rect 27246 41080 27252 41132
rect 27304 41080 27310 41132
rect 29917 41123 29975 41129
rect 29917 41089 29929 41123
rect 29963 41120 29975 41123
rect 32582 41120 32588 41132
rect 29963 41092 32588 41120
rect 29963 41089 29975 41092
rect 29917 41083 29975 41089
rect 32582 41080 32588 41092
rect 32640 41080 32646 41132
rect 1820 41024 19334 41052
rect 22465 41055 22523 41061
rect 1820 41012 1826 41024
rect 22465 41021 22477 41055
rect 22511 41021 22523 41055
rect 22465 41015 22523 41021
rect 22649 41055 22707 41061
rect 22649 41021 22661 41055
rect 22695 41052 22707 41055
rect 22738 41052 22744 41064
rect 22695 41024 22744 41052
rect 22695 41021 22707 41024
rect 22649 41015 22707 41021
rect 22480 40916 22508 41015
rect 22738 41012 22744 41024
rect 22796 41012 22802 41064
rect 25038 41012 25044 41064
rect 25096 41012 25102 41064
rect 26513 41055 26571 41061
rect 26513 41021 26525 41055
rect 26559 41052 26571 41055
rect 27522 41052 27528 41064
rect 26559 41024 27528 41052
rect 26559 41021 26571 41024
rect 26513 41015 26571 41021
rect 27522 41012 27528 41024
rect 27580 41012 27586 41064
rect 27982 41012 27988 41064
rect 28040 41052 28046 41064
rect 29086 41052 29092 41064
rect 28040 41024 29092 41052
rect 28040 41012 28046 41024
rect 29086 41012 29092 41024
rect 29144 41012 29150 41064
rect 30009 41055 30067 41061
rect 30009 41021 30021 41055
rect 30055 41021 30067 41055
rect 30009 41015 30067 41021
rect 29914 40944 29920 40996
rect 29972 40984 29978 40996
rect 30024 40984 30052 41015
rect 32306 41012 32312 41064
rect 32364 41052 32370 41064
rect 33137 41055 33195 41061
rect 33137 41052 33149 41055
rect 32364 41024 33149 41052
rect 32364 41012 32370 41024
rect 33137 41021 33149 41024
rect 33183 41021 33195 41055
rect 33137 41015 33195 41021
rect 29972 40956 30052 40984
rect 29972 40944 29978 40956
rect 22554 40916 22560 40928
rect 22480 40888 22560 40916
rect 22554 40876 22560 40888
rect 22612 40916 22618 40928
rect 22830 40916 22836 40928
rect 22612 40888 22836 40916
rect 22612 40876 22618 40888
rect 22830 40876 22836 40888
rect 22888 40916 22894 40928
rect 23201 40919 23259 40925
rect 23201 40916 23213 40919
rect 22888 40888 23213 40916
rect 22888 40876 22894 40888
rect 23201 40885 23213 40888
rect 23247 40885 23259 40919
rect 23201 40879 23259 40885
rect 28994 40876 29000 40928
rect 29052 40916 29058 40928
rect 29822 40916 29828 40928
rect 29052 40888 29828 40916
rect 29052 40876 29058 40888
rect 29822 40876 29828 40888
rect 29880 40876 29886 40928
rect 33042 40876 33048 40928
rect 33100 40916 33106 40928
rect 33594 40916 33600 40928
rect 33100 40888 33600 40916
rect 33100 40876 33106 40888
rect 33594 40876 33600 40888
rect 33652 40916 33658 40928
rect 34624 40916 34652 41160
rect 36998 41148 37004 41160
rect 37056 41148 37062 41200
rect 39850 41188 39856 41200
rect 39698 41160 39856 41188
rect 39850 41148 39856 41160
rect 39908 41148 39914 41200
rect 37826 41080 37832 41132
rect 37884 41120 37890 41132
rect 38197 41123 38255 41129
rect 38197 41120 38209 41123
rect 37884 41092 38209 41120
rect 37884 41080 37890 41092
rect 38197 41089 38209 41092
rect 38243 41089 38255 41123
rect 48777 41123 48835 41129
rect 48777 41120 48789 41123
rect 38197 41083 38255 41089
rect 45526 41092 48789 41120
rect 38930 41012 38936 41064
rect 38988 41052 38994 41064
rect 39942 41052 39948 41064
rect 38988 41024 39948 41052
rect 38988 41012 38994 41024
rect 39942 41012 39948 41024
rect 40000 41012 40006 41064
rect 45526 41052 45554 41092
rect 48777 41089 48789 41092
rect 48823 41089 48835 41123
rect 48777 41083 48835 41089
rect 41386 41024 45554 41052
rect 39482 40944 39488 40996
rect 39540 40984 39546 40996
rect 41386 40984 41414 41024
rect 48498 41012 48504 41064
rect 48556 41012 48562 41064
rect 39540 40956 41414 40984
rect 39540 40944 39546 40956
rect 33652 40888 34652 40916
rect 33652 40876 33658 40888
rect 34790 40876 34796 40928
rect 34848 40916 34854 40928
rect 34885 40919 34943 40925
rect 34885 40916 34897 40919
rect 34848 40888 34897 40916
rect 34848 40876 34854 40888
rect 34885 40885 34897 40888
rect 34931 40916 34943 40919
rect 35158 40916 35164 40928
rect 34931 40888 35164 40916
rect 34931 40885 34943 40888
rect 34885 40879 34943 40885
rect 35158 40876 35164 40888
rect 35216 40876 35222 40928
rect 38460 40919 38518 40925
rect 38460 40885 38472 40919
rect 38506 40916 38518 40919
rect 39206 40916 39212 40928
rect 38506 40888 39212 40916
rect 38506 40885 38518 40888
rect 38460 40879 38518 40885
rect 39206 40876 39212 40888
rect 39264 40916 39270 40928
rect 39758 40916 39764 40928
rect 39264 40888 39764 40916
rect 39264 40876 39270 40888
rect 39758 40876 39764 40888
rect 39816 40876 39822 40928
rect 39942 40876 39948 40928
rect 40000 40876 40006 40928
rect 1104 40826 49864 40848
rect 1104 40774 2950 40826
rect 3002 40774 3014 40826
rect 3066 40774 3078 40826
rect 3130 40774 3142 40826
rect 3194 40774 3206 40826
rect 3258 40774 12950 40826
rect 13002 40774 13014 40826
rect 13066 40774 13078 40826
rect 13130 40774 13142 40826
rect 13194 40774 13206 40826
rect 13258 40774 22950 40826
rect 23002 40774 23014 40826
rect 23066 40774 23078 40826
rect 23130 40774 23142 40826
rect 23194 40774 23206 40826
rect 23258 40774 32950 40826
rect 33002 40774 33014 40826
rect 33066 40774 33078 40826
rect 33130 40774 33142 40826
rect 33194 40774 33206 40826
rect 33258 40774 42950 40826
rect 43002 40774 43014 40826
rect 43066 40774 43078 40826
rect 43130 40774 43142 40826
rect 43194 40774 43206 40826
rect 43258 40774 49864 40826
rect 1104 40752 49864 40774
rect 20530 40672 20536 40724
rect 20588 40712 20594 40724
rect 23293 40715 23351 40721
rect 23293 40712 23305 40715
rect 20588 40684 23305 40712
rect 20588 40672 20594 40684
rect 23293 40681 23305 40684
rect 23339 40681 23351 40715
rect 29546 40712 29552 40724
rect 23293 40675 23351 40681
rect 25976 40684 29552 40712
rect 22002 40604 22008 40656
rect 22060 40644 22066 40656
rect 25501 40647 25559 40653
rect 25501 40644 25513 40647
rect 22060 40616 25513 40644
rect 22060 40604 22066 40616
rect 25501 40613 25513 40616
rect 25547 40613 25559 40647
rect 25501 40607 25559 40613
rect 23937 40579 23995 40585
rect 23937 40545 23949 40579
rect 23983 40576 23995 40579
rect 25038 40576 25044 40588
rect 23983 40548 25044 40576
rect 23983 40545 23995 40548
rect 23937 40539 23995 40545
rect 25038 40536 25044 40548
rect 25096 40536 25102 40588
rect 25976 40585 26004 40684
rect 29546 40672 29552 40684
rect 29604 40672 29610 40724
rect 31018 40712 31024 40724
rect 29656 40684 31024 40712
rect 28994 40644 29000 40656
rect 26160 40616 29000 40644
rect 26160 40585 26188 40616
rect 28994 40604 29000 40616
rect 29052 40604 29058 40656
rect 25961 40579 26019 40585
rect 25961 40545 25973 40579
rect 26007 40545 26019 40579
rect 25961 40539 26019 40545
rect 26145 40579 26203 40585
rect 26145 40545 26157 40579
rect 26191 40545 26203 40579
rect 26145 40539 26203 40545
rect 27246 40536 27252 40588
rect 27304 40536 27310 40588
rect 22738 40468 22744 40520
rect 22796 40508 22802 40520
rect 24302 40508 24308 40520
rect 22796 40480 24308 40508
rect 22796 40468 22802 40480
rect 24302 40468 24308 40480
rect 24360 40508 24366 40520
rect 24360 40480 26004 40508
rect 24360 40468 24366 40480
rect 23382 40400 23388 40452
rect 23440 40440 23446 40452
rect 25869 40443 25927 40449
rect 25869 40440 25881 40443
rect 23440 40412 25881 40440
rect 23440 40400 23446 40412
rect 25869 40409 25881 40412
rect 25915 40409 25927 40443
rect 25976 40440 26004 40480
rect 27062 40468 27068 40520
rect 27120 40468 27126 40520
rect 29656 40440 29684 40684
rect 31018 40672 31024 40684
rect 31076 40712 31082 40724
rect 31076 40684 31754 40712
rect 31076 40672 31082 40684
rect 31726 40644 31754 40684
rect 35066 40672 35072 40724
rect 35124 40712 35130 40724
rect 35253 40715 35311 40721
rect 35253 40712 35265 40715
rect 35124 40684 35265 40712
rect 35124 40672 35130 40684
rect 35253 40681 35265 40684
rect 35299 40681 35311 40715
rect 35253 40675 35311 40681
rect 38749 40715 38807 40721
rect 38749 40681 38761 40715
rect 38795 40712 38807 40715
rect 39574 40712 39580 40724
rect 38795 40684 39580 40712
rect 38795 40681 38807 40684
rect 38749 40675 38807 40681
rect 39574 40672 39580 40684
rect 39632 40672 39638 40724
rect 31726 40616 35848 40644
rect 30009 40579 30067 40585
rect 30009 40545 30021 40579
rect 30055 40576 30067 40579
rect 31018 40576 31024 40588
rect 30055 40548 31024 40576
rect 30055 40545 30067 40548
rect 30009 40539 30067 40545
rect 31018 40536 31024 40548
rect 31076 40536 31082 40588
rect 32674 40536 32680 40588
rect 32732 40536 32738 40588
rect 32766 40536 32772 40588
rect 32824 40536 32830 40588
rect 33502 40536 33508 40588
rect 33560 40576 33566 40588
rect 34057 40579 34115 40585
rect 34057 40576 34069 40579
rect 33560 40548 34069 40576
rect 33560 40536 33566 40548
rect 34057 40545 34069 40548
rect 34103 40545 34115 40579
rect 34057 40539 34115 40545
rect 34146 40536 34152 40588
rect 34204 40536 34210 40588
rect 35820 40585 35848 40616
rect 35805 40579 35863 40585
rect 35805 40545 35817 40579
rect 35851 40545 35863 40579
rect 35805 40539 35863 40545
rect 38746 40536 38752 40588
rect 38804 40576 38810 40588
rect 39209 40579 39267 40585
rect 39209 40576 39221 40579
rect 38804 40548 39221 40576
rect 38804 40536 38810 40548
rect 39209 40545 39221 40548
rect 39255 40545 39267 40579
rect 39209 40539 39267 40545
rect 39390 40536 39396 40588
rect 39448 40576 39454 40588
rect 39942 40576 39948 40588
rect 39448 40548 39948 40576
rect 39448 40536 39454 40548
rect 39942 40536 39948 40548
rect 40000 40536 40006 40588
rect 48774 40536 48780 40588
rect 48832 40536 48838 40588
rect 29730 40468 29736 40520
rect 29788 40468 29794 40520
rect 32585 40511 32643 40517
rect 32585 40477 32597 40511
rect 32631 40508 32643 40511
rect 35713 40511 35771 40517
rect 32631 40480 35572 40508
rect 32631 40477 32643 40480
rect 32585 40471 32643 40477
rect 31662 40440 31668 40452
rect 25976 40412 29684 40440
rect 31234 40412 31668 40440
rect 25869 40403 25927 40409
rect 31662 40400 31668 40412
rect 31720 40400 31726 40452
rect 33318 40440 33324 40452
rect 32232 40412 33324 40440
rect 22094 40332 22100 40384
rect 22152 40372 22158 40384
rect 23661 40375 23719 40381
rect 23661 40372 23673 40375
rect 22152 40344 23673 40372
rect 22152 40332 22158 40344
rect 23661 40341 23673 40344
rect 23707 40341 23719 40375
rect 23661 40335 23719 40341
rect 23753 40375 23811 40381
rect 23753 40341 23765 40375
rect 23799 40372 23811 40375
rect 26602 40372 26608 40384
rect 23799 40344 26608 40372
rect 23799 40341 23811 40344
rect 23753 40335 23811 40341
rect 26602 40332 26608 40344
rect 26660 40332 26666 40384
rect 26694 40332 26700 40384
rect 26752 40332 26758 40384
rect 27062 40332 27068 40384
rect 27120 40372 27126 40384
rect 27157 40375 27215 40381
rect 27157 40372 27169 40375
rect 27120 40344 27169 40372
rect 27120 40332 27126 40344
rect 27157 40341 27169 40344
rect 27203 40341 27215 40375
rect 27157 40335 27215 40341
rect 29914 40332 29920 40384
rect 29972 40372 29978 40384
rect 32232 40381 32260 40412
rect 33318 40400 33324 40412
rect 33376 40400 33382 40452
rect 33962 40400 33968 40452
rect 34020 40400 34026 40452
rect 31481 40375 31539 40381
rect 31481 40372 31493 40375
rect 29972 40344 31493 40372
rect 29972 40332 29978 40344
rect 31481 40341 31493 40344
rect 31527 40341 31539 40375
rect 31481 40335 31539 40341
rect 32217 40375 32275 40381
rect 32217 40341 32229 40375
rect 32263 40341 32275 40375
rect 32217 40335 32275 40341
rect 33597 40375 33655 40381
rect 33597 40341 33609 40375
rect 33643 40372 33655 40375
rect 33870 40372 33876 40384
rect 33643 40344 33876 40372
rect 33643 40341 33655 40344
rect 33597 40335 33655 40341
rect 33870 40332 33876 40344
rect 33928 40332 33934 40384
rect 35544 40372 35572 40480
rect 35713 40477 35725 40511
rect 35759 40508 35771 40511
rect 37734 40508 37740 40520
rect 35759 40480 37740 40508
rect 35759 40477 35771 40480
rect 35713 40471 35771 40477
rect 37734 40468 37740 40480
rect 37792 40508 37798 40520
rect 38562 40508 38568 40520
rect 37792 40480 38568 40508
rect 37792 40468 37798 40480
rect 38562 40468 38568 40480
rect 38620 40468 38626 40520
rect 48498 40468 48504 40520
rect 48556 40468 48562 40520
rect 35621 40443 35679 40449
rect 35621 40409 35633 40443
rect 35667 40440 35679 40443
rect 39942 40440 39948 40452
rect 35667 40412 39948 40440
rect 35667 40409 35679 40412
rect 35621 40403 35679 40409
rect 39942 40400 39948 40412
rect 40000 40400 40006 40452
rect 37366 40372 37372 40384
rect 35544 40344 37372 40372
rect 37366 40332 37372 40344
rect 37424 40332 37430 40384
rect 39114 40332 39120 40384
rect 39172 40332 39178 40384
rect 1104 40282 49864 40304
rect 1104 40230 7950 40282
rect 8002 40230 8014 40282
rect 8066 40230 8078 40282
rect 8130 40230 8142 40282
rect 8194 40230 8206 40282
rect 8258 40230 17950 40282
rect 18002 40230 18014 40282
rect 18066 40230 18078 40282
rect 18130 40230 18142 40282
rect 18194 40230 18206 40282
rect 18258 40230 27950 40282
rect 28002 40230 28014 40282
rect 28066 40230 28078 40282
rect 28130 40230 28142 40282
rect 28194 40230 28206 40282
rect 28258 40230 37950 40282
rect 38002 40230 38014 40282
rect 38066 40230 38078 40282
rect 38130 40230 38142 40282
rect 38194 40230 38206 40282
rect 38258 40230 47950 40282
rect 48002 40230 48014 40282
rect 48066 40230 48078 40282
rect 48130 40230 48142 40282
rect 48194 40230 48206 40282
rect 48258 40230 49864 40282
rect 1104 40208 49864 40230
rect 25038 40128 25044 40180
rect 25096 40128 25102 40180
rect 31662 40168 31668 40180
rect 29564 40140 31668 40168
rect 24854 40100 24860 40112
rect 24794 40072 24860 40100
rect 24854 40060 24860 40072
rect 24912 40060 24918 40112
rect 29564 40018 29592 40140
rect 31662 40128 31668 40140
rect 31720 40128 31726 40180
rect 32766 40128 32772 40180
rect 32824 40168 32830 40180
rect 35250 40168 35256 40180
rect 32824 40140 35256 40168
rect 32824 40128 32830 40140
rect 35250 40128 35256 40140
rect 35308 40168 35314 40180
rect 35618 40168 35624 40180
rect 35308 40140 35624 40168
rect 35308 40128 35314 40140
rect 35618 40128 35624 40140
rect 35676 40128 35682 40180
rect 35894 40128 35900 40180
rect 35952 40168 35958 40180
rect 36449 40171 36507 40177
rect 36449 40168 36461 40171
rect 35952 40140 36461 40168
rect 35952 40128 35958 40140
rect 36449 40137 36461 40140
rect 36495 40168 36507 40171
rect 36814 40168 36820 40180
rect 36495 40140 36820 40168
rect 36495 40137 36507 40140
rect 36449 40131 36507 40137
rect 36814 40128 36820 40140
rect 36872 40128 36878 40180
rect 39850 40128 39856 40180
rect 39908 40168 39914 40180
rect 39908 40140 39988 40168
rect 39908 40128 39914 40140
rect 29730 40060 29736 40112
rect 29788 40060 29794 40112
rect 33594 40060 33600 40112
rect 33652 40060 33658 40112
rect 34514 40100 34520 40112
rect 34072 40072 34520 40100
rect 29748 40032 29776 40060
rect 31294 40032 31300 40044
rect 29748 40004 31300 40032
rect 21082 39924 21088 39976
rect 21140 39964 21146 39976
rect 23293 39967 23351 39973
rect 23293 39964 23305 39967
rect 21140 39936 23305 39964
rect 21140 39924 21146 39936
rect 23293 39933 23305 39936
rect 23339 39933 23351 39967
rect 23293 39927 23351 39933
rect 23566 39924 23572 39976
rect 23624 39924 23630 39976
rect 28169 39967 28227 39973
rect 28169 39933 28181 39967
rect 28215 39964 28227 39967
rect 28445 39967 28503 39973
rect 28215 39936 28304 39964
rect 28215 39933 28227 39936
rect 28169 39927 28227 39933
rect 24670 39856 24676 39908
rect 24728 39896 24734 39908
rect 27706 39896 27712 39908
rect 24728 39868 27712 39896
rect 24728 39856 24734 39868
rect 27706 39856 27712 39868
rect 27764 39856 27770 39908
rect 22462 39788 22468 39840
rect 22520 39828 22526 39840
rect 26050 39828 26056 39840
rect 22520 39800 26056 39828
rect 22520 39788 22526 39800
rect 26050 39788 26056 39800
rect 26108 39788 26114 39840
rect 28276 39828 28304 39936
rect 28445 39933 28457 39967
rect 28491 39964 28503 39967
rect 28902 39964 28908 39976
rect 28491 39936 28908 39964
rect 28491 39933 28503 39936
rect 28445 39927 28503 39933
rect 28902 39924 28908 39936
rect 28960 39924 28966 39976
rect 29748 39828 29776 40004
rect 31294 39992 31300 40004
rect 31352 40032 31358 40044
rect 32306 40032 32312 40044
rect 31352 40004 32312 40032
rect 31352 39992 31358 40004
rect 32306 39992 32312 40004
rect 32364 39992 32370 40044
rect 34072 39973 34100 40072
rect 34514 40060 34520 40072
rect 34572 40060 34578 40112
rect 36998 40100 37004 40112
rect 36202 40072 37004 40100
rect 36998 40060 37004 40072
rect 37056 40060 37062 40112
rect 34698 39992 34704 40044
rect 34756 39992 34762 40044
rect 37826 39992 37832 40044
rect 37884 40032 37890 40044
rect 38562 40032 38568 40044
rect 37884 40004 38568 40032
rect 37884 39992 37890 40004
rect 38562 39992 38568 40004
rect 38620 39992 38626 40044
rect 39960 40032 39988 40140
rect 40310 40128 40316 40180
rect 40368 40128 40374 40180
rect 40773 40171 40831 40177
rect 40773 40137 40785 40171
rect 40819 40168 40831 40171
rect 42426 40168 42432 40180
rect 40819 40140 42432 40168
rect 40819 40137 40831 40140
rect 40773 40131 40831 40137
rect 42426 40128 42432 40140
rect 42484 40128 42490 40180
rect 41138 40060 41144 40112
rect 41196 40060 41202 40112
rect 39960 40018 40080 40032
rect 39974 40004 40080 40018
rect 32585 39967 32643 39973
rect 32585 39964 32597 39967
rect 32140 39936 32597 39964
rect 29822 39856 29828 39908
rect 29880 39896 29886 39908
rect 32140 39896 32168 39936
rect 32585 39933 32597 39936
rect 32631 39933 32643 39967
rect 32585 39927 32643 39933
rect 34057 39967 34115 39973
rect 34057 39933 34069 39967
rect 34103 39933 34115 39967
rect 34977 39967 35035 39973
rect 34977 39964 34989 39967
rect 34057 39927 34115 39933
rect 34808 39936 34989 39964
rect 29880 39868 32168 39896
rect 29880 39856 29886 39868
rect 33778 39856 33784 39908
rect 33836 39896 33842 39908
rect 34808 39896 34836 39936
rect 34977 39933 34989 39936
rect 35023 39964 35035 39967
rect 36446 39964 36452 39976
rect 35023 39936 36452 39964
rect 35023 39933 35035 39936
rect 34977 39927 35035 39933
rect 36446 39924 36452 39936
rect 36504 39964 36510 39976
rect 36722 39964 36728 39976
rect 36504 39936 36728 39964
rect 36504 39924 36510 39936
rect 36722 39924 36728 39936
rect 36780 39924 36786 39976
rect 38841 39967 38899 39973
rect 38841 39933 38853 39967
rect 38887 39964 38899 39967
rect 39390 39964 39396 39976
rect 38887 39936 39396 39964
rect 38887 39933 38899 39936
rect 38841 39927 38899 39933
rect 39390 39924 39396 39936
rect 39448 39924 39454 39976
rect 33836 39868 34836 39896
rect 40052 39896 40080 40004
rect 41230 39992 41236 40044
rect 41288 39992 41294 40044
rect 41417 39967 41475 39973
rect 41417 39933 41429 39967
rect 41463 39964 41475 39967
rect 41690 39964 41696 39976
rect 41463 39936 41696 39964
rect 41463 39933 41475 39936
rect 41417 39927 41475 39933
rect 41690 39924 41696 39936
rect 41748 39924 41754 39976
rect 48498 39924 48504 39976
rect 48556 39924 48562 39976
rect 48590 39924 48596 39976
rect 48648 39964 48654 39976
rect 48777 39967 48835 39973
rect 48777 39964 48789 39967
rect 48648 39936 48789 39964
rect 48648 39924 48654 39936
rect 48777 39933 48789 39936
rect 48823 39933 48835 39967
rect 48777 39927 48835 39933
rect 41874 39896 41880 39908
rect 40052 39868 41880 39896
rect 33836 39856 33842 39868
rect 41874 39856 41880 39868
rect 41932 39856 41938 39908
rect 28276 39800 29776 39828
rect 29917 39831 29975 39837
rect 29917 39797 29929 39831
rect 29963 39828 29975 39831
rect 30190 39828 30196 39840
rect 29963 39800 30196 39828
rect 29963 39797 29975 39800
rect 29917 39791 29975 39797
rect 30190 39788 30196 39800
rect 30248 39788 30254 39840
rect 30282 39788 30288 39840
rect 30340 39828 30346 39840
rect 31570 39828 31576 39840
rect 30340 39800 31576 39828
rect 30340 39788 30346 39800
rect 31570 39788 31576 39800
rect 31628 39788 31634 39840
rect 34790 39788 34796 39840
rect 34848 39828 34854 39840
rect 40954 39828 40960 39840
rect 34848 39800 40960 39828
rect 34848 39788 34854 39800
rect 40954 39788 40960 39800
rect 41012 39788 41018 39840
rect 1104 39738 49864 39760
rect 1104 39686 2950 39738
rect 3002 39686 3014 39738
rect 3066 39686 3078 39738
rect 3130 39686 3142 39738
rect 3194 39686 3206 39738
rect 3258 39686 12950 39738
rect 13002 39686 13014 39738
rect 13066 39686 13078 39738
rect 13130 39686 13142 39738
rect 13194 39686 13206 39738
rect 13258 39686 22950 39738
rect 23002 39686 23014 39738
rect 23066 39686 23078 39738
rect 23130 39686 23142 39738
rect 23194 39686 23206 39738
rect 23258 39686 32950 39738
rect 33002 39686 33014 39738
rect 33066 39686 33078 39738
rect 33130 39686 33142 39738
rect 33194 39686 33206 39738
rect 33258 39686 42950 39738
rect 43002 39686 43014 39738
rect 43066 39686 43078 39738
rect 43130 39686 43142 39738
rect 43194 39686 43206 39738
rect 43258 39686 49864 39738
rect 1104 39664 49864 39686
rect 22005 39627 22063 39633
rect 22005 39593 22017 39627
rect 22051 39624 22063 39627
rect 25958 39624 25964 39636
rect 22051 39596 25964 39624
rect 22051 39593 22063 39596
rect 22005 39587 22063 39593
rect 25958 39584 25964 39596
rect 26016 39584 26022 39636
rect 29178 39584 29184 39636
rect 29236 39624 29242 39636
rect 29638 39624 29644 39636
rect 29236 39596 29644 39624
rect 29236 39584 29242 39596
rect 29638 39584 29644 39596
rect 29696 39624 29702 39636
rect 30282 39624 30288 39636
rect 29696 39596 30288 39624
rect 29696 39584 29702 39596
rect 30282 39584 30288 39596
rect 30340 39624 30346 39636
rect 30450 39627 30508 39633
rect 30450 39624 30462 39627
rect 30340 39596 30462 39624
rect 30340 39584 30346 39596
rect 30450 39593 30462 39596
rect 30496 39593 30508 39627
rect 30450 39587 30508 39593
rect 31018 39584 31024 39636
rect 31076 39624 31082 39636
rect 31478 39624 31484 39636
rect 31076 39596 31484 39624
rect 31076 39584 31082 39596
rect 31478 39584 31484 39596
rect 31536 39624 31542 39636
rect 31536 39596 31984 39624
rect 31536 39584 31542 39596
rect 26050 39516 26056 39568
rect 26108 39556 26114 39568
rect 26108 39528 28580 39556
rect 26108 39516 26114 39528
rect 22462 39488 22468 39500
rect 22066 39460 22468 39488
rect 1854 39244 1860 39296
rect 1912 39284 1918 39296
rect 21453 39287 21511 39293
rect 21453 39284 21465 39287
rect 1912 39256 21465 39284
rect 1912 39244 1918 39256
rect 21453 39253 21465 39256
rect 21499 39284 21511 39287
rect 22066 39284 22094 39460
rect 22462 39448 22468 39460
rect 22520 39448 22526 39500
rect 22557 39491 22615 39497
rect 22557 39457 22569 39491
rect 22603 39457 22615 39491
rect 22557 39451 22615 39457
rect 22186 39380 22192 39432
rect 22244 39420 22250 39432
rect 22572 39420 22600 39451
rect 24578 39448 24584 39500
rect 24636 39448 24642 39500
rect 24857 39491 24915 39497
rect 24857 39457 24869 39491
rect 24903 39488 24915 39491
rect 25222 39488 25228 39500
rect 24903 39460 25228 39488
rect 24903 39457 24915 39460
rect 24857 39451 24915 39457
rect 25222 39448 25228 39460
rect 25280 39488 25286 39500
rect 28442 39488 28448 39500
rect 25280 39460 28448 39488
rect 25280 39448 25286 39460
rect 28442 39448 28448 39460
rect 28500 39448 28506 39500
rect 28552 39488 28580 39528
rect 31570 39516 31576 39568
rect 31628 39556 31634 39568
rect 31628 39528 31708 39556
rect 31628 39516 31634 39528
rect 31110 39488 31116 39500
rect 28552 39460 31116 39488
rect 31110 39448 31116 39460
rect 31168 39448 31174 39500
rect 22244 39392 22600 39420
rect 22244 39380 22250 39392
rect 26142 39380 26148 39432
rect 26200 39420 26206 39432
rect 28718 39420 28724 39432
rect 26200 39392 28724 39420
rect 26200 39380 26206 39392
rect 28718 39380 28724 39392
rect 28776 39380 28782 39432
rect 30098 39380 30104 39432
rect 30156 39420 30162 39432
rect 30193 39423 30251 39429
rect 30193 39420 30205 39423
rect 30156 39392 30205 39420
rect 30156 39380 30162 39392
rect 30193 39389 30205 39392
rect 30239 39389 30251 39423
rect 30193 39383 30251 39389
rect 31570 39380 31576 39432
rect 31628 39380 31634 39432
rect 31680 39420 31708 39528
rect 31956 39497 31984 39596
rect 32582 39584 32588 39636
rect 32640 39584 32646 39636
rect 34330 39584 34336 39636
rect 34388 39624 34394 39636
rect 39206 39624 39212 39636
rect 34388 39596 39212 39624
rect 34388 39584 34394 39596
rect 39206 39584 39212 39596
rect 39264 39584 39270 39636
rect 39850 39584 39856 39636
rect 39908 39624 39914 39636
rect 42613 39627 42671 39633
rect 42613 39624 42625 39627
rect 39908 39596 42625 39624
rect 39908 39584 39914 39596
rect 42613 39593 42625 39596
rect 42659 39593 42671 39627
rect 42613 39587 42671 39593
rect 32214 39516 32220 39568
rect 32272 39556 32278 39568
rect 35986 39556 35992 39568
rect 32272 39528 35992 39556
rect 32272 39516 32278 39528
rect 35986 39516 35992 39528
rect 36044 39516 36050 39568
rect 38470 39516 38476 39568
rect 38528 39556 38534 39568
rect 38838 39556 38844 39568
rect 38528 39528 38844 39556
rect 38528 39516 38534 39528
rect 38838 39516 38844 39528
rect 38896 39516 38902 39568
rect 48958 39556 48964 39568
rect 45526 39528 48964 39556
rect 31941 39491 31999 39497
rect 31941 39457 31953 39491
rect 31987 39488 31999 39491
rect 33137 39491 33195 39497
rect 33137 39488 33149 39491
rect 31987 39460 33149 39488
rect 31987 39457 31999 39460
rect 31941 39451 31999 39457
rect 33137 39457 33149 39460
rect 33183 39457 33195 39491
rect 33137 39451 33195 39457
rect 36265 39491 36323 39497
rect 36265 39457 36277 39491
rect 36311 39488 36323 39491
rect 38286 39488 38292 39500
rect 36311 39460 38292 39488
rect 36311 39457 36323 39460
rect 36265 39451 36323 39457
rect 38286 39448 38292 39460
rect 38344 39448 38350 39500
rect 41141 39491 41199 39497
rect 41141 39457 41153 39491
rect 41187 39488 41199 39491
rect 42794 39488 42800 39500
rect 41187 39460 42800 39488
rect 41187 39457 41199 39460
rect 41141 39451 41199 39457
rect 42794 39448 42800 39460
rect 42852 39448 42858 39500
rect 45526 39488 45554 39528
rect 48958 39516 48964 39528
rect 49016 39516 49022 39568
rect 42904 39460 45554 39488
rect 34330 39420 34336 39432
rect 31680 39392 34336 39420
rect 34330 39380 34336 39392
rect 34388 39380 34394 39432
rect 34698 39380 34704 39432
rect 34756 39420 34762 39432
rect 35989 39423 36047 39429
rect 35989 39420 36001 39423
rect 34756 39392 36001 39420
rect 34756 39380 34762 39392
rect 35989 39389 36001 39392
rect 36035 39389 36047 39423
rect 35989 39383 36047 39389
rect 38473 39423 38531 39429
rect 38473 39389 38485 39423
rect 38519 39420 38531 39423
rect 38838 39420 38844 39432
rect 38519 39392 38844 39420
rect 38519 39389 38531 39392
rect 38473 39383 38531 39389
rect 38838 39380 38844 39392
rect 38896 39380 38902 39432
rect 40862 39380 40868 39432
rect 40920 39380 40926 39432
rect 24854 39312 24860 39364
rect 24912 39352 24918 39364
rect 24912 39324 25346 39352
rect 24912 39312 24918 39324
rect 26970 39312 26976 39364
rect 27028 39352 27034 39364
rect 32953 39355 33011 39361
rect 27028 39324 30420 39352
rect 27028 39312 27034 39324
rect 21499 39256 22094 39284
rect 21499 39253 21511 39256
rect 21453 39247 21511 39253
rect 22370 39244 22376 39296
rect 22428 39244 22434 39296
rect 23566 39244 23572 39296
rect 23624 39284 23630 39296
rect 26329 39287 26387 39293
rect 26329 39284 26341 39287
rect 23624 39256 26341 39284
rect 23624 39244 23630 39256
rect 26329 39253 26341 39256
rect 26375 39284 26387 39287
rect 28810 39284 28816 39296
rect 26375 39256 28816 39284
rect 26375 39253 26387 39256
rect 26329 39247 26387 39253
rect 28810 39244 28816 39256
rect 28868 39244 28874 39296
rect 30392 39284 30420 39324
rect 32953 39321 32965 39355
rect 32999 39352 33011 39355
rect 32999 39324 36676 39352
rect 32999 39321 33011 39324
rect 32953 39315 33011 39321
rect 30742 39284 30748 39296
rect 30392 39256 30748 39284
rect 30742 39244 30748 39256
rect 30800 39244 30806 39296
rect 33045 39287 33103 39293
rect 33045 39253 33057 39287
rect 33091 39284 33103 39287
rect 33594 39284 33600 39296
rect 33091 39256 33600 39284
rect 33091 39253 33103 39256
rect 33045 39247 33103 39253
rect 33594 39244 33600 39256
rect 33652 39244 33658 39296
rect 36648 39284 36676 39324
rect 36998 39312 37004 39364
rect 37056 39312 37062 39364
rect 37550 39312 37556 39364
rect 37608 39352 37614 39364
rect 41414 39352 41420 39364
rect 37608 39324 41420 39352
rect 37608 39312 37614 39324
rect 41414 39312 41420 39324
rect 41472 39312 41478 39364
rect 42610 39352 42616 39364
rect 42366 39324 42616 39352
rect 42610 39312 42616 39324
rect 42668 39312 42674 39364
rect 37642 39284 37648 39296
rect 36648 39256 37648 39284
rect 37642 39244 37648 39256
rect 37700 39244 37706 39296
rect 37737 39287 37795 39293
rect 37737 39253 37749 39287
rect 37783 39284 37795 39287
rect 37826 39284 37832 39296
rect 37783 39256 37832 39284
rect 37783 39253 37795 39256
rect 37737 39247 37795 39253
rect 37826 39244 37832 39256
rect 37884 39244 37890 39296
rect 39666 39244 39672 39296
rect 39724 39284 39730 39296
rect 42904 39284 42932 39460
rect 48774 39448 48780 39500
rect 48832 39448 48838 39500
rect 43990 39380 43996 39432
rect 44048 39420 44054 39432
rect 46934 39420 46940 39432
rect 44048 39392 46940 39420
rect 44048 39380 44054 39392
rect 46934 39380 46940 39392
rect 46992 39380 46998 39432
rect 48498 39380 48504 39432
rect 48556 39380 48562 39432
rect 39724 39256 42932 39284
rect 39724 39244 39730 39256
rect 1104 39194 49864 39216
rect 1104 39142 7950 39194
rect 8002 39142 8014 39194
rect 8066 39142 8078 39194
rect 8130 39142 8142 39194
rect 8194 39142 8206 39194
rect 8258 39142 17950 39194
rect 18002 39142 18014 39194
rect 18066 39142 18078 39194
rect 18130 39142 18142 39194
rect 18194 39142 18206 39194
rect 18258 39142 27950 39194
rect 28002 39142 28014 39194
rect 28066 39142 28078 39194
rect 28130 39142 28142 39194
rect 28194 39142 28206 39194
rect 28258 39142 37950 39194
rect 38002 39142 38014 39194
rect 38066 39142 38078 39194
rect 38130 39142 38142 39194
rect 38194 39142 38206 39194
rect 38258 39142 47950 39194
rect 48002 39142 48014 39194
rect 48066 39142 48078 39194
rect 48130 39142 48142 39194
rect 48194 39142 48206 39194
rect 48258 39142 49864 39194
rect 1104 39120 49864 39142
rect 24486 39040 24492 39092
rect 24544 39040 24550 39092
rect 24578 39040 24584 39092
rect 24636 39080 24642 39092
rect 25038 39080 25044 39092
rect 24636 39052 25044 39080
rect 24636 39040 24642 39052
rect 25038 39040 25044 39052
rect 25096 39040 25102 39092
rect 25866 39040 25872 39092
rect 25924 39040 25930 39092
rect 26329 39083 26387 39089
rect 26329 39049 26341 39083
rect 26375 39080 26387 39083
rect 26970 39080 26976 39092
rect 26375 39052 26976 39080
rect 26375 39049 26387 39052
rect 26329 39043 26387 39049
rect 26970 39040 26976 39052
rect 27028 39040 27034 39092
rect 27154 39040 27160 39092
rect 27212 39080 27218 39092
rect 27341 39083 27399 39089
rect 27341 39080 27353 39083
rect 27212 39052 27353 39080
rect 27212 39040 27218 39052
rect 27341 39049 27353 39052
rect 27387 39049 27399 39083
rect 27341 39043 27399 39049
rect 28905 39083 28963 39089
rect 28905 39049 28917 39083
rect 28951 39080 28963 39083
rect 32214 39080 32220 39092
rect 28951 39052 32220 39080
rect 28951 39049 28963 39052
rect 28905 39043 28963 39049
rect 32214 39040 32220 39052
rect 32272 39040 32278 39092
rect 32398 39040 32404 39092
rect 32456 39040 32462 39092
rect 33594 39040 33600 39092
rect 33652 39040 33658 39092
rect 33965 39083 34023 39089
rect 33965 39049 33977 39083
rect 34011 39080 34023 39083
rect 34790 39080 34796 39092
rect 34011 39052 34796 39080
rect 34011 39049 34023 39052
rect 33965 39043 34023 39049
rect 34790 39040 34796 39052
rect 34848 39040 34854 39092
rect 34882 39040 34888 39092
rect 34940 39080 34946 39092
rect 35437 39083 35495 39089
rect 35437 39080 35449 39083
rect 34940 39052 35449 39080
rect 34940 39040 34946 39052
rect 35437 39049 35449 39052
rect 35483 39049 35495 39083
rect 35437 39043 35495 39049
rect 36170 39040 36176 39092
rect 36228 39080 36234 39092
rect 36633 39083 36691 39089
rect 36633 39080 36645 39083
rect 36228 39052 36645 39080
rect 36228 39040 36234 39052
rect 36633 39049 36645 39052
rect 36679 39049 36691 39083
rect 36633 39043 36691 39049
rect 37274 39040 37280 39092
rect 37332 39080 37338 39092
rect 37921 39083 37979 39089
rect 37921 39080 37933 39083
rect 37332 39052 37933 39080
rect 37332 39040 37338 39052
rect 37921 39049 37933 39052
rect 37967 39049 37979 39083
rect 37921 39043 37979 39049
rect 38838 39040 38844 39092
rect 38896 39040 38902 39092
rect 39114 39040 39120 39092
rect 39172 39080 39178 39092
rect 39301 39083 39359 39089
rect 39301 39080 39313 39083
rect 39172 39052 39313 39080
rect 39172 39040 39178 39052
rect 39301 39049 39313 39052
rect 39347 39049 39359 39083
rect 39301 39043 39359 39049
rect 40034 39040 40040 39092
rect 40092 39080 40098 39092
rect 40770 39080 40776 39092
rect 40092 39052 40776 39080
rect 40092 39040 40098 39052
rect 40770 39040 40776 39052
rect 40828 39040 40834 39092
rect 41414 39040 41420 39092
rect 41472 39080 41478 39092
rect 42058 39080 42064 39092
rect 41472 39052 42064 39080
rect 41472 39040 41478 39052
rect 42058 39040 42064 39052
rect 42116 39040 42122 39092
rect 22830 38972 22836 39024
rect 22888 39012 22894 39024
rect 23293 39015 23351 39021
rect 23293 39012 23305 39015
rect 22888 38984 23305 39012
rect 22888 38972 22894 38984
rect 23293 38981 23305 38984
rect 23339 39012 23351 39015
rect 24670 39012 24676 39024
rect 23339 38984 24676 39012
rect 23339 38981 23351 38984
rect 23293 38975 23351 38981
rect 24670 38972 24676 38984
rect 24728 38972 24734 39024
rect 24854 38972 24860 39024
rect 24912 38972 24918 39024
rect 24949 39015 25007 39021
rect 24949 38981 24961 39015
rect 24995 39012 25007 39015
rect 27062 39012 27068 39024
rect 24995 38984 27068 39012
rect 24995 38981 25007 38984
rect 24949 38975 25007 38981
rect 27062 38972 27068 38984
rect 27120 38972 27126 39024
rect 27801 39015 27859 39021
rect 27801 38981 27813 39015
rect 27847 39012 27859 39015
rect 29822 39012 29828 39024
rect 27847 38984 29828 39012
rect 27847 38981 27859 38984
rect 27801 38975 27859 38981
rect 29822 38972 29828 38984
rect 29880 38972 29886 39024
rect 31573 39015 31631 39021
rect 31573 38981 31585 39015
rect 31619 39012 31631 39015
rect 32769 39015 32827 39021
rect 32769 39012 32781 39015
rect 31619 38984 32781 39012
rect 31619 38981 31631 38984
rect 31573 38975 31631 38981
rect 32769 38981 32781 38984
rect 32815 39012 32827 39015
rect 37550 39012 37556 39024
rect 32815 38984 37556 39012
rect 32815 38981 32827 38984
rect 32769 38975 32827 38981
rect 37550 38972 37556 38984
rect 37608 38972 37614 39024
rect 38562 38972 38568 39024
rect 38620 39012 38626 39024
rect 40862 39012 40868 39024
rect 38620 38984 40868 39012
rect 38620 38972 38626 38984
rect 934 38904 940 38956
rect 992 38944 998 38956
rect 1765 38947 1823 38953
rect 1765 38944 1777 38947
rect 992 38916 1777 38944
rect 992 38904 998 38916
rect 1765 38913 1777 38916
rect 1811 38913 1823 38947
rect 1765 38907 1823 38913
rect 1946 38904 1952 38956
rect 2004 38944 2010 38956
rect 22373 38947 22431 38953
rect 22373 38944 22385 38947
rect 2004 38916 22385 38944
rect 2004 38904 2010 38916
rect 22373 38913 22385 38916
rect 22419 38944 22431 38947
rect 23201 38947 23259 38953
rect 23201 38944 23213 38947
rect 22419 38916 23213 38944
rect 22419 38913 22431 38916
rect 22373 38907 22431 38913
rect 23201 38913 23213 38916
rect 23247 38944 23259 38947
rect 26142 38944 26148 38956
rect 23247 38916 26148 38944
rect 23247 38913 23259 38916
rect 23201 38907 23259 38913
rect 26142 38904 26148 38916
rect 26200 38904 26206 38956
rect 26234 38904 26240 38956
rect 26292 38904 26298 38956
rect 26786 38904 26792 38956
rect 26844 38944 26850 38956
rect 27709 38947 27767 38953
rect 27709 38944 27721 38947
rect 26844 38916 27721 38944
rect 26844 38904 26850 38916
rect 27709 38913 27721 38916
rect 27755 38913 27767 38947
rect 27709 38907 27767 38913
rect 28442 38904 28448 38956
rect 28500 38944 28506 38956
rect 28500 38916 29132 38944
rect 28500 38904 28506 38916
rect 23477 38879 23535 38885
rect 23477 38845 23489 38879
rect 23523 38876 23535 38879
rect 24578 38876 24584 38888
rect 23523 38848 24584 38876
rect 23523 38845 23535 38848
rect 23477 38839 23535 38845
rect 24578 38836 24584 38848
rect 24636 38836 24642 38888
rect 24946 38836 24952 38888
rect 25004 38876 25010 38888
rect 25041 38879 25099 38885
rect 25041 38876 25053 38879
rect 25004 38848 25053 38876
rect 25004 38836 25010 38848
rect 25041 38845 25053 38848
rect 25087 38845 25099 38879
rect 25041 38839 25099 38845
rect 26510 38836 26516 38888
rect 26568 38836 26574 38888
rect 27890 38836 27896 38888
rect 27948 38836 27954 38888
rect 27982 38836 27988 38888
rect 28040 38876 28046 38888
rect 29104 38885 29132 38916
rect 32582 38904 32588 38956
rect 32640 38944 32646 38956
rect 35345 38947 35403 38953
rect 35345 38944 35357 38947
rect 32640 38916 35357 38944
rect 32640 38904 32646 38916
rect 35345 38913 35357 38916
rect 35391 38944 35403 38947
rect 36541 38947 36599 38953
rect 35391 38916 36308 38944
rect 35391 38913 35403 38916
rect 35345 38907 35403 38913
rect 28997 38879 29055 38885
rect 28997 38876 29009 38879
rect 28040 38848 29009 38876
rect 28040 38836 28046 38848
rect 28997 38845 29009 38848
rect 29043 38845 29055 38879
rect 28997 38839 29055 38845
rect 29089 38879 29147 38885
rect 29089 38845 29101 38879
rect 29135 38845 29147 38879
rect 29089 38839 29147 38845
rect 31021 38879 31079 38885
rect 31021 38845 31033 38879
rect 31067 38876 31079 38879
rect 32861 38879 32919 38885
rect 32861 38876 32873 38879
rect 31067 38848 32873 38876
rect 31067 38845 31079 38848
rect 31021 38839 31079 38845
rect 32861 38845 32873 38848
rect 32907 38845 32919 38879
rect 32861 38839 32919 38845
rect 32953 38879 33011 38885
rect 32953 38845 32965 38879
rect 32999 38845 33011 38879
rect 32953 38839 33011 38845
rect 34057 38879 34115 38885
rect 34057 38845 34069 38879
rect 34103 38845 34115 38879
rect 34057 38839 34115 38845
rect 34241 38879 34299 38885
rect 34241 38845 34253 38879
rect 34287 38876 34299 38879
rect 34330 38876 34336 38888
rect 34287 38848 34336 38876
rect 34287 38845 34299 38848
rect 34241 38839 34299 38845
rect 26050 38768 26056 38820
rect 26108 38808 26114 38820
rect 26786 38808 26792 38820
rect 26108 38780 26792 38808
rect 26108 38768 26114 38780
rect 26786 38768 26792 38780
rect 26844 38768 26850 38820
rect 28718 38768 28724 38820
rect 28776 38808 28782 38820
rect 31036 38808 31064 38839
rect 28776 38780 31064 38808
rect 28776 38768 28782 38780
rect 31570 38768 31576 38820
rect 31628 38808 31634 38820
rect 32968 38808 32996 38839
rect 31628 38780 32996 38808
rect 31628 38768 31634 38780
rect 1581 38743 1639 38749
rect 1581 38709 1593 38743
rect 1627 38740 1639 38743
rect 7374 38740 7380 38752
rect 1627 38712 7380 38740
rect 1627 38709 1639 38712
rect 1581 38703 1639 38709
rect 7374 38700 7380 38712
rect 7432 38700 7438 38752
rect 22833 38743 22891 38749
rect 22833 38709 22845 38743
rect 22879 38740 22891 38743
rect 26970 38740 26976 38752
rect 22879 38712 26976 38740
rect 22879 38709 22891 38712
rect 22833 38703 22891 38709
rect 26970 38700 26976 38712
rect 27028 38700 27034 38752
rect 28534 38700 28540 38752
rect 28592 38700 28598 38752
rect 31110 38700 31116 38752
rect 31168 38740 31174 38752
rect 34072 38740 34100 38839
rect 34330 38836 34336 38848
rect 34388 38836 34394 38888
rect 35250 38836 35256 38888
rect 35308 38876 35314 38888
rect 35529 38879 35587 38885
rect 35529 38876 35541 38879
rect 35308 38848 35541 38876
rect 35308 38836 35314 38848
rect 35529 38845 35541 38848
rect 35575 38845 35587 38879
rect 35529 38839 35587 38845
rect 31168 38712 34100 38740
rect 31168 38700 31174 38712
rect 34974 38700 34980 38752
rect 35032 38700 35038 38752
rect 36170 38700 36176 38752
rect 36228 38700 36234 38752
rect 36280 38740 36308 38916
rect 36541 38913 36553 38947
rect 36587 38944 36599 38947
rect 36906 38944 36912 38956
rect 36587 38916 36912 38944
rect 36587 38913 36599 38916
rect 36541 38907 36599 38913
rect 36906 38904 36912 38916
rect 36964 38904 36970 38956
rect 37826 38904 37832 38956
rect 37884 38904 37890 38956
rect 39666 38904 39672 38956
rect 39724 38904 39730 38956
rect 40328 38953 40356 38984
rect 40862 38972 40868 38984
rect 40920 38972 40926 39024
rect 41874 39012 41880 39024
rect 41814 38984 41880 39012
rect 41874 38972 41880 38984
rect 41932 39012 41938 39024
rect 42610 39012 42616 39024
rect 41932 38984 42616 39012
rect 41932 38972 41938 38984
rect 42610 38972 42616 38984
rect 42668 38972 42674 39024
rect 40313 38947 40371 38953
rect 40313 38913 40325 38947
rect 40359 38913 40371 38947
rect 40313 38907 40371 38913
rect 36446 38836 36452 38888
rect 36504 38876 36510 38888
rect 36725 38879 36783 38885
rect 36725 38876 36737 38879
rect 36504 38848 36737 38876
rect 36504 38836 36510 38848
rect 36725 38845 36737 38848
rect 36771 38845 36783 38879
rect 36725 38839 36783 38845
rect 37182 38836 37188 38888
rect 37240 38876 37246 38888
rect 37918 38876 37924 38888
rect 37240 38848 37924 38876
rect 37240 38836 37246 38848
rect 37918 38836 37924 38848
rect 37976 38876 37982 38888
rect 38013 38879 38071 38885
rect 38013 38876 38025 38879
rect 37976 38848 38025 38876
rect 37976 38836 37982 38848
rect 38013 38845 38025 38848
rect 38059 38845 38071 38879
rect 38013 38839 38071 38845
rect 38654 38836 38660 38888
rect 38712 38876 38718 38888
rect 38933 38879 38991 38885
rect 38933 38876 38945 38879
rect 38712 38848 38945 38876
rect 38712 38836 38718 38848
rect 38933 38845 38945 38848
rect 38979 38845 38991 38879
rect 38933 38839 38991 38845
rect 39117 38879 39175 38885
rect 39117 38845 39129 38879
rect 39163 38876 39175 38879
rect 39390 38876 39396 38888
rect 39163 38848 39396 38876
rect 39163 38845 39175 38848
rect 39117 38839 39175 38845
rect 39390 38836 39396 38848
rect 39448 38836 39454 38888
rect 39761 38879 39819 38885
rect 39761 38845 39773 38879
rect 39807 38845 39819 38879
rect 39761 38839 39819 38845
rect 39776 38808 39804 38839
rect 39850 38836 39856 38888
rect 39908 38836 39914 38888
rect 40586 38836 40592 38888
rect 40644 38836 40650 38888
rect 40034 38808 40040 38820
rect 37384 38780 40040 38808
rect 37384 38740 37412 38780
rect 40034 38768 40040 38780
rect 40092 38768 40098 38820
rect 36280 38712 37412 38740
rect 37458 38700 37464 38752
rect 37516 38700 37522 38752
rect 38473 38743 38531 38749
rect 38473 38709 38485 38743
rect 38519 38740 38531 38743
rect 41230 38740 41236 38752
rect 38519 38712 41236 38740
rect 38519 38709 38531 38712
rect 38473 38703 38531 38709
rect 41230 38700 41236 38712
rect 41288 38700 41294 38752
rect 41690 38700 41696 38752
rect 41748 38740 41754 38752
rect 42061 38743 42119 38749
rect 42061 38740 42073 38743
rect 41748 38712 42073 38740
rect 41748 38700 41754 38712
rect 42061 38709 42073 38712
rect 42107 38709 42119 38743
rect 42061 38703 42119 38709
rect 1104 38650 49864 38672
rect 1104 38598 2950 38650
rect 3002 38598 3014 38650
rect 3066 38598 3078 38650
rect 3130 38598 3142 38650
rect 3194 38598 3206 38650
rect 3258 38598 12950 38650
rect 13002 38598 13014 38650
rect 13066 38598 13078 38650
rect 13130 38598 13142 38650
rect 13194 38598 13206 38650
rect 13258 38598 22950 38650
rect 23002 38598 23014 38650
rect 23066 38598 23078 38650
rect 23130 38598 23142 38650
rect 23194 38598 23206 38650
rect 23258 38598 32950 38650
rect 33002 38598 33014 38650
rect 33066 38598 33078 38650
rect 33130 38598 33142 38650
rect 33194 38598 33206 38650
rect 33258 38598 42950 38650
rect 43002 38598 43014 38650
rect 43066 38598 43078 38650
rect 43130 38598 43142 38650
rect 43194 38598 43206 38650
rect 43258 38598 49864 38650
rect 1104 38576 49864 38598
rect 23290 38496 23296 38548
rect 23348 38496 23354 38548
rect 27062 38496 27068 38548
rect 27120 38496 27126 38548
rect 32861 38539 32919 38545
rect 32861 38505 32873 38539
rect 32907 38536 32919 38539
rect 36262 38536 36268 38548
rect 32907 38508 36268 38536
rect 32907 38505 32919 38508
rect 32861 38499 32919 38505
rect 36262 38496 36268 38508
rect 36320 38496 36326 38548
rect 36630 38496 36636 38548
rect 36688 38496 36694 38548
rect 40037 38539 40095 38545
rect 40037 38505 40049 38539
rect 40083 38536 40095 38539
rect 41138 38536 41144 38548
rect 40083 38508 41144 38536
rect 40083 38505 40095 38508
rect 40037 38499 40095 38505
rect 41138 38496 41144 38508
rect 41196 38496 41202 38548
rect 42794 38496 42800 38548
rect 42852 38536 42858 38548
rect 43257 38539 43315 38545
rect 43257 38536 43269 38539
rect 42852 38508 43269 38536
rect 42852 38496 42858 38508
rect 43257 38505 43269 38508
rect 43303 38536 43315 38539
rect 43346 38536 43352 38548
rect 43303 38508 43352 38536
rect 43303 38505 43315 38508
rect 43257 38499 43315 38505
rect 43346 38496 43352 38508
rect 43404 38496 43410 38548
rect 22833 38471 22891 38477
rect 22833 38437 22845 38471
rect 22879 38468 22891 38471
rect 25222 38468 25228 38480
rect 22879 38440 25228 38468
rect 22879 38437 22891 38440
rect 22833 38431 22891 38437
rect 25222 38428 25228 38440
rect 25280 38428 25286 38480
rect 26602 38428 26608 38480
rect 26660 38468 26666 38480
rect 28445 38471 28503 38477
rect 28445 38468 28457 38471
rect 26660 38440 28457 38468
rect 26660 38428 26666 38440
rect 28445 38437 28457 38440
rect 28491 38437 28503 38471
rect 28445 38431 28503 38437
rect 28810 38428 28816 38480
rect 28868 38468 28874 38480
rect 28868 38440 29040 38468
rect 28868 38428 28874 38440
rect 21082 38360 21088 38412
rect 21140 38360 21146 38412
rect 23842 38360 23848 38412
rect 23900 38360 23906 38412
rect 27062 38360 27068 38412
rect 27120 38400 27126 38412
rect 27617 38403 27675 38409
rect 27617 38400 27629 38403
rect 27120 38372 27629 38400
rect 27120 38360 27126 38372
rect 27617 38369 27629 38372
rect 27663 38369 27675 38403
rect 27617 38363 27675 38369
rect 28534 38360 28540 38412
rect 28592 38400 28598 38412
rect 29012 38409 29040 38440
rect 31846 38428 31852 38480
rect 31904 38468 31910 38480
rect 31904 38440 33456 38468
rect 31904 38428 31910 38440
rect 28905 38403 28963 38409
rect 28905 38400 28917 38403
rect 28592 38372 28917 38400
rect 28592 38360 28598 38372
rect 28905 38369 28917 38372
rect 28951 38369 28963 38403
rect 28905 38363 28963 38369
rect 28997 38403 29055 38409
rect 28997 38369 29009 38403
rect 29043 38369 29055 38403
rect 28997 38363 29055 38369
rect 29733 38403 29791 38409
rect 29733 38369 29745 38403
rect 29779 38400 29791 38403
rect 30098 38400 30104 38412
rect 29779 38372 30104 38400
rect 29779 38369 29791 38372
rect 29733 38363 29791 38369
rect 27154 38292 27160 38344
rect 27212 38332 27218 38344
rect 29748 38332 29776 38363
rect 30098 38360 30104 38372
rect 30156 38400 30162 38412
rect 30156 38372 32260 38400
rect 30156 38360 30162 38372
rect 27212 38304 29776 38332
rect 27212 38292 27218 38304
rect 31662 38292 31668 38344
rect 31720 38332 31726 38344
rect 31849 38335 31907 38341
rect 31849 38332 31861 38335
rect 31720 38304 31861 38332
rect 31720 38292 31726 38304
rect 31849 38301 31861 38304
rect 31895 38301 31907 38335
rect 31849 38295 31907 38301
rect 32232 38276 32260 38372
rect 33318 38360 33324 38412
rect 33376 38360 33382 38412
rect 33428 38409 33456 38440
rect 34514 38428 34520 38480
rect 34572 38468 34578 38480
rect 34572 38440 35020 38468
rect 34572 38428 34578 38440
rect 33413 38403 33471 38409
rect 33413 38369 33425 38403
rect 33459 38369 33471 38403
rect 33413 38363 33471 38369
rect 34698 38360 34704 38412
rect 34756 38400 34762 38412
rect 34885 38403 34943 38409
rect 34885 38400 34897 38403
rect 34756 38372 34897 38400
rect 34756 38360 34762 38372
rect 34885 38369 34897 38372
rect 34931 38369 34943 38403
rect 34992 38400 35020 38440
rect 36188 38440 41414 38468
rect 35250 38400 35256 38412
rect 34992 38372 35256 38400
rect 34885 38363 34943 38369
rect 35250 38360 35256 38372
rect 35308 38400 35314 38412
rect 36188 38400 36216 38440
rect 35308 38372 36216 38400
rect 35308 38360 35314 38372
rect 37366 38360 37372 38412
rect 37424 38400 37430 38412
rect 39209 38403 39267 38409
rect 39209 38400 39221 38403
rect 37424 38372 39221 38400
rect 37424 38360 37430 38372
rect 39209 38369 39221 38372
rect 39255 38400 39267 38403
rect 40402 38400 40408 38412
rect 39255 38372 40408 38400
rect 39255 38369 39267 38372
rect 39209 38363 39267 38369
rect 40402 38360 40408 38372
rect 40460 38360 40466 38412
rect 40586 38360 40592 38412
rect 40644 38360 40650 38412
rect 41386 38400 41414 38440
rect 43162 38400 43168 38412
rect 41386 38372 43168 38400
rect 43162 38360 43168 38372
rect 43220 38360 43226 38412
rect 36906 38292 36912 38344
rect 36964 38332 36970 38344
rect 37550 38332 37556 38344
rect 36964 38304 37556 38332
rect 36964 38292 36970 38304
rect 37550 38292 37556 38304
rect 37608 38332 37614 38344
rect 40497 38335 40555 38341
rect 40497 38332 40509 38335
rect 37608 38304 40509 38332
rect 37608 38292 37614 38304
rect 40497 38301 40509 38304
rect 40543 38332 40555 38335
rect 41046 38332 41052 38344
rect 40543 38304 41052 38332
rect 40543 38301 40555 38304
rect 40497 38295 40555 38301
rect 41046 38292 41052 38304
rect 41104 38332 41110 38344
rect 41233 38335 41291 38341
rect 41233 38332 41245 38335
rect 41104 38304 41245 38332
rect 41104 38292 41110 38304
rect 41233 38301 41245 38304
rect 41279 38301 41291 38335
rect 41233 38295 41291 38301
rect 41506 38292 41512 38344
rect 41564 38292 41570 38344
rect 42794 38292 42800 38344
rect 42852 38332 42858 38344
rect 43990 38332 43996 38344
rect 42852 38304 43996 38332
rect 42852 38292 42858 38304
rect 43990 38292 43996 38304
rect 44048 38292 44054 38344
rect 49326 38292 49332 38344
rect 49384 38292 49390 38344
rect 21358 38224 21364 38276
rect 21416 38224 21422 38276
rect 24670 38264 24676 38276
rect 22586 38236 24676 38264
rect 24670 38224 24676 38236
rect 24728 38224 24734 38276
rect 26605 38267 26663 38273
rect 26605 38233 26617 38267
rect 26651 38264 26663 38267
rect 27433 38267 27491 38273
rect 27433 38264 27445 38267
rect 26651 38236 27445 38264
rect 26651 38233 26663 38236
rect 26605 38227 26663 38233
rect 27433 38233 27445 38236
rect 27479 38264 27491 38267
rect 27479 38236 28948 38264
rect 27479 38233 27491 38236
rect 27433 38227 27491 38233
rect 23658 38156 23664 38208
rect 23716 38156 23722 38208
rect 23753 38199 23811 38205
rect 23753 38165 23765 38199
rect 23799 38196 23811 38199
rect 25498 38196 25504 38208
rect 23799 38168 25504 38196
rect 23799 38165 23811 38168
rect 23753 38159 23811 38165
rect 25498 38156 25504 38168
rect 25556 38156 25562 38208
rect 26970 38156 26976 38208
rect 27028 38196 27034 38208
rect 27525 38199 27583 38205
rect 27525 38196 27537 38199
rect 27028 38168 27537 38196
rect 27028 38156 27034 38168
rect 27525 38165 27537 38168
rect 27571 38165 27583 38199
rect 27525 38159 27583 38165
rect 28810 38156 28816 38208
rect 28868 38156 28874 38208
rect 28920 38196 28948 38236
rect 29914 38224 29920 38276
rect 29972 38264 29978 38276
rect 30009 38267 30067 38273
rect 30009 38264 30021 38267
rect 29972 38236 30021 38264
rect 29972 38224 29978 38236
rect 30009 38233 30021 38236
rect 30055 38233 30067 38267
rect 30009 38227 30067 38233
rect 30466 38224 30472 38276
rect 30524 38224 30530 38276
rect 31570 38224 31576 38276
rect 31628 38264 31634 38276
rect 31757 38267 31815 38273
rect 31757 38264 31769 38267
rect 31628 38236 31769 38264
rect 31628 38224 31634 38236
rect 31757 38233 31769 38236
rect 31803 38233 31815 38267
rect 31757 38227 31815 38233
rect 32214 38224 32220 38276
rect 32272 38264 32278 38276
rect 32585 38267 32643 38273
rect 32585 38264 32597 38267
rect 32272 38236 32597 38264
rect 32272 38224 32278 38236
rect 32585 38233 32597 38236
rect 32631 38233 32643 38267
rect 35161 38267 35219 38273
rect 32585 38227 32643 38233
rect 32784 38236 35112 38264
rect 32784 38196 32812 38236
rect 28920 38168 32812 38196
rect 33226 38156 33232 38208
rect 33284 38156 33290 38208
rect 35084 38196 35112 38236
rect 35161 38233 35173 38267
rect 35207 38264 35219 38267
rect 35434 38264 35440 38276
rect 35207 38236 35440 38264
rect 35207 38233 35219 38236
rect 35161 38227 35219 38233
rect 35434 38224 35440 38236
rect 35492 38224 35498 38276
rect 36446 38264 36452 38276
rect 36386 38236 36452 38264
rect 36446 38224 36452 38236
rect 36504 38264 36510 38276
rect 36998 38264 37004 38276
rect 36504 38236 37004 38264
rect 36504 38224 36510 38236
rect 36998 38224 37004 38236
rect 37056 38224 37062 38276
rect 37090 38224 37096 38276
rect 37148 38224 37154 38276
rect 37921 38267 37979 38273
rect 37921 38233 37933 38267
rect 37967 38264 37979 38267
rect 38654 38264 38660 38276
rect 37967 38236 38660 38264
rect 37967 38233 37979 38236
rect 37921 38227 37979 38233
rect 38654 38224 38660 38236
rect 38712 38224 38718 38276
rect 38764 38236 41414 38264
rect 37274 38196 37280 38208
rect 35084 38168 37280 38196
rect 37274 38156 37280 38168
rect 37332 38156 37338 38208
rect 38562 38156 38568 38208
rect 38620 38196 38626 38208
rect 38764 38196 38792 38236
rect 38620 38168 38792 38196
rect 38620 38156 38626 38168
rect 40402 38156 40408 38208
rect 40460 38196 40466 38208
rect 40678 38196 40684 38208
rect 40460 38168 40684 38196
rect 40460 38156 40466 38168
rect 40678 38156 40684 38168
rect 40736 38156 40742 38208
rect 41386 38196 41414 38236
rect 41690 38224 41696 38276
rect 41748 38264 41754 38276
rect 41785 38267 41843 38273
rect 41785 38264 41797 38267
rect 41748 38236 41797 38264
rect 41748 38224 41754 38236
rect 41785 38233 41797 38236
rect 41831 38233 41843 38267
rect 41785 38227 41843 38233
rect 43254 38224 43260 38276
rect 43312 38264 43318 38276
rect 46198 38264 46204 38276
rect 43312 38236 46204 38264
rect 43312 38224 43318 38236
rect 46198 38224 46204 38236
rect 46256 38224 46262 38276
rect 43714 38196 43720 38208
rect 41386 38168 43720 38196
rect 43714 38156 43720 38168
rect 43772 38156 43778 38208
rect 49142 38156 49148 38208
rect 49200 38156 49206 38208
rect 1104 38106 49864 38128
rect 1104 38054 7950 38106
rect 8002 38054 8014 38106
rect 8066 38054 8078 38106
rect 8130 38054 8142 38106
rect 8194 38054 8206 38106
rect 8258 38054 17950 38106
rect 18002 38054 18014 38106
rect 18066 38054 18078 38106
rect 18130 38054 18142 38106
rect 18194 38054 18206 38106
rect 18258 38054 27950 38106
rect 28002 38054 28014 38106
rect 28066 38054 28078 38106
rect 28130 38054 28142 38106
rect 28194 38054 28206 38106
rect 28258 38054 37950 38106
rect 38002 38054 38014 38106
rect 38066 38054 38078 38106
rect 38130 38054 38142 38106
rect 38194 38054 38206 38106
rect 38258 38054 47950 38106
rect 48002 38054 48014 38106
rect 48066 38054 48078 38106
rect 48130 38054 48142 38106
rect 48194 38054 48206 38106
rect 48258 38054 49864 38106
rect 1104 38032 49864 38054
rect 27154 37992 27160 38004
rect 23124 37964 27160 37992
rect 23124 37865 23152 37964
rect 27154 37952 27160 37964
rect 27212 37952 27218 38004
rect 27522 37952 27528 38004
rect 27580 37992 27586 38004
rect 32858 37992 32864 38004
rect 27580 37964 32864 37992
rect 27580 37952 27586 37964
rect 32858 37952 32864 37964
rect 32916 37952 32922 38004
rect 33870 37952 33876 38004
rect 33928 37992 33934 38004
rect 33965 37995 34023 38001
rect 33965 37992 33977 37995
rect 33928 37964 33977 37992
rect 33928 37952 33934 37964
rect 33965 37961 33977 37964
rect 34011 37961 34023 37995
rect 33965 37955 34023 37961
rect 35342 37952 35348 38004
rect 35400 37992 35406 38004
rect 37182 37992 37188 38004
rect 35400 37964 37188 37992
rect 35400 37952 35406 37964
rect 37182 37952 37188 37964
rect 37240 37952 37246 38004
rect 37461 37995 37519 38001
rect 37461 37961 37473 37995
rect 37507 37992 37519 37995
rect 37826 37992 37832 38004
rect 37507 37964 37832 37992
rect 37507 37961 37519 37964
rect 37461 37955 37519 37961
rect 37826 37952 37832 37964
rect 37884 37952 37890 38004
rect 39574 37952 39580 38004
rect 39632 37992 39638 38004
rect 39632 37964 40264 37992
rect 39632 37952 39638 37964
rect 24670 37924 24676 37936
rect 24610 37896 24676 37924
rect 24670 37884 24676 37896
rect 24728 37884 24734 37936
rect 28166 37884 28172 37936
rect 28224 37884 28230 37936
rect 31294 37884 31300 37936
rect 31352 37884 31358 37936
rect 31662 37884 31668 37936
rect 31720 37924 31726 37936
rect 35989 37927 36047 37933
rect 35989 37924 36001 37927
rect 31720 37896 36001 37924
rect 31720 37884 31754 37896
rect 35989 37893 36001 37896
rect 36035 37924 36047 37927
rect 37090 37924 37096 37936
rect 36035 37896 37096 37924
rect 36035 37893 36047 37896
rect 35989 37887 36047 37893
rect 37090 37884 37096 37896
rect 37148 37884 37154 37936
rect 40236 37924 40264 37964
rect 41230 37952 41236 38004
rect 41288 37952 41294 38004
rect 42794 37952 42800 38004
rect 42852 37992 42858 38004
rect 43073 37995 43131 38001
rect 43073 37992 43085 37995
rect 42852 37964 43085 37992
rect 42852 37952 42858 37964
rect 43073 37961 43085 37964
rect 43119 37992 43131 37995
rect 43438 37992 43444 38004
rect 43119 37964 43444 37992
rect 43119 37961 43131 37964
rect 43073 37955 43131 37961
rect 43438 37952 43444 37964
rect 43496 37952 43502 38004
rect 43714 37952 43720 38004
rect 43772 37992 43778 38004
rect 48590 37992 48596 38004
rect 43772 37964 48596 37992
rect 43772 37952 43778 37964
rect 48590 37952 48596 37964
rect 48648 37952 48654 38004
rect 41325 37927 41383 37933
rect 41325 37924 41337 37927
rect 40236 37896 41337 37924
rect 41325 37893 41337 37896
rect 41371 37893 41383 37927
rect 43254 37924 43260 37936
rect 41325 37887 41383 37893
rect 42168 37896 43260 37924
rect 23109 37859 23167 37865
rect 23109 37825 23121 37859
rect 23155 37825 23167 37859
rect 23109 37819 23167 37825
rect 27154 37816 27160 37868
rect 27212 37816 27218 37868
rect 30374 37816 30380 37868
rect 30432 37856 30438 37868
rect 30469 37859 30527 37865
rect 30469 37856 30481 37859
rect 30432 37828 30481 37856
rect 30432 37816 30438 37828
rect 30469 37825 30481 37828
rect 30515 37856 30527 37859
rect 31726 37856 31754 37884
rect 30515 37828 31754 37856
rect 32677 37859 32735 37865
rect 30515 37825 30527 37828
rect 30469 37819 30527 37825
rect 32677 37825 32689 37859
rect 32723 37856 32735 37859
rect 33502 37856 33508 37868
rect 32723 37828 33508 37856
rect 32723 37825 32735 37828
rect 32677 37819 32735 37825
rect 33502 37816 33508 37828
rect 33560 37816 33566 37868
rect 33873 37859 33931 37865
rect 33873 37825 33885 37859
rect 33919 37825 33931 37859
rect 33873 37819 33931 37825
rect 23385 37791 23443 37797
rect 23385 37757 23397 37791
rect 23431 37788 23443 37791
rect 26326 37788 26332 37800
rect 23431 37760 26332 37788
rect 23431 37757 23443 37760
rect 23385 37751 23443 37757
rect 26326 37748 26332 37760
rect 26384 37788 26390 37800
rect 27062 37788 27068 37800
rect 26384 37760 27068 37788
rect 26384 37748 26390 37760
rect 27062 37748 27068 37760
rect 27120 37748 27126 37800
rect 27433 37791 27491 37797
rect 27433 37757 27445 37791
rect 27479 37788 27491 37791
rect 27798 37788 27804 37800
rect 27479 37760 27804 37788
rect 27479 37757 27491 37760
rect 27433 37751 27491 37757
rect 27798 37748 27804 37760
rect 27856 37748 27862 37800
rect 29181 37791 29239 37797
rect 29181 37788 29193 37791
rect 28460 37760 29193 37788
rect 22462 37612 22468 37664
rect 22520 37652 22526 37664
rect 22649 37655 22707 37661
rect 22649 37652 22661 37655
rect 22520 37624 22661 37652
rect 22520 37612 22526 37624
rect 22649 37621 22661 37624
rect 22695 37621 22707 37655
rect 22649 37615 22707 37621
rect 24857 37655 24915 37661
rect 24857 37621 24869 37655
rect 24903 37652 24915 37655
rect 24946 37652 24952 37664
rect 24903 37624 24952 37652
rect 24903 37621 24915 37624
rect 24857 37615 24915 37621
rect 24946 37612 24952 37624
rect 25004 37612 25010 37664
rect 25038 37612 25044 37664
rect 25096 37652 25102 37664
rect 28460 37652 28488 37760
rect 29181 37757 29193 37760
rect 29227 37788 29239 37791
rect 29454 37788 29460 37800
rect 29227 37760 29460 37788
rect 29227 37757 29239 37760
rect 29181 37751 29239 37757
rect 29454 37748 29460 37760
rect 29512 37748 29518 37800
rect 32769 37791 32827 37797
rect 32769 37788 32781 37791
rect 29656 37760 32781 37788
rect 28902 37680 28908 37732
rect 28960 37720 28966 37732
rect 29656 37720 29684 37760
rect 32769 37757 32781 37760
rect 32815 37757 32827 37791
rect 32769 37751 32827 37757
rect 32950 37748 32956 37800
rect 33008 37748 33014 37800
rect 28960 37692 29684 37720
rect 28960 37680 28966 37692
rect 29730 37680 29736 37732
rect 29788 37720 29794 37732
rect 33888 37720 33916 37819
rect 34698 37816 34704 37868
rect 34756 37856 34762 37868
rect 36725 37859 36783 37865
rect 36725 37856 36737 37859
rect 34756 37828 36737 37856
rect 34756 37816 34762 37828
rect 36725 37825 36737 37828
rect 36771 37825 36783 37859
rect 36725 37819 36783 37825
rect 37826 37816 37832 37868
rect 37884 37816 37890 37868
rect 40402 37856 40408 37868
rect 40066 37828 40408 37856
rect 40402 37816 40408 37828
rect 40460 37816 40466 37868
rect 40678 37816 40684 37868
rect 40736 37856 40742 37868
rect 42168 37856 42196 37896
rect 43254 37884 43260 37896
rect 43312 37884 43318 37936
rect 40736 37828 42196 37856
rect 40736 37816 40742 37828
rect 42242 37816 42248 37868
rect 42300 37856 42306 37868
rect 42981 37859 43039 37865
rect 42981 37856 42993 37859
rect 42300 37828 42993 37856
rect 42300 37816 42306 37828
rect 42981 37825 42993 37828
rect 43027 37856 43039 37859
rect 43027 37828 45554 37856
rect 43027 37825 43039 37828
rect 42981 37819 43039 37825
rect 34054 37748 34060 37800
rect 34112 37748 34118 37800
rect 37918 37748 37924 37800
rect 37976 37748 37982 37800
rect 38105 37791 38163 37797
rect 38105 37757 38117 37791
rect 38151 37788 38163 37791
rect 38286 37788 38292 37800
rect 38151 37760 38292 37788
rect 38151 37757 38163 37760
rect 38105 37751 38163 37757
rect 38286 37748 38292 37760
rect 38344 37748 38350 37800
rect 38654 37748 38660 37800
rect 38712 37748 38718 37800
rect 38933 37791 38991 37797
rect 38933 37757 38945 37791
rect 38979 37788 38991 37791
rect 40126 37788 40132 37800
rect 38979 37760 40132 37788
rect 38979 37757 38991 37760
rect 38933 37751 38991 37757
rect 40126 37748 40132 37760
rect 40184 37748 40190 37800
rect 40310 37748 40316 37800
rect 40368 37788 40374 37800
rect 41417 37791 41475 37797
rect 41417 37788 41429 37791
rect 40368 37760 41429 37788
rect 40368 37748 40374 37760
rect 41417 37757 41429 37760
rect 41463 37757 41475 37791
rect 41417 37751 41475 37757
rect 43162 37748 43168 37800
rect 43220 37748 43226 37800
rect 29788 37692 33916 37720
rect 40144 37720 40172 37748
rect 40865 37723 40923 37729
rect 40144 37692 40816 37720
rect 29788 37680 29794 37692
rect 25096 37624 28488 37652
rect 30009 37655 30067 37661
rect 25096 37612 25102 37624
rect 30009 37621 30021 37655
rect 30055 37652 30067 37655
rect 31294 37652 31300 37664
rect 30055 37624 31300 37652
rect 30055 37621 30067 37624
rect 30009 37615 30067 37621
rect 31294 37612 31300 37624
rect 31352 37612 31358 37664
rect 31386 37612 31392 37664
rect 31444 37652 31450 37664
rect 32309 37655 32367 37661
rect 32309 37652 32321 37655
rect 31444 37624 32321 37652
rect 31444 37612 31450 37624
rect 32309 37621 32321 37624
rect 32355 37621 32367 37655
rect 32309 37615 32367 37621
rect 32490 37612 32496 37664
rect 32548 37652 32554 37664
rect 32674 37652 32680 37664
rect 32548 37624 32680 37652
rect 32548 37612 32554 37624
rect 32674 37612 32680 37624
rect 32732 37652 32738 37664
rect 32950 37652 32956 37664
rect 32732 37624 32956 37652
rect 32732 37612 32738 37624
rect 32950 37612 32956 37624
rect 33008 37612 33014 37664
rect 33505 37655 33563 37661
rect 33505 37621 33517 37655
rect 33551 37652 33563 37655
rect 34330 37652 34336 37664
rect 33551 37624 34336 37652
rect 33551 37621 33563 37624
rect 33505 37615 33563 37621
rect 34330 37612 34336 37624
rect 34388 37612 34394 37664
rect 40310 37612 40316 37664
rect 40368 37652 40374 37664
rect 40405 37655 40463 37661
rect 40405 37652 40417 37655
rect 40368 37624 40417 37652
rect 40368 37612 40374 37624
rect 40405 37621 40417 37624
rect 40451 37621 40463 37655
rect 40788 37652 40816 37692
rect 40865 37689 40877 37723
rect 40911 37720 40923 37723
rect 43806 37720 43812 37732
rect 40911 37692 43812 37720
rect 40911 37689 40923 37692
rect 40865 37683 40923 37689
rect 43806 37680 43812 37692
rect 43864 37680 43870 37732
rect 45526 37720 45554 37828
rect 49326 37816 49332 37868
rect 49384 37816 49390 37868
rect 49145 37723 49203 37729
rect 49145 37720 49157 37723
rect 45526 37692 49157 37720
rect 49145 37689 49157 37692
rect 49191 37689 49203 37723
rect 49145 37683 49203 37689
rect 40954 37652 40960 37664
rect 40788 37624 40960 37652
rect 40405 37615 40463 37621
rect 40954 37612 40960 37624
rect 41012 37612 41018 37664
rect 41414 37612 41420 37664
rect 41472 37652 41478 37664
rect 42613 37655 42671 37661
rect 42613 37652 42625 37655
rect 41472 37624 42625 37652
rect 41472 37612 41478 37624
rect 42613 37621 42625 37624
rect 42659 37621 42671 37655
rect 42613 37615 42671 37621
rect 1104 37562 49864 37584
rect 1104 37510 2950 37562
rect 3002 37510 3014 37562
rect 3066 37510 3078 37562
rect 3130 37510 3142 37562
rect 3194 37510 3206 37562
rect 3258 37510 12950 37562
rect 13002 37510 13014 37562
rect 13066 37510 13078 37562
rect 13130 37510 13142 37562
rect 13194 37510 13206 37562
rect 13258 37510 22950 37562
rect 23002 37510 23014 37562
rect 23066 37510 23078 37562
rect 23130 37510 23142 37562
rect 23194 37510 23206 37562
rect 23258 37510 32950 37562
rect 33002 37510 33014 37562
rect 33066 37510 33078 37562
rect 33130 37510 33142 37562
rect 33194 37510 33206 37562
rect 33258 37510 42950 37562
rect 43002 37510 43014 37562
rect 43066 37510 43078 37562
rect 43130 37510 43142 37562
rect 43194 37510 43206 37562
rect 43258 37510 49864 37562
rect 1104 37488 49864 37510
rect 22094 37408 22100 37460
rect 22152 37408 22158 37460
rect 25498 37408 25504 37460
rect 25556 37408 25562 37460
rect 27522 37448 27528 37460
rect 25608 37420 27528 37448
rect 25608 37380 25636 37420
rect 27522 37408 27528 37420
rect 27580 37408 27586 37460
rect 27798 37408 27804 37460
rect 27856 37448 27862 37460
rect 28537 37451 28595 37457
rect 28537 37448 28549 37451
rect 27856 37420 28549 37448
rect 27856 37408 27862 37420
rect 28537 37417 28549 37420
rect 28583 37417 28595 37451
rect 28537 37411 28595 37417
rect 28810 37408 28816 37460
rect 28868 37448 28874 37460
rect 34146 37448 34152 37460
rect 28868 37420 34152 37448
rect 28868 37408 28874 37420
rect 34146 37408 34152 37420
rect 34204 37408 34210 37460
rect 49142 37448 49148 37460
rect 36096 37420 49148 37448
rect 19306 37352 23796 37380
rect 14458 37136 14464 37188
rect 14516 37176 14522 37188
rect 19306 37176 19334 37352
rect 23768 37324 23796 37352
rect 23860 37352 25636 37380
rect 22741 37315 22799 37321
rect 22741 37281 22753 37315
rect 22787 37312 22799 37315
rect 23566 37312 23572 37324
rect 22787 37284 23572 37312
rect 22787 37281 22799 37284
rect 22741 37275 22799 37281
rect 23566 37272 23572 37284
rect 23624 37272 23630 37324
rect 23750 37272 23756 37324
rect 23808 37272 23814 37324
rect 23860 37321 23888 37352
rect 29730 37340 29736 37392
rect 29788 37340 29794 37392
rect 30190 37340 30196 37392
rect 30248 37380 30254 37392
rect 30248 37352 31754 37380
rect 30248 37340 30254 37352
rect 23845 37315 23903 37321
rect 23845 37281 23857 37315
rect 23891 37281 23903 37315
rect 23845 37275 23903 37281
rect 23934 37272 23940 37324
rect 23992 37312 23998 37324
rect 26053 37315 26111 37321
rect 26053 37312 26065 37315
rect 23992 37284 26065 37312
rect 23992 37272 23998 37284
rect 26053 37281 26065 37284
rect 26099 37281 26111 37315
rect 26053 37275 26111 37281
rect 26789 37315 26847 37321
rect 26789 37281 26801 37315
rect 26835 37312 26847 37315
rect 27154 37312 27160 37324
rect 26835 37284 27160 37312
rect 26835 37281 26847 37284
rect 26789 37275 26847 37281
rect 27154 37272 27160 37284
rect 27212 37272 27218 37324
rect 27614 37272 27620 37324
rect 27672 37312 27678 37324
rect 27672 37284 28212 37312
rect 27672 37272 27678 37284
rect 28184 37256 28212 37284
rect 29086 37272 29092 37324
rect 29144 37312 29150 37324
rect 30208 37312 30236 37340
rect 29144 37284 30236 37312
rect 30285 37315 30343 37321
rect 29144 37272 29150 37284
rect 30285 37281 30297 37315
rect 30331 37312 30343 37315
rect 31202 37312 31208 37324
rect 30331 37284 31208 37312
rect 30331 37281 30343 37284
rect 30285 37275 30343 37281
rect 31202 37272 31208 37284
rect 31260 37272 31266 37324
rect 31478 37272 31484 37324
rect 31536 37272 31542 37324
rect 31726 37312 31754 37352
rect 32677 37315 32735 37321
rect 32677 37312 32689 37315
rect 31726 37284 32689 37312
rect 32677 37281 32689 37284
rect 32723 37281 32735 37315
rect 32677 37275 32735 37281
rect 32858 37272 32864 37324
rect 32916 37312 32922 37324
rect 33965 37315 34023 37321
rect 33965 37312 33977 37315
rect 32916 37284 33977 37312
rect 32916 37272 32922 37284
rect 33965 37281 33977 37284
rect 34011 37281 34023 37315
rect 33965 37275 34023 37281
rect 22462 37204 22468 37256
rect 22520 37204 22526 37256
rect 22557 37247 22615 37253
rect 22557 37213 22569 37247
rect 22603 37244 22615 37247
rect 23661 37247 23719 37253
rect 22603 37216 23612 37244
rect 22603 37213 22615 37216
rect 22557 37207 22615 37213
rect 14516 37148 19334 37176
rect 14516 37136 14522 37148
rect 14918 37068 14924 37120
rect 14976 37108 14982 37120
rect 22572 37108 22600 37207
rect 14976 37080 22600 37108
rect 23293 37111 23351 37117
rect 14976 37068 14982 37080
rect 23293 37077 23305 37111
rect 23339 37108 23351 37111
rect 23382 37108 23388 37120
rect 23339 37080 23388 37108
rect 23339 37077 23351 37080
rect 23293 37071 23351 37077
rect 23382 37068 23388 37080
rect 23440 37068 23446 37120
rect 23584 37108 23612 37216
rect 23661 37213 23673 37247
rect 23707 37244 23719 37247
rect 24765 37247 24823 37253
rect 24765 37244 24777 37247
rect 23707 37216 24777 37244
rect 23707 37213 23719 37216
rect 23661 37207 23719 37213
rect 24765 37213 24777 37216
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 28166 37204 28172 37256
rect 28224 37204 28230 37256
rect 29181 37247 29239 37253
rect 29181 37213 29193 37247
rect 29227 37244 29239 37247
rect 30101 37247 30159 37253
rect 30101 37244 30113 37247
rect 29227 37216 30113 37244
rect 29227 37213 29239 37216
rect 29181 37207 29239 37213
rect 30101 37213 30113 37216
rect 30147 37213 30159 37247
rect 30101 37207 30159 37213
rect 31294 37204 31300 37256
rect 31352 37204 31358 37256
rect 32030 37204 32036 37256
rect 32088 37244 32094 37256
rect 32585 37247 32643 37253
rect 32585 37244 32597 37247
rect 32088 37216 32597 37244
rect 32088 37204 32094 37216
rect 32585 37213 32597 37216
rect 32631 37213 32643 37247
rect 32585 37207 32643 37213
rect 25608 37148 26096 37176
rect 25608 37120 25636 37148
rect 25590 37108 25596 37120
rect 23584 37080 25596 37108
rect 25590 37068 25596 37080
rect 25648 37068 25654 37120
rect 25866 37068 25872 37120
rect 25924 37068 25930 37120
rect 25958 37068 25964 37120
rect 26016 37068 26022 37120
rect 26068 37108 26096 37148
rect 27062 37136 27068 37188
rect 27120 37136 27126 37188
rect 29270 37136 29276 37188
rect 29328 37176 29334 37188
rect 31389 37179 31447 37185
rect 31389 37176 31401 37179
rect 29328 37148 31401 37176
rect 29328 37136 29334 37148
rect 31389 37145 31401 37148
rect 31435 37145 31447 37179
rect 31389 37139 31447 37145
rect 31938 37136 31944 37188
rect 31996 37176 32002 37188
rect 31996 37148 33456 37176
rect 31996 37136 32002 37148
rect 30193 37111 30251 37117
rect 30193 37108 30205 37111
rect 26068 37080 30205 37108
rect 30193 37077 30205 37080
rect 30239 37077 30251 37111
rect 30193 37071 30251 37077
rect 30834 37068 30840 37120
rect 30892 37108 30898 37120
rect 30929 37111 30987 37117
rect 30929 37108 30941 37111
rect 30892 37080 30941 37108
rect 30892 37068 30898 37080
rect 30929 37077 30941 37080
rect 30975 37077 30987 37111
rect 30929 37071 30987 37077
rect 31478 37068 31484 37120
rect 31536 37108 31542 37120
rect 32125 37111 32183 37117
rect 32125 37108 32137 37111
rect 31536 37080 32137 37108
rect 31536 37068 31542 37080
rect 32125 37077 32137 37080
rect 32171 37077 32183 37111
rect 32125 37071 32183 37077
rect 32490 37068 32496 37120
rect 32548 37068 32554 37120
rect 33428 37117 33456 37148
rect 33502 37136 33508 37188
rect 33560 37176 33566 37188
rect 33873 37179 33931 37185
rect 33873 37176 33885 37179
rect 33560 37148 33885 37176
rect 33560 37136 33566 37148
rect 33873 37145 33885 37148
rect 33919 37176 33931 37179
rect 36096 37176 36124 37420
rect 49142 37408 49148 37420
rect 49200 37408 49206 37460
rect 38654 37340 38660 37392
rect 38712 37380 38718 37392
rect 38712 37352 41552 37380
rect 38712 37340 38718 37352
rect 41524 37324 41552 37352
rect 39209 37315 39267 37321
rect 39209 37281 39221 37315
rect 39255 37312 39267 37315
rect 40126 37312 40132 37324
rect 39255 37284 40132 37312
rect 39255 37281 39267 37284
rect 39209 37275 39267 37281
rect 40126 37272 40132 37284
rect 40184 37272 40190 37324
rect 40310 37272 40316 37324
rect 40368 37312 40374 37324
rect 40589 37315 40647 37321
rect 40589 37312 40601 37315
rect 40368 37284 40601 37312
rect 40368 37272 40374 37284
rect 40589 37281 40601 37284
rect 40635 37281 40647 37315
rect 40589 37275 40647 37281
rect 40678 37272 40684 37324
rect 40736 37312 40742 37324
rect 41417 37315 41475 37321
rect 41417 37312 41429 37315
rect 40736 37284 41429 37312
rect 40736 37272 40742 37284
rect 41417 37281 41429 37284
rect 41463 37281 41475 37315
rect 41417 37275 41475 37281
rect 41506 37272 41512 37324
rect 41564 37312 41570 37324
rect 42153 37315 42211 37321
rect 42153 37312 42165 37315
rect 41564 37284 42165 37312
rect 41564 37272 41570 37284
rect 42153 37281 42165 37284
rect 42199 37312 42211 37315
rect 42518 37312 42524 37324
rect 42199 37284 42524 37312
rect 42199 37281 42211 37284
rect 42153 37275 42211 37281
rect 42518 37272 42524 37284
rect 42576 37272 42582 37324
rect 48041 37315 48099 37321
rect 48041 37281 48053 37315
rect 48087 37312 48099 37315
rect 48498 37312 48504 37324
rect 48087 37284 48504 37312
rect 48087 37281 48099 37284
rect 48041 37275 48099 37281
rect 48498 37272 48504 37284
rect 48556 37272 48562 37324
rect 36998 37204 37004 37256
rect 37056 37244 37062 37256
rect 37826 37244 37832 37256
rect 37056 37216 37832 37244
rect 37056 37204 37062 37216
rect 37826 37204 37832 37216
rect 37884 37244 37890 37256
rect 38470 37244 38476 37256
rect 37884 37216 38476 37244
rect 37884 37204 37890 37216
rect 38470 37204 38476 37216
rect 38528 37244 38534 37256
rect 38933 37247 38991 37253
rect 38933 37244 38945 37247
rect 38528 37216 38945 37244
rect 38528 37204 38534 37216
rect 38933 37213 38945 37216
rect 38979 37213 38991 37247
rect 38933 37207 38991 37213
rect 40218 37204 40224 37256
rect 40276 37244 40282 37256
rect 40497 37247 40555 37253
rect 40497 37244 40509 37247
rect 40276 37216 40509 37244
rect 40276 37204 40282 37216
rect 40497 37213 40509 37216
rect 40543 37213 40555 37247
rect 40497 37207 40555 37213
rect 48774 37204 48780 37256
rect 48832 37204 48838 37256
rect 40405 37179 40463 37185
rect 40405 37176 40417 37179
rect 33919 37148 36124 37176
rect 38580 37148 40417 37176
rect 33919 37145 33931 37148
rect 33873 37139 33931 37145
rect 33413 37111 33471 37117
rect 33413 37077 33425 37111
rect 33459 37077 33471 37111
rect 33413 37071 33471 37077
rect 33781 37111 33839 37117
rect 33781 37077 33793 37111
rect 33827 37108 33839 37111
rect 34514 37108 34520 37120
rect 33827 37080 34520 37108
rect 33827 37077 33839 37080
rect 33781 37071 33839 37077
rect 34514 37068 34520 37080
rect 34572 37108 34578 37120
rect 35434 37108 35440 37120
rect 34572 37080 35440 37108
rect 34572 37068 34578 37080
rect 35434 37068 35440 37080
rect 35492 37068 35498 37120
rect 35710 37068 35716 37120
rect 35768 37108 35774 37120
rect 36446 37108 36452 37120
rect 35768 37080 36452 37108
rect 35768 37068 35774 37080
rect 36446 37068 36452 37080
rect 36504 37068 36510 37120
rect 38580 37117 38608 37148
rect 40405 37145 40417 37148
rect 40451 37145 40463 37179
rect 40405 37139 40463 37145
rect 42429 37179 42487 37185
rect 42429 37145 42441 37179
rect 42475 37176 42487 37179
rect 43990 37176 43996 37188
rect 42475 37148 42840 37176
rect 43654 37148 43996 37176
rect 42475 37145 42487 37148
rect 42429 37139 42487 37145
rect 38565 37111 38623 37117
rect 38565 37077 38577 37111
rect 38611 37077 38623 37111
rect 38565 37071 38623 37077
rect 39025 37111 39083 37117
rect 39025 37077 39037 37111
rect 39071 37108 39083 37111
rect 39114 37108 39120 37120
rect 39071 37080 39120 37108
rect 39071 37077 39083 37080
rect 39025 37071 39083 37077
rect 39114 37068 39120 37080
rect 39172 37068 39178 37120
rect 39482 37068 39488 37120
rect 39540 37108 39546 37120
rect 40037 37111 40095 37117
rect 40037 37108 40049 37111
rect 39540 37080 40049 37108
rect 39540 37068 39546 37080
rect 40037 37077 40049 37080
rect 40083 37077 40095 37111
rect 42812 37108 42840 37148
rect 43990 37136 43996 37148
rect 44048 37136 44054 37188
rect 43438 37108 43444 37120
rect 42812 37080 43444 37108
rect 40037 37071 40095 37077
rect 43438 37068 43444 37080
rect 43496 37068 43502 37120
rect 43714 37068 43720 37120
rect 43772 37108 43778 37120
rect 43901 37111 43959 37117
rect 43901 37108 43913 37111
rect 43772 37080 43913 37108
rect 43772 37068 43778 37080
rect 43901 37077 43913 37080
rect 43947 37077 43959 37111
rect 43901 37071 43959 37077
rect 1104 37018 49864 37040
rect 1104 36966 7950 37018
rect 8002 36966 8014 37018
rect 8066 36966 8078 37018
rect 8130 36966 8142 37018
rect 8194 36966 8206 37018
rect 8258 36966 17950 37018
rect 18002 36966 18014 37018
rect 18066 36966 18078 37018
rect 18130 36966 18142 37018
rect 18194 36966 18206 37018
rect 18258 36966 27950 37018
rect 28002 36966 28014 37018
rect 28066 36966 28078 37018
rect 28130 36966 28142 37018
rect 28194 36966 28206 37018
rect 28258 36966 37950 37018
rect 38002 36966 38014 37018
rect 38066 36966 38078 37018
rect 38130 36966 38142 37018
rect 38194 36966 38206 37018
rect 38258 36966 47950 37018
rect 48002 36966 48014 37018
rect 48066 36966 48078 37018
rect 48130 36966 48142 37018
rect 48194 36966 48206 37018
rect 48258 36966 49864 37018
rect 1104 36944 49864 36966
rect 19426 36864 19432 36916
rect 19484 36864 19490 36916
rect 23750 36864 23756 36916
rect 23808 36904 23814 36916
rect 27617 36907 27675 36913
rect 27617 36904 27629 36907
rect 23808 36876 27629 36904
rect 23808 36864 23814 36876
rect 27617 36873 27629 36876
rect 27663 36873 27675 36907
rect 27617 36867 27675 36873
rect 29822 36864 29828 36916
rect 29880 36904 29886 36916
rect 32309 36907 32367 36913
rect 32309 36904 32321 36907
rect 29880 36876 32321 36904
rect 29880 36864 29886 36876
rect 32309 36873 32321 36876
rect 32355 36873 32367 36907
rect 32309 36867 32367 36873
rect 32398 36864 32404 36916
rect 32456 36904 32462 36916
rect 32769 36907 32827 36913
rect 32769 36904 32781 36907
rect 32456 36876 32781 36904
rect 32456 36864 32462 36876
rect 32769 36873 32781 36876
rect 32815 36873 32827 36907
rect 32769 36867 32827 36873
rect 34348 36876 37688 36904
rect 24670 36796 24676 36848
rect 24728 36796 24734 36848
rect 26329 36839 26387 36845
rect 26329 36805 26341 36839
rect 26375 36836 26387 36839
rect 30377 36839 30435 36845
rect 26375 36808 27936 36836
rect 26375 36805 26387 36808
rect 26329 36799 26387 36805
rect 934 36728 940 36780
rect 992 36768 998 36780
rect 1765 36771 1823 36777
rect 1765 36768 1777 36771
rect 992 36740 1777 36768
rect 992 36728 998 36740
rect 1765 36737 1777 36740
rect 1811 36737 1823 36771
rect 1765 36731 1823 36737
rect 17218 36728 17224 36780
rect 17276 36768 17282 36780
rect 19797 36771 19855 36777
rect 19797 36768 19809 36771
rect 17276 36740 19809 36768
rect 17276 36728 17282 36740
rect 19797 36737 19809 36740
rect 19843 36737 19855 36771
rect 19797 36731 19855 36737
rect 19889 36771 19947 36777
rect 19889 36737 19901 36771
rect 19935 36768 19947 36771
rect 21818 36768 21824 36780
rect 19935 36740 21824 36768
rect 19935 36737 19947 36740
rect 19889 36731 19947 36737
rect 21818 36728 21824 36740
rect 21876 36728 21882 36780
rect 26237 36771 26295 36777
rect 26237 36737 26249 36771
rect 26283 36768 26295 36771
rect 26283 36740 27292 36768
rect 26283 36737 26295 36740
rect 26237 36731 26295 36737
rect 20073 36703 20131 36709
rect 20073 36669 20085 36703
rect 20119 36700 20131 36703
rect 21358 36700 21364 36712
rect 20119 36672 21364 36700
rect 20119 36669 20131 36672
rect 20073 36663 20131 36669
rect 21358 36660 21364 36672
rect 21416 36660 21422 36712
rect 22554 36660 22560 36712
rect 22612 36700 22618 36712
rect 23385 36703 23443 36709
rect 23385 36700 23397 36703
rect 22612 36672 23397 36700
rect 22612 36660 22618 36672
rect 23385 36669 23397 36672
rect 23431 36669 23443 36703
rect 23385 36663 23443 36669
rect 23661 36703 23719 36709
rect 23661 36669 23673 36703
rect 23707 36700 23719 36703
rect 24946 36700 24952 36712
rect 23707 36672 24952 36700
rect 23707 36669 23719 36672
rect 23661 36663 23719 36669
rect 24946 36660 24952 36672
rect 25004 36660 25010 36712
rect 25409 36703 25467 36709
rect 25409 36669 25421 36703
rect 25455 36700 25467 36703
rect 25774 36700 25780 36712
rect 25455 36672 25780 36700
rect 25455 36669 25467 36672
rect 25409 36663 25467 36669
rect 25774 36660 25780 36672
rect 25832 36660 25838 36712
rect 26418 36660 26424 36712
rect 26476 36660 26482 36712
rect 27264 36700 27292 36740
rect 27338 36728 27344 36780
rect 27396 36768 27402 36780
rect 27525 36771 27583 36777
rect 27525 36768 27537 36771
rect 27396 36740 27537 36768
rect 27396 36728 27402 36740
rect 27525 36737 27537 36740
rect 27571 36737 27583 36771
rect 27798 36768 27804 36780
rect 27525 36731 27583 36737
rect 27724 36740 27804 36768
rect 27430 36700 27436 36712
rect 27264 36672 27436 36700
rect 27430 36660 27436 36672
rect 27488 36660 27494 36712
rect 27724 36709 27752 36740
rect 27798 36728 27804 36740
rect 27856 36728 27862 36780
rect 27709 36703 27767 36709
rect 27709 36669 27721 36703
rect 27755 36669 27767 36703
rect 27908 36700 27936 36808
rect 30377 36805 30389 36839
rect 30423 36836 30435 36839
rect 34238 36836 34244 36848
rect 30423 36808 34244 36836
rect 30423 36805 30435 36808
rect 30377 36799 30435 36805
rect 34238 36796 34244 36808
rect 34296 36796 34302 36848
rect 28994 36728 29000 36780
rect 29052 36768 29058 36780
rect 30285 36771 30343 36777
rect 30285 36768 30297 36771
rect 29052 36740 30297 36768
rect 29052 36728 29058 36740
rect 30285 36737 30297 36740
rect 30331 36737 30343 36771
rect 31386 36768 31392 36780
rect 30285 36731 30343 36737
rect 30392 36740 31392 36768
rect 30392 36700 30420 36740
rect 31386 36728 31392 36740
rect 31444 36728 31450 36780
rect 31754 36728 31760 36780
rect 31812 36728 31818 36780
rect 32677 36771 32735 36777
rect 32677 36737 32689 36771
rect 32723 36768 32735 36771
rect 34348 36768 34376 36876
rect 37660 36836 37688 36876
rect 37734 36864 37740 36916
rect 37792 36904 37798 36916
rect 37829 36907 37887 36913
rect 37829 36904 37841 36907
rect 37792 36876 37841 36904
rect 37792 36864 37798 36876
rect 37829 36873 37841 36876
rect 37875 36873 37887 36907
rect 37829 36867 37887 36873
rect 40586 36864 40592 36916
rect 40644 36904 40650 36916
rect 41417 36907 41475 36913
rect 41417 36904 41429 36907
rect 40644 36876 41429 36904
rect 40644 36864 40650 36876
rect 41417 36873 41429 36876
rect 41463 36873 41475 36907
rect 41417 36867 41475 36873
rect 42426 36864 42432 36916
rect 42484 36904 42490 36916
rect 43073 36907 43131 36913
rect 43073 36904 43085 36907
rect 42484 36876 43085 36904
rect 42484 36864 42490 36876
rect 43073 36873 43085 36876
rect 43119 36873 43131 36907
rect 43073 36867 43131 36873
rect 39022 36836 39028 36848
rect 37660 36808 39028 36836
rect 39022 36796 39028 36808
rect 39080 36796 39086 36848
rect 39574 36796 39580 36848
rect 39632 36836 39638 36848
rect 40402 36836 40408 36848
rect 39632 36808 40408 36836
rect 39632 36796 39638 36808
rect 40402 36796 40408 36808
rect 40460 36796 40466 36848
rect 42334 36796 42340 36848
rect 42392 36836 42398 36848
rect 48774 36836 48780 36848
rect 42392 36808 48780 36836
rect 42392 36796 42398 36808
rect 48774 36796 48780 36808
rect 48832 36796 48838 36848
rect 32723 36740 34376 36768
rect 32723 36737 32735 36740
rect 32677 36731 32735 36737
rect 35710 36728 35716 36780
rect 35768 36728 35774 36780
rect 41230 36728 41236 36780
rect 41288 36768 41294 36780
rect 42981 36771 43039 36777
rect 42981 36768 42993 36771
rect 41288 36740 42993 36768
rect 41288 36728 41294 36740
rect 42981 36737 42993 36740
rect 43027 36737 43039 36771
rect 43714 36768 43720 36780
rect 42981 36731 43039 36737
rect 43088 36740 43720 36768
rect 27908 36672 30420 36700
rect 30561 36703 30619 36709
rect 27709 36663 27767 36669
rect 30561 36669 30573 36703
rect 30607 36669 30619 36703
rect 30561 36663 30619 36669
rect 30576 36632 30604 36663
rect 30834 36660 30840 36712
rect 30892 36700 30898 36712
rect 32953 36703 33011 36709
rect 30892 36672 32352 36700
rect 30892 36660 30898 36672
rect 32122 36632 32128 36644
rect 30576 36604 32128 36632
rect 32122 36592 32128 36604
rect 32180 36592 32186 36644
rect 32324 36632 32352 36672
rect 32953 36669 32965 36703
rect 32999 36669 33011 36703
rect 32953 36663 33011 36669
rect 32968 36632 32996 36663
rect 33962 36660 33968 36712
rect 34020 36700 34026 36712
rect 34333 36703 34391 36709
rect 34333 36700 34345 36703
rect 34020 36672 34345 36700
rect 34020 36660 34026 36672
rect 34333 36669 34345 36672
rect 34379 36669 34391 36703
rect 34333 36663 34391 36669
rect 34609 36703 34667 36709
rect 34609 36669 34621 36703
rect 34655 36700 34667 36703
rect 35250 36700 35256 36712
rect 34655 36672 35256 36700
rect 34655 36669 34667 36672
rect 34609 36663 34667 36669
rect 35250 36660 35256 36672
rect 35308 36660 35314 36712
rect 37921 36703 37979 36709
rect 37921 36700 37933 36703
rect 35636 36672 37933 36700
rect 32324 36604 32996 36632
rect 1581 36567 1639 36573
rect 1581 36533 1593 36567
rect 1627 36564 1639 36567
rect 7558 36564 7564 36576
rect 1627 36536 7564 36564
rect 1627 36533 1639 36536
rect 1581 36527 1639 36533
rect 7558 36524 7564 36536
rect 7616 36524 7622 36576
rect 22830 36524 22836 36576
rect 22888 36564 22894 36576
rect 22925 36567 22983 36573
rect 22925 36564 22937 36567
rect 22888 36536 22937 36564
rect 22888 36524 22894 36536
rect 22925 36533 22937 36536
rect 22971 36533 22983 36567
rect 22925 36527 22983 36533
rect 25498 36524 25504 36576
rect 25556 36564 25562 36576
rect 25869 36567 25927 36573
rect 25869 36564 25881 36567
rect 25556 36536 25881 36564
rect 25556 36524 25562 36536
rect 25869 36533 25881 36536
rect 25915 36533 25927 36567
rect 25869 36527 25927 36533
rect 27157 36567 27215 36573
rect 27157 36533 27169 36567
rect 27203 36564 27215 36567
rect 29638 36564 29644 36576
rect 27203 36536 29644 36564
rect 27203 36533 27215 36536
rect 27157 36527 27215 36533
rect 29638 36524 29644 36536
rect 29696 36524 29702 36576
rect 29914 36524 29920 36576
rect 29972 36524 29978 36576
rect 34054 36524 34060 36576
rect 34112 36564 34118 36576
rect 35636 36564 35664 36672
rect 37921 36669 37933 36672
rect 37967 36669 37979 36703
rect 37921 36663 37979 36669
rect 38105 36703 38163 36709
rect 38105 36669 38117 36703
rect 38151 36700 38163 36703
rect 38470 36700 38476 36712
rect 38151 36672 38476 36700
rect 38151 36669 38163 36672
rect 38105 36663 38163 36669
rect 38470 36660 38476 36672
rect 38528 36660 38534 36712
rect 38654 36660 38660 36712
rect 38712 36700 38718 36712
rect 39669 36703 39727 36709
rect 39669 36700 39681 36703
rect 38712 36672 39681 36700
rect 38712 36660 38718 36672
rect 39669 36669 39681 36672
rect 39715 36669 39727 36703
rect 39669 36663 39727 36669
rect 39942 36660 39948 36712
rect 40000 36660 40006 36712
rect 40954 36660 40960 36712
rect 41012 36700 41018 36712
rect 43088 36700 43116 36740
rect 43714 36728 43720 36740
rect 43772 36728 43778 36780
rect 49326 36728 49332 36780
rect 49384 36728 49390 36780
rect 41012 36672 43116 36700
rect 43257 36703 43315 36709
rect 41012 36660 41018 36672
rect 43257 36669 43269 36703
rect 43303 36700 43315 36703
rect 43346 36700 43352 36712
rect 43303 36672 43352 36700
rect 43303 36669 43315 36672
rect 43257 36663 43315 36669
rect 43346 36660 43352 36672
rect 43404 36660 43410 36712
rect 35802 36592 35808 36644
rect 35860 36632 35866 36644
rect 37461 36635 37519 36641
rect 37461 36632 37473 36635
rect 35860 36604 37473 36632
rect 35860 36592 35866 36604
rect 37461 36601 37473 36604
rect 37507 36601 37519 36635
rect 37461 36595 37519 36601
rect 34112 36536 35664 36564
rect 34112 36524 34118 36536
rect 36078 36524 36084 36576
rect 36136 36524 36142 36576
rect 36538 36524 36544 36576
rect 36596 36564 36602 36576
rect 36906 36564 36912 36576
rect 36596 36536 36912 36564
rect 36596 36524 36602 36536
rect 36906 36524 36912 36536
rect 36964 36524 36970 36576
rect 40402 36524 40408 36576
rect 40460 36564 40466 36576
rect 40586 36564 40592 36576
rect 40460 36536 40592 36564
rect 40460 36524 40466 36536
rect 40586 36524 40592 36536
rect 40644 36524 40650 36576
rect 42613 36567 42671 36573
rect 42613 36533 42625 36567
rect 42659 36564 42671 36567
rect 44082 36564 44088 36576
rect 42659 36536 44088 36564
rect 42659 36533 42671 36536
rect 42613 36527 42671 36533
rect 44082 36524 44088 36536
rect 44140 36524 44146 36576
rect 49142 36524 49148 36576
rect 49200 36524 49206 36576
rect 1104 36474 49864 36496
rect 1104 36422 2950 36474
rect 3002 36422 3014 36474
rect 3066 36422 3078 36474
rect 3130 36422 3142 36474
rect 3194 36422 3206 36474
rect 3258 36422 12950 36474
rect 13002 36422 13014 36474
rect 13066 36422 13078 36474
rect 13130 36422 13142 36474
rect 13194 36422 13206 36474
rect 13258 36422 22950 36474
rect 23002 36422 23014 36474
rect 23066 36422 23078 36474
rect 23130 36422 23142 36474
rect 23194 36422 23206 36474
rect 23258 36422 32950 36474
rect 33002 36422 33014 36474
rect 33066 36422 33078 36474
rect 33130 36422 33142 36474
rect 33194 36422 33206 36474
rect 33258 36422 42950 36474
rect 43002 36422 43014 36474
rect 43066 36422 43078 36474
rect 43130 36422 43142 36474
rect 43194 36422 43206 36474
rect 43258 36422 49864 36474
rect 1104 36400 49864 36422
rect 21910 36320 21916 36372
rect 21968 36320 21974 36372
rect 22465 36363 22523 36369
rect 22465 36329 22477 36363
rect 22511 36360 22523 36363
rect 26234 36360 26240 36372
rect 22511 36332 26240 36360
rect 22511 36329 22523 36332
rect 22465 36323 22523 36329
rect 26234 36320 26240 36332
rect 26292 36320 26298 36372
rect 27338 36320 27344 36372
rect 27396 36320 27402 36372
rect 27430 36320 27436 36372
rect 27488 36360 27494 36372
rect 32033 36363 32091 36369
rect 32033 36360 32045 36363
rect 27488 36332 32045 36360
rect 27488 36320 27494 36332
rect 32033 36329 32045 36332
rect 32079 36329 32091 36363
rect 32033 36323 32091 36329
rect 32122 36320 32128 36372
rect 32180 36360 32186 36372
rect 33870 36360 33876 36372
rect 32180 36332 33876 36360
rect 32180 36320 32186 36332
rect 33870 36320 33876 36332
rect 33928 36320 33934 36372
rect 34422 36320 34428 36372
rect 34480 36360 34486 36372
rect 36354 36360 36360 36372
rect 34480 36332 36360 36360
rect 34480 36320 34486 36332
rect 36354 36320 36360 36332
rect 36412 36320 36418 36372
rect 37274 36320 37280 36372
rect 37332 36360 37338 36372
rect 37461 36363 37519 36369
rect 37461 36360 37473 36363
rect 37332 36332 37473 36360
rect 37332 36320 37338 36332
rect 37461 36329 37473 36332
rect 37507 36329 37519 36363
rect 37461 36323 37519 36329
rect 40129 36363 40187 36369
rect 40129 36329 40141 36363
rect 40175 36360 40187 36363
rect 41230 36360 41236 36372
rect 40175 36332 41236 36360
rect 40175 36329 40187 36332
rect 40129 36323 40187 36329
rect 41230 36320 41236 36332
rect 41288 36320 41294 36372
rect 21928 36224 21956 36320
rect 25866 36252 25872 36304
rect 25924 36292 25930 36304
rect 36265 36295 36323 36301
rect 25924 36264 28856 36292
rect 25924 36252 25930 36264
rect 22646 36224 22652 36236
rect 21928 36196 22652 36224
rect 22646 36184 22652 36196
rect 22704 36184 22710 36236
rect 22738 36184 22744 36236
rect 22796 36224 22802 36236
rect 23017 36227 23075 36233
rect 23017 36224 23029 36227
rect 22796 36196 23029 36224
rect 22796 36184 22802 36196
rect 23017 36193 23029 36196
rect 23063 36193 23075 36227
rect 23017 36187 23075 36193
rect 28445 36227 28503 36233
rect 28445 36193 28457 36227
rect 28491 36224 28503 36227
rect 28626 36224 28632 36236
rect 28491 36196 28632 36224
rect 28491 36193 28503 36196
rect 28445 36187 28503 36193
rect 28626 36184 28632 36196
rect 28684 36184 28690 36236
rect 28828 36224 28856 36264
rect 36265 36261 36277 36295
rect 36311 36261 36323 36295
rect 36265 36255 36323 36261
rect 28828 36196 32536 36224
rect 22830 36116 22836 36168
rect 22888 36116 22894 36168
rect 28166 36116 28172 36168
rect 28224 36116 28230 36168
rect 28261 36159 28319 36165
rect 28261 36125 28273 36159
rect 28307 36156 28319 36159
rect 28718 36156 28724 36168
rect 28307 36128 28724 36156
rect 28307 36125 28319 36128
rect 28261 36119 28319 36125
rect 28718 36116 28724 36128
rect 28776 36116 28782 36168
rect 31754 36116 31760 36168
rect 31812 36156 31818 36168
rect 32401 36159 32459 36165
rect 32401 36156 32413 36159
rect 31812 36128 32413 36156
rect 31812 36116 31818 36128
rect 32401 36125 32413 36128
rect 32447 36125 32459 36159
rect 32508 36156 32536 36196
rect 32674 36184 32680 36236
rect 32732 36224 32738 36236
rect 34606 36224 34612 36236
rect 32732 36196 34612 36224
rect 32732 36184 32738 36196
rect 34606 36184 34612 36196
rect 34664 36184 34670 36236
rect 34974 36184 34980 36236
rect 35032 36224 35038 36236
rect 35529 36227 35587 36233
rect 35529 36224 35541 36227
rect 35032 36196 35541 36224
rect 35032 36184 35038 36196
rect 35529 36193 35541 36196
rect 35575 36193 35587 36227
rect 35529 36187 35587 36193
rect 35621 36227 35679 36233
rect 35621 36193 35633 36227
rect 35667 36193 35679 36227
rect 35621 36187 35679 36193
rect 35066 36156 35072 36168
rect 32508 36128 35072 36156
rect 32401 36119 32459 36125
rect 35066 36116 35072 36128
rect 35124 36116 35130 36168
rect 35158 36116 35164 36168
rect 35216 36156 35222 36168
rect 35636 36156 35664 36187
rect 35216 36128 35664 36156
rect 36280 36156 36308 36255
rect 40586 36252 40592 36304
rect 40644 36292 40650 36304
rect 49142 36292 49148 36304
rect 40644 36264 49148 36292
rect 40644 36252 40650 36264
rect 49142 36252 49148 36264
rect 49200 36252 49206 36304
rect 36446 36184 36452 36236
rect 36504 36224 36510 36236
rect 36725 36227 36783 36233
rect 36725 36224 36737 36227
rect 36504 36196 36737 36224
rect 36504 36184 36510 36196
rect 36725 36193 36737 36196
rect 36771 36193 36783 36227
rect 36725 36187 36783 36193
rect 36814 36184 36820 36236
rect 36872 36184 36878 36236
rect 38010 36184 38016 36236
rect 38068 36184 38074 36236
rect 38102 36184 38108 36236
rect 38160 36224 38166 36236
rect 40494 36224 40500 36236
rect 38160 36196 40500 36224
rect 38160 36184 38166 36196
rect 40494 36184 40500 36196
rect 40552 36184 40558 36236
rect 40773 36227 40831 36233
rect 40773 36193 40785 36227
rect 40819 36224 40831 36227
rect 41690 36224 41696 36236
rect 40819 36196 41696 36224
rect 40819 36193 40831 36196
rect 40773 36187 40831 36193
rect 41690 36184 41696 36196
rect 41748 36184 41754 36236
rect 41782 36184 41788 36236
rect 41840 36184 41846 36236
rect 41874 36184 41880 36236
rect 41932 36184 41938 36236
rect 43165 36227 43223 36233
rect 43165 36193 43177 36227
rect 43211 36224 43223 36227
rect 43346 36224 43352 36236
rect 43211 36196 43352 36224
rect 43211 36193 43223 36196
rect 43165 36187 43223 36193
rect 43346 36184 43352 36196
rect 43404 36184 43410 36236
rect 41598 36156 41604 36168
rect 36280 36128 41604 36156
rect 35216 36116 35222 36128
rect 41598 36116 41604 36128
rect 41656 36116 41662 36168
rect 42794 36156 42800 36168
rect 41708 36128 42800 36156
rect 21726 36048 21732 36100
rect 21784 36088 21790 36100
rect 29914 36088 29920 36100
rect 21784 36060 29920 36088
rect 21784 36048 21790 36060
rect 29914 36048 29920 36060
rect 29972 36048 29978 36100
rect 33134 36048 33140 36100
rect 33192 36088 33198 36100
rect 35437 36091 35495 36097
rect 35437 36088 35449 36091
rect 33192 36060 35449 36088
rect 33192 36048 33198 36060
rect 35437 36057 35449 36060
rect 35483 36057 35495 36091
rect 35437 36051 35495 36057
rect 35618 36048 35624 36100
rect 35676 36088 35682 36100
rect 35802 36088 35808 36100
rect 35676 36060 35808 36088
rect 35676 36048 35682 36060
rect 35802 36048 35808 36060
rect 35860 36048 35866 36100
rect 36354 36048 36360 36100
rect 36412 36088 36418 36100
rect 36633 36091 36691 36097
rect 36633 36088 36645 36091
rect 36412 36060 36645 36088
rect 36412 36048 36418 36060
rect 36633 36057 36645 36060
rect 36679 36057 36691 36091
rect 36633 36051 36691 36057
rect 37829 36091 37887 36097
rect 37829 36057 37841 36091
rect 37875 36088 37887 36091
rect 40218 36088 40224 36100
rect 37875 36060 40224 36088
rect 37875 36057 37887 36060
rect 37829 36051 37887 36057
rect 40218 36048 40224 36060
rect 40276 36048 40282 36100
rect 40497 36091 40555 36097
rect 40497 36057 40509 36091
rect 40543 36088 40555 36091
rect 40678 36088 40684 36100
rect 40543 36060 40684 36088
rect 40543 36057 40555 36060
rect 40497 36051 40555 36057
rect 40678 36048 40684 36060
rect 40736 36048 40742 36100
rect 41708 36097 41736 36128
rect 42794 36116 42800 36128
rect 42852 36116 42858 36168
rect 42981 36159 43039 36165
rect 42981 36125 42993 36159
rect 43027 36156 43039 36159
rect 43530 36156 43536 36168
rect 43027 36128 43536 36156
rect 43027 36125 43039 36128
rect 42981 36119 43039 36125
rect 43530 36116 43536 36128
rect 43588 36116 43594 36168
rect 41693 36091 41751 36097
rect 41693 36057 41705 36091
rect 41739 36057 41751 36091
rect 41693 36051 41751 36057
rect 22646 35980 22652 36032
rect 22704 36020 22710 36032
rect 22925 36023 22983 36029
rect 22925 36020 22937 36023
rect 22704 35992 22937 36020
rect 22704 35980 22710 35992
rect 22925 35989 22937 35992
rect 22971 35989 22983 36023
rect 22925 35983 22983 35989
rect 26234 35980 26240 36032
rect 26292 36020 26298 36032
rect 27801 36023 27859 36029
rect 27801 36020 27813 36023
rect 26292 35992 27813 36020
rect 26292 35980 26298 35992
rect 27801 35989 27813 35992
rect 27847 35989 27859 36023
rect 27801 35983 27859 35989
rect 32493 36023 32551 36029
rect 32493 35989 32505 36023
rect 32539 36020 32551 36023
rect 34514 36020 34520 36032
rect 32539 35992 34520 36020
rect 32539 35989 32551 35992
rect 32493 35983 32551 35989
rect 34514 35980 34520 35992
rect 34572 35980 34578 36032
rect 35069 36023 35127 36029
rect 35069 35989 35081 36023
rect 35115 36020 35127 36023
rect 36814 36020 36820 36032
rect 35115 35992 36820 36020
rect 35115 35989 35127 35992
rect 35069 35983 35127 35989
rect 36814 35980 36820 35992
rect 36872 35980 36878 36032
rect 37921 36023 37979 36029
rect 37921 35989 37933 36023
rect 37967 36020 37979 36023
rect 38102 36020 38108 36032
rect 37967 35992 38108 36020
rect 37967 35989 37979 35992
rect 37921 35983 37979 35989
rect 38102 35980 38108 35992
rect 38160 35980 38166 36032
rect 38746 35980 38752 36032
rect 38804 36020 38810 36032
rect 40589 36023 40647 36029
rect 40589 36020 40601 36023
rect 38804 35992 40601 36020
rect 38804 35980 38810 35992
rect 40589 35989 40601 35992
rect 40635 35989 40647 36023
rect 40589 35983 40647 35989
rect 41322 35980 41328 36032
rect 41380 35980 41386 36032
rect 42521 36023 42579 36029
rect 42521 35989 42533 36023
rect 42567 36020 42579 36023
rect 42794 36020 42800 36032
rect 42567 35992 42800 36020
rect 42567 35989 42579 35992
rect 42521 35983 42579 35989
rect 42794 35980 42800 35992
rect 42852 35980 42858 36032
rect 42886 35980 42892 36032
rect 42944 35980 42950 36032
rect 43254 35980 43260 36032
rect 43312 36020 43318 36032
rect 43898 36020 43904 36032
rect 43312 35992 43904 36020
rect 43312 35980 43318 35992
rect 43898 35980 43904 35992
rect 43956 35980 43962 36032
rect 1104 35930 49864 35952
rect 1104 35878 7950 35930
rect 8002 35878 8014 35930
rect 8066 35878 8078 35930
rect 8130 35878 8142 35930
rect 8194 35878 8206 35930
rect 8258 35878 17950 35930
rect 18002 35878 18014 35930
rect 18066 35878 18078 35930
rect 18130 35878 18142 35930
rect 18194 35878 18206 35930
rect 18258 35878 27950 35930
rect 28002 35878 28014 35930
rect 28066 35878 28078 35930
rect 28130 35878 28142 35930
rect 28194 35878 28206 35930
rect 28258 35878 37950 35930
rect 38002 35878 38014 35930
rect 38066 35878 38078 35930
rect 38130 35878 38142 35930
rect 38194 35878 38206 35930
rect 38258 35878 47950 35930
rect 48002 35878 48014 35930
rect 48066 35878 48078 35930
rect 48130 35878 48142 35930
rect 48194 35878 48206 35930
rect 48258 35878 49864 35930
rect 1104 35856 49864 35878
rect 21082 35816 21088 35828
rect 19536 35788 21088 35816
rect 19536 35689 19564 35788
rect 21082 35776 21088 35788
rect 21140 35776 21146 35828
rect 21269 35819 21327 35825
rect 21269 35785 21281 35819
rect 21315 35816 21327 35819
rect 21358 35816 21364 35828
rect 21315 35788 21364 35816
rect 21315 35785 21327 35788
rect 21269 35779 21327 35785
rect 21358 35776 21364 35788
rect 21416 35776 21422 35828
rect 23753 35819 23811 35825
rect 22066 35788 23428 35816
rect 22066 35748 22094 35788
rect 21022 35720 22094 35748
rect 19521 35683 19579 35689
rect 19521 35649 19533 35683
rect 19567 35649 19579 35683
rect 19521 35643 19579 35649
rect 23290 35640 23296 35692
rect 23348 35680 23354 35692
rect 23400 35680 23428 35788
rect 23753 35785 23765 35819
rect 23799 35816 23811 35819
rect 23842 35816 23848 35828
rect 23799 35788 23848 35816
rect 23799 35785 23811 35788
rect 23753 35779 23811 35785
rect 23842 35776 23848 35788
rect 23900 35776 23906 35828
rect 27154 35816 27160 35828
rect 24688 35788 27160 35816
rect 24688 35689 24716 35788
rect 27154 35776 27160 35788
rect 27212 35776 27218 35828
rect 30834 35816 30840 35828
rect 29104 35788 30840 35816
rect 24949 35751 25007 35757
rect 24949 35717 24961 35751
rect 24995 35748 25007 35751
rect 25038 35748 25044 35760
rect 24995 35720 25044 35748
rect 24995 35717 25007 35720
rect 24949 35711 25007 35717
rect 25038 35708 25044 35720
rect 25096 35708 25102 35760
rect 27062 35708 27068 35760
rect 27120 35748 27126 35760
rect 29104 35748 29132 35788
rect 30834 35776 30840 35788
rect 30892 35776 30898 35828
rect 32309 35819 32367 35825
rect 32309 35785 32321 35819
rect 32355 35816 32367 35819
rect 33134 35816 33140 35828
rect 32355 35788 33140 35816
rect 32355 35785 32367 35788
rect 32309 35779 32367 35785
rect 33134 35776 33140 35788
rect 33192 35776 33198 35828
rect 35066 35776 35072 35828
rect 35124 35816 35130 35828
rect 35621 35819 35679 35825
rect 35621 35816 35633 35819
rect 35124 35788 35633 35816
rect 35124 35776 35130 35788
rect 35621 35785 35633 35788
rect 35667 35785 35679 35819
rect 35621 35779 35679 35785
rect 36081 35819 36139 35825
rect 36081 35785 36093 35819
rect 36127 35816 36139 35819
rect 39298 35816 39304 35828
rect 36127 35788 39304 35816
rect 36127 35785 36139 35788
rect 36081 35779 36139 35785
rect 39298 35776 39304 35788
rect 39356 35776 39362 35828
rect 39942 35776 39948 35828
rect 40000 35776 40006 35828
rect 49050 35816 49056 35828
rect 40052 35788 49056 35816
rect 27120 35720 29132 35748
rect 27120 35708 27126 35720
rect 33962 35708 33968 35760
rect 34020 35748 34026 35760
rect 38562 35748 38568 35760
rect 34020 35720 38568 35748
rect 34020 35708 34026 35720
rect 24673 35683 24731 35689
rect 23348 35652 24440 35680
rect 23348 35640 23354 35652
rect 17862 35572 17868 35624
rect 17920 35612 17926 35624
rect 19797 35615 19855 35621
rect 19797 35612 19809 35615
rect 17920 35584 19809 35612
rect 17920 35572 17926 35584
rect 19797 35581 19809 35584
rect 19843 35612 19855 35615
rect 19843 35584 21036 35612
rect 19843 35581 19855 35584
rect 19797 35575 19855 35581
rect 21008 35476 21036 35584
rect 21082 35572 21088 35624
rect 21140 35612 21146 35624
rect 22002 35612 22008 35624
rect 21140 35584 22008 35612
rect 21140 35572 21146 35584
rect 22002 35572 22008 35584
rect 22060 35572 22066 35624
rect 22281 35615 22339 35621
rect 22281 35581 22293 35615
rect 22327 35612 22339 35615
rect 23934 35612 23940 35624
rect 22327 35584 23940 35612
rect 22327 35581 22339 35584
rect 22281 35575 22339 35581
rect 23934 35572 23940 35584
rect 23992 35572 23998 35624
rect 24412 35612 24440 35652
rect 24673 35649 24685 35683
rect 24719 35649 24731 35683
rect 26082 35666 26556 35680
rect 24673 35643 24731 35649
rect 26068 35652 26556 35666
rect 26068 35612 26096 35652
rect 24412 35584 26096 35612
rect 24688 35556 24716 35584
rect 26326 35572 26332 35624
rect 26384 35612 26390 35624
rect 26421 35615 26479 35621
rect 26421 35612 26433 35615
rect 26384 35584 26433 35612
rect 26384 35572 26390 35584
rect 26421 35581 26433 35584
rect 26467 35581 26479 35615
rect 26528 35612 26556 35652
rect 27154 35640 27160 35692
rect 27212 35680 27218 35692
rect 29089 35683 29147 35689
rect 29089 35680 29101 35683
rect 27212 35652 29101 35680
rect 27212 35640 27218 35652
rect 29089 35649 29101 35652
rect 29135 35649 29147 35683
rect 29089 35643 29147 35649
rect 30466 35640 30472 35692
rect 30524 35640 30530 35692
rect 31757 35683 31815 35689
rect 31757 35649 31769 35683
rect 31803 35680 31815 35683
rect 32677 35683 32735 35689
rect 32677 35680 32689 35683
rect 31803 35652 32689 35680
rect 31803 35649 31815 35652
rect 31757 35643 31815 35649
rect 32677 35649 32689 35652
rect 32723 35649 32735 35683
rect 32677 35643 32735 35649
rect 34514 35640 34520 35692
rect 34572 35680 34578 35692
rect 38212 35689 38240 35720
rect 38562 35708 38568 35720
rect 38620 35708 38626 35760
rect 34793 35683 34851 35689
rect 34793 35680 34805 35683
rect 34572 35652 34805 35680
rect 34572 35640 34578 35652
rect 34793 35649 34805 35652
rect 34839 35649 34851 35683
rect 34793 35643 34851 35649
rect 34885 35683 34943 35689
rect 34885 35649 34897 35683
rect 34931 35680 34943 35683
rect 35989 35683 36047 35689
rect 34931 35652 35940 35680
rect 34931 35649 34943 35652
rect 34885 35643 34943 35649
rect 27614 35612 27620 35624
rect 26528 35584 27620 35612
rect 26421 35575 26479 35581
rect 27614 35572 27620 35584
rect 27672 35572 27678 35624
rect 29365 35615 29423 35621
rect 29365 35581 29377 35615
rect 29411 35612 29423 35615
rect 29454 35612 29460 35624
rect 29411 35584 29460 35612
rect 29411 35581 29423 35584
rect 29365 35575 29423 35581
rect 29454 35572 29460 35584
rect 29512 35612 29518 35624
rect 31570 35612 31576 35624
rect 29512 35584 31576 35612
rect 29512 35572 29518 35584
rect 31570 35572 31576 35584
rect 31628 35572 31634 35624
rect 32766 35572 32772 35624
rect 32824 35572 32830 35624
rect 32858 35572 32864 35624
rect 32916 35572 32922 35624
rect 35069 35615 35127 35621
rect 35069 35581 35081 35615
rect 35115 35612 35127 35615
rect 35802 35612 35808 35624
rect 35115 35584 35808 35612
rect 35115 35581 35127 35584
rect 35069 35575 35127 35581
rect 35802 35572 35808 35584
rect 35860 35572 35866 35624
rect 35912 35612 35940 35652
rect 35989 35649 36001 35683
rect 36035 35680 36047 35683
rect 38197 35683 38255 35689
rect 36035 35652 38148 35680
rect 36035 35649 36047 35652
rect 35989 35643 36047 35649
rect 35912 35584 36124 35612
rect 24670 35504 24676 35556
rect 24728 35504 24734 35556
rect 32784 35544 32812 35572
rect 33505 35547 33563 35553
rect 33505 35544 33517 35547
rect 32784 35516 33517 35544
rect 33505 35513 33517 35516
rect 33551 35513 33563 35547
rect 33505 35507 33563 35513
rect 34425 35547 34483 35553
rect 34425 35513 34437 35547
rect 34471 35544 34483 35547
rect 35894 35544 35900 35556
rect 34471 35516 35900 35544
rect 34471 35513 34483 35516
rect 34425 35507 34483 35513
rect 35894 35504 35900 35516
rect 35952 35504 35958 35556
rect 36096 35544 36124 35584
rect 36170 35572 36176 35624
rect 36228 35572 36234 35624
rect 38120 35612 38148 35652
rect 38197 35649 38209 35683
rect 38243 35649 38255 35683
rect 38197 35643 38255 35649
rect 39574 35640 39580 35692
rect 39632 35640 39638 35692
rect 39114 35612 39120 35624
rect 38120 35584 39120 35612
rect 39114 35572 39120 35584
rect 39172 35612 39178 35624
rect 40052 35612 40080 35788
rect 49050 35776 49056 35788
rect 49108 35776 49114 35828
rect 40770 35708 40776 35760
rect 40828 35708 40834 35760
rect 42889 35751 42947 35757
rect 42889 35748 42901 35751
rect 41386 35720 42901 35748
rect 40678 35640 40684 35692
rect 40736 35680 40742 35692
rect 40865 35683 40923 35689
rect 40865 35680 40877 35683
rect 40736 35652 40877 35680
rect 40736 35640 40742 35652
rect 40865 35649 40877 35652
rect 40911 35649 40923 35683
rect 40865 35643 40923 35649
rect 39172 35584 40080 35612
rect 39172 35572 39178 35584
rect 40954 35572 40960 35624
rect 41012 35612 41018 35624
rect 41386 35612 41414 35720
rect 42889 35717 42901 35720
rect 42935 35748 42947 35751
rect 43162 35748 43168 35760
rect 42935 35720 43168 35748
rect 42935 35717 42947 35720
rect 42889 35711 42947 35717
rect 43162 35708 43168 35720
rect 43220 35708 43226 35760
rect 42518 35640 42524 35692
rect 42576 35680 42582 35692
rect 42613 35683 42671 35689
rect 42613 35680 42625 35683
rect 42576 35652 42625 35680
rect 42576 35640 42582 35652
rect 42613 35649 42625 35652
rect 42659 35649 42671 35683
rect 42613 35643 42671 35649
rect 43990 35640 43996 35692
rect 44048 35640 44054 35692
rect 49326 35640 49332 35692
rect 49384 35640 49390 35692
rect 41012 35584 41414 35612
rect 41012 35572 41018 35584
rect 41966 35572 41972 35624
rect 42024 35612 42030 35624
rect 42024 35584 45554 35612
rect 42024 35572 42030 35584
rect 38194 35544 38200 35556
rect 36096 35516 38200 35544
rect 38194 35504 38200 35516
rect 38252 35504 38258 35556
rect 45526 35544 45554 35584
rect 49145 35547 49203 35553
rect 49145 35544 49157 35547
rect 45526 35516 49157 35544
rect 49145 35513 49157 35516
rect 49191 35513 49203 35547
rect 49145 35507 49203 35513
rect 23382 35476 23388 35488
rect 21008 35448 23388 35476
rect 23382 35436 23388 35448
rect 23440 35436 23446 35488
rect 26510 35436 26516 35488
rect 26568 35476 26574 35488
rect 27341 35479 27399 35485
rect 27341 35476 27353 35479
rect 26568 35448 27353 35476
rect 26568 35436 26574 35448
rect 27341 35445 27353 35448
rect 27387 35445 27399 35479
rect 27341 35439 27399 35445
rect 27706 35436 27712 35488
rect 27764 35476 27770 35488
rect 30098 35476 30104 35488
rect 27764 35448 30104 35476
rect 27764 35436 27770 35448
rect 30098 35436 30104 35448
rect 30156 35436 30162 35488
rect 30466 35436 30472 35488
rect 30524 35476 30530 35488
rect 33594 35476 33600 35488
rect 30524 35448 33600 35476
rect 30524 35436 30530 35448
rect 33594 35436 33600 35448
rect 33652 35436 33658 35488
rect 37274 35436 37280 35488
rect 37332 35476 37338 35488
rect 38454 35479 38512 35485
rect 38454 35476 38466 35479
rect 37332 35448 38466 35476
rect 37332 35436 37338 35448
rect 38454 35445 38466 35448
rect 38500 35476 38512 35479
rect 40310 35476 40316 35488
rect 38500 35448 40316 35476
rect 38500 35445 38512 35448
rect 38454 35439 38512 35445
rect 40310 35436 40316 35448
rect 40368 35436 40374 35488
rect 40405 35479 40463 35485
rect 40405 35445 40417 35479
rect 40451 35476 40463 35479
rect 42886 35476 42892 35488
rect 40451 35448 42892 35476
rect 40451 35445 40463 35448
rect 40405 35439 40463 35445
rect 42886 35436 42892 35448
rect 42944 35436 42950 35488
rect 43346 35436 43352 35488
rect 43404 35476 43410 35488
rect 44361 35479 44419 35485
rect 44361 35476 44373 35479
rect 43404 35448 44373 35476
rect 43404 35436 43410 35448
rect 44361 35445 44373 35448
rect 44407 35445 44419 35479
rect 44361 35439 44419 35445
rect 1104 35386 49864 35408
rect 1104 35334 2950 35386
rect 3002 35334 3014 35386
rect 3066 35334 3078 35386
rect 3130 35334 3142 35386
rect 3194 35334 3206 35386
rect 3258 35334 12950 35386
rect 13002 35334 13014 35386
rect 13066 35334 13078 35386
rect 13130 35334 13142 35386
rect 13194 35334 13206 35386
rect 13258 35334 22950 35386
rect 23002 35334 23014 35386
rect 23066 35334 23078 35386
rect 23130 35334 23142 35386
rect 23194 35334 23206 35386
rect 23258 35334 32950 35386
rect 33002 35334 33014 35386
rect 33066 35334 33078 35386
rect 33130 35334 33142 35386
rect 33194 35334 33206 35386
rect 33258 35334 42950 35386
rect 43002 35334 43014 35386
rect 43066 35334 43078 35386
rect 43130 35334 43142 35386
rect 43194 35334 43206 35386
rect 43258 35334 49864 35386
rect 1104 35312 49864 35334
rect 21818 35232 21824 35284
rect 21876 35272 21882 35284
rect 24581 35275 24639 35281
rect 24581 35272 24593 35275
rect 21876 35244 24593 35272
rect 21876 35232 21882 35244
rect 24581 35241 24593 35244
rect 24627 35241 24639 35275
rect 24581 35235 24639 35241
rect 26050 35232 26056 35284
rect 26108 35232 26114 35284
rect 26602 35232 26608 35284
rect 26660 35272 26666 35284
rect 27246 35272 27252 35284
rect 26660 35244 27252 35272
rect 26660 35232 26666 35244
rect 27246 35232 27252 35244
rect 27304 35272 27310 35284
rect 28997 35275 29055 35281
rect 28997 35272 29009 35275
rect 27304 35244 29009 35272
rect 27304 35232 27310 35244
rect 28997 35241 29009 35244
rect 29043 35241 29055 35275
rect 28997 35235 29055 35241
rect 30466 35232 30472 35284
rect 30524 35272 30530 35284
rect 30524 35244 33824 35272
rect 30524 35232 30530 35244
rect 23477 35207 23535 35213
rect 23477 35173 23489 35207
rect 23523 35204 23535 35207
rect 23934 35204 23940 35216
rect 23523 35176 23940 35204
rect 23523 35173 23535 35176
rect 23477 35167 23535 35173
rect 23934 35164 23940 35176
rect 23992 35204 23998 35216
rect 24210 35204 24216 35216
rect 23992 35176 24216 35204
rect 23992 35164 23998 35176
rect 24210 35164 24216 35176
rect 24268 35164 24274 35216
rect 29454 35164 29460 35216
rect 29512 35204 29518 35216
rect 33796 35204 33824 35244
rect 33870 35232 33876 35284
rect 33928 35272 33934 35284
rect 33965 35275 34023 35281
rect 33965 35272 33977 35275
rect 33928 35244 33977 35272
rect 33928 35232 33934 35244
rect 33965 35241 33977 35244
rect 34011 35241 34023 35275
rect 33965 35235 34023 35241
rect 38010 35232 38016 35284
rect 38068 35272 38074 35284
rect 38068 35244 38654 35272
rect 38068 35232 38074 35244
rect 38626 35204 38654 35244
rect 41414 35204 41420 35216
rect 29512 35176 32352 35204
rect 33796 35176 37596 35204
rect 38626 35176 41420 35204
rect 29512 35164 29518 35176
rect 21729 35139 21787 35145
rect 21729 35105 21741 35139
rect 21775 35136 21787 35139
rect 22002 35136 22008 35148
rect 21775 35108 22008 35136
rect 21775 35105 21787 35108
rect 21729 35099 21787 35105
rect 22002 35096 22008 35108
rect 22060 35136 22066 35148
rect 22554 35136 22560 35148
rect 22060 35108 22560 35136
rect 22060 35096 22066 35108
rect 22554 35096 22560 35108
rect 22612 35096 22618 35148
rect 23382 35096 23388 35148
rect 23440 35136 23446 35148
rect 25133 35139 25191 35145
rect 25133 35136 25145 35139
rect 23440 35108 25145 35136
rect 23440 35096 23446 35108
rect 25133 35105 25145 35108
rect 25179 35105 25191 35139
rect 25133 35099 25191 35105
rect 26697 35139 26755 35145
rect 26697 35105 26709 35139
rect 26743 35136 26755 35139
rect 27062 35136 27068 35148
rect 26743 35108 27068 35136
rect 26743 35105 26755 35108
rect 26697 35099 26755 35105
rect 27062 35096 27068 35108
rect 27120 35096 27126 35148
rect 27154 35096 27160 35148
rect 27212 35136 27218 35148
rect 27249 35139 27307 35145
rect 27249 35136 27261 35139
rect 27212 35108 27261 35136
rect 27212 35096 27218 35108
rect 27249 35105 27261 35108
rect 27295 35105 27307 35139
rect 27249 35099 27307 35105
rect 27525 35139 27583 35145
rect 27525 35105 27537 35139
rect 27571 35136 27583 35139
rect 29914 35136 29920 35148
rect 27571 35108 29920 35136
rect 27571 35105 27583 35108
rect 27525 35099 27583 35105
rect 29914 35096 29920 35108
rect 29972 35096 29978 35148
rect 30558 35096 30564 35148
rect 30616 35096 30622 35148
rect 31110 35096 31116 35148
rect 31168 35136 31174 35148
rect 31481 35139 31539 35145
rect 31481 35136 31493 35139
rect 31168 35108 31493 35136
rect 31168 35096 31174 35108
rect 31481 35105 31493 35108
rect 31527 35105 31539 35139
rect 31481 35099 31539 35105
rect 31662 35096 31668 35148
rect 31720 35096 31726 35148
rect 32214 35096 32220 35148
rect 32272 35096 32278 35148
rect 32324 35136 32352 35176
rect 32493 35139 32551 35145
rect 32493 35136 32505 35139
rect 32324 35108 32505 35136
rect 32493 35105 32505 35108
rect 32539 35136 32551 35139
rect 36078 35136 36084 35148
rect 32539 35108 36084 35136
rect 32539 35105 32551 35108
rect 32493 35099 32551 35105
rect 36078 35096 36084 35108
rect 36136 35096 36142 35148
rect 36630 35096 36636 35148
rect 36688 35096 36694 35148
rect 25041 35071 25099 35077
rect 25041 35037 25053 35071
rect 25087 35068 25099 35071
rect 26234 35068 26240 35080
rect 25087 35040 26240 35068
rect 25087 35037 25099 35040
rect 25041 35031 25099 35037
rect 26234 35028 26240 35040
rect 26292 35028 26298 35080
rect 26421 35071 26479 35077
rect 26421 35037 26433 35071
rect 26467 35068 26479 35071
rect 26510 35068 26516 35080
rect 26467 35040 26516 35068
rect 26467 35037 26479 35040
rect 26421 35031 26479 35037
rect 26510 35028 26516 35040
rect 26568 35028 26574 35080
rect 30576 35068 30604 35096
rect 28658 35040 30604 35068
rect 33594 35028 33600 35080
rect 33652 35068 33658 35080
rect 35710 35068 35716 35080
rect 33652 35040 35716 35068
rect 33652 35028 33658 35040
rect 35710 35028 35716 35040
rect 35768 35028 35774 35080
rect 36449 35071 36507 35077
rect 36449 35037 36461 35071
rect 36495 35068 36507 35071
rect 37458 35068 37464 35080
rect 36495 35040 37464 35068
rect 36495 35037 36507 35040
rect 36449 35031 36507 35037
rect 37458 35028 37464 35040
rect 37516 35028 37522 35080
rect 22005 35003 22063 35009
rect 22005 34969 22017 35003
rect 22051 35000 22063 35003
rect 22094 35000 22100 35012
rect 22051 34972 22100 35000
rect 22051 34969 22063 34972
rect 22005 34963 22063 34969
rect 22094 34960 22100 34972
rect 22152 34960 22158 35012
rect 23290 35000 23296 35012
rect 23230 34972 23296 35000
rect 23290 34960 23296 34972
rect 23348 34960 23354 35012
rect 24949 35003 25007 35009
rect 24949 34969 24961 35003
rect 24995 35000 25007 35003
rect 30561 35003 30619 35009
rect 24995 34972 27476 35000
rect 24995 34969 25007 34972
rect 24949 34963 25007 34969
rect 24578 34892 24584 34944
rect 24636 34932 24642 34944
rect 26513 34935 26571 34941
rect 26513 34932 26525 34935
rect 24636 34904 26525 34932
rect 24636 34892 24642 34904
rect 26513 34901 26525 34904
rect 26559 34901 26571 34935
rect 27448 34932 27476 34972
rect 30561 34969 30573 35003
rect 30607 35000 30619 35003
rect 31389 35003 31447 35009
rect 31389 35000 31401 35003
rect 30607 34972 31401 35000
rect 30607 34969 30619 34972
rect 30561 34963 30619 34969
rect 31389 34969 31401 34972
rect 31435 35000 31447 35003
rect 31435 34972 31754 35000
rect 31435 34969 31447 34972
rect 31389 34963 31447 34969
rect 28442 34932 28448 34944
rect 27448 34904 28448 34932
rect 26513 34895 26571 34901
rect 28442 34892 28448 34904
rect 28500 34892 28506 34944
rect 28534 34892 28540 34944
rect 28592 34932 28598 34944
rect 29822 34932 29828 34944
rect 28592 34904 29828 34932
rect 28592 34892 28598 34904
rect 29822 34892 29828 34904
rect 29880 34892 29886 34944
rect 30190 34892 30196 34944
rect 30248 34932 30254 34944
rect 31021 34935 31079 34941
rect 31021 34932 31033 34935
rect 30248 34904 31033 34932
rect 30248 34892 30254 34904
rect 31021 34901 31033 34904
rect 31067 34901 31079 34935
rect 31726 34932 31754 34972
rect 34238 34960 34244 35012
rect 34296 35000 34302 35012
rect 37568 35000 37596 35176
rect 41414 35164 41420 35176
rect 41472 35164 41478 35216
rect 42076 35176 42840 35204
rect 37826 35096 37832 35148
rect 37884 35096 37890 35148
rect 37918 35096 37924 35148
rect 37976 35096 37982 35148
rect 39206 35096 39212 35148
rect 39264 35096 39270 35148
rect 42076 35145 42104 35176
rect 42061 35139 42119 35145
rect 42061 35105 42073 35139
rect 42107 35105 42119 35139
rect 42061 35099 42119 35105
rect 42518 35096 42524 35148
rect 42576 35136 42582 35148
rect 42705 35139 42763 35145
rect 42705 35136 42717 35139
rect 42576 35108 42717 35136
rect 42576 35096 42582 35108
rect 42705 35105 42717 35108
rect 42751 35105 42763 35139
rect 42812 35136 42840 35176
rect 42981 35139 43039 35145
rect 42981 35136 42993 35139
rect 42812 35108 42993 35136
rect 42705 35099 42763 35105
rect 42981 35105 42993 35108
rect 43027 35136 43039 35139
rect 43346 35136 43352 35148
rect 43027 35108 43352 35136
rect 43027 35105 43039 35108
rect 42981 35099 43039 35105
rect 43346 35096 43352 35108
rect 43404 35096 43410 35148
rect 43530 35096 43536 35148
rect 43588 35136 43594 35148
rect 44453 35139 44511 35145
rect 44453 35136 44465 35139
rect 43588 35108 44465 35136
rect 43588 35096 43594 35108
rect 44453 35105 44465 35108
rect 44499 35105 44511 35139
rect 44453 35099 44511 35105
rect 37737 35071 37795 35077
rect 37737 35037 37749 35071
rect 37783 35068 37795 35071
rect 39574 35068 39580 35080
rect 37783 35040 39580 35068
rect 37783 35037 37795 35040
rect 37737 35031 37795 35037
rect 39574 35028 39580 35040
rect 39632 35028 39638 35080
rect 40218 35028 40224 35080
rect 40276 35068 40282 35080
rect 40678 35068 40684 35080
rect 40276 35040 40684 35068
rect 40276 35028 40282 35040
rect 40678 35028 40684 35040
rect 40736 35068 40742 35080
rect 40736 35040 42748 35068
rect 40736 35028 40742 35040
rect 38654 35000 38660 35012
rect 34296 34972 37412 35000
rect 37568 34972 38660 35000
rect 34296 34960 34302 34972
rect 35894 34932 35900 34944
rect 31726 34904 35900 34932
rect 31021 34895 31079 34901
rect 35894 34892 35900 34904
rect 35952 34892 35958 34944
rect 35986 34892 35992 34944
rect 36044 34892 36050 34944
rect 36354 34892 36360 34944
rect 36412 34892 36418 34944
rect 37384 34941 37412 34972
rect 38654 34960 38660 34972
rect 38712 34960 38718 35012
rect 38933 35003 38991 35009
rect 38933 34969 38945 35003
rect 38979 35000 38991 35003
rect 39206 35000 39212 35012
rect 38979 34972 39212 35000
rect 38979 34969 38991 34972
rect 38933 34963 38991 34969
rect 39206 34960 39212 34972
rect 39264 34960 39270 35012
rect 40126 34960 40132 35012
rect 40184 35000 40190 35012
rect 41877 35003 41935 35009
rect 41877 35000 41889 35003
rect 40184 34972 41889 35000
rect 40184 34960 40190 34972
rect 41877 34969 41889 34972
rect 41923 34969 41935 35003
rect 41877 34963 41935 34969
rect 37369 34935 37427 34941
rect 37369 34901 37381 34935
rect 37415 34901 37427 34935
rect 37369 34895 37427 34901
rect 37642 34892 37648 34944
rect 37700 34932 37706 34944
rect 38565 34935 38623 34941
rect 38565 34932 38577 34935
rect 37700 34904 38577 34932
rect 37700 34892 37706 34904
rect 38565 34901 38577 34904
rect 38611 34901 38623 34935
rect 38565 34895 38623 34901
rect 39025 34935 39083 34941
rect 39025 34901 39037 34935
rect 39071 34932 39083 34935
rect 40586 34932 40592 34944
rect 39071 34904 40592 34932
rect 39071 34901 39083 34904
rect 39025 34895 39083 34901
rect 40586 34892 40592 34904
rect 40644 34892 40650 34944
rect 41414 34892 41420 34944
rect 41472 34892 41478 34944
rect 41782 34892 41788 34944
rect 41840 34892 41846 34944
rect 42720 34932 42748 35040
rect 49326 35028 49332 35080
rect 49384 35028 49390 35080
rect 43990 34960 43996 35012
rect 44048 34960 44054 35012
rect 43622 34932 43628 34944
rect 42720 34904 43628 34932
rect 43622 34892 43628 34904
rect 43680 34892 43686 34944
rect 49142 34892 49148 34944
rect 49200 34892 49206 34944
rect 1104 34842 49864 34864
rect 1104 34790 7950 34842
rect 8002 34790 8014 34842
rect 8066 34790 8078 34842
rect 8130 34790 8142 34842
rect 8194 34790 8206 34842
rect 8258 34790 17950 34842
rect 18002 34790 18014 34842
rect 18066 34790 18078 34842
rect 18130 34790 18142 34842
rect 18194 34790 18206 34842
rect 18258 34790 27950 34842
rect 28002 34790 28014 34842
rect 28066 34790 28078 34842
rect 28130 34790 28142 34842
rect 28194 34790 28206 34842
rect 28258 34790 37950 34842
rect 38002 34790 38014 34842
rect 38066 34790 38078 34842
rect 38130 34790 38142 34842
rect 38194 34790 38206 34842
rect 38258 34790 47950 34842
rect 48002 34790 48014 34842
rect 48066 34790 48078 34842
rect 48130 34790 48142 34842
rect 48194 34790 48206 34842
rect 48258 34790 49864 34842
rect 1104 34768 49864 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34728 1639 34731
rect 7834 34728 7840 34740
rect 1627 34700 7840 34728
rect 1627 34697 1639 34700
rect 1581 34691 1639 34697
rect 7834 34688 7840 34700
rect 7892 34688 7898 34740
rect 19978 34688 19984 34740
rect 20036 34728 20042 34740
rect 22186 34728 22192 34740
rect 20036 34700 22192 34728
rect 20036 34688 20042 34700
rect 22186 34688 22192 34700
rect 22244 34728 22250 34740
rect 22244 34700 24808 34728
rect 22244 34688 22250 34700
rect 24670 34660 24676 34672
rect 24610 34632 24676 34660
rect 24670 34620 24676 34632
rect 24728 34620 24734 34672
rect 24780 34660 24808 34700
rect 24854 34688 24860 34740
rect 24912 34728 24918 34740
rect 25409 34731 25467 34737
rect 25409 34728 25421 34731
rect 24912 34700 25421 34728
rect 24912 34688 24918 34700
rect 25409 34697 25421 34700
rect 25455 34697 25467 34731
rect 25409 34691 25467 34697
rect 28718 34688 28724 34740
rect 28776 34728 28782 34740
rect 30101 34731 30159 34737
rect 30101 34728 30113 34731
rect 28776 34700 30113 34728
rect 28776 34688 28782 34700
rect 30101 34697 30113 34700
rect 30147 34697 30159 34731
rect 30101 34691 30159 34697
rect 30466 34688 30472 34740
rect 30524 34688 30530 34740
rect 30650 34688 30656 34740
rect 30708 34728 30714 34740
rect 31386 34728 31392 34740
rect 30708 34700 31392 34728
rect 30708 34688 30714 34700
rect 31386 34688 31392 34700
rect 31444 34688 31450 34740
rect 32309 34731 32367 34737
rect 32309 34697 32321 34731
rect 32355 34728 32367 34731
rect 34422 34728 34428 34740
rect 32355 34700 34428 34728
rect 32355 34697 32367 34700
rect 32309 34691 32367 34697
rect 34422 34688 34428 34700
rect 34480 34688 34486 34740
rect 34606 34688 34612 34740
rect 34664 34728 34670 34740
rect 35805 34731 35863 34737
rect 35805 34728 35817 34731
rect 34664 34700 35817 34728
rect 34664 34688 34670 34700
rect 35805 34697 35817 34700
rect 35851 34697 35863 34731
rect 35805 34691 35863 34697
rect 35894 34688 35900 34740
rect 35952 34728 35958 34740
rect 38930 34728 38936 34740
rect 35952 34700 38936 34728
rect 35952 34688 35958 34700
rect 38930 34688 38936 34700
rect 38988 34688 38994 34740
rect 39025 34731 39083 34737
rect 39025 34697 39037 34731
rect 39071 34697 39083 34731
rect 39025 34691 39083 34697
rect 28534 34660 28540 34672
rect 24780 34632 28540 34660
rect 28534 34620 28540 34632
rect 28592 34620 28598 34672
rect 30558 34660 30564 34672
rect 29762 34632 30564 34660
rect 30558 34620 30564 34632
rect 30616 34620 30622 34672
rect 31481 34663 31539 34669
rect 31481 34629 31493 34663
rect 31527 34660 31539 34663
rect 35710 34660 35716 34672
rect 31527 34632 33916 34660
rect 35558 34632 35716 34660
rect 31527 34629 31539 34632
rect 31481 34623 31539 34629
rect 1762 34552 1768 34604
rect 1820 34552 1826 34604
rect 24946 34552 24952 34604
rect 25004 34592 25010 34604
rect 25777 34595 25835 34601
rect 25777 34592 25789 34595
rect 25004 34564 25789 34592
rect 25004 34552 25010 34564
rect 25777 34561 25789 34564
rect 25823 34561 25835 34595
rect 25777 34555 25835 34561
rect 27154 34552 27160 34604
rect 27212 34592 27218 34604
rect 28261 34595 28319 34601
rect 28261 34592 28273 34595
rect 27212 34564 28273 34592
rect 27212 34552 27218 34564
rect 28261 34561 28273 34564
rect 28307 34561 28319 34595
rect 28261 34555 28319 34561
rect 29822 34552 29828 34604
rect 29880 34592 29886 34604
rect 29880 34564 31754 34592
rect 29880 34552 29886 34564
rect 22554 34484 22560 34536
rect 22612 34524 22618 34536
rect 23109 34527 23167 34533
rect 23109 34524 23121 34527
rect 22612 34496 23121 34524
rect 22612 34484 22618 34496
rect 23109 34493 23121 34496
rect 23155 34493 23167 34527
rect 23109 34487 23167 34493
rect 23385 34527 23443 34533
rect 23385 34493 23397 34527
rect 23431 34524 23443 34527
rect 23842 34524 23848 34536
rect 23431 34496 23848 34524
rect 23431 34493 23443 34496
rect 23385 34487 23443 34493
rect 23842 34484 23848 34496
rect 23900 34484 23906 34536
rect 24857 34527 24915 34533
rect 24857 34493 24869 34527
rect 24903 34524 24915 34527
rect 25130 34524 25136 34536
rect 24903 34496 25136 34524
rect 24903 34493 24915 34496
rect 24857 34487 24915 34493
rect 25130 34484 25136 34496
rect 25188 34484 25194 34536
rect 25866 34484 25872 34536
rect 25924 34484 25930 34536
rect 26053 34527 26111 34533
rect 26053 34493 26065 34527
rect 26099 34524 26111 34527
rect 26326 34524 26332 34536
rect 26099 34496 26332 34524
rect 26099 34493 26111 34496
rect 26053 34487 26111 34493
rect 26326 34484 26332 34496
rect 26384 34484 26390 34536
rect 28534 34484 28540 34536
rect 28592 34524 28598 34536
rect 29086 34524 29092 34536
rect 28592 34496 29092 34524
rect 28592 34484 28598 34496
rect 29086 34484 29092 34496
rect 29144 34484 29150 34536
rect 29914 34484 29920 34536
rect 29972 34524 29978 34536
rect 30009 34527 30067 34533
rect 30009 34524 30021 34527
rect 29972 34496 30021 34524
rect 29972 34484 29978 34496
rect 30009 34493 30021 34496
rect 30055 34524 30067 34527
rect 30282 34524 30288 34536
rect 30055 34496 30288 34524
rect 30055 34493 30067 34496
rect 30009 34487 30067 34493
rect 30282 34484 30288 34496
rect 30340 34484 30346 34536
rect 30561 34527 30619 34533
rect 30561 34524 30573 34527
rect 30392 34496 30573 34524
rect 28166 34456 28172 34468
rect 25056 34428 28172 34456
rect 20438 34348 20444 34400
rect 20496 34388 20502 34400
rect 25056 34388 25084 34428
rect 28166 34416 28172 34428
rect 28224 34416 28230 34468
rect 30098 34416 30104 34468
rect 30156 34456 30162 34468
rect 30392 34456 30420 34496
rect 30561 34493 30573 34496
rect 30607 34493 30619 34527
rect 30561 34487 30619 34493
rect 30653 34527 30711 34533
rect 30653 34493 30665 34527
rect 30699 34493 30711 34527
rect 30653 34487 30711 34493
rect 30668 34456 30696 34487
rect 30742 34484 30748 34536
rect 30800 34524 30806 34536
rect 31573 34527 31631 34533
rect 30800 34496 31064 34524
rect 30800 34484 30806 34496
rect 31036 34465 31064 34496
rect 31573 34493 31585 34527
rect 31619 34493 31631 34527
rect 31726 34524 31754 34564
rect 32674 34552 32680 34604
rect 32732 34552 32738 34604
rect 32769 34595 32827 34601
rect 32769 34561 32781 34595
rect 32815 34592 32827 34595
rect 33505 34595 33563 34601
rect 33505 34592 33517 34595
rect 32815 34564 33517 34592
rect 32815 34561 32827 34564
rect 32769 34555 32827 34561
rect 33505 34561 33517 34564
rect 33551 34561 33563 34595
rect 33505 34555 33563 34561
rect 32784 34524 32812 34555
rect 31726 34496 32812 34524
rect 32953 34527 33011 34533
rect 31573 34487 31631 34493
rect 32953 34493 32965 34527
rect 32999 34493 33011 34527
rect 32953 34487 33011 34493
rect 30156 34428 30420 34456
rect 30576 34428 30696 34456
rect 31021 34459 31079 34465
rect 30156 34416 30162 34428
rect 30576 34400 30604 34428
rect 31021 34425 31033 34459
rect 31067 34425 31079 34459
rect 31021 34419 31079 34425
rect 20496 34360 25084 34388
rect 20496 34348 20502 34360
rect 25130 34348 25136 34400
rect 25188 34388 25194 34400
rect 30558 34388 30564 34400
rect 25188 34360 30564 34388
rect 25188 34348 25194 34360
rect 30558 34348 30564 34360
rect 30616 34348 30622 34400
rect 30926 34348 30932 34400
rect 30984 34388 30990 34400
rect 31588 34388 31616 34487
rect 32968 34456 32996 34487
rect 33778 34456 33784 34468
rect 32968 34428 33784 34456
rect 33778 34416 33784 34428
rect 33836 34416 33842 34468
rect 33888 34456 33916 34632
rect 35710 34620 35716 34632
rect 35768 34620 35774 34672
rect 39040 34660 39068 34691
rect 39482 34688 39488 34740
rect 39540 34688 39546 34740
rect 39574 34688 39580 34740
rect 39632 34728 39638 34740
rect 39632 34700 41368 34728
rect 39632 34688 39638 34700
rect 39040 34632 41276 34660
rect 35802 34552 35808 34604
rect 35860 34592 35866 34604
rect 35860 34564 37412 34592
rect 35860 34552 35866 34564
rect 33962 34484 33968 34536
rect 34020 34524 34026 34536
rect 34057 34527 34115 34533
rect 34057 34524 34069 34527
rect 34020 34496 34069 34524
rect 34020 34484 34026 34496
rect 34057 34493 34069 34496
rect 34103 34493 34115 34527
rect 37182 34524 37188 34536
rect 34057 34487 34115 34493
rect 34164 34496 37188 34524
rect 34164 34456 34192 34496
rect 37182 34484 37188 34496
rect 37240 34484 37246 34536
rect 37384 34524 37412 34564
rect 37826 34552 37832 34604
rect 37884 34592 37890 34604
rect 39393 34595 39451 34601
rect 39393 34592 39405 34595
rect 37884 34564 39405 34592
rect 37884 34552 37890 34564
rect 39393 34561 39405 34564
rect 39439 34561 39451 34595
rect 39850 34592 39856 34604
rect 39393 34555 39451 34561
rect 39592 34564 39856 34592
rect 39592 34524 39620 34564
rect 39850 34552 39856 34564
rect 39908 34552 39914 34604
rect 40586 34552 40592 34604
rect 40644 34552 40650 34604
rect 40681 34595 40739 34601
rect 40681 34561 40693 34595
rect 40727 34592 40739 34595
rect 40862 34592 40868 34604
rect 40727 34564 40868 34592
rect 40727 34561 40739 34564
rect 40681 34555 40739 34561
rect 40862 34552 40868 34564
rect 40920 34552 40926 34604
rect 37384 34496 39620 34524
rect 39669 34527 39727 34533
rect 39669 34493 39681 34527
rect 39715 34524 39727 34527
rect 39942 34524 39948 34536
rect 39715 34496 39948 34524
rect 39715 34493 39727 34496
rect 39669 34487 39727 34493
rect 39942 34484 39948 34496
rect 40000 34484 40006 34536
rect 40773 34527 40831 34533
rect 40773 34493 40785 34527
rect 40819 34493 40831 34527
rect 40773 34487 40831 34493
rect 33888 34428 34192 34456
rect 36078 34416 36084 34468
rect 36136 34456 36142 34468
rect 40402 34456 40408 34468
rect 36136 34428 40408 34456
rect 36136 34416 36142 34428
rect 40402 34416 40408 34428
rect 40460 34416 40466 34468
rect 40788 34400 40816 34487
rect 30984 34360 31616 34388
rect 34320 34391 34378 34397
rect 30984 34348 30990 34360
rect 34320 34357 34332 34391
rect 34366 34388 34378 34391
rect 39942 34388 39948 34400
rect 34366 34360 39948 34388
rect 34366 34357 34378 34360
rect 34320 34351 34378 34357
rect 39942 34348 39948 34360
rect 40000 34348 40006 34400
rect 40218 34348 40224 34400
rect 40276 34348 40282 34400
rect 40770 34348 40776 34400
rect 40828 34348 40834 34400
rect 41248 34388 41276 34632
rect 41340 34524 41368 34700
rect 41414 34688 41420 34740
rect 41472 34728 41478 34740
rect 43349 34731 43407 34737
rect 43349 34728 43361 34731
rect 41472 34700 43361 34728
rect 41472 34688 41478 34700
rect 43349 34697 43361 34700
rect 43395 34697 43407 34731
rect 43349 34691 43407 34697
rect 41616 34632 42748 34660
rect 41616 34524 41644 34632
rect 41782 34552 41788 34604
rect 41840 34592 41846 34604
rect 41969 34595 42027 34601
rect 41969 34592 41981 34595
rect 41840 34564 41981 34592
rect 41840 34552 41846 34564
rect 41969 34561 41981 34564
rect 42015 34561 42027 34595
rect 42720 34592 42748 34632
rect 42794 34620 42800 34672
rect 42852 34660 42858 34672
rect 43441 34663 43499 34669
rect 43441 34660 43453 34663
rect 42852 34632 43453 34660
rect 42852 34620 42858 34632
rect 43441 34629 43453 34632
rect 43487 34629 43499 34663
rect 43441 34623 43499 34629
rect 43622 34620 43628 34672
rect 43680 34660 43686 34672
rect 49142 34660 49148 34672
rect 43680 34632 49148 34660
rect 43680 34620 43686 34632
rect 49142 34620 49148 34632
rect 49200 34620 49206 34672
rect 42720 34564 43484 34592
rect 41969 34555 42027 34561
rect 43456 34536 43484 34564
rect 49326 34552 49332 34604
rect 49384 34552 49390 34604
rect 43346 34524 43352 34536
rect 41340 34496 41644 34524
rect 41708 34496 43352 34524
rect 41708 34388 41736 34496
rect 43346 34484 43352 34496
rect 43404 34484 43410 34536
rect 43438 34484 43444 34536
rect 43496 34484 43502 34536
rect 43530 34484 43536 34536
rect 43588 34484 43594 34536
rect 44266 34524 44272 34536
rect 43640 34496 44272 34524
rect 42981 34459 43039 34465
rect 42981 34425 42993 34459
rect 43027 34456 43039 34459
rect 43640 34456 43668 34496
rect 44266 34484 44272 34496
rect 44324 34484 44330 34536
rect 49050 34484 49056 34536
rect 49108 34524 49114 34536
rect 49108 34496 49188 34524
rect 49108 34484 49114 34496
rect 49160 34465 49188 34496
rect 43027 34428 43668 34456
rect 49145 34459 49203 34465
rect 43027 34425 43039 34428
rect 42981 34419 43039 34425
rect 49145 34425 49157 34459
rect 49191 34425 49203 34459
rect 49145 34419 49203 34425
rect 41248 34360 41736 34388
rect 1104 34298 49864 34320
rect 1104 34246 2950 34298
rect 3002 34246 3014 34298
rect 3066 34246 3078 34298
rect 3130 34246 3142 34298
rect 3194 34246 3206 34298
rect 3258 34246 12950 34298
rect 13002 34246 13014 34298
rect 13066 34246 13078 34298
rect 13130 34246 13142 34298
rect 13194 34246 13206 34298
rect 13258 34246 22950 34298
rect 23002 34246 23014 34298
rect 23066 34246 23078 34298
rect 23130 34246 23142 34298
rect 23194 34246 23206 34298
rect 23258 34246 32950 34298
rect 33002 34246 33014 34298
rect 33066 34246 33078 34298
rect 33130 34246 33142 34298
rect 33194 34246 33206 34298
rect 33258 34246 42950 34298
rect 43002 34246 43014 34298
rect 43066 34246 43078 34298
rect 43130 34246 43142 34298
rect 43194 34246 43206 34298
rect 43258 34246 49864 34298
rect 1104 34224 49864 34246
rect 20806 34144 20812 34196
rect 20864 34184 20870 34196
rect 23293 34187 23351 34193
rect 23293 34184 23305 34187
rect 20864 34156 23305 34184
rect 20864 34144 20870 34156
rect 23293 34153 23305 34156
rect 23339 34153 23351 34187
rect 23293 34147 23351 34153
rect 28166 34144 28172 34196
rect 28224 34184 28230 34196
rect 30650 34184 30656 34196
rect 28224 34156 30656 34184
rect 28224 34144 28230 34156
rect 30650 34144 30656 34156
rect 30708 34144 30714 34196
rect 32493 34187 32551 34193
rect 32493 34153 32505 34187
rect 32539 34184 32551 34187
rect 32674 34184 32680 34196
rect 32539 34156 32680 34184
rect 32539 34153 32551 34156
rect 32493 34147 32551 34153
rect 32674 34144 32680 34156
rect 32732 34144 32738 34196
rect 34606 34144 34612 34196
rect 34664 34184 34670 34196
rect 35342 34184 35348 34196
rect 34664 34156 35348 34184
rect 34664 34144 34670 34156
rect 35342 34144 35348 34156
rect 35400 34144 35406 34196
rect 35434 34144 35440 34196
rect 35492 34184 35498 34196
rect 36817 34187 36875 34193
rect 35492 34156 36584 34184
rect 35492 34144 35498 34156
rect 22833 34119 22891 34125
rect 22833 34085 22845 34119
rect 22879 34116 22891 34119
rect 23382 34116 23388 34128
rect 22879 34088 23388 34116
rect 22879 34085 22891 34088
rect 22833 34079 22891 34085
rect 23382 34076 23388 34088
rect 23440 34076 23446 34128
rect 24581 34119 24639 34125
rect 24581 34116 24593 34119
rect 23492 34088 24593 34116
rect 21085 34051 21143 34057
rect 21085 34017 21097 34051
rect 21131 34048 21143 34051
rect 22002 34048 22008 34060
rect 21131 34020 22008 34048
rect 21131 34017 21143 34020
rect 21085 34011 21143 34017
rect 22002 34008 22008 34020
rect 22060 34008 22066 34060
rect 22370 34008 22376 34060
rect 22428 34048 22434 34060
rect 23492 34048 23520 34088
rect 24581 34085 24593 34088
rect 24627 34085 24639 34119
rect 24581 34079 24639 34085
rect 30745 34119 30803 34125
rect 30745 34085 30757 34119
rect 30791 34116 30803 34119
rect 36354 34116 36360 34128
rect 30791 34088 36360 34116
rect 30791 34085 30803 34088
rect 30745 34079 30803 34085
rect 36354 34076 36360 34088
rect 36412 34076 36418 34128
rect 22428 34020 23520 34048
rect 22428 34008 22434 34020
rect 23934 34008 23940 34060
rect 23992 34008 23998 34060
rect 25222 34008 25228 34060
rect 25280 34008 25286 34060
rect 26237 34051 26295 34057
rect 26237 34017 26249 34051
rect 26283 34048 26295 34051
rect 27154 34048 27160 34060
rect 26283 34020 27160 34048
rect 26283 34017 26295 34020
rect 26237 34011 26295 34017
rect 27154 34008 27160 34020
rect 27212 34008 27218 34060
rect 31389 34051 31447 34057
rect 31389 34017 31401 34051
rect 31435 34048 31447 34051
rect 34606 34048 34612 34060
rect 31435 34020 34612 34048
rect 31435 34017 31447 34020
rect 31389 34011 31447 34017
rect 34606 34008 34612 34020
rect 34664 34008 34670 34060
rect 36078 34008 36084 34060
rect 36136 34048 36142 34060
rect 36173 34051 36231 34057
rect 36173 34048 36185 34051
rect 36136 34020 36185 34048
rect 36136 34008 36142 34020
rect 36173 34017 36185 34020
rect 36219 34017 36231 34051
rect 36173 34011 36231 34017
rect 22830 33980 22836 33992
rect 22494 33952 22836 33980
rect 22830 33940 22836 33952
rect 22888 33980 22894 33992
rect 23290 33980 23296 33992
rect 22888 33952 23296 33980
rect 22888 33940 22894 33952
rect 23290 33940 23296 33952
rect 23348 33940 23354 33992
rect 23842 33980 23848 33992
rect 23400 33952 23848 33980
rect 21361 33915 21419 33921
rect 21361 33881 21373 33915
rect 21407 33881 21419 33915
rect 23400 33912 23428 33952
rect 23842 33940 23848 33952
rect 23900 33940 23906 33992
rect 27614 33940 27620 33992
rect 27672 33940 27678 33992
rect 29086 33940 29092 33992
rect 29144 33980 29150 33992
rect 29917 33983 29975 33989
rect 29917 33980 29929 33983
rect 29144 33952 29929 33980
rect 29144 33940 29150 33952
rect 29917 33949 29929 33952
rect 29963 33949 29975 33983
rect 29917 33943 29975 33949
rect 30558 33940 30564 33992
rect 30616 33980 30622 33992
rect 35802 33980 35808 33992
rect 30616 33952 35808 33980
rect 30616 33940 30622 33952
rect 35802 33940 35808 33952
rect 35860 33940 35866 33992
rect 36556 33980 36584 34156
rect 36817 34153 36829 34187
rect 36863 34184 36875 34187
rect 38608 34184 38614 34196
rect 36863 34156 38614 34184
rect 36863 34153 36875 34156
rect 36817 34147 36875 34153
rect 38608 34144 38614 34156
rect 38666 34144 38672 34196
rect 38930 34144 38936 34196
rect 38988 34184 38994 34196
rect 38988 34156 48314 34184
rect 38988 34144 38994 34156
rect 36630 34076 36636 34128
rect 36688 34116 36694 34128
rect 38289 34119 38347 34125
rect 38289 34116 38301 34119
rect 36688 34088 38301 34116
rect 36688 34076 36694 34088
rect 38289 34085 38301 34088
rect 38335 34085 38347 34119
rect 39574 34116 39580 34128
rect 38289 34079 38347 34085
rect 38948 34088 39580 34116
rect 37182 34008 37188 34060
rect 37240 34048 37246 34060
rect 37734 34048 37740 34060
rect 37240 34020 37740 34048
rect 37240 34008 37246 34020
rect 37734 34008 37740 34020
rect 37792 34008 37798 34060
rect 38470 34008 38476 34060
rect 38528 34048 38534 34060
rect 38654 34048 38660 34060
rect 38528 34020 38660 34048
rect 38528 34008 38534 34020
rect 38654 34008 38660 34020
rect 38712 34008 38718 34060
rect 38746 34008 38752 34060
rect 38804 34008 38810 34060
rect 38948 34057 38976 34088
rect 39574 34076 39580 34088
rect 39632 34076 39638 34128
rect 42150 34076 42156 34128
rect 42208 34116 42214 34128
rect 42208 34088 42380 34116
rect 42208 34076 42214 34088
rect 42352 34057 42380 34088
rect 38933 34051 38991 34057
rect 38933 34017 38945 34051
rect 38979 34017 38991 34051
rect 38933 34011 38991 34017
rect 42337 34051 42395 34057
rect 42337 34017 42349 34051
rect 42383 34017 42395 34051
rect 42337 34011 42395 34017
rect 38838 33980 38844 33992
rect 36556 33952 38844 33980
rect 38838 33940 38844 33952
rect 38896 33940 38902 33992
rect 41322 33940 41328 33992
rect 41380 33980 41386 33992
rect 42153 33983 42211 33989
rect 41380 33952 41920 33980
rect 41380 33940 41386 33952
rect 21361 33875 21419 33881
rect 22664 33884 23428 33912
rect 21376 33844 21404 33875
rect 22664 33844 22692 33884
rect 23474 33872 23480 33924
rect 23532 33912 23538 33924
rect 24949 33915 25007 33921
rect 24949 33912 24961 33915
rect 23532 33884 24961 33912
rect 23532 33872 23538 33884
rect 24949 33881 24961 33884
rect 24995 33881 25007 33915
rect 24949 33875 25007 33881
rect 26513 33915 26571 33921
rect 26513 33881 26525 33915
rect 26559 33912 26571 33915
rect 26602 33912 26608 33924
rect 26559 33884 26608 33912
rect 26559 33881 26571 33884
rect 26513 33875 26571 33881
rect 26602 33872 26608 33884
rect 26660 33872 26666 33924
rect 36446 33872 36452 33924
rect 36504 33872 36510 33924
rect 36538 33872 36544 33924
rect 36596 33912 36602 33924
rect 39390 33912 39396 33924
rect 36596 33884 39396 33912
rect 36596 33872 36602 33884
rect 39390 33872 39396 33884
rect 39448 33872 39454 33924
rect 21376 33816 22692 33844
rect 23382 33804 23388 33856
rect 23440 33844 23446 33856
rect 23661 33847 23719 33853
rect 23661 33844 23673 33847
rect 23440 33816 23673 33844
rect 23440 33804 23446 33816
rect 23661 33813 23673 33816
rect 23707 33813 23719 33847
rect 23661 33807 23719 33813
rect 23750 33804 23756 33856
rect 23808 33804 23814 33856
rect 25041 33847 25099 33853
rect 25041 33813 25053 33847
rect 25087 33844 25099 33847
rect 27798 33844 27804 33856
rect 25087 33816 27804 33844
rect 25087 33813 25099 33816
rect 25041 33807 25099 33813
rect 27798 33804 27804 33816
rect 27856 33804 27862 33856
rect 27982 33804 27988 33856
rect 28040 33804 28046 33856
rect 31110 33804 31116 33856
rect 31168 33804 31174 33856
rect 31202 33804 31208 33856
rect 31260 33804 31266 33856
rect 33778 33804 33784 33856
rect 33836 33844 33842 33856
rect 35529 33847 35587 33853
rect 35529 33844 35541 33847
rect 33836 33816 35541 33844
rect 33836 33804 33842 33816
rect 35529 33813 35541 33816
rect 35575 33844 35587 33847
rect 36357 33847 36415 33853
rect 36357 33844 36369 33847
rect 35575 33816 36369 33844
rect 35575 33813 35587 33816
rect 35529 33807 35587 33813
rect 36357 33813 36369 33816
rect 36403 33844 36415 33847
rect 37090 33844 37096 33856
rect 36403 33816 37096 33844
rect 36403 33813 36415 33816
rect 36357 33807 36415 33813
rect 37090 33804 37096 33816
rect 37148 33804 37154 33856
rect 37734 33804 37740 33856
rect 37792 33844 37798 33856
rect 38608 33844 38614 33856
rect 37792 33816 38614 33844
rect 37792 33804 37798 33816
rect 38608 33804 38614 33816
rect 38666 33853 38672 33856
rect 38666 33847 38715 33853
rect 38666 33813 38669 33847
rect 38703 33813 38715 33847
rect 38666 33807 38715 33813
rect 38666 33804 38672 33807
rect 39758 33804 39764 33856
rect 39816 33844 39822 33856
rect 41785 33847 41843 33853
rect 41785 33844 41797 33847
rect 39816 33816 41797 33844
rect 39816 33804 39822 33816
rect 41785 33813 41797 33816
rect 41831 33813 41843 33847
rect 41892 33844 41920 33952
rect 42153 33949 42165 33983
rect 42199 33980 42211 33983
rect 42242 33980 42248 33992
rect 42199 33952 42248 33980
rect 42199 33949 42211 33952
rect 42153 33943 42211 33949
rect 42242 33940 42248 33952
rect 42300 33940 42306 33992
rect 48286 33924 48314 34156
rect 49326 33940 49332 33992
rect 49384 33940 49390 33992
rect 48286 33884 48320 33924
rect 48314 33872 48320 33884
rect 48372 33872 48378 33924
rect 42245 33847 42303 33853
rect 42245 33844 42257 33847
rect 41892 33816 42257 33844
rect 41785 33807 41843 33813
rect 42245 33813 42257 33816
rect 42291 33813 42303 33847
rect 42245 33807 42303 33813
rect 48590 33804 48596 33856
rect 48648 33844 48654 33856
rect 49145 33847 49203 33853
rect 49145 33844 49157 33847
rect 48648 33816 49157 33844
rect 48648 33804 48654 33816
rect 49145 33813 49157 33816
rect 49191 33813 49203 33847
rect 49145 33807 49203 33813
rect 1104 33754 49864 33776
rect 1104 33702 7950 33754
rect 8002 33702 8014 33754
rect 8066 33702 8078 33754
rect 8130 33702 8142 33754
rect 8194 33702 8206 33754
rect 8258 33702 17950 33754
rect 18002 33702 18014 33754
rect 18066 33702 18078 33754
rect 18130 33702 18142 33754
rect 18194 33702 18206 33754
rect 18258 33702 27950 33754
rect 28002 33702 28014 33754
rect 28066 33702 28078 33754
rect 28130 33702 28142 33754
rect 28194 33702 28206 33754
rect 28258 33702 37950 33754
rect 38002 33702 38014 33754
rect 38066 33702 38078 33754
rect 38130 33702 38142 33754
rect 38194 33702 38206 33754
rect 38258 33702 47950 33754
rect 48002 33702 48014 33754
rect 48066 33702 48078 33754
rect 48130 33702 48142 33754
rect 48194 33702 48206 33754
rect 48258 33702 49864 33754
rect 1104 33680 49864 33702
rect 23658 33600 23664 33652
rect 23716 33600 23722 33652
rect 28721 33643 28779 33649
rect 28721 33609 28733 33643
rect 28767 33640 28779 33643
rect 28994 33640 29000 33652
rect 28767 33612 29000 33640
rect 28767 33609 28779 33612
rect 28721 33603 28779 33609
rect 28994 33600 29000 33612
rect 29052 33600 29058 33652
rect 29086 33600 29092 33652
rect 29144 33600 29150 33652
rect 36998 33640 37004 33652
rect 30300 33612 37004 33640
rect 21450 33464 21456 33516
rect 21508 33504 21514 33516
rect 24029 33507 24087 33513
rect 24029 33504 24041 33507
rect 21508 33476 24041 33504
rect 21508 33464 21514 33476
rect 24029 33473 24041 33476
rect 24075 33473 24087 33507
rect 24029 33467 24087 33473
rect 24121 33507 24179 33513
rect 24121 33473 24133 33507
rect 24167 33504 24179 33507
rect 25774 33504 25780 33516
rect 24167 33476 25780 33504
rect 24167 33473 24179 33476
rect 24121 33467 24179 33473
rect 25774 33464 25780 33476
rect 25832 33464 25838 33516
rect 26694 33464 26700 33516
rect 26752 33504 26758 33516
rect 26752 33476 29592 33504
rect 26752 33464 26758 33476
rect 24210 33396 24216 33448
rect 24268 33396 24274 33448
rect 27338 33396 27344 33448
rect 27396 33436 27402 33448
rect 27396 33408 28994 33436
rect 27396 33396 27402 33408
rect 27246 33328 27252 33380
rect 27304 33368 27310 33380
rect 28966 33368 28994 33408
rect 29086 33396 29092 33448
rect 29144 33436 29150 33448
rect 29181 33439 29239 33445
rect 29181 33436 29193 33439
rect 29144 33408 29193 33436
rect 29144 33396 29150 33408
rect 29181 33405 29193 33408
rect 29227 33405 29239 33439
rect 29181 33399 29239 33405
rect 29365 33439 29423 33445
rect 29365 33405 29377 33439
rect 29411 33436 29423 33439
rect 29454 33436 29460 33448
rect 29411 33408 29460 33436
rect 29411 33405 29423 33408
rect 29365 33399 29423 33405
rect 29454 33396 29460 33408
rect 29512 33396 29518 33448
rect 29564 33436 29592 33476
rect 29638 33464 29644 33516
rect 29696 33504 29702 33516
rect 30300 33513 30328 33612
rect 36998 33600 37004 33612
rect 37056 33600 37062 33652
rect 37461 33643 37519 33649
rect 37461 33609 37473 33643
rect 37507 33640 37519 33643
rect 40126 33640 40132 33652
rect 37507 33612 38700 33640
rect 37507 33609 37519 33612
rect 37461 33603 37519 33609
rect 33870 33532 33876 33584
rect 33928 33572 33934 33584
rect 34241 33575 34299 33581
rect 34241 33572 34253 33575
rect 33928 33544 34253 33572
rect 33928 33532 33934 33544
rect 34241 33541 34253 33544
rect 34287 33541 34299 33575
rect 35710 33572 35716 33584
rect 35466 33558 35716 33572
rect 34241 33535 34299 33541
rect 35452 33544 35716 33558
rect 30285 33507 30343 33513
rect 30285 33504 30297 33507
rect 29696 33476 30297 33504
rect 29696 33464 29702 33476
rect 30285 33473 30297 33476
rect 30331 33473 30343 33507
rect 30285 33467 30343 33473
rect 31110 33464 31116 33516
rect 31168 33504 31174 33516
rect 31297 33507 31355 33513
rect 31297 33504 31309 33507
rect 31168 33476 31309 33504
rect 31168 33464 31174 33476
rect 31297 33473 31309 33476
rect 31343 33473 31355 33507
rect 31297 33467 31355 33473
rect 33962 33464 33968 33516
rect 34020 33464 34026 33516
rect 30377 33439 30435 33445
rect 30377 33436 30389 33439
rect 29564 33408 30389 33436
rect 30377 33405 30389 33408
rect 30423 33405 30435 33439
rect 30377 33399 30435 33405
rect 30469 33439 30527 33445
rect 30469 33405 30481 33439
rect 30515 33405 30527 33439
rect 30469 33399 30527 33405
rect 30484 33368 30512 33399
rect 34698 33396 34704 33448
rect 34756 33436 34762 33448
rect 35452 33436 35480 33544
rect 35710 33532 35716 33544
rect 35768 33572 35774 33584
rect 36630 33572 36636 33584
rect 35768 33544 36636 33572
rect 35768 33532 35774 33544
rect 36630 33532 36636 33544
rect 36688 33532 36694 33584
rect 37366 33532 37372 33584
rect 37424 33572 37430 33584
rect 37921 33575 37979 33581
rect 37921 33572 37933 33575
rect 37424 33544 37933 33572
rect 37424 33532 37430 33544
rect 37921 33541 37933 33544
rect 37967 33572 37979 33575
rect 38286 33572 38292 33584
rect 37967 33544 38292 33572
rect 37967 33541 37979 33544
rect 37921 33535 37979 33541
rect 38286 33532 38292 33544
rect 38344 33532 38350 33584
rect 38672 33572 38700 33612
rect 38856 33612 40132 33640
rect 38856 33572 38884 33612
rect 40126 33600 40132 33612
rect 40184 33600 40190 33652
rect 41966 33640 41972 33652
rect 40328 33612 41972 33640
rect 38672 33544 38884 33572
rect 39209 33575 39267 33581
rect 39209 33541 39221 33575
rect 39255 33572 39267 33575
rect 39298 33572 39304 33584
rect 39255 33544 39304 33572
rect 39255 33541 39267 33544
rect 39209 33535 39267 33541
rect 39298 33532 39304 33544
rect 39356 33532 39362 33584
rect 37826 33464 37832 33516
rect 37884 33504 37890 33516
rect 38749 33507 38807 33513
rect 38749 33504 38761 33507
rect 37884 33476 38761 33504
rect 37884 33464 37890 33476
rect 38749 33473 38761 33476
rect 38795 33473 38807 33507
rect 40328 33504 40356 33612
rect 41966 33600 41972 33612
rect 42024 33600 42030 33652
rect 42610 33572 42616 33584
rect 41814 33544 42616 33572
rect 42610 33532 42616 33544
rect 42668 33572 42674 33584
rect 43990 33572 43996 33584
rect 42668 33544 43996 33572
rect 42668 33532 42674 33544
rect 43990 33532 43996 33544
rect 44048 33532 44054 33584
rect 38749 33467 38807 33473
rect 39316 33476 40356 33504
rect 34756 33408 35480 33436
rect 34756 33396 34762 33408
rect 35710 33396 35716 33448
rect 35768 33436 35774 33448
rect 37274 33436 37280 33448
rect 35768 33408 37280 33436
rect 35768 33396 35774 33408
rect 37274 33396 37280 33408
rect 37332 33396 37338 33448
rect 39316 33445 39344 33476
rect 38105 33439 38163 33445
rect 38105 33405 38117 33439
rect 38151 33405 38163 33439
rect 38105 33399 38163 33405
rect 39301 33439 39359 33445
rect 39301 33405 39313 33439
rect 39347 33405 39359 33439
rect 39301 33399 39359 33405
rect 36173 33371 36231 33377
rect 36173 33368 36185 33371
rect 27304 33340 28856 33368
rect 28966 33340 30512 33368
rect 35268 33340 36185 33368
rect 27304 33328 27310 33340
rect 28828 33312 28856 33340
rect 28810 33260 28816 33312
rect 28868 33260 28874 33312
rect 28948 33260 28954 33312
rect 29006 33300 29012 33312
rect 29178 33300 29184 33312
rect 29006 33272 29184 33300
rect 29006 33260 29012 33272
rect 29178 33260 29184 33272
rect 29236 33260 29242 33312
rect 29917 33303 29975 33309
rect 29917 33269 29929 33303
rect 29963 33300 29975 33303
rect 30098 33300 30104 33312
rect 29963 33272 30104 33300
rect 29963 33269 29975 33272
rect 29917 33263 29975 33269
rect 30098 33260 30104 33272
rect 30156 33260 30162 33312
rect 30650 33260 30656 33312
rect 30708 33300 30714 33312
rect 35268 33300 35296 33340
rect 36173 33337 36185 33340
rect 36219 33368 36231 33371
rect 36446 33368 36452 33380
rect 36219 33340 36452 33368
rect 36219 33337 36231 33340
rect 36173 33331 36231 33337
rect 36446 33328 36452 33340
rect 36504 33328 36510 33380
rect 38120 33368 38148 33399
rect 39390 33396 39396 33448
rect 39448 33396 39454 33448
rect 40310 33396 40316 33448
rect 40368 33396 40374 33448
rect 40586 33396 40592 33448
rect 40644 33436 40650 33448
rect 41874 33436 41880 33448
rect 40644 33408 41880 33436
rect 40644 33396 40650 33408
rect 41874 33396 41880 33408
rect 41932 33396 41938 33448
rect 38120 33340 40448 33368
rect 30708 33272 35296 33300
rect 35713 33303 35771 33309
rect 30708 33260 30714 33272
rect 35713 33269 35725 33303
rect 35759 33300 35771 33303
rect 38378 33300 38384 33312
rect 35759 33272 38384 33300
rect 35759 33269 35771 33272
rect 35713 33263 35771 33269
rect 38378 33260 38384 33272
rect 38436 33260 38442 33312
rect 38841 33303 38899 33309
rect 38841 33269 38853 33303
rect 38887 33300 38899 33303
rect 39022 33300 39028 33312
rect 38887 33272 39028 33300
rect 38887 33269 38899 33272
rect 38841 33263 38899 33269
rect 39022 33260 39028 33272
rect 39080 33260 39086 33312
rect 40420 33300 40448 33340
rect 40954 33300 40960 33312
rect 40420 33272 40960 33300
rect 40954 33260 40960 33272
rect 41012 33260 41018 33312
rect 42061 33303 42119 33309
rect 42061 33269 42073 33303
rect 42107 33300 42119 33303
rect 42150 33300 42156 33312
rect 42107 33272 42156 33300
rect 42107 33269 42119 33272
rect 42061 33263 42119 33269
rect 42150 33260 42156 33272
rect 42208 33260 42214 33312
rect 1104 33210 49864 33232
rect 1104 33158 2950 33210
rect 3002 33158 3014 33210
rect 3066 33158 3078 33210
rect 3130 33158 3142 33210
rect 3194 33158 3206 33210
rect 3258 33158 12950 33210
rect 13002 33158 13014 33210
rect 13066 33158 13078 33210
rect 13130 33158 13142 33210
rect 13194 33158 13206 33210
rect 13258 33158 22950 33210
rect 23002 33158 23014 33210
rect 23066 33158 23078 33210
rect 23130 33158 23142 33210
rect 23194 33158 23206 33210
rect 23258 33158 32950 33210
rect 33002 33158 33014 33210
rect 33066 33158 33078 33210
rect 33130 33158 33142 33210
rect 33194 33158 33206 33210
rect 33258 33158 42950 33210
rect 43002 33158 43014 33210
rect 43066 33158 43078 33210
rect 43130 33158 43142 33210
rect 43194 33158 43206 33210
rect 43258 33158 49864 33210
rect 1104 33136 49864 33158
rect 27798 33056 27804 33108
rect 27856 33096 27862 33108
rect 28445 33099 28503 33105
rect 28445 33096 28457 33099
rect 27856 33068 28457 33096
rect 27856 33056 27862 33068
rect 28445 33065 28457 33068
rect 28491 33065 28503 33099
rect 28445 33059 28503 33065
rect 30282 33056 30288 33108
rect 30340 33096 30346 33108
rect 31478 33096 31484 33108
rect 30340 33068 31484 33096
rect 30340 33056 30346 33068
rect 31478 33056 31484 33068
rect 31536 33056 31542 33108
rect 34790 33056 34796 33108
rect 34848 33096 34854 33108
rect 37645 33099 37703 33105
rect 34848 33068 37228 33096
rect 34848 33056 34854 33068
rect 23750 32988 23756 33040
rect 23808 33028 23814 33040
rect 29733 33031 29791 33037
rect 29733 33028 29745 33031
rect 23808 33000 29745 33028
rect 23808 32988 23814 33000
rect 29733 32997 29745 33000
rect 29779 32997 29791 33031
rect 34885 33031 34943 33037
rect 29733 32991 29791 32997
rect 30116 33000 34836 33028
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 23934 32960 23940 32972
rect 22603 32932 23940 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 23934 32920 23940 32932
rect 23992 32920 23998 32972
rect 24029 32963 24087 32969
rect 24029 32929 24041 32963
rect 24075 32929 24087 32963
rect 24029 32923 24087 32929
rect 22278 32852 22284 32904
rect 22336 32852 22342 32904
rect 23842 32852 23848 32904
rect 23900 32892 23906 32904
rect 24044 32892 24072 32923
rect 24302 32920 24308 32972
rect 24360 32960 24366 32972
rect 26970 32960 26976 32972
rect 24360 32932 26976 32960
rect 24360 32920 24366 32932
rect 26970 32920 26976 32932
rect 27028 32960 27034 32972
rect 27065 32963 27123 32969
rect 27065 32960 27077 32963
rect 27028 32932 27077 32960
rect 27028 32920 27034 32932
rect 27065 32929 27077 32932
rect 27111 32929 27123 32963
rect 27065 32923 27123 32929
rect 27246 32920 27252 32972
rect 27304 32920 27310 32972
rect 28626 32960 28632 32972
rect 27356 32932 28632 32960
rect 27356 32892 27384 32932
rect 28626 32920 28632 32932
rect 28684 32920 28690 32972
rect 28997 32963 29055 32969
rect 28997 32960 29009 32963
rect 28736 32932 29009 32960
rect 28736 32904 28764 32932
rect 28997 32929 29009 32932
rect 29043 32929 29055 32963
rect 28997 32923 29055 32929
rect 23900 32864 27384 32892
rect 23900 32852 23906 32864
rect 28718 32852 28724 32904
rect 28776 32852 28782 32904
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 30116 32892 30144 33000
rect 30190 32920 30196 32972
rect 30248 32920 30254 32972
rect 30285 32963 30343 32969
rect 30285 32929 30297 32963
rect 30331 32929 30343 32963
rect 30285 32923 30343 32929
rect 28859 32864 30144 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 22830 32784 22836 32836
rect 22888 32824 22894 32836
rect 26053 32827 26111 32833
rect 26053 32824 26065 32827
rect 22888 32796 23046 32824
rect 23952 32796 26065 32824
rect 22888 32784 22894 32796
rect 21542 32716 21548 32768
rect 21600 32756 21606 32768
rect 23952 32756 23980 32796
rect 26053 32793 26065 32796
rect 26099 32824 26111 32827
rect 26418 32824 26424 32836
rect 26099 32796 26424 32824
rect 26099 32793 26111 32796
rect 26053 32787 26111 32793
rect 26418 32784 26424 32796
rect 26476 32824 26482 32836
rect 26973 32827 27031 32833
rect 26973 32824 26985 32827
rect 26476 32796 26985 32824
rect 26476 32784 26482 32796
rect 26973 32793 26985 32796
rect 27019 32793 27031 32827
rect 26973 32787 27031 32793
rect 28902 32784 28908 32836
rect 28960 32784 28966 32836
rect 28994 32784 29000 32836
rect 29052 32824 29058 32836
rect 30300 32824 30328 32923
rect 31294 32920 31300 32972
rect 31352 32960 31358 32972
rect 31389 32963 31447 32969
rect 31389 32960 31401 32963
rect 31352 32932 31401 32960
rect 31352 32920 31358 32932
rect 31389 32929 31401 32932
rect 31435 32929 31447 32963
rect 31389 32923 31447 32929
rect 31478 32920 31484 32972
rect 31536 32920 31542 32972
rect 34808 32960 34836 33000
rect 34885 32997 34897 33031
rect 34931 33028 34943 33031
rect 37200 33028 37228 33068
rect 37645 33065 37657 33099
rect 37691 33096 37703 33099
rect 40586 33096 40592 33108
rect 37691 33068 40592 33096
rect 37691 33065 37703 33068
rect 37645 33059 37703 33065
rect 40586 33056 40592 33068
rect 40644 33056 40650 33108
rect 40862 33056 40868 33108
rect 40920 33096 40926 33108
rect 48774 33096 48780 33108
rect 40920 33068 48780 33096
rect 40920 33056 40926 33068
rect 48774 33056 48780 33068
rect 48832 33056 48838 33108
rect 38381 33031 38439 33037
rect 38381 33028 38393 33031
rect 34931 33000 36032 33028
rect 37200 33000 38393 33028
rect 34931 32997 34943 33000
rect 34885 32991 34943 32997
rect 35434 32960 35440 32972
rect 34808 32932 35440 32960
rect 35434 32920 35440 32932
rect 35492 32920 35498 32972
rect 35529 32963 35587 32969
rect 35529 32929 35541 32963
rect 35575 32960 35587 32963
rect 35710 32960 35716 32972
rect 35575 32932 35716 32960
rect 35575 32929 35587 32932
rect 35529 32923 35587 32929
rect 35710 32920 35716 32932
rect 35768 32920 35774 32972
rect 36004 32960 36032 33000
rect 38381 32997 38393 33000
rect 38427 32997 38439 33031
rect 38381 32991 38439 32997
rect 38562 32988 38568 33040
rect 38620 33028 38626 33040
rect 43714 33028 43720 33040
rect 38620 33000 40448 33028
rect 38620 32988 38626 33000
rect 37734 32960 37740 32972
rect 36004 32932 37740 32960
rect 37734 32920 37740 32932
rect 37792 32920 37798 32972
rect 38746 32920 38752 32972
rect 38804 32960 38810 32972
rect 38841 32963 38899 32969
rect 38841 32960 38853 32963
rect 38804 32932 38853 32960
rect 38804 32920 38810 32932
rect 38841 32929 38853 32932
rect 38887 32929 38899 32963
rect 38841 32923 38899 32929
rect 38930 32920 38936 32972
rect 38988 32920 38994 32972
rect 40420 32960 40448 33000
rect 40696 33000 43720 33028
rect 40696 32960 40724 33000
rect 43714 32988 43720 33000
rect 43772 32988 43778 33040
rect 40420 32932 40724 32960
rect 40957 32963 41015 32969
rect 40957 32929 40969 32963
rect 41003 32929 41015 32963
rect 40957 32923 41015 32929
rect 29052 32796 30328 32824
rect 30852 32864 31616 32892
rect 29052 32784 29058 32796
rect 21600 32728 23980 32756
rect 21600 32716 21606 32728
rect 24026 32716 24032 32768
rect 24084 32756 24090 32768
rect 24486 32756 24492 32768
rect 24084 32728 24492 32756
rect 24084 32716 24090 32728
rect 24486 32716 24492 32728
rect 24544 32756 24550 32768
rect 26510 32756 26516 32768
rect 24544 32728 26516 32756
rect 24544 32716 24550 32728
rect 26510 32716 26516 32728
rect 26568 32716 26574 32768
rect 26602 32716 26608 32768
rect 26660 32716 26666 32768
rect 28718 32716 28724 32768
rect 28776 32756 28782 32768
rect 29270 32756 29276 32768
rect 28776 32728 29276 32756
rect 28776 32716 28782 32728
rect 29270 32716 29276 32728
rect 29328 32716 29334 32768
rect 30101 32759 30159 32765
rect 30101 32725 30113 32759
rect 30147 32756 30159 32759
rect 30852 32756 30880 32864
rect 31588 32824 31616 32864
rect 31754 32852 31760 32904
rect 31812 32892 31818 32904
rect 32306 32892 32312 32904
rect 31812 32864 32312 32892
rect 31812 32852 31818 32864
rect 32306 32852 32312 32864
rect 32364 32852 32370 32904
rect 34517 32895 34575 32901
rect 34517 32861 34529 32895
rect 34563 32892 34575 32895
rect 35253 32895 35311 32901
rect 35253 32892 35265 32895
rect 34563 32864 35265 32892
rect 34563 32861 34575 32864
rect 34517 32855 34575 32861
rect 35253 32861 35265 32864
rect 35299 32861 35311 32895
rect 35253 32855 35311 32861
rect 35894 32852 35900 32904
rect 35952 32852 35958 32904
rect 37826 32852 37832 32904
rect 37884 32892 37890 32904
rect 40586 32892 40592 32904
rect 37884 32864 40592 32892
rect 37884 32852 37890 32864
rect 40586 32852 40592 32864
rect 40644 32852 40650 32904
rect 40678 32852 40684 32904
rect 40736 32892 40742 32904
rect 40773 32895 40831 32901
rect 40773 32892 40785 32895
rect 40736 32864 40785 32892
rect 40736 32852 40742 32864
rect 40773 32861 40785 32864
rect 40819 32861 40831 32895
rect 40773 32855 40831 32861
rect 30944 32796 31524 32824
rect 31588 32796 32812 32824
rect 30944 32765 30972 32796
rect 30147 32728 30880 32756
rect 30929 32759 30987 32765
rect 30147 32725 30159 32728
rect 30101 32719 30159 32725
rect 30929 32725 30941 32759
rect 30975 32725 30987 32759
rect 30929 32719 30987 32725
rect 31294 32716 31300 32768
rect 31352 32716 31358 32768
rect 31496 32756 31524 32796
rect 32214 32756 32220 32768
rect 31496 32728 32220 32756
rect 32214 32716 32220 32728
rect 32272 32716 32278 32768
rect 32784 32756 32812 32796
rect 35710 32784 35716 32836
rect 35768 32824 35774 32836
rect 36173 32827 36231 32833
rect 36173 32824 36185 32827
rect 35768 32796 36185 32824
rect 35768 32784 35774 32796
rect 36173 32793 36185 32796
rect 36219 32793 36231 32827
rect 36173 32787 36231 32793
rect 36630 32784 36636 32836
rect 36688 32784 36694 32836
rect 40972 32824 41000 32923
rect 42058 32920 42064 32972
rect 42116 32920 42122 32972
rect 42242 32920 42248 32972
rect 42300 32920 42306 32972
rect 41966 32852 41972 32904
rect 42024 32852 42030 32904
rect 43806 32852 43812 32904
rect 43864 32852 43870 32904
rect 49326 32852 49332 32904
rect 49384 32852 49390 32904
rect 37752 32796 41000 32824
rect 34606 32756 34612 32768
rect 32784 32728 34612 32756
rect 34606 32716 34612 32728
rect 34664 32716 34670 32768
rect 35342 32716 35348 32768
rect 35400 32716 35406 32768
rect 37182 32716 37188 32768
rect 37240 32756 37246 32768
rect 37752 32756 37780 32796
rect 41322 32784 41328 32836
rect 41380 32824 41386 32836
rect 41414 32824 41420 32836
rect 41380 32796 41420 32824
rect 41380 32784 41386 32796
rect 41414 32784 41420 32796
rect 41472 32784 41478 32836
rect 37240 32728 37780 32756
rect 38749 32759 38807 32765
rect 37240 32716 37246 32728
rect 38749 32725 38761 32759
rect 38795 32756 38807 32759
rect 39114 32756 39120 32768
rect 38795 32728 39120 32756
rect 38795 32725 38807 32728
rect 38749 32719 38807 32725
rect 39114 32716 39120 32728
rect 39172 32716 39178 32768
rect 40126 32716 40132 32768
rect 40184 32756 40190 32768
rect 40405 32759 40463 32765
rect 40405 32756 40417 32759
rect 40184 32728 40417 32756
rect 40184 32716 40190 32728
rect 40405 32725 40417 32728
rect 40451 32725 40463 32759
rect 40405 32719 40463 32725
rect 40494 32716 40500 32768
rect 40552 32756 40558 32768
rect 40865 32759 40923 32765
rect 40865 32756 40877 32759
rect 40552 32728 40877 32756
rect 40552 32716 40558 32728
rect 40865 32725 40877 32728
rect 40911 32725 40923 32759
rect 40865 32719 40923 32725
rect 40954 32716 40960 32768
rect 41012 32756 41018 32768
rect 41601 32759 41659 32765
rect 41601 32756 41613 32759
rect 41012 32728 41613 32756
rect 41012 32716 41018 32728
rect 41601 32725 41613 32728
rect 41647 32725 41659 32759
rect 41601 32719 41659 32725
rect 43625 32759 43683 32765
rect 43625 32725 43637 32759
rect 43671 32756 43683 32759
rect 46382 32756 46388 32768
rect 43671 32728 46388 32756
rect 43671 32725 43683 32728
rect 43625 32719 43683 32725
rect 46382 32716 46388 32728
rect 46440 32716 46446 32768
rect 49142 32716 49148 32768
rect 49200 32716 49206 32768
rect 1104 32666 49864 32688
rect 1104 32614 7950 32666
rect 8002 32614 8014 32666
rect 8066 32614 8078 32666
rect 8130 32614 8142 32666
rect 8194 32614 8206 32666
rect 8258 32614 17950 32666
rect 18002 32614 18014 32666
rect 18066 32614 18078 32666
rect 18130 32614 18142 32666
rect 18194 32614 18206 32666
rect 18258 32614 27950 32666
rect 28002 32614 28014 32666
rect 28066 32614 28078 32666
rect 28130 32614 28142 32666
rect 28194 32614 28206 32666
rect 28258 32614 37950 32666
rect 38002 32614 38014 32666
rect 38066 32614 38078 32666
rect 38130 32614 38142 32666
rect 38194 32614 38206 32666
rect 38258 32614 47950 32666
rect 48002 32614 48014 32666
rect 48066 32614 48078 32666
rect 48130 32614 48142 32666
rect 48194 32614 48206 32666
rect 48258 32614 49864 32666
rect 1104 32592 49864 32614
rect 17218 32512 17224 32564
rect 17276 32512 17282 32564
rect 25222 32512 25228 32564
rect 25280 32552 25286 32564
rect 25685 32555 25743 32561
rect 25685 32552 25697 32555
rect 25280 32524 25697 32552
rect 25280 32512 25286 32524
rect 25685 32521 25697 32524
rect 25731 32552 25743 32555
rect 26050 32552 26056 32564
rect 25731 32524 26056 32552
rect 25731 32521 25743 32524
rect 25685 32515 25743 32521
rect 26050 32512 26056 32524
rect 26108 32512 26114 32564
rect 27249 32555 27307 32561
rect 27249 32521 27261 32555
rect 27295 32552 27307 32555
rect 31294 32552 31300 32564
rect 27295 32524 31300 32552
rect 27295 32521 27307 32524
rect 27249 32515 27307 32521
rect 31294 32512 31300 32524
rect 31352 32512 31358 32564
rect 35069 32555 35127 32561
rect 35069 32521 35081 32555
rect 35115 32552 35127 32555
rect 36538 32552 36544 32564
rect 35115 32524 36544 32552
rect 35115 32521 35127 32524
rect 35069 32515 35127 32521
rect 36538 32512 36544 32524
rect 36596 32512 36602 32564
rect 39574 32512 39580 32564
rect 39632 32552 39638 32564
rect 41322 32552 41328 32564
rect 39632 32524 41328 32552
rect 39632 32512 39638 32524
rect 41322 32512 41328 32524
rect 41380 32512 41386 32564
rect 41506 32512 41512 32564
rect 41564 32552 41570 32564
rect 47118 32552 47124 32564
rect 41564 32524 47124 32552
rect 41564 32512 41570 32524
rect 47118 32512 47124 32524
rect 47176 32512 47182 32564
rect 22830 32444 22836 32496
rect 22888 32484 22894 32496
rect 24670 32484 24676 32496
rect 22888 32456 24676 32484
rect 22888 32444 22894 32456
rect 24670 32444 24676 32456
rect 24728 32444 24734 32496
rect 26510 32444 26516 32496
rect 26568 32484 26574 32496
rect 27709 32487 27767 32493
rect 27709 32484 27721 32487
rect 26568 32456 27721 32484
rect 26568 32444 26574 32456
rect 27709 32453 27721 32456
rect 27755 32484 27767 32487
rect 28445 32487 28503 32493
rect 28445 32484 28457 32487
rect 27755 32456 28457 32484
rect 27755 32453 27767 32456
rect 27709 32447 27767 32453
rect 28445 32453 28457 32456
rect 28491 32484 28503 32487
rect 29086 32484 29092 32496
rect 28491 32456 28856 32484
rect 28491 32453 28503 32456
rect 28445 32447 28503 32453
rect 934 32376 940 32428
rect 992 32416 998 32428
rect 1765 32419 1823 32425
rect 1765 32416 1777 32419
rect 992 32388 1777 32416
rect 992 32376 998 32388
rect 1765 32385 1777 32388
rect 1811 32385 1823 32419
rect 1765 32379 1823 32385
rect 17589 32419 17647 32425
rect 17589 32385 17601 32419
rect 17635 32416 17647 32419
rect 18785 32419 18843 32425
rect 18785 32416 18797 32419
rect 17635 32388 18797 32416
rect 17635 32385 17647 32388
rect 17589 32379 17647 32385
rect 18785 32385 18797 32388
rect 18831 32385 18843 32419
rect 18785 32379 18843 32385
rect 27617 32419 27675 32425
rect 27617 32385 27629 32419
rect 27663 32416 27675 32419
rect 28828 32416 28856 32456
rect 28966 32456 29092 32484
rect 28966 32416 28994 32456
rect 29086 32444 29092 32456
rect 29144 32444 29150 32496
rect 34698 32484 34704 32496
rect 33994 32456 34704 32484
rect 34698 32444 34704 32456
rect 34756 32444 34762 32496
rect 35161 32487 35219 32493
rect 35161 32453 35173 32487
rect 35207 32484 35219 32487
rect 35618 32484 35624 32496
rect 35207 32456 35624 32484
rect 35207 32453 35219 32456
rect 35161 32447 35219 32453
rect 35618 32444 35624 32456
rect 35676 32444 35682 32496
rect 36630 32444 36636 32496
rect 36688 32484 36694 32496
rect 40034 32484 40040 32496
rect 36688 32456 40040 32484
rect 36688 32444 36694 32456
rect 40034 32444 40040 32456
rect 40092 32444 40098 32496
rect 41414 32484 41420 32496
rect 40986 32456 41420 32484
rect 41414 32444 41420 32456
rect 41472 32484 41478 32496
rect 42610 32484 42616 32496
rect 41472 32456 42616 32484
rect 41472 32444 41478 32456
rect 42610 32444 42616 32456
rect 42668 32444 42674 32496
rect 27663 32388 28672 32416
rect 28828 32388 28994 32416
rect 27663 32385 27675 32388
rect 27617 32379 27675 32385
rect 5718 32308 5724 32360
rect 5776 32348 5782 32360
rect 17681 32351 17739 32357
rect 17681 32348 17693 32351
rect 5776 32320 17693 32348
rect 5776 32308 5782 32320
rect 17681 32317 17693 32320
rect 17727 32317 17739 32351
rect 17681 32311 17739 32317
rect 1581 32215 1639 32221
rect 1581 32181 1593 32215
rect 1627 32212 1639 32215
rect 7466 32212 7472 32224
rect 1627 32184 7472 32212
rect 1627 32181 1639 32184
rect 1581 32175 1639 32181
rect 7466 32172 7472 32184
rect 7524 32172 7530 32224
rect 17696 32212 17724 32311
rect 17862 32308 17868 32360
rect 17920 32308 17926 32360
rect 23937 32351 23995 32357
rect 23937 32317 23949 32351
rect 23983 32317 23995 32351
rect 23937 32311 23995 32317
rect 18506 32212 18512 32224
rect 17696 32184 18512 32212
rect 18506 32172 18512 32184
rect 18564 32172 18570 32224
rect 22554 32172 22560 32224
rect 22612 32212 22618 32224
rect 23952 32212 23980 32311
rect 24210 32308 24216 32360
rect 24268 32308 24274 32360
rect 24670 32308 24676 32360
rect 24728 32348 24734 32360
rect 26234 32348 26240 32360
rect 24728 32320 26240 32348
rect 24728 32308 24734 32320
rect 26234 32308 26240 32320
rect 26292 32308 26298 32360
rect 27893 32351 27951 32357
rect 27893 32317 27905 32351
rect 27939 32348 27951 32351
rect 28534 32348 28540 32360
rect 27939 32320 28540 32348
rect 27939 32317 27951 32320
rect 27893 32311 27951 32317
rect 28534 32308 28540 32320
rect 28592 32308 28598 32360
rect 28644 32348 28672 32388
rect 34606 32376 34612 32428
rect 34664 32416 34670 32428
rect 37458 32416 37464 32428
rect 34664 32388 37464 32416
rect 34664 32376 34670 32388
rect 37458 32376 37464 32388
rect 37516 32376 37522 32428
rect 44082 32376 44088 32428
rect 44140 32416 44146 32428
rect 44821 32419 44879 32425
rect 44821 32416 44833 32419
rect 44140 32388 44833 32416
rect 44140 32376 44146 32388
rect 44821 32385 44833 32388
rect 44867 32385 44879 32419
rect 44821 32379 44879 32385
rect 48774 32376 48780 32428
rect 48832 32376 48838 32428
rect 28813 32351 28871 32357
rect 28813 32348 28825 32351
rect 28644 32320 28825 32348
rect 28813 32317 28825 32320
rect 28859 32317 28871 32351
rect 28813 32311 28871 32317
rect 31938 32308 31944 32360
rect 31996 32348 32002 32360
rect 32493 32351 32551 32357
rect 32493 32348 32505 32351
rect 31996 32320 32505 32348
rect 31996 32308 32002 32320
rect 32493 32317 32505 32320
rect 32539 32317 32551 32351
rect 32493 32311 32551 32317
rect 32769 32351 32827 32357
rect 32769 32317 32781 32351
rect 32815 32348 32827 32351
rect 32815 32320 35112 32348
rect 32815 32317 32827 32320
rect 32769 32311 32827 32317
rect 26602 32240 26608 32292
rect 26660 32280 26666 32292
rect 28718 32280 28724 32292
rect 26660 32252 28724 32280
rect 26660 32240 26666 32252
rect 28718 32240 28724 32252
rect 28776 32240 28782 32292
rect 34238 32240 34244 32292
rect 34296 32280 34302 32292
rect 34974 32280 34980 32292
rect 34296 32252 34980 32280
rect 34296 32240 34302 32252
rect 34974 32240 34980 32252
rect 35032 32240 35038 32292
rect 35084 32280 35112 32320
rect 35158 32308 35164 32360
rect 35216 32348 35222 32360
rect 35253 32351 35311 32357
rect 35253 32348 35265 32351
rect 35216 32320 35265 32348
rect 35216 32308 35222 32320
rect 35253 32317 35265 32320
rect 35299 32317 35311 32351
rect 35253 32311 35311 32317
rect 39022 32308 39028 32360
rect 39080 32348 39086 32360
rect 39485 32351 39543 32357
rect 39485 32348 39497 32351
rect 39080 32320 39497 32348
rect 39080 32308 39086 32320
rect 39485 32317 39497 32320
rect 39531 32317 39543 32351
rect 39485 32311 39543 32317
rect 39761 32351 39819 32357
rect 39761 32317 39773 32351
rect 39807 32348 39819 32351
rect 42150 32348 42156 32360
rect 39807 32320 42156 32348
rect 39807 32317 39819 32320
rect 39761 32311 39819 32317
rect 42150 32308 42156 32320
rect 42208 32308 42214 32360
rect 48498 32308 48504 32360
rect 48556 32308 48562 32360
rect 36078 32280 36084 32292
rect 35084 32252 36084 32280
rect 36078 32240 36084 32252
rect 36136 32280 36142 32292
rect 38470 32280 38476 32292
rect 36136 32252 38476 32280
rect 36136 32240 36142 32252
rect 38470 32240 38476 32252
rect 38528 32240 38534 32292
rect 41322 32240 41328 32292
rect 41380 32280 41386 32292
rect 49142 32280 49148 32292
rect 41380 32252 49148 32280
rect 41380 32240 41386 32252
rect 49142 32240 49148 32252
rect 49200 32240 49206 32292
rect 24854 32212 24860 32224
rect 22612 32184 24860 32212
rect 22612 32172 22618 32184
rect 24854 32172 24860 32184
rect 24912 32172 24918 32224
rect 32122 32172 32128 32224
rect 32180 32212 32186 32224
rect 34701 32215 34759 32221
rect 34701 32212 34713 32215
rect 32180 32184 34713 32212
rect 32180 32172 32186 32184
rect 34701 32181 34713 32184
rect 34747 32181 34759 32215
rect 34701 32175 34759 32181
rect 34882 32172 34888 32224
rect 34940 32212 34946 32224
rect 35710 32212 35716 32224
rect 34940 32184 35716 32212
rect 34940 32172 34946 32184
rect 35710 32172 35716 32184
rect 35768 32172 35774 32224
rect 39942 32172 39948 32224
rect 40000 32212 40006 32224
rect 41233 32215 41291 32221
rect 41233 32212 41245 32215
rect 40000 32184 41245 32212
rect 40000 32172 40006 32184
rect 41233 32181 41245 32184
rect 41279 32181 41291 32215
rect 41233 32175 41291 32181
rect 42794 32172 42800 32224
rect 42852 32172 42858 32224
rect 44634 32172 44640 32224
rect 44692 32172 44698 32224
rect 1104 32122 49864 32144
rect 1104 32070 2950 32122
rect 3002 32070 3014 32122
rect 3066 32070 3078 32122
rect 3130 32070 3142 32122
rect 3194 32070 3206 32122
rect 3258 32070 12950 32122
rect 13002 32070 13014 32122
rect 13066 32070 13078 32122
rect 13130 32070 13142 32122
rect 13194 32070 13206 32122
rect 13258 32070 22950 32122
rect 23002 32070 23014 32122
rect 23066 32070 23078 32122
rect 23130 32070 23142 32122
rect 23194 32070 23206 32122
rect 23258 32070 32950 32122
rect 33002 32070 33014 32122
rect 33066 32070 33078 32122
rect 33130 32070 33142 32122
rect 33194 32070 33206 32122
rect 33258 32070 42950 32122
rect 43002 32070 43014 32122
rect 43066 32070 43078 32122
rect 43130 32070 43142 32122
rect 43194 32070 43206 32122
rect 43258 32070 49864 32122
rect 1104 32048 49864 32070
rect 22554 32008 22560 32020
rect 22388 31980 22560 32008
rect 22281 31875 22339 31881
rect 22281 31841 22293 31875
rect 22327 31872 22339 31875
rect 22388 31872 22416 31980
rect 22554 31968 22560 31980
rect 22612 31968 22618 32020
rect 23934 31968 23940 32020
rect 23992 32008 23998 32020
rect 24029 32011 24087 32017
rect 24029 32008 24041 32011
rect 23992 31980 24041 32008
rect 23992 31968 23998 31980
rect 24029 31977 24041 31980
rect 24075 31977 24087 32011
rect 27062 32008 27068 32020
rect 24029 31971 24087 31977
rect 25792 31980 27068 32008
rect 22327 31844 22416 31872
rect 22557 31875 22615 31881
rect 22327 31841 22339 31844
rect 22281 31835 22339 31841
rect 22557 31841 22569 31875
rect 22603 31872 22615 31875
rect 23842 31872 23848 31884
rect 22603 31844 23848 31872
rect 22603 31841 22615 31844
rect 22557 31835 22615 31841
rect 23842 31832 23848 31844
rect 23900 31832 23906 31884
rect 25792 31881 25820 31980
rect 27062 31968 27068 31980
rect 27120 31968 27126 32020
rect 28442 31968 28448 32020
rect 28500 31968 28506 32020
rect 34330 31968 34336 32020
rect 34388 32008 34394 32020
rect 39301 32011 39359 32017
rect 34388 31980 38976 32008
rect 34388 31968 34394 31980
rect 31662 31940 31668 31952
rect 27816 31912 31668 31940
rect 25777 31875 25835 31881
rect 25777 31841 25789 31875
rect 25823 31841 25835 31875
rect 25777 31835 25835 31841
rect 26050 31832 26056 31884
rect 26108 31832 26114 31884
rect 27246 31832 27252 31884
rect 27304 31872 27310 31884
rect 27816 31881 27844 31912
rect 31662 31900 31668 31912
rect 31720 31940 31726 31952
rect 32030 31940 32036 31952
rect 31720 31912 32036 31940
rect 31720 31900 31726 31912
rect 32030 31900 32036 31912
rect 32088 31900 32094 31952
rect 32309 31943 32367 31949
rect 32309 31909 32321 31943
rect 32355 31940 32367 31943
rect 32355 31912 34100 31940
rect 32355 31909 32367 31912
rect 32309 31903 32367 31909
rect 27801 31875 27859 31881
rect 27801 31872 27813 31875
rect 27304 31844 27813 31872
rect 27304 31832 27310 31844
rect 27801 31841 27813 31844
rect 27847 31841 27859 31875
rect 27801 31835 27859 31841
rect 28626 31832 28632 31884
rect 28684 31872 28690 31884
rect 28997 31875 29055 31881
rect 28997 31872 29009 31875
rect 28684 31844 29009 31872
rect 28684 31832 28690 31844
rect 28997 31841 29009 31844
rect 29043 31841 29055 31875
rect 28997 31835 29055 31841
rect 31754 31832 31760 31884
rect 31812 31872 31818 31884
rect 32769 31875 32827 31881
rect 32769 31872 32781 31875
rect 31812 31844 32781 31872
rect 31812 31832 31818 31844
rect 32769 31841 32781 31844
rect 32815 31841 32827 31875
rect 32769 31835 32827 31841
rect 32953 31875 33011 31881
rect 32953 31841 32965 31875
rect 32999 31872 33011 31875
rect 33686 31872 33692 31884
rect 32999 31844 33692 31872
rect 32999 31841 33011 31844
rect 32953 31835 33011 31841
rect 33686 31832 33692 31844
rect 33744 31832 33750 31884
rect 34072 31872 34100 31912
rect 35250 31900 35256 31952
rect 35308 31940 35314 31952
rect 35345 31943 35403 31949
rect 35345 31940 35357 31943
rect 35308 31912 35357 31940
rect 35308 31900 35314 31912
rect 35345 31909 35357 31912
rect 35391 31909 35403 31943
rect 35345 31903 35403 31909
rect 36262 31900 36268 31952
rect 36320 31940 36326 31952
rect 36722 31940 36728 31952
rect 36320 31912 36728 31940
rect 36320 31900 36326 31912
rect 36722 31900 36728 31912
rect 36780 31900 36786 31952
rect 37921 31943 37979 31949
rect 37921 31909 37933 31943
rect 37967 31940 37979 31943
rect 38654 31940 38660 31952
rect 37967 31912 38660 31940
rect 37967 31909 37979 31912
rect 37921 31903 37979 31909
rect 38654 31900 38660 31912
rect 38712 31900 38718 31952
rect 35805 31875 35863 31881
rect 35805 31872 35817 31875
rect 34072 31844 35817 31872
rect 35805 31841 35817 31844
rect 35851 31841 35863 31875
rect 35805 31835 35863 31841
rect 35989 31875 36047 31881
rect 35989 31841 36001 31875
rect 36035 31872 36047 31875
rect 36170 31872 36176 31884
rect 36035 31844 36176 31872
rect 36035 31841 36047 31844
rect 35989 31835 36047 31841
rect 36170 31832 36176 31844
rect 36228 31832 36234 31884
rect 37274 31832 37280 31884
rect 37332 31872 37338 31884
rect 37642 31872 37648 31884
rect 37332 31844 37648 31872
rect 37332 31832 37338 31844
rect 37642 31832 37648 31844
rect 37700 31872 37706 31884
rect 37700 31844 37964 31872
rect 37700 31832 37706 31844
rect 21818 31764 21824 31816
rect 21876 31764 21882 31816
rect 24762 31764 24768 31816
rect 24820 31764 24826 31816
rect 28905 31807 28963 31813
rect 28905 31773 28917 31807
rect 28951 31804 28963 31807
rect 37826 31804 37832 31816
rect 28951 31776 37832 31804
rect 28951 31773 28963 31776
rect 28905 31767 28963 31773
rect 37826 31764 37832 31776
rect 37884 31764 37890 31816
rect 37936 31804 37964 31844
rect 38470 31832 38476 31884
rect 38528 31832 38534 31884
rect 38562 31832 38568 31884
rect 38620 31832 38626 31884
rect 38289 31807 38347 31813
rect 38289 31804 38301 31807
rect 37936 31776 38301 31804
rect 38289 31773 38301 31776
rect 38335 31773 38347 31807
rect 38289 31767 38347 31773
rect 38381 31807 38439 31813
rect 38381 31773 38393 31807
rect 38427 31804 38439 31807
rect 38580 31804 38608 31832
rect 38427 31776 38608 31804
rect 38948 31804 38976 31980
rect 39301 31977 39313 32011
rect 39347 32008 39359 32011
rect 43438 32008 43444 32020
rect 39347 31980 43444 32008
rect 39347 31977 39359 31980
rect 39301 31971 39359 31977
rect 43438 31968 43444 31980
rect 43496 31968 43502 32020
rect 43625 32011 43683 32017
rect 43625 31977 43637 32011
rect 43671 32008 43683 32011
rect 43898 32008 43904 32020
rect 43671 31980 43904 32008
rect 43671 31977 43683 31980
rect 43625 31971 43683 31977
rect 43898 31968 43904 31980
rect 43956 31968 43962 32020
rect 39022 31832 39028 31884
rect 39080 31872 39086 31884
rect 40310 31872 40316 31884
rect 39080 31844 40316 31872
rect 39080 31832 39086 31844
rect 40310 31832 40316 31844
rect 40368 31872 40374 31884
rect 41877 31875 41935 31881
rect 41877 31872 41889 31875
rect 40368 31844 41889 31872
rect 40368 31832 40374 31844
rect 41877 31841 41889 31844
rect 41923 31841 41935 31875
rect 41877 31835 41935 31841
rect 42153 31875 42211 31881
rect 42153 31841 42165 31875
rect 42199 31872 42211 31875
rect 42702 31872 42708 31884
rect 42199 31844 42708 31872
rect 42199 31841 42211 31844
rect 42153 31835 42211 31841
rect 42702 31832 42708 31844
rect 42760 31832 42766 31884
rect 47118 31832 47124 31884
rect 47176 31872 47182 31884
rect 48777 31875 48835 31881
rect 48777 31872 48789 31875
rect 47176 31844 48789 31872
rect 47176 31832 47182 31844
rect 48777 31841 48789 31844
rect 48823 31841 48835 31875
rect 48777 31835 48835 31841
rect 39485 31807 39543 31813
rect 39485 31804 39497 31807
rect 38948 31776 39497 31804
rect 38427 31773 38439 31776
rect 38381 31767 38439 31773
rect 39485 31773 39497 31776
rect 39531 31773 39543 31807
rect 39485 31767 39543 31773
rect 40034 31764 40040 31816
rect 40092 31804 40098 31816
rect 41506 31804 41512 31816
rect 40092 31776 41512 31804
rect 40092 31764 40098 31776
rect 41506 31764 41512 31776
rect 41564 31764 41570 31816
rect 48041 31807 48099 31813
rect 48041 31773 48053 31807
rect 48087 31804 48099 31807
rect 48498 31804 48504 31816
rect 48087 31776 48504 31804
rect 48087 31773 48099 31776
rect 48041 31767 48099 31773
rect 48498 31764 48504 31776
rect 48556 31764 48562 31816
rect 22830 31696 22836 31748
rect 22888 31736 22894 31748
rect 27522 31736 27528 31748
rect 22888 31708 23046 31736
rect 27278 31708 27528 31736
rect 22888 31696 22894 31708
rect 27522 31696 27528 31708
rect 27580 31696 27586 31748
rect 27798 31696 27804 31748
rect 27856 31736 27862 31748
rect 35713 31739 35771 31745
rect 27856 31708 31892 31736
rect 27856 31696 27862 31708
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 31864 31677 31892 31708
rect 35713 31705 35725 31739
rect 35759 31736 35771 31739
rect 40218 31736 40224 31748
rect 35759 31708 40224 31736
rect 35759 31705 35771 31708
rect 35713 31699 35771 31705
rect 40218 31696 40224 31708
rect 40276 31696 40282 31748
rect 42610 31696 42616 31748
rect 42668 31696 42674 31748
rect 28813 31671 28871 31677
rect 28813 31668 28825 31671
rect 27764 31640 28825 31668
rect 27764 31628 27770 31640
rect 28813 31637 28825 31640
rect 28859 31637 28871 31671
rect 28813 31631 28871 31637
rect 31849 31671 31907 31677
rect 31849 31637 31861 31671
rect 31895 31668 31907 31671
rect 32677 31671 32735 31677
rect 32677 31668 32689 31671
rect 31895 31640 32689 31668
rect 31895 31637 31907 31640
rect 31849 31631 31907 31637
rect 32677 31637 32689 31640
rect 32723 31637 32735 31671
rect 32677 31631 32735 31637
rect 34146 31628 34152 31680
rect 34204 31668 34210 31680
rect 35802 31668 35808 31680
rect 34204 31640 35808 31668
rect 34204 31628 34210 31640
rect 35802 31628 35808 31640
rect 35860 31668 35866 31680
rect 36630 31668 36636 31680
rect 35860 31640 36636 31668
rect 35860 31628 35866 31640
rect 36630 31628 36636 31640
rect 36688 31628 36694 31680
rect 38470 31628 38476 31680
rect 38528 31668 38534 31680
rect 41506 31668 41512 31680
rect 38528 31640 41512 31668
rect 38528 31628 38534 31640
rect 41506 31628 41512 31640
rect 41564 31628 41570 31680
rect 1104 31578 49864 31600
rect 1104 31526 7950 31578
rect 8002 31526 8014 31578
rect 8066 31526 8078 31578
rect 8130 31526 8142 31578
rect 8194 31526 8206 31578
rect 8258 31526 17950 31578
rect 18002 31526 18014 31578
rect 18066 31526 18078 31578
rect 18130 31526 18142 31578
rect 18194 31526 18206 31578
rect 18258 31526 27950 31578
rect 28002 31526 28014 31578
rect 28066 31526 28078 31578
rect 28130 31526 28142 31578
rect 28194 31526 28206 31578
rect 28258 31526 37950 31578
rect 38002 31526 38014 31578
rect 38066 31526 38078 31578
rect 38130 31526 38142 31578
rect 38194 31526 38206 31578
rect 38258 31526 47950 31578
rect 48002 31526 48014 31578
rect 48066 31526 48078 31578
rect 48130 31526 48142 31578
rect 48194 31526 48206 31578
rect 48258 31526 49864 31578
rect 1104 31504 49864 31526
rect 23474 31424 23480 31476
rect 23532 31424 23538 31476
rect 23845 31467 23903 31473
rect 23845 31433 23857 31467
rect 23891 31464 23903 31467
rect 24762 31464 24768 31476
rect 23891 31436 24768 31464
rect 23891 31433 23903 31436
rect 23845 31427 23903 31433
rect 24762 31424 24768 31436
rect 24820 31424 24826 31476
rect 25406 31424 25412 31476
rect 25464 31464 25470 31476
rect 26605 31467 26663 31473
rect 25464 31436 26556 31464
rect 25464 31424 25470 31436
rect 25038 31396 25044 31408
rect 22756 31368 25044 31396
rect 21453 31331 21511 31337
rect 21453 31297 21465 31331
rect 21499 31328 21511 31331
rect 22373 31331 22431 31337
rect 22373 31328 22385 31331
rect 21499 31300 22385 31328
rect 21499 31297 21511 31300
rect 21453 31291 21511 31297
rect 22373 31297 22385 31300
rect 22419 31297 22431 31331
rect 22373 31291 22431 31297
rect 22462 31220 22468 31272
rect 22520 31220 22526 31272
rect 22649 31263 22707 31269
rect 22649 31229 22661 31263
rect 22695 31260 22707 31263
rect 22756 31260 22784 31368
rect 25038 31356 25044 31368
rect 25096 31356 25102 31408
rect 24854 31288 24860 31340
rect 24912 31288 24918 31340
rect 26234 31288 26240 31340
rect 26292 31288 26298 31340
rect 26528 31328 26556 31436
rect 26605 31433 26617 31467
rect 26651 31464 26663 31467
rect 26694 31464 26700 31476
rect 26651 31436 26700 31464
rect 26651 31433 26663 31436
rect 26605 31427 26663 31433
rect 26694 31424 26700 31436
rect 26752 31424 26758 31476
rect 32030 31424 32036 31476
rect 32088 31464 32094 31476
rect 32088 31436 36032 31464
rect 32088 31424 32094 31436
rect 27154 31356 27160 31408
rect 27212 31396 27218 31408
rect 27212 31368 31754 31396
rect 27212 31356 27218 31368
rect 27798 31328 27804 31340
rect 26528 31300 27804 31328
rect 27798 31288 27804 31300
rect 27856 31288 27862 31340
rect 31726 31328 31754 31368
rect 34606 31356 34612 31408
rect 34664 31396 34670 31408
rect 36004 31396 36032 31436
rect 36078 31424 36084 31476
rect 36136 31464 36142 31476
rect 36173 31467 36231 31473
rect 36173 31464 36185 31467
rect 36136 31436 36185 31464
rect 36136 31424 36142 31436
rect 36173 31433 36185 31436
rect 36219 31433 36231 31467
rect 36173 31427 36231 31433
rect 36814 31424 36820 31476
rect 36872 31464 36878 31476
rect 36872 31436 38056 31464
rect 36872 31424 36878 31436
rect 37918 31396 37924 31408
rect 34664 31368 35190 31396
rect 36004 31368 37924 31396
rect 34664 31356 34670 31368
rect 37918 31356 37924 31368
rect 37976 31356 37982 31408
rect 38028 31396 38056 31436
rect 38562 31424 38568 31476
rect 38620 31424 38626 31476
rect 38654 31424 38660 31476
rect 38712 31464 38718 31476
rect 40034 31464 40040 31476
rect 38712 31436 40040 31464
rect 38712 31424 38718 31436
rect 40034 31424 40040 31436
rect 40092 31424 40098 31476
rect 40218 31424 40224 31476
rect 40276 31464 40282 31476
rect 41322 31464 41328 31476
rect 40276 31436 41328 31464
rect 40276 31424 40282 31436
rect 41322 31424 41328 31436
rect 41380 31424 41386 31476
rect 42794 31424 42800 31476
rect 42852 31464 42858 31476
rect 42981 31467 43039 31473
rect 42981 31464 42993 31467
rect 42852 31436 42993 31464
rect 42852 31424 42858 31436
rect 42981 31433 42993 31436
rect 43027 31433 43039 31467
rect 42981 31427 43039 31433
rect 43073 31399 43131 31405
rect 38028 31368 40816 31396
rect 33321 31331 33379 31337
rect 33321 31328 33333 31331
rect 31726 31300 33333 31328
rect 33321 31297 33333 31300
rect 33367 31297 33379 31331
rect 33321 31291 33379 31297
rect 33413 31331 33471 31337
rect 33413 31297 33425 31331
rect 33459 31328 33471 31331
rect 33594 31328 33600 31340
rect 33459 31300 33600 31328
rect 33459 31297 33471 31300
rect 33413 31291 33471 31297
rect 33594 31288 33600 31300
rect 33652 31288 33658 31340
rect 36538 31288 36544 31340
rect 36596 31328 36602 31340
rect 37737 31331 37795 31337
rect 37737 31328 37749 31331
rect 36596 31300 37749 31328
rect 36596 31288 36602 31300
rect 37737 31297 37749 31300
rect 37783 31297 37795 31331
rect 37737 31291 37795 31297
rect 38378 31288 38384 31340
rect 38436 31328 38442 31340
rect 38562 31328 38568 31340
rect 38436 31300 38568 31328
rect 38436 31288 38442 31300
rect 38562 31288 38568 31300
rect 38620 31328 38626 31340
rect 40788 31337 40816 31368
rect 43073 31365 43085 31399
rect 43119 31396 43131 31399
rect 43530 31396 43536 31408
rect 43119 31368 43536 31396
rect 43119 31365 43131 31368
rect 43073 31359 43131 31365
rect 43530 31356 43536 31368
rect 43588 31356 43594 31408
rect 40773 31331 40831 31337
rect 38620 31300 38792 31328
rect 38620 31288 38626 31300
rect 22695 31232 22784 31260
rect 22695 31229 22707 31232
rect 22649 31223 22707 31229
rect 22830 31220 22836 31272
rect 22888 31260 22894 31272
rect 23937 31263 23995 31269
rect 23937 31260 23949 31263
rect 22888 31232 23949 31260
rect 22888 31220 22894 31232
rect 23937 31229 23949 31232
rect 23983 31229 23995 31263
rect 23937 31223 23995 31229
rect 24121 31263 24179 31269
rect 24121 31229 24133 31263
rect 24167 31260 24179 31263
rect 24210 31260 24216 31272
rect 24167 31232 24216 31260
rect 24167 31229 24179 31232
rect 24121 31223 24179 31229
rect 24210 31220 24216 31232
rect 24268 31220 24274 31272
rect 25130 31220 25136 31272
rect 25188 31220 25194 31272
rect 22005 31127 22063 31133
rect 22005 31093 22017 31127
rect 22051 31124 22063 31127
rect 24946 31124 24952 31136
rect 22051 31096 24952 31124
rect 22051 31093 22063 31096
rect 22005 31087 22063 31093
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 26252 31124 26280 31288
rect 32030 31220 32036 31272
rect 32088 31260 32094 31272
rect 32398 31260 32404 31272
rect 32088 31232 32404 31260
rect 32088 31220 32094 31232
rect 32398 31220 32404 31232
rect 32456 31220 32462 31272
rect 32674 31220 32680 31272
rect 32732 31260 32738 31272
rect 33505 31263 33563 31269
rect 33505 31260 33517 31263
rect 32732 31232 33517 31260
rect 32732 31220 32738 31232
rect 33505 31229 33517 31232
rect 33551 31260 33563 31263
rect 34330 31260 34336 31272
rect 33551 31232 34336 31260
rect 33551 31229 33563 31232
rect 33505 31223 33563 31229
rect 34330 31220 34336 31232
rect 34388 31220 34394 31272
rect 34425 31263 34483 31269
rect 34425 31229 34437 31263
rect 34471 31229 34483 31263
rect 34425 31223 34483 31229
rect 34701 31263 34759 31269
rect 34701 31229 34713 31263
rect 34747 31260 34759 31263
rect 35158 31260 35164 31272
rect 34747 31232 35164 31260
rect 34747 31229 34759 31232
rect 34701 31223 34759 31229
rect 26878 31124 26884 31136
rect 26252 31096 26884 31124
rect 26878 31084 26884 31096
rect 26936 31124 26942 31136
rect 27522 31124 27528 31136
rect 26936 31096 27528 31124
rect 26936 31084 26942 31096
rect 27522 31084 27528 31096
rect 27580 31124 27586 31136
rect 29270 31124 29276 31136
rect 27580 31096 29276 31124
rect 27580 31084 27586 31096
rect 29270 31084 29276 31096
rect 29328 31084 29334 31136
rect 32858 31084 32864 31136
rect 32916 31124 32922 31136
rect 32953 31127 33011 31133
rect 32953 31124 32965 31127
rect 32916 31096 32965 31124
rect 32916 31084 32922 31096
rect 32953 31093 32965 31096
rect 32999 31093 33011 31127
rect 34440 31124 34468 31223
rect 35158 31220 35164 31232
rect 35216 31220 35222 31272
rect 38470 31220 38476 31272
rect 38528 31260 38534 31272
rect 38764 31269 38792 31300
rect 40773 31297 40785 31331
rect 40819 31297 40831 31331
rect 40773 31291 40831 31297
rect 42150 31288 42156 31340
rect 42208 31328 42214 31340
rect 42208 31300 43208 31328
rect 42208 31288 42214 31300
rect 43180 31269 43208 31300
rect 44266 31288 44272 31340
rect 44324 31328 44330 31340
rect 45557 31331 45615 31337
rect 45557 31328 45569 31331
rect 44324 31300 45569 31328
rect 44324 31288 44330 31300
rect 45557 31297 45569 31300
rect 45603 31297 45615 31331
rect 45557 31291 45615 31297
rect 48314 31288 48320 31340
rect 48372 31328 48378 31340
rect 48777 31331 48835 31337
rect 48777 31328 48789 31331
rect 48372 31300 48789 31328
rect 48372 31288 48378 31300
rect 48777 31297 48789 31300
rect 48823 31297 48835 31331
rect 48777 31291 48835 31297
rect 38657 31263 38715 31269
rect 38657 31260 38669 31263
rect 38528 31232 38669 31260
rect 38528 31220 38534 31232
rect 38657 31229 38669 31232
rect 38703 31229 38715 31263
rect 38657 31223 38715 31229
rect 38749 31263 38807 31269
rect 38749 31229 38761 31263
rect 38795 31229 38807 31263
rect 43165 31263 43223 31269
rect 38749 31223 38807 31229
rect 39684 31232 42932 31260
rect 37553 31195 37611 31201
rect 37553 31161 37565 31195
rect 37599 31192 37611 31195
rect 39684 31192 39712 31232
rect 37599 31164 39712 31192
rect 40589 31195 40647 31201
rect 37599 31161 37611 31164
rect 37553 31155 37611 31161
rect 40589 31161 40601 31195
rect 40635 31192 40647 31195
rect 42904 31192 42932 31232
rect 43165 31229 43177 31263
rect 43211 31229 43223 31263
rect 43165 31223 43223 31229
rect 48498 31220 48504 31272
rect 48556 31220 48562 31272
rect 44358 31192 44364 31204
rect 40635 31164 42840 31192
rect 42904 31164 44364 31192
rect 40635 31161 40647 31164
rect 40589 31155 40647 31161
rect 35894 31124 35900 31136
rect 34440 31096 35900 31124
rect 32953 31087 33011 31093
rect 35894 31084 35900 31096
rect 35952 31084 35958 31136
rect 38197 31127 38255 31133
rect 38197 31093 38209 31127
rect 38243 31124 38255 31127
rect 40402 31124 40408 31136
rect 38243 31096 40408 31124
rect 38243 31093 38255 31096
rect 38197 31087 38255 31093
rect 40402 31084 40408 31096
rect 40460 31084 40466 31136
rect 40494 31084 40500 31136
rect 40552 31124 40558 31136
rect 42613 31127 42671 31133
rect 42613 31124 42625 31127
rect 40552 31096 42625 31124
rect 40552 31084 40558 31096
rect 42613 31093 42625 31096
rect 42659 31093 42671 31127
rect 42812 31124 42840 31164
rect 44358 31152 44364 31164
rect 44416 31152 44422 31204
rect 45554 31192 45560 31204
rect 44468 31164 45560 31192
rect 44468 31124 44496 31164
rect 45554 31152 45560 31164
rect 45612 31152 45618 31204
rect 42812 31096 44496 31124
rect 45373 31127 45431 31133
rect 42613 31087 42671 31093
rect 45373 31093 45385 31127
rect 45419 31124 45431 31127
rect 47854 31124 47860 31136
rect 45419 31096 47860 31124
rect 45419 31093 45431 31096
rect 45373 31087 45431 31093
rect 47854 31084 47860 31096
rect 47912 31084 47918 31136
rect 1104 31034 49864 31056
rect 1104 30982 2950 31034
rect 3002 30982 3014 31034
rect 3066 30982 3078 31034
rect 3130 30982 3142 31034
rect 3194 30982 3206 31034
rect 3258 30982 12950 31034
rect 13002 30982 13014 31034
rect 13066 30982 13078 31034
rect 13130 30982 13142 31034
rect 13194 30982 13206 31034
rect 13258 30982 22950 31034
rect 23002 30982 23014 31034
rect 23066 30982 23078 31034
rect 23130 30982 23142 31034
rect 23194 30982 23206 31034
rect 23258 30982 32950 31034
rect 33002 30982 33014 31034
rect 33066 30982 33078 31034
rect 33130 30982 33142 31034
rect 33194 30982 33206 31034
rect 33258 30982 42950 31034
rect 43002 30982 43014 31034
rect 43066 30982 43078 31034
rect 43130 30982 43142 31034
rect 43194 30982 43206 31034
rect 43258 30982 49864 31034
rect 1104 30960 49864 30982
rect 21450 30880 21456 30932
rect 21508 30880 21514 30932
rect 23201 30923 23259 30929
rect 23201 30889 23213 30923
rect 23247 30920 23259 30923
rect 23382 30920 23388 30932
rect 23247 30892 23388 30920
rect 23247 30889 23259 30892
rect 23201 30883 23259 30889
rect 23382 30880 23388 30892
rect 23440 30880 23446 30932
rect 27522 30880 27528 30932
rect 27580 30920 27586 30932
rect 29733 30923 29791 30929
rect 29733 30920 29745 30923
rect 27580 30892 29745 30920
rect 27580 30880 27586 30892
rect 29733 30889 29745 30892
rect 29779 30889 29791 30923
rect 29733 30883 29791 30889
rect 30190 30880 30196 30932
rect 30248 30920 30254 30932
rect 30248 30892 35388 30920
rect 30248 30880 30254 30892
rect 26605 30855 26663 30861
rect 26605 30821 26617 30855
rect 26651 30852 26663 30855
rect 28902 30852 28908 30864
rect 26651 30824 27200 30852
rect 26651 30821 26663 30824
rect 26605 30815 26663 30821
rect 22094 30744 22100 30796
rect 22152 30744 22158 30796
rect 23842 30744 23848 30796
rect 23900 30784 23906 30796
rect 26620 30784 26648 30815
rect 23900 30756 26648 30784
rect 23900 30744 23906 30756
rect 27062 30744 27068 30796
rect 27120 30744 27126 30796
rect 27172 30784 27200 30824
rect 28368 30824 28908 30852
rect 28368 30784 28396 30824
rect 28902 30812 28908 30824
rect 28960 30812 28966 30864
rect 32582 30812 32588 30864
rect 32640 30852 32646 30864
rect 33045 30855 33103 30861
rect 33045 30852 33057 30855
rect 32640 30824 33057 30852
rect 32640 30812 32646 30824
rect 33045 30821 33057 30824
rect 33091 30852 33103 30855
rect 34882 30852 34888 30864
rect 33091 30824 34888 30852
rect 33091 30821 33103 30824
rect 33045 30815 33103 30821
rect 34882 30812 34888 30824
rect 34940 30812 34946 30864
rect 29270 30784 29276 30796
rect 27172 30756 28396 30784
rect 28644 30756 29276 30784
rect 21818 30676 21824 30728
rect 21876 30676 21882 30728
rect 23382 30676 23388 30728
rect 23440 30716 23446 30728
rect 23440 30688 23796 30716
rect 23440 30676 23446 30688
rect 9122 30608 9128 30660
rect 9180 30648 9186 30660
rect 20901 30651 20959 30657
rect 20901 30648 20913 30651
rect 9180 30620 20913 30648
rect 9180 30608 9186 30620
rect 20901 30617 20913 30620
rect 20947 30648 20959 30651
rect 21910 30648 21916 30660
rect 20947 30620 21916 30648
rect 20947 30617 20959 30620
rect 20901 30611 20959 30617
rect 21910 30608 21916 30620
rect 21968 30608 21974 30660
rect 23290 30608 23296 30660
rect 23348 30648 23354 30660
rect 23661 30651 23719 30657
rect 23661 30648 23673 30651
rect 23348 30620 23673 30648
rect 23348 30608 23354 30620
rect 23661 30617 23673 30620
rect 23707 30617 23719 30651
rect 23768 30648 23796 30688
rect 24854 30676 24860 30728
rect 24912 30676 24918 30728
rect 28644 30716 28672 30756
rect 29270 30744 29276 30756
rect 29328 30744 29334 30796
rect 30285 30787 30343 30793
rect 30285 30753 30297 30787
rect 30331 30753 30343 30787
rect 31938 30784 31944 30796
rect 30285 30747 30343 30753
rect 31312 30756 31944 30784
rect 30300 30716 30328 30747
rect 28474 30688 28672 30716
rect 28736 30688 30328 30716
rect 25133 30651 25191 30657
rect 25133 30648 25145 30651
rect 23768 30620 25145 30648
rect 23661 30611 23719 30617
rect 25133 30617 25145 30620
rect 25179 30617 25191 30651
rect 26878 30648 26884 30660
rect 26358 30620 26884 30648
rect 25133 30611 25191 30617
rect 23566 30540 23572 30592
rect 23624 30540 23630 30592
rect 25148 30580 25176 30611
rect 26878 30608 26884 30620
rect 26936 30608 26942 30660
rect 27338 30608 27344 30660
rect 27396 30608 27402 30660
rect 27246 30580 27252 30592
rect 25148 30552 27252 30580
rect 27246 30540 27252 30552
rect 27304 30540 27310 30592
rect 27430 30540 27436 30592
rect 27488 30580 27494 30592
rect 28736 30580 28764 30688
rect 30558 30676 30564 30728
rect 30616 30716 30622 30728
rect 31312 30725 31340 30756
rect 31938 30744 31944 30756
rect 31996 30784 32002 30796
rect 32306 30784 32312 30796
rect 31996 30756 32312 30784
rect 31996 30744 32002 30756
rect 32306 30744 32312 30756
rect 32364 30744 32370 30796
rect 31297 30719 31355 30725
rect 31297 30716 31309 30719
rect 30616 30688 31309 30716
rect 30616 30676 30622 30688
rect 31297 30685 31309 30688
rect 31343 30685 31355 30719
rect 33318 30716 33324 30728
rect 32706 30688 33324 30716
rect 31297 30679 31355 30685
rect 33318 30676 33324 30688
rect 33376 30676 33382 30728
rect 35360 30725 35388 30892
rect 35434 30880 35440 30932
rect 35492 30920 35498 30932
rect 36173 30923 36231 30929
rect 36173 30920 36185 30923
rect 35492 30892 36185 30920
rect 35492 30880 35498 30892
rect 36173 30889 36185 30892
rect 36219 30889 36231 30923
rect 36173 30883 36231 30889
rect 37369 30923 37427 30929
rect 37369 30889 37381 30923
rect 37415 30920 37427 30923
rect 37458 30920 37464 30932
rect 37415 30892 37464 30920
rect 37415 30889 37427 30892
rect 37369 30883 37427 30889
rect 37458 30880 37464 30892
rect 37516 30880 37522 30932
rect 37550 30880 37556 30932
rect 37608 30920 37614 30932
rect 38470 30920 38476 30932
rect 37608 30892 38476 30920
rect 37608 30880 37614 30892
rect 38470 30880 38476 30892
rect 38528 30880 38534 30932
rect 39666 30880 39672 30932
rect 39724 30920 39730 30932
rect 40494 30920 40500 30932
rect 39724 30892 40500 30920
rect 39724 30880 39730 30892
rect 40494 30880 40500 30892
rect 40552 30880 40558 30932
rect 37568 30852 37596 30880
rect 40218 30852 40224 30864
rect 35452 30824 37596 30852
rect 37844 30824 40224 30852
rect 35345 30719 35403 30725
rect 35345 30685 35357 30719
rect 35391 30685 35403 30719
rect 35345 30679 35403 30685
rect 30101 30651 30159 30657
rect 30101 30617 30113 30651
rect 30147 30648 30159 30651
rect 30147 30620 30972 30648
rect 30147 30617 30159 30620
rect 30101 30611 30159 30617
rect 27488 30552 28764 30580
rect 27488 30540 27494 30552
rect 28810 30540 28816 30592
rect 28868 30540 28874 30592
rect 30190 30540 30196 30592
rect 30248 30540 30254 30592
rect 30944 30580 30972 30620
rect 31570 30608 31576 30660
rect 31628 30608 31634 30660
rect 35452 30648 35480 30824
rect 35621 30787 35679 30793
rect 35621 30753 35633 30787
rect 35667 30753 35679 30787
rect 35621 30747 35679 30753
rect 35636 30716 35664 30747
rect 35710 30744 35716 30796
rect 35768 30784 35774 30796
rect 37844 30793 37872 30824
rect 40218 30812 40224 30824
rect 40276 30812 40282 30864
rect 40310 30812 40316 30864
rect 40368 30852 40374 30864
rect 40368 30824 40632 30852
rect 40368 30812 40374 30824
rect 36725 30787 36783 30793
rect 36725 30784 36737 30787
rect 35768 30756 36737 30784
rect 35768 30744 35774 30756
rect 36725 30753 36737 30756
rect 36771 30753 36783 30787
rect 36725 30747 36783 30753
rect 37829 30787 37887 30793
rect 37829 30753 37841 30787
rect 37875 30753 37887 30787
rect 37829 30747 37887 30753
rect 37918 30744 37924 30796
rect 37976 30744 37982 30796
rect 38654 30744 38660 30796
rect 38712 30784 38718 30796
rect 39209 30787 39267 30793
rect 39209 30784 39221 30787
rect 38712 30756 39221 30784
rect 38712 30744 38718 30756
rect 39209 30753 39221 30756
rect 39255 30753 39267 30787
rect 39209 30747 39267 30753
rect 40034 30744 40040 30796
rect 40092 30784 40098 30796
rect 40604 30793 40632 30824
rect 40497 30787 40555 30793
rect 40497 30784 40509 30787
rect 40092 30756 40509 30784
rect 40092 30744 40098 30756
rect 40497 30753 40509 30756
rect 40543 30753 40555 30787
rect 40497 30747 40555 30753
rect 40589 30787 40647 30793
rect 40589 30753 40601 30787
rect 40635 30753 40647 30787
rect 48590 30784 48596 30796
rect 40589 30747 40647 30753
rect 41386 30756 48596 30784
rect 37550 30716 37556 30728
rect 35636 30688 37556 30716
rect 37550 30676 37556 30688
rect 37608 30676 37614 30728
rect 39117 30719 39175 30725
rect 39117 30685 39129 30719
rect 39163 30716 39175 30719
rect 39482 30716 39488 30728
rect 39163 30688 39488 30716
rect 39163 30685 39175 30688
rect 39117 30679 39175 30685
rect 39482 30676 39488 30688
rect 39540 30676 39546 30728
rect 40402 30676 40408 30728
rect 40460 30676 40466 30728
rect 41386 30716 41414 30756
rect 48590 30744 48596 30756
rect 48648 30744 48654 30796
rect 40512 30688 41414 30716
rect 32876 30620 35480 30648
rect 36633 30651 36691 30657
rect 32876 30580 32904 30620
rect 36633 30617 36645 30651
rect 36679 30648 36691 30651
rect 39025 30651 39083 30657
rect 39025 30648 39037 30651
rect 36679 30620 39037 30648
rect 36679 30617 36691 30620
rect 36633 30611 36691 30617
rect 39025 30617 39037 30620
rect 39071 30648 39083 30651
rect 40512 30648 40540 30688
rect 41506 30676 41512 30728
rect 41564 30676 41570 30728
rect 41598 30676 41604 30728
rect 41656 30716 41662 30728
rect 42153 30719 42211 30725
rect 42153 30716 42165 30719
rect 41656 30688 42165 30716
rect 41656 30676 41662 30688
rect 42153 30685 42165 30688
rect 42199 30685 42211 30719
rect 42153 30679 42211 30685
rect 43165 30719 43223 30725
rect 43165 30685 43177 30719
rect 43211 30716 43223 30719
rect 43346 30716 43352 30728
rect 43211 30688 43352 30716
rect 43211 30685 43223 30688
rect 43165 30679 43223 30685
rect 43346 30676 43352 30688
rect 43404 30676 43410 30728
rect 46014 30648 46020 30660
rect 39071 30620 40540 30648
rect 41340 30620 46020 30648
rect 39071 30617 39083 30620
rect 39025 30611 39083 30617
rect 30944 30552 32904 30580
rect 34974 30540 34980 30592
rect 35032 30540 35038 30592
rect 35437 30583 35495 30589
rect 35437 30549 35449 30583
rect 35483 30580 35495 30583
rect 35526 30580 35532 30592
rect 35483 30552 35532 30580
rect 35483 30549 35495 30552
rect 35437 30543 35495 30549
rect 35526 30540 35532 30552
rect 35584 30540 35590 30592
rect 36538 30540 36544 30592
rect 36596 30540 36602 30592
rect 37734 30540 37740 30592
rect 37792 30540 37798 30592
rect 38657 30583 38715 30589
rect 38657 30549 38669 30583
rect 38703 30580 38715 30583
rect 38746 30580 38752 30592
rect 38703 30552 38752 30580
rect 38703 30549 38715 30552
rect 38657 30543 38715 30549
rect 38746 30540 38752 30552
rect 38804 30540 38810 30592
rect 40037 30583 40095 30589
rect 40037 30549 40049 30583
rect 40083 30580 40095 30583
rect 41230 30580 41236 30592
rect 40083 30552 41236 30580
rect 40083 30549 40095 30552
rect 40037 30543 40095 30549
rect 41230 30540 41236 30552
rect 41288 30540 41294 30592
rect 41340 30589 41368 30620
rect 46014 30608 46020 30620
rect 46072 30608 46078 30660
rect 41325 30583 41383 30589
rect 41325 30549 41337 30583
rect 41371 30549 41383 30583
rect 41325 30543 41383 30549
rect 41969 30583 42027 30589
rect 41969 30549 41981 30583
rect 42015 30580 42027 30583
rect 42794 30580 42800 30592
rect 42015 30552 42800 30580
rect 42015 30549 42027 30552
rect 41969 30543 42027 30549
rect 42794 30540 42800 30552
rect 42852 30540 42858 30592
rect 42981 30583 43039 30589
rect 42981 30549 42993 30583
rect 43027 30580 43039 30583
rect 45462 30580 45468 30592
rect 43027 30552 45468 30580
rect 43027 30549 43039 30552
rect 42981 30543 43039 30549
rect 45462 30540 45468 30552
rect 45520 30540 45526 30592
rect 1104 30490 49864 30512
rect 1104 30438 7950 30490
rect 8002 30438 8014 30490
rect 8066 30438 8078 30490
rect 8130 30438 8142 30490
rect 8194 30438 8206 30490
rect 8258 30438 17950 30490
rect 18002 30438 18014 30490
rect 18066 30438 18078 30490
rect 18130 30438 18142 30490
rect 18194 30438 18206 30490
rect 18258 30438 27950 30490
rect 28002 30438 28014 30490
rect 28066 30438 28078 30490
rect 28130 30438 28142 30490
rect 28194 30438 28206 30490
rect 28258 30438 37950 30490
rect 38002 30438 38014 30490
rect 38066 30438 38078 30490
rect 38130 30438 38142 30490
rect 38194 30438 38206 30490
rect 38258 30438 47950 30490
rect 48002 30438 48014 30490
rect 48066 30438 48078 30490
rect 48130 30438 48142 30490
rect 48194 30438 48206 30490
rect 48258 30438 49864 30490
rect 1104 30416 49864 30438
rect 20254 30336 20260 30388
rect 20312 30376 20318 30388
rect 23845 30379 23903 30385
rect 23845 30376 23857 30379
rect 20312 30348 23857 30376
rect 20312 30336 20318 30348
rect 23845 30345 23857 30348
rect 23891 30376 23903 30379
rect 24857 30379 24915 30385
rect 24857 30376 24869 30379
rect 23891 30348 24869 30376
rect 23891 30345 23903 30348
rect 23845 30339 23903 30345
rect 24857 30345 24869 30348
rect 24903 30376 24915 30379
rect 27614 30376 27620 30388
rect 24903 30348 27620 30376
rect 24903 30345 24915 30348
rect 24857 30339 24915 30345
rect 27614 30336 27620 30348
rect 27672 30336 27678 30388
rect 28258 30336 28264 30388
rect 28316 30376 28322 30388
rect 28721 30379 28779 30385
rect 28721 30376 28733 30379
rect 28316 30348 28733 30376
rect 28316 30336 28322 30348
rect 28721 30345 28733 30348
rect 28767 30345 28779 30379
rect 28721 30339 28779 30345
rect 30282 30336 30288 30388
rect 30340 30376 30346 30388
rect 31570 30376 31576 30388
rect 30340 30348 31576 30376
rect 30340 30336 30346 30348
rect 31570 30336 31576 30348
rect 31628 30376 31634 30388
rect 34238 30376 34244 30388
rect 31628 30348 34244 30376
rect 31628 30336 31634 30348
rect 34238 30336 34244 30348
rect 34296 30336 34302 30388
rect 34422 30336 34428 30388
rect 34480 30376 34486 30388
rect 38930 30376 38936 30388
rect 34480 30348 38936 30376
rect 34480 30336 34486 30348
rect 38930 30336 38936 30348
rect 38988 30336 38994 30388
rect 10686 30268 10692 30320
rect 10744 30308 10750 30320
rect 24765 30311 24823 30317
rect 24765 30308 24777 30311
rect 10744 30280 24777 30308
rect 10744 30268 10750 30280
rect 24765 30277 24777 30280
rect 24811 30308 24823 30311
rect 25590 30308 25596 30320
rect 24811 30280 25596 30308
rect 24811 30277 24823 30280
rect 24765 30271 24823 30277
rect 25590 30268 25596 30280
rect 25648 30268 25654 30320
rect 27062 30268 27068 30320
rect 27120 30308 27126 30320
rect 30558 30308 30564 30320
rect 27120 30280 30564 30308
rect 27120 30268 27126 30280
rect 30558 30268 30564 30280
rect 30616 30268 30622 30320
rect 30650 30268 30656 30320
rect 30708 30308 30714 30320
rect 30745 30311 30803 30317
rect 30745 30308 30757 30311
rect 30708 30280 30757 30308
rect 30708 30268 30714 30280
rect 30745 30277 30757 30280
rect 30791 30277 30803 30311
rect 30745 30271 30803 30277
rect 33410 30268 33416 30320
rect 33468 30308 33474 30320
rect 34149 30311 34207 30317
rect 34149 30308 34161 30311
rect 33468 30280 34161 30308
rect 33468 30268 33474 30280
rect 34149 30277 34161 30280
rect 34195 30308 34207 30311
rect 34330 30308 34336 30320
rect 34195 30280 34336 30308
rect 34195 30277 34207 30280
rect 34149 30271 34207 30277
rect 34330 30268 34336 30280
rect 34388 30268 34394 30320
rect 35802 30268 35808 30320
rect 35860 30308 35866 30320
rect 35897 30311 35955 30317
rect 35897 30308 35909 30311
rect 35860 30280 35909 30308
rect 35860 30268 35866 30280
rect 35897 30277 35909 30280
rect 35943 30277 35955 30311
rect 35897 30271 35955 30277
rect 35989 30311 36047 30317
rect 35989 30277 36001 30311
rect 36035 30308 36047 30311
rect 36262 30308 36268 30320
rect 36035 30280 36268 30308
rect 36035 30277 36047 30280
rect 35989 30271 36047 30277
rect 36262 30268 36268 30280
rect 36320 30268 36326 30320
rect 37826 30268 37832 30320
rect 37884 30268 37890 30320
rect 37918 30268 37924 30320
rect 37976 30268 37982 30320
rect 39022 30308 39028 30320
rect 38672 30280 39028 30308
rect 7374 30200 7380 30252
rect 7432 30200 7438 30252
rect 23566 30200 23572 30252
rect 23624 30240 23630 30252
rect 24213 30243 24271 30249
rect 24213 30240 24225 30243
rect 23624 30212 24225 30240
rect 23624 30200 23630 30212
rect 24213 30209 24225 30212
rect 24259 30209 24271 30243
rect 24213 30203 24271 30209
rect 28994 30200 29000 30252
rect 29052 30240 29058 30252
rect 30006 30240 30012 30252
rect 29052 30212 30012 30240
rect 29052 30200 29058 30212
rect 30006 30200 30012 30212
rect 30064 30200 30070 30252
rect 34057 30243 34115 30249
rect 34057 30240 34069 30243
rect 30760 30212 34069 30240
rect 7561 30175 7619 30181
rect 7561 30141 7573 30175
rect 7607 30172 7619 30175
rect 7650 30172 7656 30184
rect 7607 30144 7656 30172
rect 7607 30141 7619 30144
rect 7561 30135 7619 30141
rect 7650 30132 7656 30144
rect 7708 30132 7714 30184
rect 9122 30132 9128 30184
rect 9180 30132 9186 30184
rect 25038 30132 25044 30184
rect 25096 30132 25102 30184
rect 25866 30132 25872 30184
rect 25924 30172 25930 30184
rect 28813 30175 28871 30181
rect 25924 30144 28488 30172
rect 25924 30132 25930 30144
rect 24397 30107 24455 30113
rect 24397 30073 24409 30107
rect 24443 30104 24455 30107
rect 24578 30104 24584 30116
rect 24443 30076 24584 30104
rect 24443 30073 24455 30076
rect 24397 30067 24455 30073
rect 24578 30064 24584 30076
rect 24636 30064 24642 30116
rect 27801 30107 27859 30113
rect 27801 30104 27813 30107
rect 25516 30076 27813 30104
rect 18690 29996 18696 30048
rect 18748 30036 18754 30048
rect 25516 30036 25544 30076
rect 27801 30073 27813 30076
rect 27847 30104 27859 30107
rect 28258 30104 28264 30116
rect 27847 30076 28264 30104
rect 27847 30073 27859 30076
rect 27801 30067 27859 30073
rect 28258 30064 28264 30076
rect 28316 30064 28322 30116
rect 18748 30008 25544 30036
rect 18748 29996 18754 30008
rect 25774 29996 25780 30048
rect 25832 30036 25838 30048
rect 28353 30039 28411 30045
rect 28353 30036 28365 30039
rect 25832 30008 28365 30036
rect 25832 29996 25838 30008
rect 28353 30005 28365 30008
rect 28399 30005 28411 30039
rect 28460 30036 28488 30144
rect 28813 30141 28825 30175
rect 28859 30141 28871 30175
rect 28813 30135 28871 30141
rect 28828 30104 28856 30135
rect 28902 30132 28908 30184
rect 28960 30132 28966 30184
rect 29822 30132 29828 30184
rect 29880 30172 29886 30184
rect 30760 30172 30788 30212
rect 34057 30209 34069 30212
rect 34103 30209 34115 30243
rect 34698 30240 34704 30252
rect 34057 30203 34115 30209
rect 34256 30212 34704 30240
rect 29880 30144 30788 30172
rect 30837 30175 30895 30181
rect 29880 30132 29886 30144
rect 30837 30141 30849 30175
rect 30883 30141 30895 30175
rect 30837 30135 30895 30141
rect 30742 30104 30748 30116
rect 28828 30076 30748 30104
rect 30742 30064 30748 30076
rect 30800 30064 30806 30116
rect 30377 30039 30435 30045
rect 30377 30036 30389 30039
rect 28460 30008 30389 30036
rect 28353 29999 28411 30005
rect 30377 30005 30389 30008
rect 30423 30005 30435 30039
rect 30852 30036 30880 30135
rect 31018 30132 31024 30184
rect 31076 30132 31082 30184
rect 34256 30172 34284 30212
rect 34698 30200 34704 30212
rect 34756 30200 34762 30252
rect 33612 30144 34284 30172
rect 34333 30175 34391 30181
rect 30926 30064 30932 30116
rect 30984 30104 30990 30116
rect 32766 30104 32772 30116
rect 30984 30076 32772 30104
rect 30984 30064 30990 30076
rect 32766 30064 32772 30076
rect 32824 30064 32830 30116
rect 33612 30036 33640 30144
rect 34333 30141 34345 30175
rect 34379 30172 34391 30175
rect 35986 30172 35992 30184
rect 34379 30144 35992 30172
rect 34379 30141 34391 30144
rect 34333 30135 34391 30141
rect 35986 30132 35992 30144
rect 36044 30132 36050 30184
rect 36078 30132 36084 30184
rect 36136 30132 36142 30184
rect 38010 30132 38016 30184
rect 38068 30132 38074 30184
rect 38672 30181 38700 30280
rect 39022 30268 39028 30280
rect 39080 30268 39086 30320
rect 39574 30268 39580 30320
rect 39632 30268 39638 30320
rect 41138 30268 41144 30320
rect 41196 30308 41202 30320
rect 41325 30311 41383 30317
rect 41325 30308 41337 30311
rect 41196 30280 41337 30308
rect 41196 30268 41202 30280
rect 41325 30277 41337 30280
rect 41371 30277 41383 30311
rect 41325 30271 41383 30277
rect 40218 30200 40224 30252
rect 40276 30240 40282 30252
rect 41233 30243 41291 30249
rect 41233 30240 41245 30243
rect 40276 30212 41245 30240
rect 40276 30200 40282 30212
rect 41233 30209 41245 30212
rect 41279 30209 41291 30243
rect 41233 30203 41291 30209
rect 41340 30212 41460 30240
rect 38657 30175 38715 30181
rect 38657 30141 38669 30175
rect 38703 30141 38715 30175
rect 38933 30175 38991 30181
rect 38933 30172 38945 30175
rect 38657 30135 38715 30141
rect 38764 30144 38945 30172
rect 33689 30107 33747 30113
rect 33689 30073 33701 30107
rect 33735 30104 33747 30107
rect 33735 30076 35848 30104
rect 33735 30073 33747 30076
rect 33689 30067 33747 30073
rect 30852 30008 33640 30036
rect 30377 29999 30435 30005
rect 34514 29996 34520 30048
rect 34572 30036 34578 30048
rect 35529 30039 35587 30045
rect 35529 30036 35541 30039
rect 34572 30008 35541 30036
rect 34572 29996 34578 30008
rect 35529 30005 35541 30008
rect 35575 30005 35587 30039
rect 35820 30036 35848 30076
rect 35894 30064 35900 30116
rect 35952 30104 35958 30116
rect 38378 30104 38384 30116
rect 35952 30076 38384 30104
rect 35952 30064 35958 30076
rect 38378 30064 38384 30076
rect 38436 30104 38442 30116
rect 38672 30104 38700 30135
rect 38436 30076 38700 30104
rect 38436 30064 38442 30076
rect 37366 30036 37372 30048
rect 35820 30008 37372 30036
rect 35529 29999 35587 30005
rect 37366 29996 37372 30008
rect 37424 29996 37430 30048
rect 37458 29996 37464 30048
rect 37516 29996 37522 30048
rect 38562 29996 38568 30048
rect 38620 30036 38626 30048
rect 38764 30036 38792 30144
rect 38933 30141 38945 30144
rect 38979 30141 38991 30175
rect 38933 30135 38991 30141
rect 39022 30132 39028 30184
rect 39080 30172 39086 30184
rect 41340 30172 41368 30212
rect 41432 30181 41460 30212
rect 49326 30200 49332 30252
rect 49384 30200 49390 30252
rect 39080 30144 41368 30172
rect 41417 30175 41475 30181
rect 39080 30132 39086 30144
rect 41417 30141 41429 30175
rect 41463 30141 41475 30175
rect 41417 30135 41475 30141
rect 39942 30064 39948 30116
rect 40000 30104 40006 30116
rect 40865 30107 40923 30113
rect 40865 30104 40877 30107
rect 40000 30076 40877 30104
rect 40000 30064 40006 30076
rect 40865 30073 40877 30076
rect 40911 30073 40923 30107
rect 40865 30067 40923 30073
rect 43530 30064 43536 30116
rect 43588 30104 43594 30116
rect 49145 30107 49203 30113
rect 49145 30104 49157 30107
rect 43588 30076 49157 30104
rect 43588 30064 43594 30076
rect 49145 30073 49157 30076
rect 49191 30073 49203 30107
rect 49145 30067 49203 30073
rect 38620 30008 38792 30036
rect 38620 29996 38626 30008
rect 40310 29996 40316 30048
rect 40368 30036 40374 30048
rect 40405 30039 40463 30045
rect 40405 30036 40417 30039
rect 40368 30008 40417 30036
rect 40368 29996 40374 30008
rect 40405 30005 40417 30008
rect 40451 30005 40463 30039
rect 40405 29999 40463 30005
rect 1104 29946 49864 29968
rect 1104 29894 2950 29946
rect 3002 29894 3014 29946
rect 3066 29894 3078 29946
rect 3130 29894 3142 29946
rect 3194 29894 3206 29946
rect 3258 29894 12950 29946
rect 13002 29894 13014 29946
rect 13066 29894 13078 29946
rect 13130 29894 13142 29946
rect 13194 29894 13206 29946
rect 13258 29894 22950 29946
rect 23002 29894 23014 29946
rect 23066 29894 23078 29946
rect 23130 29894 23142 29946
rect 23194 29894 23206 29946
rect 23258 29894 32950 29946
rect 33002 29894 33014 29946
rect 33066 29894 33078 29946
rect 33130 29894 33142 29946
rect 33194 29894 33206 29946
rect 33258 29894 42950 29946
rect 43002 29894 43014 29946
rect 43066 29894 43078 29946
rect 43130 29894 43142 29946
rect 43194 29894 43206 29946
rect 43258 29894 49864 29946
rect 1104 29872 49864 29894
rect 25038 29792 25044 29844
rect 25096 29832 25102 29844
rect 29546 29832 29552 29844
rect 25096 29804 29552 29832
rect 25096 29792 25102 29804
rect 29546 29792 29552 29804
rect 29604 29792 29610 29844
rect 35342 29832 35348 29844
rect 29656 29804 35348 29832
rect 22646 29724 22652 29776
rect 22704 29764 22710 29776
rect 22704 29736 25820 29764
rect 22704 29724 22710 29736
rect 1302 29656 1308 29708
rect 1360 29696 1366 29708
rect 2041 29699 2099 29705
rect 2041 29696 2053 29699
rect 1360 29668 2053 29696
rect 1360 29656 1366 29668
rect 2041 29665 2053 29668
rect 2087 29665 2099 29699
rect 2041 29659 2099 29665
rect 22554 29656 22560 29708
rect 22612 29696 22618 29708
rect 25792 29705 25820 29736
rect 25866 29724 25872 29776
rect 25924 29764 25930 29776
rect 25924 29736 27568 29764
rect 25924 29724 25930 29736
rect 23201 29699 23259 29705
rect 23201 29696 23213 29699
rect 22612 29668 23213 29696
rect 22612 29656 22618 29668
rect 23201 29665 23213 29668
rect 23247 29665 23259 29699
rect 23201 29659 23259 29665
rect 25777 29699 25835 29705
rect 25777 29665 25789 29699
rect 25823 29665 25835 29699
rect 25777 29659 25835 29665
rect 25961 29699 26019 29705
rect 25961 29665 25973 29699
rect 26007 29696 26019 29699
rect 27338 29696 27344 29708
rect 26007 29668 27344 29696
rect 26007 29665 26019 29668
rect 25961 29659 26019 29665
rect 27338 29656 27344 29668
rect 27396 29656 27402 29708
rect 1765 29631 1823 29637
rect 1765 29597 1777 29631
rect 1811 29628 1823 29631
rect 4890 29628 4896 29640
rect 1811 29600 4896 29628
rect 1811 29597 1823 29600
rect 1765 29591 1823 29597
rect 4890 29588 4896 29600
rect 4948 29588 4954 29640
rect 25685 29631 25743 29637
rect 25685 29597 25697 29631
rect 25731 29628 25743 29631
rect 26697 29631 26755 29637
rect 26697 29628 26709 29631
rect 25731 29600 26709 29628
rect 25731 29597 25743 29600
rect 25685 29591 25743 29597
rect 26697 29597 26709 29600
rect 26743 29597 26755 29631
rect 27540 29628 27568 29736
rect 27614 29656 27620 29708
rect 27672 29696 27678 29708
rect 28902 29696 28908 29708
rect 27672 29668 28908 29696
rect 27672 29656 27678 29668
rect 28902 29656 28908 29668
rect 28960 29696 28966 29708
rect 29656 29696 29684 29804
rect 35342 29792 35348 29804
rect 35400 29792 35406 29844
rect 38010 29832 38016 29844
rect 35452 29804 38016 29832
rect 29733 29767 29791 29773
rect 29733 29733 29745 29767
rect 29779 29733 29791 29767
rect 29733 29727 29791 29733
rect 28960 29668 29684 29696
rect 29748 29696 29776 29727
rect 30006 29724 30012 29776
rect 30064 29764 30070 29776
rect 30064 29736 30328 29764
rect 30064 29724 30070 29736
rect 29748 29668 29960 29696
rect 28960 29656 28966 29668
rect 29822 29628 29828 29640
rect 27540 29600 29828 29628
rect 26697 29591 26755 29597
rect 29822 29588 29828 29600
rect 29880 29588 29886 29640
rect 29932 29628 29960 29668
rect 30098 29656 30104 29708
rect 30156 29696 30162 29708
rect 30300 29705 30328 29736
rect 31938 29724 31944 29776
rect 31996 29764 32002 29776
rect 32674 29764 32680 29776
rect 31996 29736 32680 29764
rect 31996 29724 32002 29736
rect 32674 29724 32680 29736
rect 32732 29724 32738 29776
rect 34054 29724 34060 29776
rect 34112 29764 34118 29776
rect 35452 29764 35480 29804
rect 38010 29792 38016 29804
rect 38068 29792 38074 29844
rect 38286 29792 38292 29844
rect 38344 29832 38350 29844
rect 39022 29832 39028 29844
rect 38344 29804 39028 29832
rect 38344 29792 38350 29804
rect 39022 29792 39028 29804
rect 39080 29792 39086 29844
rect 39114 29792 39120 29844
rect 39172 29832 39178 29844
rect 39172 29804 42288 29832
rect 39172 29792 39178 29804
rect 34112 29736 35480 29764
rect 35820 29736 36492 29764
rect 34112 29724 34118 29736
rect 30193 29699 30251 29705
rect 30193 29696 30205 29699
rect 30156 29668 30205 29696
rect 30156 29656 30162 29668
rect 30193 29665 30205 29668
rect 30239 29665 30251 29699
rect 30193 29659 30251 29665
rect 30285 29699 30343 29705
rect 30285 29665 30297 29699
rect 30331 29665 30343 29699
rect 32493 29699 32551 29705
rect 32493 29696 32505 29699
rect 30285 29659 30343 29665
rect 31726 29668 32505 29696
rect 30006 29628 30012 29640
rect 29932 29600 30012 29628
rect 30006 29588 30012 29600
rect 30064 29588 30070 29640
rect 31726 29628 31754 29668
rect 32493 29665 32505 29668
rect 32539 29665 32551 29699
rect 32493 29659 32551 29665
rect 30208 29600 31754 29628
rect 32309 29631 32367 29637
rect 30208 29572 30236 29600
rect 32309 29597 32321 29631
rect 32355 29628 32367 29631
rect 35820 29628 35848 29736
rect 35894 29656 35900 29708
rect 35952 29696 35958 29708
rect 36357 29699 36415 29705
rect 36357 29696 36369 29699
rect 35952 29668 36369 29696
rect 35952 29656 35958 29668
rect 36357 29665 36369 29668
rect 36403 29665 36415 29699
rect 36464 29696 36492 29736
rect 37642 29696 37648 29708
rect 36464 29668 37648 29696
rect 36357 29659 36415 29665
rect 37642 29656 37648 29668
rect 37700 29656 37706 29708
rect 40310 29656 40316 29708
rect 40368 29696 40374 29708
rect 41233 29699 41291 29705
rect 41233 29696 41245 29699
rect 40368 29668 41245 29696
rect 40368 29656 40374 29668
rect 41233 29665 41245 29668
rect 41279 29665 41291 29699
rect 42260 29696 42288 29804
rect 42702 29792 42708 29844
rect 42760 29792 42766 29844
rect 48777 29699 48835 29705
rect 48777 29696 48789 29699
rect 42260 29668 48789 29696
rect 41233 29659 41291 29665
rect 48777 29665 48789 29668
rect 48823 29665 48835 29699
rect 48777 29659 48835 29665
rect 32355 29600 35848 29628
rect 32355 29597 32367 29600
rect 32309 29591 32367 29597
rect 40034 29588 40040 29640
rect 40092 29628 40098 29640
rect 40957 29631 41015 29637
rect 40957 29628 40969 29631
rect 40092 29600 40969 29628
rect 40092 29588 40098 29600
rect 40957 29597 40969 29600
rect 41003 29597 41015 29631
rect 40957 29591 41015 29597
rect 48498 29588 48504 29640
rect 48556 29588 48562 29640
rect 22462 29520 22468 29572
rect 22520 29520 22526 29572
rect 30101 29563 30159 29569
rect 30101 29560 30113 29563
rect 25332 29532 30113 29560
rect 25332 29501 25360 29532
rect 30101 29529 30113 29532
rect 30147 29529 30159 29563
rect 30101 29523 30159 29529
rect 30190 29520 30196 29572
rect 30248 29520 30254 29572
rect 32214 29520 32220 29572
rect 32272 29560 32278 29572
rect 32674 29560 32680 29572
rect 32272 29532 32680 29560
rect 32272 29520 32278 29532
rect 32674 29520 32680 29532
rect 32732 29520 32738 29572
rect 33686 29520 33692 29572
rect 33744 29560 33750 29572
rect 36630 29560 36636 29572
rect 33744 29532 36636 29560
rect 33744 29520 33750 29532
rect 36630 29520 36636 29532
rect 36688 29520 36694 29572
rect 37090 29520 37096 29572
rect 37148 29520 37154 29572
rect 42610 29560 42616 29572
rect 42458 29532 42616 29560
rect 42610 29520 42616 29532
rect 42668 29520 42674 29572
rect 25317 29495 25375 29501
rect 25317 29461 25329 29495
rect 25363 29461 25375 29495
rect 25317 29455 25375 29461
rect 29362 29452 29368 29504
rect 29420 29492 29426 29504
rect 31294 29492 31300 29504
rect 29420 29464 31300 29492
rect 29420 29452 29426 29464
rect 31294 29452 31300 29464
rect 31352 29452 31358 29504
rect 31754 29452 31760 29504
rect 31812 29492 31818 29504
rect 31941 29495 31999 29501
rect 31941 29492 31953 29495
rect 31812 29464 31953 29492
rect 31812 29452 31818 29464
rect 31941 29461 31953 29464
rect 31987 29461 31999 29495
rect 31941 29455 31999 29461
rect 32398 29452 32404 29504
rect 32456 29492 32462 29504
rect 35894 29492 35900 29504
rect 32456 29464 35900 29492
rect 32456 29452 32462 29464
rect 35894 29452 35900 29464
rect 35952 29452 35958 29504
rect 36262 29452 36268 29504
rect 36320 29492 36326 29504
rect 38105 29495 38163 29501
rect 38105 29492 38117 29495
rect 36320 29464 38117 29492
rect 36320 29452 36326 29464
rect 38105 29461 38117 29464
rect 38151 29461 38163 29495
rect 38105 29455 38163 29461
rect 1104 29402 49864 29424
rect 1104 29350 7950 29402
rect 8002 29350 8014 29402
rect 8066 29350 8078 29402
rect 8130 29350 8142 29402
rect 8194 29350 8206 29402
rect 8258 29350 17950 29402
rect 18002 29350 18014 29402
rect 18066 29350 18078 29402
rect 18130 29350 18142 29402
rect 18194 29350 18206 29402
rect 18258 29350 27950 29402
rect 28002 29350 28014 29402
rect 28066 29350 28078 29402
rect 28130 29350 28142 29402
rect 28194 29350 28206 29402
rect 28258 29350 37950 29402
rect 38002 29350 38014 29402
rect 38066 29350 38078 29402
rect 38130 29350 38142 29402
rect 38194 29350 38206 29402
rect 38258 29350 47950 29402
rect 48002 29350 48014 29402
rect 48066 29350 48078 29402
rect 48130 29350 48142 29402
rect 48194 29350 48206 29402
rect 48258 29350 49864 29402
rect 1104 29328 49864 29350
rect 17310 29248 17316 29300
rect 17368 29288 17374 29300
rect 21177 29291 21235 29297
rect 21177 29288 21189 29291
rect 17368 29260 21189 29288
rect 17368 29248 17374 29260
rect 21177 29257 21189 29260
rect 21223 29257 21235 29291
rect 21177 29251 21235 29257
rect 22005 29291 22063 29297
rect 22005 29257 22017 29291
rect 22051 29288 22063 29291
rect 22830 29288 22836 29300
rect 22051 29260 22836 29288
rect 22051 29257 22063 29260
rect 22005 29251 22063 29257
rect 21192 29220 21220 29251
rect 22830 29248 22836 29260
rect 22888 29248 22894 29300
rect 28810 29288 28816 29300
rect 28000 29260 28816 29288
rect 22094 29220 22100 29232
rect 21192 29192 22100 29220
rect 22094 29180 22100 29192
rect 22152 29220 22158 29232
rect 28000 29229 28028 29260
rect 28810 29248 28816 29260
rect 28868 29248 28874 29300
rect 31202 29288 31208 29300
rect 29656 29260 31208 29288
rect 22465 29223 22523 29229
rect 22152 29192 22416 29220
rect 22152 29180 22158 29192
rect 17402 29112 17408 29164
rect 17460 29152 17466 29164
rect 22388 29161 22416 29192
rect 22465 29189 22477 29223
rect 22511 29189 22523 29223
rect 22465 29183 22523 29189
rect 27985 29223 28043 29229
rect 27985 29189 27997 29223
rect 28031 29189 28043 29223
rect 29270 29220 29276 29232
rect 29210 29192 29276 29220
rect 27985 29183 28043 29189
rect 22373 29155 22431 29161
rect 17460 29124 22094 29152
rect 17460 29112 17466 29124
rect 22066 29084 22094 29124
rect 22373 29121 22385 29155
rect 22419 29121 22431 29155
rect 22373 29115 22431 29121
rect 22480 29152 22508 29183
rect 29270 29180 29276 29192
rect 29328 29180 29334 29232
rect 23293 29155 23351 29161
rect 23293 29152 23305 29155
rect 22480 29124 23305 29152
rect 22480 29084 22508 29124
rect 23293 29121 23305 29124
rect 23339 29152 23351 29155
rect 23339 29124 25268 29152
rect 23339 29121 23351 29124
rect 23293 29115 23351 29121
rect 22066 29056 22508 29084
rect 22649 29087 22707 29093
rect 22649 29053 22661 29087
rect 22695 29084 22707 29087
rect 25130 29084 25136 29096
rect 22695 29056 25136 29084
rect 22695 29053 22707 29056
rect 22649 29047 22707 29053
rect 25130 29044 25136 29056
rect 25188 29044 25194 29096
rect 25240 29084 25268 29124
rect 27062 29112 27068 29164
rect 27120 29152 27126 29164
rect 27709 29155 27767 29161
rect 27709 29152 27721 29155
rect 27120 29124 27721 29152
rect 27120 29112 27126 29124
rect 27709 29121 27721 29124
rect 27755 29121 27767 29155
rect 29656 29152 29684 29260
rect 31202 29248 31208 29260
rect 31260 29248 31266 29300
rect 31294 29248 31300 29300
rect 31352 29288 31358 29300
rect 32398 29288 32404 29300
rect 31352 29260 32404 29288
rect 31352 29248 31358 29260
rect 32398 29248 32404 29260
rect 32456 29248 32462 29300
rect 34606 29248 34612 29300
rect 34664 29248 34670 29300
rect 35158 29248 35164 29300
rect 35216 29288 35222 29300
rect 35713 29291 35771 29297
rect 35713 29288 35725 29291
rect 35216 29260 35725 29288
rect 35216 29248 35222 29260
rect 35713 29257 35725 29260
rect 35759 29257 35771 29291
rect 35713 29251 35771 29257
rect 36722 29248 36728 29300
rect 36780 29288 36786 29300
rect 39301 29291 39359 29297
rect 39301 29288 39313 29291
rect 36780 29260 39313 29288
rect 36780 29248 36786 29260
rect 39301 29257 39313 29260
rect 39347 29257 39359 29291
rect 39301 29251 39359 29257
rect 39666 29248 39672 29300
rect 39724 29248 39730 29300
rect 39758 29248 39764 29300
rect 39816 29248 39822 29300
rect 41230 29248 41236 29300
rect 41288 29248 41294 29300
rect 49145 29291 49203 29297
rect 49145 29288 49157 29291
rect 41386 29260 49157 29288
rect 30006 29180 30012 29232
rect 30064 29220 30070 29232
rect 33778 29220 33784 29232
rect 30064 29192 33784 29220
rect 30064 29180 30070 29192
rect 33778 29180 33784 29192
rect 33836 29180 33842 29232
rect 34624 29220 34652 29248
rect 34624 29192 34730 29220
rect 35986 29180 35992 29232
rect 36044 29220 36050 29232
rect 37182 29220 37188 29232
rect 36044 29192 37188 29220
rect 36044 29180 36050 29192
rect 37182 29180 37188 29192
rect 37240 29180 37246 29232
rect 39206 29180 39212 29232
rect 39264 29220 39270 29232
rect 41386 29220 41414 29260
rect 49145 29257 49157 29260
rect 49191 29257 49203 29291
rect 49145 29251 49203 29257
rect 39264 29192 41414 29220
rect 39264 29180 39270 29192
rect 27709 29115 27767 29121
rect 29196 29124 29684 29152
rect 30285 29155 30343 29161
rect 29196 29084 29224 29124
rect 30285 29121 30297 29155
rect 30331 29152 30343 29155
rect 30331 29124 31754 29152
rect 30331 29121 30343 29124
rect 30285 29115 30343 29121
rect 25240 29056 29224 29084
rect 29454 29044 29460 29096
rect 29512 29044 29518 29096
rect 29822 29044 29828 29096
rect 29880 29084 29886 29096
rect 30377 29087 30435 29093
rect 30377 29084 30389 29087
rect 29880 29056 30389 29084
rect 29880 29044 29886 29056
rect 30377 29053 30389 29056
rect 30423 29053 30435 29087
rect 30377 29047 30435 29053
rect 30469 29087 30527 29093
rect 30469 29053 30481 29087
rect 30515 29053 30527 29087
rect 30469 29047 30527 29053
rect 28994 28976 29000 29028
rect 29052 29016 29058 29028
rect 29917 29019 29975 29025
rect 29917 29016 29929 29019
rect 29052 28988 29929 29016
rect 29052 28976 29058 28988
rect 29917 28985 29929 28988
rect 29963 28985 29975 29019
rect 29917 28979 29975 28985
rect 30006 28976 30012 29028
rect 30064 29016 30070 29028
rect 30484 29016 30512 29047
rect 30064 28988 30512 29016
rect 31726 29016 31754 29124
rect 36630 29112 36636 29164
rect 36688 29152 36694 29164
rect 39666 29152 39672 29164
rect 36688 29124 39672 29152
rect 36688 29112 36694 29124
rect 39666 29112 39672 29124
rect 39724 29152 39730 29164
rect 40770 29152 40776 29164
rect 39724 29124 40776 29152
rect 39724 29112 39730 29124
rect 40770 29112 40776 29124
rect 40828 29112 40834 29164
rect 41138 29112 41144 29164
rect 41196 29112 41202 29164
rect 49326 29112 49332 29164
rect 49384 29112 49390 29164
rect 33962 29044 33968 29096
rect 34020 29044 34026 29096
rect 34606 29044 34612 29096
rect 34664 29084 34670 29096
rect 37090 29084 37096 29096
rect 34664 29056 37096 29084
rect 34664 29044 34670 29056
rect 37090 29044 37096 29056
rect 37148 29084 37154 29096
rect 37826 29084 37832 29096
rect 37148 29056 37832 29084
rect 37148 29044 37154 29056
rect 37826 29044 37832 29056
rect 37884 29044 37890 29096
rect 39850 29044 39856 29096
rect 39908 29044 39914 29096
rect 41417 29087 41475 29093
rect 41417 29053 41429 29087
rect 41463 29084 41475 29087
rect 42702 29084 42708 29096
rect 41463 29056 42708 29084
rect 41463 29053 41475 29056
rect 41417 29047 41475 29053
rect 42702 29044 42708 29056
rect 42760 29044 42766 29096
rect 33410 29016 33416 29028
rect 31726 28988 33416 29016
rect 30064 28976 30070 28988
rect 33410 28976 33416 28988
rect 33468 29016 33474 29028
rect 33686 29016 33692 29028
rect 33468 28988 33692 29016
rect 33468 28976 33474 28988
rect 33686 28976 33692 28988
rect 33744 28976 33750 29028
rect 38378 28976 38384 29028
rect 38436 29016 38442 29028
rect 40034 29016 40040 29028
rect 38436 28988 40040 29016
rect 38436 28976 38442 28988
rect 40034 28976 40040 28988
rect 40092 28976 40098 29028
rect 40773 29019 40831 29025
rect 40773 28985 40785 29019
rect 40819 29016 40831 29019
rect 43990 29016 43996 29028
rect 40819 28988 43996 29016
rect 40819 28985 40831 28988
rect 40773 28979 40831 28985
rect 43990 28976 43996 28988
rect 44048 28976 44054 29028
rect 32306 28908 32312 28960
rect 32364 28948 32370 28960
rect 33962 28948 33968 28960
rect 32364 28920 33968 28948
rect 32364 28908 32370 28920
rect 33962 28908 33968 28920
rect 34020 28908 34026 28960
rect 34228 28951 34286 28957
rect 34228 28917 34240 28951
rect 34274 28948 34286 28951
rect 36262 28948 36268 28960
rect 34274 28920 36268 28948
rect 34274 28917 34286 28920
rect 34228 28911 34286 28917
rect 36262 28908 36268 28920
rect 36320 28908 36326 28960
rect 36354 28908 36360 28960
rect 36412 28908 36418 28960
rect 38654 28908 38660 28960
rect 38712 28908 38718 28960
rect 1104 28858 49864 28880
rect 1104 28806 2950 28858
rect 3002 28806 3014 28858
rect 3066 28806 3078 28858
rect 3130 28806 3142 28858
rect 3194 28806 3206 28858
rect 3258 28806 12950 28858
rect 13002 28806 13014 28858
rect 13066 28806 13078 28858
rect 13130 28806 13142 28858
rect 13194 28806 13206 28858
rect 13258 28806 22950 28858
rect 23002 28806 23014 28858
rect 23066 28806 23078 28858
rect 23130 28806 23142 28858
rect 23194 28806 23206 28858
rect 23258 28806 32950 28858
rect 33002 28806 33014 28858
rect 33066 28806 33078 28858
rect 33130 28806 33142 28858
rect 33194 28806 33206 28858
rect 33258 28806 42950 28858
rect 43002 28806 43014 28858
rect 43066 28806 43078 28858
rect 43130 28806 43142 28858
rect 43194 28806 43206 28858
rect 43258 28806 49864 28858
rect 1104 28784 49864 28806
rect 22925 28747 22983 28753
rect 22925 28713 22937 28747
rect 22971 28744 22983 28747
rect 23290 28744 23296 28756
rect 22971 28716 23296 28744
rect 22971 28713 22983 28716
rect 22925 28707 22983 28713
rect 23290 28704 23296 28716
rect 23348 28704 23354 28756
rect 33318 28704 33324 28756
rect 33376 28744 33382 28756
rect 34606 28744 34612 28756
rect 33376 28716 34612 28744
rect 33376 28704 33382 28716
rect 34606 28704 34612 28716
rect 34664 28704 34670 28756
rect 35618 28704 35624 28756
rect 35676 28744 35682 28756
rect 38562 28744 38568 28756
rect 35676 28716 38568 28744
rect 35676 28704 35682 28716
rect 38562 28704 38568 28716
rect 38620 28704 38626 28756
rect 38657 28747 38715 28753
rect 38657 28713 38669 28747
rect 38703 28744 38715 28747
rect 41138 28744 41144 28756
rect 38703 28716 41144 28744
rect 38703 28713 38715 28716
rect 38657 28707 38715 28713
rect 41138 28704 41144 28716
rect 41196 28704 41202 28756
rect 22186 28636 22192 28688
rect 22244 28676 22250 28688
rect 22244 28648 22600 28676
rect 22244 28636 22250 28648
rect 19518 28608 19524 28620
rect 12406 28580 19524 28608
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 12406 28540 12434 28580
rect 19518 28568 19524 28580
rect 19576 28608 19582 28620
rect 19576 28580 21864 28608
rect 19576 28568 19582 28580
rect 7248 28512 12434 28540
rect 20993 28543 21051 28549
rect 7248 28500 7254 28512
rect 20993 28509 21005 28543
rect 21039 28540 21051 28543
rect 21634 28540 21640 28552
rect 21039 28512 21640 28540
rect 21039 28509 21051 28512
rect 20993 28503 21051 28509
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 21836 28540 21864 28580
rect 22002 28568 22008 28620
rect 22060 28608 22066 28620
rect 22278 28608 22284 28620
rect 22060 28580 22284 28608
rect 22060 28568 22066 28580
rect 22278 28568 22284 28580
rect 22336 28568 22342 28620
rect 22572 28552 22600 28648
rect 23198 28636 23204 28688
rect 23256 28676 23262 28688
rect 27614 28676 27620 28688
rect 23256 28648 27620 28676
rect 23256 28636 23262 28648
rect 27614 28636 27620 28648
rect 27672 28676 27678 28688
rect 28353 28679 28411 28685
rect 28353 28676 28365 28679
rect 27672 28648 28365 28676
rect 27672 28636 27678 28648
rect 28353 28645 28365 28648
rect 28399 28676 28411 28679
rect 30374 28676 30380 28688
rect 28399 28648 30380 28676
rect 28399 28645 28411 28648
rect 28353 28639 28411 28645
rect 30374 28636 30380 28648
rect 30432 28636 30438 28688
rect 31938 28636 31944 28688
rect 31996 28676 32002 28688
rect 32950 28676 32956 28688
rect 31996 28648 32956 28676
rect 31996 28636 32002 28648
rect 32950 28636 32956 28648
rect 33008 28636 33014 28688
rect 34974 28636 34980 28688
rect 35032 28676 35038 28688
rect 35032 28648 40540 28676
rect 35032 28636 35038 28648
rect 23382 28568 23388 28620
rect 23440 28608 23446 28620
rect 23477 28611 23535 28617
rect 23477 28608 23489 28611
rect 23440 28580 23489 28608
rect 23440 28568 23446 28580
rect 23477 28577 23489 28580
rect 23523 28577 23535 28611
rect 23477 28571 23535 28577
rect 29454 28568 29460 28620
rect 29512 28608 29518 28620
rect 31205 28611 31263 28617
rect 31205 28608 31217 28611
rect 29512 28580 31217 28608
rect 29512 28568 29518 28580
rect 31205 28577 31217 28580
rect 31251 28577 31263 28611
rect 31205 28571 31263 28577
rect 32858 28568 32864 28620
rect 32916 28608 32922 28620
rect 34057 28611 34115 28617
rect 34057 28608 34069 28611
rect 32916 28580 34069 28608
rect 32916 28568 32922 28580
rect 34057 28577 34069 28580
rect 34103 28577 34115 28611
rect 34057 28571 34115 28577
rect 34146 28568 34152 28620
rect 34204 28568 34210 28620
rect 35529 28611 35587 28617
rect 35529 28577 35541 28611
rect 35575 28608 35587 28611
rect 35618 28608 35624 28620
rect 35575 28580 35624 28608
rect 35575 28577 35587 28580
rect 35529 28571 35587 28577
rect 35618 28568 35624 28580
rect 35676 28568 35682 28620
rect 36262 28568 36268 28620
rect 36320 28608 36326 28620
rect 36633 28611 36691 28617
rect 36633 28608 36645 28611
rect 36320 28580 36645 28608
rect 36320 28568 36326 28580
rect 36633 28577 36645 28580
rect 36679 28577 36691 28611
rect 36633 28571 36691 28577
rect 37366 28568 37372 28620
rect 37424 28568 37430 28620
rect 37553 28611 37611 28617
rect 37553 28577 37565 28611
rect 37599 28608 37611 28611
rect 38562 28608 38568 28620
rect 37599 28580 38568 28608
rect 37599 28577 37611 28580
rect 37553 28571 37611 28577
rect 38562 28568 38568 28580
rect 38620 28568 38626 28620
rect 39301 28611 39359 28617
rect 39301 28577 39313 28611
rect 39347 28608 39359 28611
rect 40310 28608 40316 28620
rect 39347 28580 40316 28608
rect 39347 28577 39359 28580
rect 39301 28571 39359 28577
rect 40310 28568 40316 28580
rect 40368 28568 40374 28620
rect 40512 28617 40540 28648
rect 40497 28611 40555 28617
rect 40497 28577 40509 28611
rect 40543 28577 40555 28611
rect 40497 28571 40555 28577
rect 40678 28568 40684 28620
rect 40736 28568 40742 28620
rect 22370 28540 22376 28552
rect 21836 28512 22376 28540
rect 22370 28500 22376 28512
rect 22428 28500 22434 28552
rect 22554 28500 22560 28552
rect 22612 28540 22618 28552
rect 22612 28512 23336 28540
rect 22612 28500 22618 28512
rect 21729 28475 21787 28481
rect 21729 28441 21741 28475
rect 21775 28441 21787 28475
rect 21729 28435 21787 28441
rect 21744 28404 21772 28435
rect 21818 28432 21824 28484
rect 21876 28472 21882 28484
rect 22462 28472 22468 28484
rect 21876 28444 22468 28472
rect 21876 28432 21882 28444
rect 22462 28432 22468 28444
rect 22520 28472 22526 28484
rect 23198 28472 23204 28484
rect 22520 28444 23204 28472
rect 22520 28432 22526 28444
rect 23198 28432 23204 28444
rect 23256 28432 23262 28484
rect 23308 28472 23336 28512
rect 29914 28500 29920 28552
rect 29972 28500 29978 28552
rect 31021 28543 31079 28549
rect 31021 28509 31033 28543
rect 31067 28540 31079 28543
rect 33594 28540 33600 28552
rect 31067 28512 33600 28540
rect 31067 28509 31079 28512
rect 31021 28503 31079 28509
rect 33594 28500 33600 28512
rect 33652 28500 33658 28552
rect 33965 28543 34023 28549
rect 33965 28509 33977 28543
rect 34011 28540 34023 28543
rect 34790 28540 34796 28552
rect 34011 28512 34796 28540
rect 34011 28509 34023 28512
rect 33965 28503 34023 28509
rect 34790 28500 34796 28512
rect 34848 28500 34854 28552
rect 36354 28500 36360 28552
rect 36412 28540 36418 28552
rect 36449 28543 36507 28549
rect 36449 28540 36461 28543
rect 36412 28512 36461 28540
rect 36412 28500 36418 28512
rect 36449 28509 36461 28512
rect 36495 28509 36507 28543
rect 36449 28503 36507 28509
rect 38654 28500 38660 28552
rect 38712 28540 38718 28552
rect 39025 28543 39083 28549
rect 39025 28540 39037 28543
rect 38712 28512 39037 28540
rect 38712 28500 38718 28512
rect 39025 28509 39037 28512
rect 39071 28509 39083 28543
rect 39025 28503 39083 28509
rect 40405 28543 40463 28549
rect 40405 28509 40417 28543
rect 40451 28540 40463 28543
rect 40954 28540 40960 28552
rect 40451 28512 40960 28540
rect 40451 28509 40463 28512
rect 40405 28503 40463 28509
rect 40954 28500 40960 28512
rect 41012 28500 41018 28552
rect 49326 28500 49332 28552
rect 49384 28500 49390 28552
rect 23308 28444 23428 28472
rect 22002 28404 22008 28416
rect 21744 28376 22008 28404
rect 22002 28364 22008 28376
rect 22060 28364 22066 28416
rect 22370 28364 22376 28416
rect 22428 28404 22434 28416
rect 23290 28404 23296 28416
rect 22428 28376 23296 28404
rect 22428 28364 22434 28376
rect 23290 28364 23296 28376
rect 23348 28364 23354 28416
rect 23400 28413 23428 28444
rect 27062 28432 27068 28484
rect 27120 28432 27126 28484
rect 29730 28432 29736 28484
rect 29788 28472 29794 28484
rect 29788 28444 31156 28472
rect 29788 28432 29794 28444
rect 23385 28407 23443 28413
rect 23385 28373 23397 28407
rect 23431 28373 23443 28407
rect 23385 28367 23443 28373
rect 30650 28364 30656 28416
rect 30708 28364 30714 28416
rect 31128 28413 31156 28444
rect 32214 28432 32220 28484
rect 32272 28472 32278 28484
rect 38105 28475 38163 28481
rect 38105 28472 38117 28475
rect 32272 28444 38117 28472
rect 32272 28432 32278 28444
rect 38105 28441 38117 28444
rect 38151 28472 38163 28475
rect 39117 28475 39175 28481
rect 39117 28472 39129 28475
rect 38151 28444 39129 28472
rect 38151 28441 38163 28444
rect 38105 28435 38163 28441
rect 39117 28441 39129 28444
rect 39163 28441 39175 28475
rect 40126 28472 40132 28484
rect 39117 28435 39175 28441
rect 39224 28444 40132 28472
rect 31113 28407 31171 28413
rect 31113 28373 31125 28407
rect 31159 28404 31171 28407
rect 31294 28404 31300 28416
rect 31159 28376 31300 28404
rect 31159 28373 31171 28376
rect 31113 28367 31171 28373
rect 31294 28364 31300 28376
rect 31352 28364 31358 28416
rect 32766 28364 32772 28416
rect 32824 28404 32830 28416
rect 33597 28407 33655 28413
rect 33597 28404 33609 28407
rect 32824 28376 33609 28404
rect 32824 28364 32830 28376
rect 33597 28373 33609 28376
rect 33643 28373 33655 28407
rect 33597 28367 33655 28373
rect 34790 28364 34796 28416
rect 34848 28404 34854 28416
rect 34885 28407 34943 28413
rect 34885 28404 34897 28407
rect 34848 28376 34897 28404
rect 34848 28364 34854 28376
rect 34885 28373 34897 28376
rect 34931 28373 34943 28407
rect 34885 28367 34943 28373
rect 34974 28364 34980 28416
rect 35032 28404 35038 28416
rect 35253 28407 35311 28413
rect 35253 28404 35265 28407
rect 35032 28376 35265 28404
rect 35032 28364 35038 28376
rect 35253 28373 35265 28376
rect 35299 28373 35311 28407
rect 35253 28367 35311 28373
rect 35342 28364 35348 28416
rect 35400 28364 35406 28416
rect 35434 28364 35440 28416
rect 35492 28404 35498 28416
rect 36081 28407 36139 28413
rect 36081 28404 36093 28407
rect 35492 28376 36093 28404
rect 35492 28364 35498 28376
rect 36081 28373 36093 28376
rect 36127 28373 36139 28407
rect 36081 28367 36139 28373
rect 36538 28364 36544 28416
rect 36596 28364 36602 28416
rect 36909 28407 36967 28413
rect 36909 28373 36921 28407
rect 36955 28404 36967 28407
rect 37182 28404 37188 28416
rect 36955 28376 37188 28404
rect 36955 28373 36967 28376
rect 36909 28367 36967 28373
rect 37182 28364 37188 28376
rect 37240 28364 37246 28416
rect 37277 28407 37335 28413
rect 37277 28373 37289 28407
rect 37323 28404 37335 28407
rect 39224 28404 39252 28444
rect 40126 28432 40132 28444
rect 40184 28432 40190 28484
rect 37323 28376 39252 28404
rect 40037 28407 40095 28413
rect 37323 28373 37335 28376
rect 37277 28367 37335 28373
rect 40037 28373 40049 28407
rect 40083 28404 40095 28407
rect 40310 28404 40316 28416
rect 40083 28376 40316 28404
rect 40083 28373 40095 28376
rect 40037 28367 40095 28373
rect 40310 28364 40316 28376
rect 40368 28364 40374 28416
rect 49142 28364 49148 28416
rect 49200 28364 49206 28416
rect 1104 28314 49864 28336
rect 1104 28262 7950 28314
rect 8002 28262 8014 28314
rect 8066 28262 8078 28314
rect 8130 28262 8142 28314
rect 8194 28262 8206 28314
rect 8258 28262 17950 28314
rect 18002 28262 18014 28314
rect 18066 28262 18078 28314
rect 18130 28262 18142 28314
rect 18194 28262 18206 28314
rect 18258 28262 27950 28314
rect 28002 28262 28014 28314
rect 28066 28262 28078 28314
rect 28130 28262 28142 28314
rect 28194 28262 28206 28314
rect 28258 28262 37950 28314
rect 38002 28262 38014 28314
rect 38066 28262 38078 28314
rect 38130 28262 38142 28314
rect 38194 28262 38206 28314
rect 38258 28262 47950 28314
rect 48002 28262 48014 28314
rect 48066 28262 48078 28314
rect 48130 28262 48142 28314
rect 48194 28262 48206 28314
rect 48258 28262 49864 28314
rect 1104 28240 49864 28262
rect 4890 28160 4896 28212
rect 4948 28160 4954 28212
rect 23382 28200 23388 28212
rect 22664 28172 23388 28200
rect 22664 28141 22692 28172
rect 23382 28160 23388 28172
rect 23440 28200 23446 28212
rect 26329 28203 26387 28209
rect 26329 28200 26341 28203
rect 23440 28172 26341 28200
rect 23440 28160 23446 28172
rect 26329 28169 26341 28172
rect 26375 28200 26387 28203
rect 27430 28200 27436 28212
rect 26375 28172 27436 28200
rect 26375 28169 26387 28172
rect 26329 28163 26387 28169
rect 27430 28160 27436 28172
rect 27488 28160 27494 28212
rect 29454 28200 29460 28212
rect 28184 28172 29460 28200
rect 22649 28135 22707 28141
rect 22649 28101 22661 28135
rect 22695 28101 22707 28135
rect 22649 28095 22707 28101
rect 24946 28092 24952 28144
rect 25004 28132 25010 28144
rect 25004 28104 25346 28132
rect 25004 28092 25010 28104
rect 27706 28092 27712 28144
rect 27764 28132 27770 28144
rect 28184 28141 28212 28172
rect 29454 28160 29460 28172
rect 29512 28160 29518 28212
rect 31297 28203 31355 28209
rect 31297 28169 31309 28203
rect 31343 28200 31355 28203
rect 32122 28200 32128 28212
rect 31343 28172 32128 28200
rect 31343 28169 31355 28172
rect 31297 28163 31355 28169
rect 32122 28160 32128 28172
rect 32180 28160 32186 28212
rect 32398 28160 32404 28212
rect 32456 28200 32462 28212
rect 34057 28203 34115 28209
rect 34057 28200 34069 28203
rect 32456 28172 34069 28200
rect 32456 28160 32462 28172
rect 34057 28169 34069 28172
rect 34103 28200 34115 28203
rect 34146 28200 34152 28212
rect 34103 28172 34152 28200
rect 34103 28169 34115 28172
rect 34057 28163 34115 28169
rect 34146 28160 34152 28172
rect 34204 28160 34210 28212
rect 35894 28160 35900 28212
rect 35952 28200 35958 28212
rect 36357 28203 36415 28209
rect 36357 28200 36369 28203
rect 35952 28172 36369 28200
rect 35952 28160 35958 28172
rect 36357 28169 36369 28172
rect 36403 28169 36415 28203
rect 36357 28163 36415 28169
rect 36446 28160 36452 28212
rect 36504 28160 36510 28212
rect 36538 28160 36544 28212
rect 36596 28200 36602 28212
rect 39025 28203 39083 28209
rect 39025 28200 39037 28203
rect 36596 28172 39037 28200
rect 36596 28160 36602 28172
rect 39025 28169 39037 28172
rect 39071 28169 39083 28203
rect 39025 28163 39083 28169
rect 39206 28160 39212 28212
rect 39264 28200 39270 28212
rect 39485 28203 39543 28209
rect 39485 28200 39497 28203
rect 39264 28172 39497 28200
rect 39264 28160 39270 28172
rect 39485 28169 39497 28172
rect 39531 28169 39543 28203
rect 39485 28163 39543 28169
rect 28169 28135 28227 28141
rect 28169 28132 28181 28135
rect 27764 28104 28181 28132
rect 27764 28092 27770 28104
rect 28169 28101 28181 28104
rect 28215 28101 28227 28135
rect 28169 28095 28227 28101
rect 35342 28092 35348 28144
rect 35400 28132 35406 28144
rect 35400 28104 38332 28132
rect 35400 28092 35406 28104
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5123 28036 6914 28064
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 6886 27928 6914 28036
rect 7558 28024 7564 28076
rect 7616 28024 7622 28076
rect 22002 28024 22008 28076
rect 22060 28064 22066 28076
rect 22278 28064 22284 28076
rect 22060 28036 22284 28064
rect 22060 28024 22066 28036
rect 22278 28024 22284 28036
rect 22336 28064 22342 28076
rect 22373 28067 22431 28073
rect 22373 28064 22385 28067
rect 22336 28036 22385 28064
rect 22336 28024 22342 28036
rect 22373 28033 22385 28036
rect 22419 28033 22431 28067
rect 22373 28027 22431 28033
rect 23750 28024 23756 28076
rect 23808 28024 23814 28076
rect 29270 28024 29276 28076
rect 29328 28024 29334 28076
rect 29454 28024 29460 28076
rect 29512 28064 29518 28076
rect 31205 28067 31263 28073
rect 31205 28064 31217 28067
rect 29512 28036 31217 28064
rect 29512 28024 29518 28036
rect 31205 28033 31217 28036
rect 31251 28033 31263 28067
rect 31205 28027 31263 28033
rect 32306 28024 32312 28076
rect 32364 28024 32370 28076
rect 34146 28064 34152 28076
rect 33718 28036 34152 28064
rect 34146 28024 34152 28036
rect 34204 28064 34210 28076
rect 34606 28064 34612 28076
rect 34204 28036 34612 28064
rect 34204 28024 34210 28036
rect 34606 28024 34612 28036
rect 34664 28024 34670 28076
rect 37458 28024 37464 28076
rect 37516 28064 37522 28076
rect 37645 28067 37703 28073
rect 37645 28064 37657 28067
rect 37516 28036 37657 28064
rect 37516 28024 37522 28036
rect 37645 28033 37657 28036
rect 37691 28033 37703 28067
rect 38304 28064 38332 28104
rect 38378 28092 38384 28144
rect 38436 28092 38442 28144
rect 39298 28092 39304 28144
rect 39356 28132 39362 28144
rect 39574 28132 39580 28144
rect 39356 28104 39580 28132
rect 39356 28092 39362 28104
rect 39574 28092 39580 28104
rect 39632 28132 39638 28144
rect 49142 28132 49148 28144
rect 39632 28104 49148 28132
rect 39632 28092 39638 28104
rect 49142 28092 49148 28104
rect 49200 28092 49206 28144
rect 38838 28064 38844 28076
rect 38304 28036 38844 28064
rect 37645 28027 37703 28033
rect 38838 28024 38844 28036
rect 38896 28024 38902 28076
rect 39206 28024 39212 28076
rect 39264 28064 39270 28076
rect 39393 28067 39451 28073
rect 39393 28064 39405 28067
rect 39264 28036 39405 28064
rect 39264 28024 39270 28036
rect 39393 28033 39405 28036
rect 39439 28033 39451 28067
rect 39393 28027 39451 28033
rect 47854 28024 47860 28076
rect 47912 28064 47918 28076
rect 48133 28067 48191 28073
rect 48133 28064 48145 28067
rect 47912 28036 48145 28064
rect 47912 28024 47918 28036
rect 48133 28033 48145 28036
rect 48179 28033 48191 28067
rect 48133 28027 48191 28033
rect 7742 27956 7748 28008
rect 7800 27956 7806 28008
rect 9401 27999 9459 28005
rect 9401 27965 9413 27999
rect 9447 27996 9459 27999
rect 9582 27996 9588 28008
rect 9447 27968 9588 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 9582 27956 9588 27968
rect 9640 27956 9646 28008
rect 24581 27999 24639 28005
rect 24581 27965 24593 27999
rect 24627 27965 24639 27999
rect 24581 27959 24639 27965
rect 24857 27999 24915 28005
rect 24857 27965 24869 27999
rect 24903 27996 24915 27999
rect 26602 27996 26608 28008
rect 24903 27968 26608 27996
rect 24903 27965 24915 27968
rect 24857 27959 24915 27965
rect 9674 27928 9680 27940
rect 6886 27900 9680 27928
rect 9674 27888 9680 27900
rect 9732 27888 9738 27940
rect 24121 27863 24179 27869
rect 24121 27829 24133 27863
rect 24167 27860 24179 27863
rect 24394 27860 24400 27872
rect 24167 27832 24400 27860
rect 24167 27829 24179 27832
rect 24121 27823 24179 27829
rect 24394 27820 24400 27832
rect 24452 27820 24458 27872
rect 24596 27860 24624 27959
rect 26602 27956 26608 27968
rect 26660 27956 26666 28008
rect 27798 27956 27804 28008
rect 27856 27996 27862 28008
rect 27893 27999 27951 28005
rect 27893 27996 27905 27999
rect 27856 27968 27905 27996
rect 27856 27956 27862 27968
rect 27893 27965 27905 27968
rect 27939 27965 27951 27999
rect 29288 27996 29316 28024
rect 30098 27996 30104 28008
rect 29288 27968 30104 27996
rect 27893 27959 27951 27965
rect 30098 27956 30104 27968
rect 30156 27956 30162 28008
rect 31481 27999 31539 28005
rect 31481 27965 31493 27999
rect 31527 27965 31539 27999
rect 31481 27959 31539 27965
rect 32585 27999 32643 28005
rect 32585 27965 32597 27999
rect 32631 27996 32643 27999
rect 32950 27996 32956 28008
rect 32631 27968 32956 27996
rect 32631 27965 32643 27968
rect 32585 27959 32643 27965
rect 24854 27860 24860 27872
rect 24596 27832 24860 27860
rect 24854 27820 24860 27832
rect 24912 27820 24918 27872
rect 29178 27820 29184 27872
rect 29236 27860 29242 27872
rect 29641 27863 29699 27869
rect 29641 27860 29653 27863
rect 29236 27832 29653 27860
rect 29236 27820 29242 27832
rect 29641 27829 29653 27832
rect 29687 27829 29699 27863
rect 29641 27823 29699 27829
rect 30834 27820 30840 27872
rect 30892 27820 30898 27872
rect 31496 27860 31524 27959
rect 32950 27956 32956 27968
rect 33008 27996 33014 28008
rect 33318 27996 33324 28008
rect 33008 27968 33324 27996
rect 33008 27956 33014 27968
rect 33318 27956 33324 27968
rect 33376 27956 33382 28008
rect 36633 27999 36691 28005
rect 36633 27965 36645 27999
rect 36679 27996 36691 27999
rect 37274 27996 37280 28008
rect 36679 27968 37280 27996
rect 36679 27965 36691 27968
rect 36633 27959 36691 27965
rect 37274 27956 37280 27968
rect 37332 27996 37338 28008
rect 38286 27996 38292 28008
rect 37332 27968 38292 27996
rect 37332 27956 37338 27968
rect 38286 27956 38292 27968
rect 38344 27956 38350 28008
rect 39666 27956 39672 28008
rect 39724 27956 39730 28008
rect 31570 27888 31576 27940
rect 31628 27928 31634 27940
rect 32214 27928 32220 27940
rect 31628 27900 32220 27928
rect 31628 27888 31634 27900
rect 32214 27888 32220 27900
rect 32272 27888 32278 27940
rect 32582 27860 32588 27872
rect 31496 27832 32588 27860
rect 32582 27820 32588 27832
rect 32640 27820 32646 27872
rect 35989 27863 36047 27869
rect 35989 27829 36001 27863
rect 36035 27860 36047 27863
rect 39390 27860 39396 27872
rect 36035 27832 39396 27860
rect 36035 27829 36047 27832
rect 35989 27823 36047 27829
rect 39390 27820 39396 27832
rect 39448 27820 39454 27872
rect 47854 27820 47860 27872
rect 47912 27860 47918 27872
rect 48225 27863 48283 27869
rect 48225 27860 48237 27863
rect 47912 27832 48237 27860
rect 47912 27820 47918 27832
rect 48225 27829 48237 27832
rect 48271 27829 48283 27863
rect 48225 27823 48283 27829
rect 1104 27770 49864 27792
rect 1104 27718 2950 27770
rect 3002 27718 3014 27770
rect 3066 27718 3078 27770
rect 3130 27718 3142 27770
rect 3194 27718 3206 27770
rect 3258 27718 12950 27770
rect 13002 27718 13014 27770
rect 13066 27718 13078 27770
rect 13130 27718 13142 27770
rect 13194 27718 13206 27770
rect 13258 27718 22950 27770
rect 23002 27718 23014 27770
rect 23066 27718 23078 27770
rect 23130 27718 23142 27770
rect 23194 27718 23206 27770
rect 23258 27718 32950 27770
rect 33002 27718 33014 27770
rect 33066 27718 33078 27770
rect 33130 27718 33142 27770
rect 33194 27718 33206 27770
rect 33258 27718 42950 27770
rect 43002 27718 43014 27770
rect 43066 27718 43078 27770
rect 43130 27718 43142 27770
rect 43194 27718 43206 27770
rect 43258 27718 49864 27770
rect 1104 27696 49864 27718
rect 35084 27628 35572 27656
rect 7650 27548 7656 27600
rect 7708 27588 7714 27600
rect 7791 27591 7849 27597
rect 7791 27588 7803 27591
rect 7708 27560 7803 27588
rect 7708 27548 7714 27560
rect 7791 27557 7803 27560
rect 7837 27557 7849 27591
rect 7791 27551 7849 27557
rect 27709 27591 27767 27597
rect 27709 27557 27721 27591
rect 27755 27588 27767 27591
rect 29454 27588 29460 27600
rect 27755 27560 29460 27588
rect 27755 27557 27767 27560
rect 27709 27551 27767 27557
rect 29454 27548 29460 27560
rect 29512 27548 29518 27600
rect 35084 27588 35112 27628
rect 32232 27560 35112 27588
rect 32232 27532 32260 27560
rect 35158 27548 35164 27600
rect 35216 27588 35222 27600
rect 35544 27588 35572 27628
rect 41340 27628 41552 27656
rect 36078 27588 36084 27600
rect 35216 27560 35480 27588
rect 35544 27560 36084 27588
rect 35216 27548 35222 27560
rect 1302 27480 1308 27532
rect 1360 27520 1366 27532
rect 2041 27523 2099 27529
rect 2041 27520 2053 27523
rect 1360 27492 2053 27520
rect 1360 27480 1366 27492
rect 2041 27489 2053 27492
rect 2087 27489 2099 27523
rect 2041 27483 2099 27489
rect 28353 27523 28411 27529
rect 28353 27489 28365 27523
rect 28399 27520 28411 27523
rect 30282 27520 30288 27532
rect 28399 27492 30288 27520
rect 28399 27489 28411 27492
rect 28353 27483 28411 27489
rect 30282 27480 30288 27492
rect 30340 27480 30346 27532
rect 30745 27523 30803 27529
rect 30745 27489 30757 27523
rect 30791 27489 30803 27523
rect 30745 27483 30803 27489
rect 1765 27455 1823 27461
rect 1765 27421 1777 27455
rect 1811 27452 1823 27455
rect 4890 27452 4896 27464
rect 1811 27424 4896 27452
rect 1811 27421 1823 27424
rect 1765 27415 1823 27421
rect 4890 27412 4896 27424
rect 4948 27412 4954 27464
rect 5442 27412 5448 27464
rect 5500 27452 5506 27464
rect 7688 27455 7746 27461
rect 7688 27452 7700 27455
rect 5500 27424 7700 27452
rect 5500 27412 5506 27424
rect 7688 27421 7700 27424
rect 7734 27421 7746 27455
rect 7688 27415 7746 27421
rect 23106 27412 23112 27464
rect 23164 27452 23170 27464
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 23164 27424 23397 27452
rect 23164 27412 23170 27424
rect 23385 27421 23397 27424
rect 23431 27421 23443 27455
rect 23385 27415 23443 27421
rect 24854 27412 24860 27464
rect 24912 27412 24918 27464
rect 28077 27455 28135 27461
rect 28077 27421 28089 27455
rect 28123 27452 28135 27455
rect 29914 27452 29920 27464
rect 28123 27424 29920 27452
rect 28123 27421 28135 27424
rect 28077 27415 28135 27421
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 30374 27412 30380 27464
rect 30432 27452 30438 27464
rect 30653 27455 30711 27461
rect 30653 27452 30665 27455
rect 30432 27424 30665 27452
rect 30432 27412 30438 27424
rect 30653 27421 30665 27424
rect 30699 27421 30711 27455
rect 30653 27415 30711 27421
rect 25130 27344 25136 27396
rect 25188 27344 25194 27396
rect 26694 27384 26700 27396
rect 25240 27356 25622 27384
rect 26528 27356 26700 27384
rect 23474 27276 23480 27328
rect 23532 27316 23538 27328
rect 23750 27316 23756 27328
rect 23532 27288 23756 27316
rect 23532 27276 23538 27288
rect 23750 27276 23756 27288
rect 23808 27316 23814 27328
rect 24946 27316 24952 27328
rect 23808 27288 24952 27316
rect 23808 27276 23814 27288
rect 24946 27276 24952 27288
rect 25004 27316 25010 27328
rect 25240 27316 25268 27356
rect 25004 27288 25268 27316
rect 25516 27316 25544 27356
rect 26528 27316 26556 27356
rect 26694 27344 26700 27356
rect 26752 27344 26758 27396
rect 28718 27344 28724 27396
rect 28776 27384 28782 27396
rect 30760 27384 30788 27483
rect 32214 27480 32220 27532
rect 32272 27480 32278 27532
rect 35250 27480 35256 27532
rect 35308 27520 35314 27532
rect 35452 27529 35480 27560
rect 36078 27548 36084 27560
rect 36136 27548 36142 27600
rect 38562 27548 38568 27600
rect 38620 27588 38626 27600
rect 38657 27591 38715 27597
rect 38657 27588 38669 27591
rect 38620 27560 38669 27588
rect 38620 27548 38626 27560
rect 38657 27557 38669 27560
rect 38703 27557 38715 27591
rect 38657 27551 38715 27557
rect 39666 27548 39672 27600
rect 39724 27588 39730 27600
rect 39724 27560 40172 27588
rect 39724 27548 39730 27560
rect 35345 27523 35403 27529
rect 35345 27520 35357 27523
rect 35308 27492 35357 27520
rect 35308 27480 35314 27492
rect 35345 27489 35357 27492
rect 35391 27489 35403 27523
rect 35345 27483 35403 27489
rect 35437 27523 35495 27529
rect 35437 27489 35449 27523
rect 35483 27489 35495 27523
rect 35437 27483 35495 27489
rect 40034 27480 40040 27532
rect 40092 27480 40098 27532
rect 40144 27520 40172 27560
rect 41340 27520 41368 27628
rect 41524 27588 41552 27628
rect 41785 27591 41843 27597
rect 41785 27588 41797 27591
rect 41524 27560 41797 27588
rect 41785 27557 41797 27560
rect 41831 27557 41843 27591
rect 41785 27551 41843 27557
rect 40144 27492 41368 27520
rect 31662 27412 31668 27464
rect 31720 27452 31726 27464
rect 32861 27455 32919 27461
rect 32861 27452 32873 27455
rect 31720 27424 32873 27452
rect 31720 27412 31726 27424
rect 32861 27421 32873 27424
rect 32907 27421 32919 27455
rect 32861 27415 32919 27421
rect 33689 27455 33747 27461
rect 33689 27421 33701 27455
rect 33735 27452 33747 27455
rect 33962 27452 33968 27464
rect 33735 27424 33968 27452
rect 33735 27421 33747 27424
rect 33689 27415 33747 27421
rect 33962 27412 33968 27424
rect 34020 27452 34026 27464
rect 36909 27455 36967 27461
rect 36909 27452 36921 27455
rect 34020 27424 36921 27452
rect 34020 27412 34026 27424
rect 36909 27421 36921 27424
rect 36955 27421 36967 27455
rect 36909 27415 36967 27421
rect 43990 27412 43996 27464
rect 44048 27412 44054 27464
rect 46382 27412 46388 27464
rect 46440 27452 46446 27464
rect 47213 27455 47271 27461
rect 47213 27452 47225 27455
rect 46440 27424 47225 27452
rect 46440 27412 46446 27424
rect 47213 27421 47225 27424
rect 47259 27421 47271 27455
rect 47213 27415 47271 27421
rect 48498 27412 48504 27464
rect 48556 27412 48562 27464
rect 48590 27412 48596 27464
rect 48648 27452 48654 27464
rect 48777 27455 48835 27461
rect 48777 27452 48789 27455
rect 48648 27424 48789 27452
rect 48648 27412 48654 27424
rect 48777 27421 48789 27424
rect 48823 27421 48835 27455
rect 48777 27415 48835 27421
rect 28776 27356 30788 27384
rect 28776 27344 28782 27356
rect 30926 27344 30932 27396
rect 30984 27384 30990 27396
rect 32033 27387 32091 27393
rect 32033 27384 32045 27387
rect 30984 27356 32045 27384
rect 30984 27344 30990 27356
rect 32033 27353 32045 27356
rect 32079 27353 32091 27387
rect 32033 27347 32091 27353
rect 32950 27344 32956 27396
rect 33008 27384 33014 27396
rect 35253 27387 35311 27393
rect 33008 27356 35204 27384
rect 33008 27344 33014 27356
rect 25516 27288 26556 27316
rect 25004 27276 25010 27288
rect 26602 27276 26608 27328
rect 26660 27316 26666 27328
rect 27246 27316 27252 27328
rect 26660 27288 27252 27316
rect 26660 27276 26666 27288
rect 27246 27276 27252 27288
rect 27304 27276 27310 27328
rect 28169 27319 28227 27325
rect 28169 27285 28181 27319
rect 28215 27316 28227 27319
rect 28442 27316 28448 27328
rect 28215 27288 28448 27316
rect 28215 27285 28227 27288
rect 28169 27279 28227 27285
rect 28442 27276 28448 27288
rect 28500 27276 28506 27328
rect 30190 27276 30196 27328
rect 30248 27276 30254 27328
rect 30558 27276 30564 27328
rect 30616 27276 30622 27328
rect 31665 27319 31723 27325
rect 31665 27285 31677 27319
rect 31711 27316 31723 27319
rect 31938 27316 31944 27328
rect 31711 27288 31944 27316
rect 31711 27285 31723 27288
rect 31665 27279 31723 27285
rect 31938 27276 31944 27288
rect 31996 27276 32002 27328
rect 32125 27319 32183 27325
rect 32125 27285 32137 27319
rect 32171 27316 32183 27319
rect 34606 27316 34612 27328
rect 32171 27288 34612 27316
rect 32171 27285 32183 27288
rect 32125 27279 32183 27285
rect 34606 27276 34612 27288
rect 34664 27276 34670 27328
rect 34885 27319 34943 27325
rect 34885 27285 34897 27319
rect 34931 27316 34943 27319
rect 35066 27316 35072 27328
rect 34931 27288 35072 27316
rect 34931 27285 34943 27288
rect 34885 27279 34943 27285
rect 35066 27276 35072 27288
rect 35124 27276 35130 27328
rect 35176 27316 35204 27356
rect 35253 27353 35265 27387
rect 35299 27384 35311 27387
rect 35434 27384 35440 27396
rect 35299 27356 35440 27384
rect 35299 27353 35311 27356
rect 35253 27347 35311 27353
rect 35434 27344 35440 27356
rect 35492 27344 35498 27396
rect 37090 27344 37096 27396
rect 37148 27384 37154 27396
rect 37185 27387 37243 27393
rect 37185 27384 37197 27387
rect 37148 27356 37197 27384
rect 37148 27344 37154 27356
rect 37185 27353 37197 27356
rect 37231 27353 37243 27387
rect 37185 27347 37243 27353
rect 37826 27344 37832 27396
rect 37884 27344 37890 27396
rect 40313 27387 40371 27393
rect 40313 27353 40325 27387
rect 40359 27384 40371 27387
rect 40402 27384 40408 27396
rect 40359 27356 40408 27384
rect 40359 27353 40371 27356
rect 40313 27347 40371 27353
rect 40402 27344 40408 27356
rect 40460 27344 40466 27396
rect 41598 27384 41604 27396
rect 41538 27356 41604 27384
rect 41598 27344 41604 27356
rect 41656 27384 41662 27396
rect 42610 27384 42616 27396
rect 41656 27356 42616 27384
rect 41656 27344 41662 27356
rect 42610 27344 42616 27356
rect 42668 27344 42674 27396
rect 47397 27387 47455 27393
rect 47397 27353 47409 27387
rect 47443 27384 47455 27387
rect 47578 27384 47584 27396
rect 47443 27356 47584 27384
rect 47443 27353 47455 27356
rect 47397 27347 47455 27353
rect 47578 27344 47584 27356
rect 47636 27344 47642 27396
rect 40954 27316 40960 27328
rect 35176 27288 40960 27316
rect 40954 27276 40960 27288
rect 41012 27276 41018 27328
rect 41046 27276 41052 27328
rect 41104 27316 41110 27328
rect 43714 27316 43720 27328
rect 41104 27288 43720 27316
rect 41104 27276 41110 27288
rect 43714 27276 43720 27288
rect 43772 27276 43778 27328
rect 43806 27276 43812 27328
rect 43864 27276 43870 27328
rect 1104 27226 49864 27248
rect 1104 27174 7950 27226
rect 8002 27174 8014 27226
rect 8066 27174 8078 27226
rect 8130 27174 8142 27226
rect 8194 27174 8206 27226
rect 8258 27174 17950 27226
rect 18002 27174 18014 27226
rect 18066 27174 18078 27226
rect 18130 27174 18142 27226
rect 18194 27174 18206 27226
rect 18258 27174 27950 27226
rect 28002 27174 28014 27226
rect 28066 27174 28078 27226
rect 28130 27174 28142 27226
rect 28194 27174 28206 27226
rect 28258 27174 37950 27226
rect 38002 27174 38014 27226
rect 38066 27174 38078 27226
rect 38130 27174 38142 27226
rect 38194 27174 38206 27226
rect 38258 27174 47950 27226
rect 48002 27174 48014 27226
rect 48066 27174 48078 27226
rect 48130 27174 48142 27226
rect 48194 27174 48206 27226
rect 48258 27174 49864 27226
rect 1104 27152 49864 27174
rect 23106 27072 23112 27124
rect 23164 27072 23170 27124
rect 23201 27115 23259 27121
rect 23201 27081 23213 27115
rect 23247 27112 23259 27115
rect 23290 27112 23296 27124
rect 23247 27084 23296 27112
rect 23247 27081 23259 27084
rect 23201 27075 23259 27081
rect 23290 27072 23296 27084
rect 23348 27072 23354 27124
rect 30282 27072 30288 27124
rect 30340 27072 30346 27124
rect 30558 27072 30564 27124
rect 30616 27112 30622 27124
rect 31386 27112 31392 27124
rect 30616 27084 31392 27112
rect 30616 27072 30622 27084
rect 31386 27072 31392 27084
rect 31444 27112 31450 27124
rect 32490 27112 32496 27124
rect 31444 27084 32496 27112
rect 31444 27072 31450 27084
rect 32490 27072 32496 27084
rect 32548 27072 32554 27124
rect 32674 27072 32680 27124
rect 32732 27112 32738 27124
rect 32732 27084 35756 27112
rect 32732 27072 32738 27084
rect 24854 27004 24860 27056
rect 24912 27044 24918 27056
rect 27798 27044 27804 27056
rect 24912 27016 27804 27044
rect 24912 27004 24918 27016
rect 27798 27004 27804 27016
rect 27856 27044 27862 27056
rect 27893 27047 27951 27053
rect 27893 27044 27905 27047
rect 27856 27016 27905 27044
rect 27856 27004 27862 27016
rect 27893 27013 27905 27016
rect 27939 27044 27951 27047
rect 30098 27044 30104 27056
rect 27939 27016 28580 27044
rect 30038 27016 30104 27044
rect 27939 27013 27951 27016
rect 27893 27007 27951 27013
rect 7834 26936 7840 26988
rect 7892 26936 7898 26988
rect 24121 26979 24179 26985
rect 24121 26945 24133 26979
rect 24167 26976 24179 26979
rect 25498 26976 25504 26988
rect 24167 26948 25504 26976
rect 24167 26945 24179 26948
rect 24121 26939 24179 26945
rect 25498 26936 25504 26948
rect 25556 26936 25562 26988
rect 27157 26979 27215 26985
rect 27157 26945 27169 26979
rect 27203 26976 27215 26979
rect 27614 26976 27620 26988
rect 27203 26948 27620 26976
rect 27203 26945 27215 26948
rect 27157 26939 27215 26945
rect 27614 26936 27620 26948
rect 27672 26936 27678 26988
rect 28552 26985 28580 27016
rect 30098 27004 30104 27016
rect 30156 27044 30162 27056
rect 30742 27044 30748 27056
rect 30156 27016 30748 27044
rect 30156 27004 30162 27016
rect 30742 27004 30748 27016
rect 30800 27004 30806 27056
rect 31113 27047 31171 27053
rect 31113 27013 31125 27047
rect 31159 27044 31171 27047
rect 31202 27044 31208 27056
rect 31159 27016 31208 27044
rect 31159 27013 31171 27016
rect 31113 27007 31171 27013
rect 31202 27004 31208 27016
rect 31260 27004 31266 27056
rect 31294 27004 31300 27056
rect 31352 27044 31358 27056
rect 33321 27047 33379 27053
rect 33321 27044 33333 27047
rect 31352 27016 33333 27044
rect 31352 27004 31358 27016
rect 33321 27013 33333 27016
rect 33367 27013 33379 27047
rect 33321 27007 33379 27013
rect 34146 27004 34152 27056
rect 34204 27044 34210 27056
rect 34204 27016 34914 27044
rect 34204 27004 34210 27016
rect 28537 26979 28595 26985
rect 28537 26945 28549 26979
rect 28583 26945 28595 26979
rect 31570 26976 31576 26988
rect 28537 26939 28595 26945
rect 31220 26948 31576 26976
rect 8021 26911 8079 26917
rect 8021 26877 8033 26911
rect 8067 26908 8079 26911
rect 8294 26908 8300 26920
rect 8067 26880 8300 26908
rect 8067 26877 8079 26880
rect 8021 26871 8079 26877
rect 8294 26868 8300 26880
rect 8352 26868 8358 26920
rect 8938 26868 8944 26920
rect 8996 26868 9002 26920
rect 23382 26868 23388 26920
rect 23440 26868 23446 26920
rect 28813 26911 28871 26917
rect 28813 26877 28825 26911
rect 28859 26908 28871 26911
rect 29178 26908 29184 26920
rect 28859 26880 29184 26908
rect 28859 26877 28871 26880
rect 28813 26871 28871 26877
rect 29178 26868 29184 26880
rect 29236 26868 29242 26920
rect 30558 26868 30564 26920
rect 30616 26908 30622 26920
rect 31220 26917 31248 26948
rect 31570 26936 31576 26948
rect 31628 26936 31634 26988
rect 33413 26979 33471 26985
rect 33413 26945 33425 26979
rect 33459 26976 33471 26979
rect 33686 26976 33692 26988
rect 33459 26948 33692 26976
rect 33459 26945 33471 26948
rect 33413 26939 33471 26945
rect 33686 26936 33692 26948
rect 33744 26936 33750 26988
rect 35728 26976 35756 27084
rect 35894 27072 35900 27124
rect 35952 27112 35958 27124
rect 37090 27112 37096 27124
rect 35952 27084 37096 27112
rect 35952 27072 35958 27084
rect 37090 27072 37096 27084
rect 37148 27072 37154 27124
rect 40678 27072 40684 27124
rect 40736 27112 40742 27124
rect 42061 27115 42119 27121
rect 42061 27112 42073 27115
rect 40736 27084 42073 27112
rect 40736 27072 40742 27084
rect 42061 27081 42073 27084
rect 42107 27081 42119 27115
rect 42061 27075 42119 27081
rect 37550 27004 37556 27056
rect 37608 27044 37614 27056
rect 40589 27047 40647 27053
rect 40589 27044 40601 27047
rect 37608 27016 40601 27044
rect 37608 27004 37614 27016
rect 36909 26979 36967 26985
rect 36909 26976 36921 26979
rect 35728 26948 36921 26976
rect 36909 26945 36921 26948
rect 36955 26945 36967 26979
rect 36909 26939 36967 26945
rect 37458 26936 37464 26988
rect 37516 26936 37522 26988
rect 31205 26911 31263 26917
rect 31205 26908 31217 26911
rect 30616 26880 31217 26908
rect 30616 26868 30622 26880
rect 31205 26877 31217 26880
rect 31251 26877 31263 26911
rect 31205 26871 31263 26877
rect 31297 26911 31355 26917
rect 31297 26877 31309 26911
rect 31343 26877 31355 26911
rect 31297 26871 31355 26877
rect 33597 26911 33655 26917
rect 33597 26877 33609 26911
rect 33643 26908 33655 26911
rect 34054 26908 34060 26920
rect 33643 26880 34060 26908
rect 33643 26877 33655 26880
rect 33597 26871 33655 26877
rect 31110 26800 31116 26852
rect 31168 26840 31174 26852
rect 31312 26840 31340 26871
rect 34054 26868 34060 26880
rect 34112 26868 34118 26920
rect 34149 26911 34207 26917
rect 34149 26877 34161 26911
rect 34195 26908 34207 26911
rect 34195 26880 34284 26908
rect 34195 26877 34207 26880
rect 34149 26871 34207 26877
rect 31168 26812 31340 26840
rect 31168 26800 31174 26812
rect 22741 26775 22799 26781
rect 22741 26741 22753 26775
rect 22787 26772 22799 26775
rect 24118 26772 24124 26784
rect 22787 26744 24124 26772
rect 22787 26741 22799 26744
rect 22741 26735 22799 26741
rect 24118 26732 24124 26744
rect 24176 26732 24182 26784
rect 24210 26732 24216 26784
rect 24268 26732 24274 26784
rect 26510 26732 26516 26784
rect 26568 26772 26574 26784
rect 27338 26772 27344 26784
rect 26568 26744 27344 26772
rect 26568 26732 26574 26744
rect 27338 26732 27344 26744
rect 27396 26772 27402 26784
rect 30374 26772 30380 26784
rect 27396 26744 30380 26772
rect 27396 26732 27402 26744
rect 30374 26732 30380 26744
rect 30432 26732 30438 26784
rect 30466 26732 30472 26784
rect 30524 26772 30530 26784
rect 30745 26775 30803 26781
rect 30745 26772 30757 26775
rect 30524 26744 30757 26772
rect 30524 26732 30530 26744
rect 30745 26741 30757 26744
rect 30791 26741 30803 26775
rect 30745 26735 30803 26741
rect 32953 26775 33011 26781
rect 32953 26741 32965 26775
rect 32999 26772 33011 26775
rect 33962 26772 33968 26784
rect 32999 26744 33968 26772
rect 32999 26741 33011 26744
rect 32953 26735 33011 26741
rect 33962 26732 33968 26744
rect 34020 26732 34026 26784
rect 34256 26772 34284 26880
rect 34422 26868 34428 26920
rect 34480 26868 34486 26920
rect 38286 26868 38292 26920
rect 38344 26868 38350 26920
rect 39960 26908 39988 27016
rect 40589 27013 40601 27016
rect 40635 27013 40647 27047
rect 40589 27007 40647 27013
rect 41598 27004 41604 27056
rect 41656 27004 41662 27056
rect 44634 27004 44640 27056
rect 44692 27044 44698 27056
rect 47857 27047 47915 27053
rect 47857 27044 47869 27047
rect 44692 27016 47869 27044
rect 44692 27004 44698 27016
rect 47857 27013 47869 27016
rect 47903 27013 47915 27047
rect 47857 27007 47915 27013
rect 40034 26936 40040 26988
rect 40092 26976 40098 26988
rect 40313 26979 40371 26985
rect 40313 26976 40325 26979
rect 40092 26948 40325 26976
rect 40092 26936 40098 26948
rect 40313 26945 40325 26948
rect 40359 26945 40371 26979
rect 40313 26939 40371 26945
rect 45462 26936 45468 26988
rect 45520 26976 45526 26988
rect 47029 26979 47087 26985
rect 47029 26976 47041 26979
rect 45520 26948 47041 26976
rect 45520 26936 45526 26948
rect 47029 26945 47041 26948
rect 47075 26945 47087 26979
rect 47029 26939 47087 26945
rect 41782 26908 41788 26920
rect 39960 26880 41788 26908
rect 41782 26868 41788 26880
rect 41840 26908 41846 26920
rect 42242 26908 42248 26920
rect 41840 26880 42248 26908
rect 41840 26868 41846 26880
rect 42242 26868 42248 26880
rect 42300 26868 42306 26920
rect 48498 26868 48504 26920
rect 48556 26868 48562 26920
rect 48774 26868 48780 26920
rect 48832 26868 48838 26920
rect 36630 26800 36636 26852
rect 36688 26840 36694 26852
rect 36688 26812 40448 26840
rect 36688 26800 36694 26812
rect 34882 26772 34888 26784
rect 34256 26744 34888 26772
rect 34882 26732 34888 26744
rect 34940 26732 34946 26784
rect 36725 26775 36783 26781
rect 36725 26741 36737 26775
rect 36771 26772 36783 26775
rect 38378 26772 38384 26784
rect 36771 26744 38384 26772
rect 36771 26741 36783 26744
rect 36725 26735 36783 26741
rect 38378 26732 38384 26744
rect 38436 26732 38442 26784
rect 40420 26772 40448 26812
rect 41046 26772 41052 26784
rect 40420 26744 41052 26772
rect 41046 26732 41052 26744
rect 41104 26732 41110 26784
rect 46842 26732 46848 26784
rect 46900 26732 46906 26784
rect 47670 26732 47676 26784
rect 47728 26772 47734 26784
rect 47949 26775 48007 26781
rect 47949 26772 47961 26775
rect 47728 26744 47961 26772
rect 47728 26732 47734 26744
rect 47949 26741 47961 26744
rect 47995 26741 48007 26775
rect 47949 26735 48007 26741
rect 1104 26682 49864 26704
rect 1104 26630 2950 26682
rect 3002 26630 3014 26682
rect 3066 26630 3078 26682
rect 3130 26630 3142 26682
rect 3194 26630 3206 26682
rect 3258 26630 12950 26682
rect 13002 26630 13014 26682
rect 13066 26630 13078 26682
rect 13130 26630 13142 26682
rect 13194 26630 13206 26682
rect 13258 26630 22950 26682
rect 23002 26630 23014 26682
rect 23066 26630 23078 26682
rect 23130 26630 23142 26682
rect 23194 26630 23206 26682
rect 23258 26630 32950 26682
rect 33002 26630 33014 26682
rect 33066 26630 33078 26682
rect 33130 26630 33142 26682
rect 33194 26630 33206 26682
rect 33258 26630 42950 26682
rect 43002 26630 43014 26682
rect 43066 26630 43078 26682
rect 43130 26630 43142 26682
rect 43194 26630 43206 26682
rect 43258 26630 49864 26682
rect 1104 26608 49864 26630
rect 7742 26528 7748 26580
rect 7800 26568 7806 26580
rect 7883 26571 7941 26577
rect 7883 26568 7895 26571
rect 7800 26540 7895 26568
rect 7800 26528 7806 26540
rect 7883 26537 7895 26540
rect 7929 26537 7941 26571
rect 7883 26531 7941 26537
rect 9674 26528 9680 26580
rect 9732 26528 9738 26580
rect 22360 26571 22418 26577
rect 22360 26537 22372 26571
rect 22406 26568 22418 26571
rect 24394 26568 24400 26580
rect 22406 26540 24400 26568
rect 22406 26537 22418 26540
rect 22360 26531 22418 26537
rect 24394 26528 24400 26540
rect 24452 26528 24458 26580
rect 25038 26528 25044 26580
rect 25096 26568 25102 26580
rect 25222 26568 25228 26580
rect 25096 26540 25228 26568
rect 25096 26528 25102 26540
rect 25222 26528 25228 26540
rect 25280 26528 25286 26580
rect 29178 26528 29184 26580
rect 29236 26568 29242 26580
rect 29236 26540 31248 26568
rect 29236 26528 29242 26540
rect 23566 26460 23572 26512
rect 23624 26500 23630 26512
rect 23845 26503 23903 26509
rect 23845 26500 23857 26503
rect 23624 26472 23857 26500
rect 23624 26460 23630 26472
rect 23845 26469 23857 26472
rect 23891 26469 23903 26503
rect 23845 26463 23903 26469
rect 23934 26460 23940 26512
rect 23992 26500 23998 26512
rect 24581 26503 24639 26509
rect 24581 26500 24593 26503
rect 23992 26472 24593 26500
rect 23992 26460 23998 26472
rect 24581 26469 24593 26472
rect 24627 26469 24639 26503
rect 31018 26500 31024 26512
rect 24581 26463 24639 26469
rect 24964 26472 31024 26500
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 10870 26432 10876 26444
rect 9171 26404 10876 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 10870 26392 10876 26404
rect 10928 26392 10934 26444
rect 22097 26435 22155 26441
rect 22097 26401 22109 26435
rect 22143 26432 22155 26435
rect 24854 26432 24860 26444
rect 22143 26404 24860 26432
rect 22143 26401 22155 26404
rect 22097 26395 22155 26401
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 7742 26324 7748 26376
rect 7800 26373 7806 26376
rect 7800 26367 7838 26373
rect 7826 26333 7838 26367
rect 7800 26327 7838 26333
rect 9309 26367 9367 26373
rect 9309 26333 9321 26367
rect 9355 26364 9367 26367
rect 10962 26364 10968 26376
rect 9355 26336 10968 26364
rect 9355 26333 9367 26336
rect 9309 26327 9367 26333
rect 7800 26324 7806 26327
rect 4982 26256 4988 26308
rect 5040 26296 5046 26308
rect 5442 26296 5448 26308
rect 5040 26268 5448 26296
rect 5040 26256 5046 26268
rect 5442 26256 5448 26268
rect 5500 26296 5506 26308
rect 9324 26296 9352 26327
rect 10962 26324 10968 26336
rect 11020 26324 11026 26376
rect 23474 26324 23480 26376
rect 23532 26324 23538 26376
rect 24964 26373 24992 26472
rect 31018 26460 31024 26472
rect 31076 26460 31082 26512
rect 25038 26392 25044 26444
rect 25096 26392 25102 26444
rect 25133 26435 25191 26441
rect 25133 26401 25145 26435
rect 25179 26401 25191 26435
rect 25133 26395 25191 26401
rect 24949 26367 25007 26373
rect 24949 26333 24961 26367
rect 24995 26333 25007 26367
rect 24949 26327 25007 26333
rect 5500 26268 9352 26296
rect 5500 26256 5506 26268
rect 23658 26256 23664 26308
rect 23716 26296 23722 26308
rect 25148 26296 25176 26395
rect 26418 26392 26424 26444
rect 26476 26432 26482 26444
rect 26513 26435 26571 26441
rect 26513 26432 26525 26435
rect 26476 26404 26525 26432
rect 26476 26392 26482 26404
rect 26513 26401 26525 26404
rect 26559 26401 26571 26435
rect 26513 26395 26571 26401
rect 26697 26435 26755 26441
rect 26697 26401 26709 26435
rect 26743 26432 26755 26435
rect 27706 26432 27712 26444
rect 26743 26404 27712 26432
rect 26743 26401 26755 26404
rect 26697 26395 26755 26401
rect 27706 26392 27712 26404
rect 27764 26392 27770 26444
rect 28350 26392 28356 26444
rect 28408 26432 28414 26444
rect 28810 26432 28816 26444
rect 28408 26404 28816 26432
rect 28408 26392 28414 26404
rect 28810 26392 28816 26404
rect 28868 26432 28874 26444
rect 30558 26432 30564 26444
rect 28868 26404 30564 26432
rect 28868 26392 28874 26404
rect 30558 26392 30564 26404
rect 30616 26392 30622 26444
rect 30650 26392 30656 26444
rect 30708 26432 30714 26444
rect 31220 26441 31248 26540
rect 32582 26528 32588 26580
rect 32640 26568 32646 26580
rect 33873 26571 33931 26577
rect 33873 26568 33885 26571
rect 32640 26540 33885 26568
rect 32640 26528 32646 26540
rect 33873 26537 33885 26540
rect 33919 26568 33931 26571
rect 34422 26568 34428 26580
rect 33919 26540 34428 26568
rect 33919 26537 33931 26540
rect 33873 26531 33931 26537
rect 34422 26528 34428 26540
rect 34480 26528 34486 26580
rect 37090 26568 37096 26580
rect 34532 26540 37096 26568
rect 33686 26460 33692 26512
rect 33744 26500 33750 26512
rect 34532 26500 34560 26540
rect 37090 26528 37096 26540
rect 37148 26528 37154 26580
rect 37369 26571 37427 26577
rect 37369 26537 37381 26571
rect 37415 26568 37427 26571
rect 40494 26568 40500 26580
rect 37415 26540 40500 26568
rect 37415 26537 37427 26540
rect 37369 26531 37427 26537
rect 40494 26528 40500 26540
rect 40552 26528 40558 26580
rect 40954 26528 40960 26580
rect 41012 26568 41018 26580
rect 48774 26568 48780 26580
rect 41012 26540 48780 26568
rect 41012 26528 41018 26540
rect 48774 26528 48780 26540
rect 48832 26528 48838 26580
rect 33744 26472 34560 26500
rect 33744 26460 33750 26472
rect 34698 26460 34704 26512
rect 34756 26500 34762 26512
rect 48590 26500 48596 26512
rect 34756 26472 40172 26500
rect 34756 26460 34762 26472
rect 31113 26435 31171 26441
rect 31113 26432 31125 26435
rect 30708 26404 31125 26432
rect 30708 26392 30714 26404
rect 31113 26401 31125 26404
rect 31159 26401 31171 26435
rect 31113 26395 31171 26401
rect 31205 26435 31263 26441
rect 31205 26401 31217 26435
rect 31251 26401 31263 26435
rect 31205 26395 31263 26401
rect 31662 26392 31668 26444
rect 31720 26432 31726 26444
rect 37458 26432 37464 26444
rect 31720 26404 37464 26432
rect 31720 26392 31754 26404
rect 27249 26367 27307 26373
rect 27249 26333 27261 26367
rect 27295 26364 27307 26367
rect 27614 26364 27620 26376
rect 27295 26336 27620 26364
rect 27295 26333 27307 26336
rect 27249 26327 27307 26333
rect 27614 26324 27620 26336
rect 27672 26364 27678 26376
rect 28626 26364 28632 26376
rect 27672 26336 28632 26364
rect 27672 26324 27678 26336
rect 28626 26324 28632 26336
rect 28684 26364 28690 26376
rect 31726 26364 31754 26392
rect 34900 26373 34928 26404
rect 37458 26392 37464 26404
rect 37516 26392 37522 26444
rect 37550 26392 37556 26444
rect 37608 26432 37614 26444
rect 37921 26435 37979 26441
rect 37921 26432 37933 26435
rect 37608 26404 37933 26432
rect 37608 26392 37614 26404
rect 37921 26401 37933 26404
rect 37967 26401 37979 26435
rect 37921 26395 37979 26401
rect 40034 26392 40040 26444
rect 40092 26392 40098 26444
rect 40144 26432 40172 26472
rect 41386 26472 48596 26500
rect 41386 26432 41414 26472
rect 48590 26460 48596 26472
rect 48648 26460 48654 26512
rect 40144 26404 41414 26432
rect 41782 26392 41788 26444
rect 41840 26392 41846 26444
rect 43714 26392 43720 26444
rect 43772 26432 43778 26444
rect 48777 26435 48835 26441
rect 48777 26432 48789 26435
rect 43772 26404 48789 26432
rect 43772 26392 43778 26404
rect 48777 26401 48789 26404
rect 48823 26401 48835 26435
rect 48777 26395 48835 26401
rect 28684 26336 31754 26364
rect 32125 26367 32183 26373
rect 28684 26324 28690 26336
rect 32125 26333 32137 26367
rect 32171 26333 32183 26367
rect 32125 26327 32183 26333
rect 34885 26367 34943 26373
rect 34885 26333 34897 26367
rect 34931 26333 34943 26367
rect 34885 26327 34943 26333
rect 37829 26367 37887 26373
rect 37829 26333 37841 26367
rect 37875 26364 37887 26367
rect 39574 26364 39580 26376
rect 37875 26336 39580 26364
rect 37875 26333 37887 26336
rect 37829 26327 37887 26333
rect 28077 26299 28135 26305
rect 23716 26268 25176 26296
rect 26068 26268 28028 26296
rect 23716 26256 23722 26268
rect 25406 26188 25412 26240
rect 25464 26228 25470 26240
rect 25682 26228 25688 26240
rect 25464 26200 25688 26228
rect 25464 26188 25470 26200
rect 25682 26188 25688 26200
rect 25740 26188 25746 26240
rect 26068 26237 26096 26268
rect 26053 26231 26111 26237
rect 26053 26197 26065 26231
rect 26099 26197 26111 26231
rect 26053 26191 26111 26197
rect 26418 26188 26424 26240
rect 26476 26188 26482 26240
rect 28000 26228 28028 26268
rect 28077 26265 28089 26299
rect 28123 26296 28135 26299
rect 28350 26296 28356 26308
rect 28123 26268 28356 26296
rect 28123 26265 28135 26268
rect 28077 26259 28135 26265
rect 28350 26256 28356 26268
rect 28408 26256 28414 26308
rect 31021 26299 31079 26305
rect 31021 26296 31033 26299
rect 28460 26268 31033 26296
rect 28460 26228 28488 26268
rect 31021 26265 31033 26268
rect 31067 26265 31079 26299
rect 32140 26296 32168 26327
rect 39574 26324 39580 26336
rect 39632 26324 39638 26376
rect 43806 26324 43812 26376
rect 43864 26364 43870 26376
rect 47397 26367 47455 26373
rect 47397 26364 47409 26367
rect 43864 26336 47409 26364
rect 43864 26324 43870 26336
rect 47397 26333 47409 26336
rect 47443 26333 47455 26367
rect 47397 26327 47455 26333
rect 48041 26367 48099 26373
rect 48041 26333 48053 26367
rect 48087 26364 48099 26367
rect 48498 26364 48504 26376
rect 48087 26336 48504 26364
rect 48087 26333 48099 26336
rect 48041 26327 48099 26333
rect 48498 26324 48504 26336
rect 48556 26324 48562 26376
rect 32306 26296 32312 26308
rect 32140 26268 32312 26296
rect 31021 26259 31079 26265
rect 32306 26256 32312 26268
rect 32364 26256 32370 26308
rect 32398 26256 32404 26308
rect 32456 26256 32462 26308
rect 34238 26296 34244 26308
rect 33626 26268 34244 26296
rect 34238 26256 34244 26268
rect 34296 26256 34302 26308
rect 35621 26299 35679 26305
rect 35621 26296 35633 26299
rect 34900 26268 35633 26296
rect 34900 26240 34928 26268
rect 35621 26265 35633 26268
rect 35667 26265 35679 26299
rect 35621 26259 35679 26265
rect 39482 26256 39488 26308
rect 39540 26296 39546 26308
rect 40313 26299 40371 26305
rect 40313 26296 40325 26299
rect 39540 26268 40325 26296
rect 39540 26256 39546 26268
rect 40313 26265 40325 26268
rect 40359 26265 40371 26299
rect 41598 26296 41604 26308
rect 41538 26268 41604 26296
rect 40313 26259 40371 26265
rect 41598 26256 41604 26268
rect 41656 26256 41662 26308
rect 28000 26200 28488 26228
rect 30650 26188 30656 26240
rect 30708 26188 30714 26240
rect 34882 26188 34888 26240
rect 34940 26188 34946 26240
rect 37734 26188 37740 26240
rect 37792 26188 37798 26240
rect 47210 26188 47216 26240
rect 47268 26188 47274 26240
rect 1104 26138 49864 26160
rect 1104 26086 7950 26138
rect 8002 26086 8014 26138
rect 8066 26086 8078 26138
rect 8130 26086 8142 26138
rect 8194 26086 8206 26138
rect 8258 26086 17950 26138
rect 18002 26086 18014 26138
rect 18066 26086 18078 26138
rect 18130 26086 18142 26138
rect 18194 26086 18206 26138
rect 18258 26086 27950 26138
rect 28002 26086 28014 26138
rect 28066 26086 28078 26138
rect 28130 26086 28142 26138
rect 28194 26086 28206 26138
rect 28258 26086 37950 26138
rect 38002 26086 38014 26138
rect 38066 26086 38078 26138
rect 38130 26086 38142 26138
rect 38194 26086 38206 26138
rect 38258 26086 47950 26138
rect 48002 26086 48014 26138
rect 48066 26086 48078 26138
rect 48130 26086 48142 26138
rect 48194 26086 48206 26138
rect 48258 26086 49864 26138
rect 1104 26064 49864 26086
rect 24118 25984 24124 26036
rect 24176 26024 24182 26036
rect 27525 26027 27583 26033
rect 27525 26024 27537 26027
rect 24176 25996 27537 26024
rect 24176 25984 24182 25996
rect 27525 25993 27537 25996
rect 27571 25993 27583 26027
rect 27525 25987 27583 25993
rect 27798 25984 27804 26036
rect 27856 26024 27862 26036
rect 28442 26024 28448 26036
rect 27856 25996 28448 26024
rect 27856 25984 27862 25996
rect 28442 25984 28448 25996
rect 28500 25984 28506 26036
rect 29546 25984 29552 26036
rect 29604 26024 29610 26036
rect 31297 26027 31355 26033
rect 31297 26024 31309 26027
rect 29604 25996 31309 26024
rect 29604 25984 29610 25996
rect 31297 25993 31309 25996
rect 31343 25993 31355 26027
rect 31297 25987 31355 25993
rect 31389 26027 31447 26033
rect 31389 25993 31401 26027
rect 31435 26024 31447 26027
rect 32309 26027 32367 26033
rect 32309 26024 32321 26027
rect 31435 25996 32321 26024
rect 31435 25993 31447 25996
rect 31389 25987 31447 25993
rect 32309 25993 32321 25996
rect 32355 25993 32367 26027
rect 32309 25987 32367 25993
rect 32674 25984 32680 26036
rect 32732 26024 32738 26036
rect 37734 26024 37740 26036
rect 32732 25996 37740 26024
rect 32732 25984 32738 25996
rect 37734 25984 37740 25996
rect 37792 25984 37798 26036
rect 39025 26027 39083 26033
rect 39025 26024 39037 26027
rect 37844 25996 39037 26024
rect 24136 25928 24440 25956
rect 7650 25848 7656 25900
rect 7708 25848 7714 25900
rect 24136 25897 24164 25928
rect 24121 25891 24179 25897
rect 24121 25857 24133 25891
rect 24167 25857 24179 25891
rect 24412 25888 24440 25928
rect 25682 25916 25688 25968
rect 25740 25956 25746 25968
rect 27816 25956 27844 25984
rect 30742 25956 30748 25968
rect 25740 25928 27844 25956
rect 29854 25928 30748 25956
rect 25740 25916 25746 25928
rect 30742 25916 30748 25928
rect 30800 25916 30806 25968
rect 32769 25959 32827 25965
rect 32769 25925 32781 25959
rect 32815 25956 32827 25959
rect 32950 25956 32956 25968
rect 32815 25928 32956 25956
rect 32815 25925 32827 25928
rect 32769 25919 32827 25925
rect 32950 25916 32956 25928
rect 33008 25916 33014 25968
rect 33778 25916 33784 25968
rect 33836 25956 33842 25968
rect 33836 25928 36308 25956
rect 33836 25916 33842 25928
rect 25133 25891 25191 25897
rect 25133 25888 25145 25891
rect 24412 25860 25145 25888
rect 24121 25851 24179 25857
rect 25133 25857 25145 25860
rect 25179 25857 25191 25891
rect 25133 25851 25191 25857
rect 26418 25848 26424 25900
rect 26476 25888 26482 25900
rect 26605 25891 26663 25897
rect 26605 25888 26617 25891
rect 26476 25860 26617 25888
rect 26476 25848 26482 25860
rect 26605 25857 26617 25860
rect 26651 25857 26663 25891
rect 26605 25851 26663 25857
rect 27522 25848 27528 25900
rect 27580 25888 27586 25900
rect 27617 25891 27675 25897
rect 27617 25888 27629 25891
rect 27580 25860 27629 25888
rect 27580 25848 27586 25860
rect 27617 25857 27629 25860
rect 27663 25857 27675 25891
rect 27617 25851 27675 25857
rect 34330 25848 34336 25900
rect 34388 25888 34394 25900
rect 36280 25897 36308 25928
rect 37642 25916 37648 25968
rect 37700 25956 37706 25968
rect 37844 25956 37872 25996
rect 39025 25993 39037 25996
rect 39071 25993 39083 26027
rect 39025 25987 39083 25993
rect 39393 26027 39451 26033
rect 39393 25993 39405 26027
rect 39439 26024 39451 26027
rect 39942 26024 39948 26036
rect 39439 25996 39948 26024
rect 39439 25993 39451 25996
rect 39393 25987 39451 25993
rect 39942 25984 39948 25996
rect 40000 25984 40006 26036
rect 40402 25984 40408 26036
rect 40460 26024 40466 26036
rect 40770 26024 40776 26036
rect 40460 25996 40776 26024
rect 40460 25984 40466 25996
rect 40770 25984 40776 25996
rect 40828 26024 40834 26036
rect 42061 26027 42119 26033
rect 42061 26024 42073 26027
rect 40828 25996 42073 26024
rect 40828 25984 40834 25996
rect 42061 25993 42073 25996
rect 42107 25993 42119 26027
rect 42061 25987 42119 25993
rect 37700 25928 37872 25956
rect 37700 25916 37706 25928
rect 38286 25916 38292 25968
rect 38344 25956 38350 25968
rect 40589 25959 40647 25965
rect 38344 25928 40356 25956
rect 38344 25916 38350 25928
rect 35253 25891 35311 25897
rect 35253 25888 35265 25891
rect 34388 25860 35265 25888
rect 34388 25848 34394 25860
rect 35253 25857 35265 25860
rect 35299 25857 35311 25891
rect 35253 25851 35311 25857
rect 36265 25891 36323 25897
rect 36265 25857 36277 25891
rect 36311 25857 36323 25891
rect 36265 25851 36323 25857
rect 37550 25848 37556 25900
rect 37608 25888 37614 25900
rect 38197 25891 38255 25897
rect 38197 25888 38209 25891
rect 37608 25860 38209 25888
rect 37608 25848 37614 25860
rect 38197 25857 38209 25860
rect 38243 25857 38255 25891
rect 38470 25888 38476 25900
rect 38197 25851 38255 25857
rect 38304 25860 38476 25888
rect 7837 25823 7895 25829
rect 7837 25789 7849 25823
rect 7883 25820 7895 25823
rect 9030 25820 9036 25832
rect 7883 25792 9036 25820
rect 7883 25789 7895 25792
rect 7837 25783 7895 25789
rect 9030 25780 9036 25792
rect 9088 25780 9094 25832
rect 9490 25780 9496 25832
rect 9548 25820 9554 25832
rect 9548 25792 12434 25820
rect 9548 25780 9554 25792
rect 12406 25752 12434 25792
rect 22094 25780 22100 25832
rect 22152 25820 22158 25832
rect 22370 25820 22376 25832
rect 22152 25792 22376 25820
rect 22152 25780 22158 25792
rect 22370 25780 22376 25792
rect 22428 25820 22434 25832
rect 24213 25823 24271 25829
rect 24213 25820 24225 25823
rect 22428 25792 24225 25820
rect 22428 25780 22434 25792
rect 24213 25789 24225 25792
rect 24259 25789 24271 25823
rect 24213 25783 24271 25789
rect 24302 25780 24308 25832
rect 24360 25780 24366 25832
rect 24394 25780 24400 25832
rect 24452 25820 24458 25832
rect 27709 25823 27767 25829
rect 27709 25820 27721 25823
rect 24452 25792 27721 25820
rect 24452 25780 24458 25792
rect 27709 25789 27721 25792
rect 27755 25789 27767 25823
rect 27709 25783 27767 25789
rect 28350 25780 28356 25832
rect 28408 25780 28414 25832
rect 28629 25823 28687 25829
rect 28629 25820 28641 25823
rect 28460 25792 28641 25820
rect 23753 25755 23811 25761
rect 12406 25724 23704 25752
rect 22646 25644 22652 25696
rect 22704 25684 22710 25696
rect 22833 25687 22891 25693
rect 22833 25684 22845 25687
rect 22704 25656 22845 25684
rect 22704 25644 22710 25656
rect 22833 25653 22845 25656
rect 22879 25653 22891 25687
rect 23676 25684 23704 25724
rect 23753 25721 23765 25755
rect 23799 25752 23811 25755
rect 28258 25752 28264 25764
rect 23799 25724 28264 25752
rect 23799 25721 23811 25724
rect 23753 25715 23811 25721
rect 28258 25712 28264 25724
rect 28316 25712 28322 25764
rect 25682 25684 25688 25696
rect 23676 25656 25688 25684
rect 22833 25647 22891 25653
rect 25682 25644 25688 25656
rect 25740 25644 25746 25696
rect 25774 25644 25780 25696
rect 25832 25684 25838 25696
rect 25961 25687 26019 25693
rect 25961 25684 25973 25687
rect 25832 25656 25973 25684
rect 25832 25644 25838 25656
rect 25961 25653 25973 25656
rect 26007 25653 26019 25687
rect 25961 25647 26019 25653
rect 27157 25687 27215 25693
rect 27157 25653 27169 25687
rect 27203 25684 27215 25687
rect 27338 25684 27344 25696
rect 27203 25656 27344 25684
rect 27203 25653 27215 25656
rect 27157 25647 27215 25653
rect 27338 25644 27344 25656
rect 27396 25644 27402 25696
rect 27430 25644 27436 25696
rect 27488 25684 27494 25696
rect 28460 25684 28488 25792
rect 28629 25789 28641 25792
rect 28675 25820 28687 25823
rect 30282 25820 30288 25832
rect 28675 25792 30288 25820
rect 28675 25789 28687 25792
rect 28629 25783 28687 25789
rect 30282 25780 30288 25792
rect 30340 25780 30346 25832
rect 31573 25823 31631 25829
rect 31573 25789 31585 25823
rect 31619 25820 31631 25823
rect 32398 25820 32404 25832
rect 31619 25792 32404 25820
rect 31619 25789 31631 25792
rect 31573 25783 31631 25789
rect 32398 25780 32404 25792
rect 32456 25780 32462 25832
rect 32861 25823 32919 25829
rect 32861 25789 32873 25823
rect 32907 25820 32919 25823
rect 33318 25820 33324 25832
rect 32907 25792 33324 25820
rect 32907 25789 32919 25792
rect 32861 25783 32919 25789
rect 29822 25712 29828 25764
rect 29880 25752 29886 25764
rect 32876 25752 32904 25783
rect 33318 25780 33324 25792
rect 33376 25780 33382 25832
rect 34698 25780 34704 25832
rect 34756 25820 34762 25832
rect 35345 25823 35403 25829
rect 35345 25820 35357 25823
rect 34756 25792 35357 25820
rect 34756 25780 34762 25792
rect 35345 25789 35357 25792
rect 35391 25789 35403 25823
rect 35345 25783 35403 25789
rect 35529 25823 35587 25829
rect 35529 25789 35541 25823
rect 35575 25820 35587 25823
rect 35894 25820 35900 25832
rect 35575 25792 35900 25820
rect 35575 25789 35587 25792
rect 35529 25783 35587 25789
rect 35894 25780 35900 25792
rect 35952 25780 35958 25832
rect 38304 25829 38332 25860
rect 38470 25848 38476 25860
rect 38528 25848 38534 25900
rect 39390 25848 39396 25900
rect 39448 25888 39454 25900
rect 40328 25897 40356 25928
rect 40589 25925 40601 25959
rect 40635 25956 40647 25959
rect 40678 25956 40684 25968
rect 40635 25928 40684 25956
rect 40635 25925 40647 25928
rect 40589 25919 40647 25925
rect 40678 25916 40684 25928
rect 40736 25916 40742 25968
rect 41598 25916 41604 25968
rect 41656 25916 41662 25968
rect 42794 25916 42800 25968
rect 42852 25956 42858 25968
rect 46753 25959 46811 25965
rect 46753 25956 46765 25959
rect 42852 25928 46765 25956
rect 42852 25916 42858 25928
rect 46753 25925 46765 25928
rect 46799 25925 46811 25959
rect 46753 25919 46811 25925
rect 39485 25891 39543 25897
rect 39485 25888 39497 25891
rect 39448 25860 39497 25888
rect 39448 25848 39454 25860
rect 39485 25857 39497 25860
rect 39531 25857 39543 25891
rect 39485 25851 39543 25857
rect 40313 25891 40371 25897
rect 40313 25857 40325 25891
rect 40359 25857 40371 25891
rect 40313 25851 40371 25857
rect 38289 25823 38347 25829
rect 38289 25789 38301 25823
rect 38335 25789 38347 25823
rect 38289 25783 38347 25789
rect 38381 25823 38439 25829
rect 38381 25789 38393 25823
rect 38427 25789 38439 25823
rect 38381 25783 38439 25789
rect 29880 25724 32904 25752
rect 36081 25755 36139 25761
rect 29880 25712 29886 25724
rect 36081 25721 36093 25755
rect 36127 25752 36139 25755
rect 37458 25752 37464 25764
rect 36127 25724 37464 25752
rect 36127 25721 36139 25724
rect 36081 25715 36139 25721
rect 37458 25712 37464 25724
rect 37516 25712 37522 25764
rect 37550 25712 37556 25764
rect 37608 25752 37614 25764
rect 38396 25752 38424 25783
rect 39574 25780 39580 25832
rect 39632 25780 39638 25832
rect 39666 25780 39672 25832
rect 39724 25820 39730 25832
rect 41616 25820 41644 25916
rect 46014 25848 46020 25900
rect 46072 25848 46078 25900
rect 49326 25848 49332 25900
rect 49384 25848 49390 25900
rect 39724 25792 41644 25820
rect 39724 25780 39730 25792
rect 37608 25724 38424 25752
rect 37608 25712 37614 25724
rect 46198 25712 46204 25764
rect 46256 25712 46262 25764
rect 46934 25712 46940 25764
rect 46992 25712 46998 25764
rect 27488 25656 28488 25684
rect 27488 25644 27494 25656
rect 29914 25644 29920 25696
rect 29972 25684 29978 25696
rect 30101 25687 30159 25693
rect 30101 25684 30113 25687
rect 29972 25656 30113 25684
rect 29972 25644 29978 25656
rect 30101 25653 30113 25656
rect 30147 25653 30159 25687
rect 30101 25647 30159 25653
rect 30926 25644 30932 25696
rect 30984 25644 30990 25696
rect 34885 25687 34943 25693
rect 34885 25653 34897 25687
rect 34931 25684 34943 25687
rect 35986 25684 35992 25696
rect 34931 25656 35992 25684
rect 34931 25653 34943 25656
rect 34885 25647 34943 25653
rect 35986 25644 35992 25656
rect 36044 25644 36050 25696
rect 36906 25644 36912 25696
rect 36964 25644 36970 25696
rect 37734 25644 37740 25696
rect 37792 25684 37798 25696
rect 37829 25687 37887 25693
rect 37829 25684 37841 25687
rect 37792 25656 37841 25684
rect 37792 25644 37798 25656
rect 37829 25653 37841 25656
rect 37875 25653 37887 25687
rect 37829 25647 37887 25653
rect 49142 25644 49148 25696
rect 49200 25644 49206 25696
rect 1104 25594 49864 25616
rect 1104 25542 2950 25594
rect 3002 25542 3014 25594
rect 3066 25542 3078 25594
rect 3130 25542 3142 25594
rect 3194 25542 3206 25594
rect 3258 25542 12950 25594
rect 13002 25542 13014 25594
rect 13066 25542 13078 25594
rect 13130 25542 13142 25594
rect 13194 25542 13206 25594
rect 13258 25542 22950 25594
rect 23002 25542 23014 25594
rect 23066 25542 23078 25594
rect 23130 25542 23142 25594
rect 23194 25542 23206 25594
rect 23258 25542 32950 25594
rect 33002 25542 33014 25594
rect 33066 25542 33078 25594
rect 33130 25542 33142 25594
rect 33194 25542 33206 25594
rect 33258 25542 42950 25594
rect 43002 25542 43014 25594
rect 43066 25542 43078 25594
rect 43130 25542 43142 25594
rect 43194 25542 43206 25594
rect 43258 25542 49864 25594
rect 1104 25520 49864 25542
rect 4890 25440 4896 25492
rect 4948 25440 4954 25492
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25449 10839 25483
rect 10781 25443 10839 25449
rect 1302 25304 1308 25356
rect 1360 25344 1366 25356
rect 2041 25347 2099 25353
rect 2041 25344 2053 25347
rect 1360 25316 2053 25344
rect 1360 25304 1366 25316
rect 2041 25313 2053 25316
rect 2087 25313 2099 25347
rect 10796 25344 10824 25443
rect 10962 25440 10968 25492
rect 11020 25480 11026 25492
rect 11057 25483 11115 25489
rect 11057 25480 11069 25483
rect 11020 25452 11069 25480
rect 11020 25440 11026 25452
rect 11057 25449 11069 25452
rect 11103 25449 11115 25483
rect 11057 25443 11115 25449
rect 24302 25440 24308 25492
rect 24360 25480 24366 25492
rect 25130 25480 25136 25492
rect 24360 25452 25136 25480
rect 24360 25440 24366 25452
rect 25130 25440 25136 25452
rect 25188 25480 25194 25492
rect 27709 25483 27767 25489
rect 27709 25480 27721 25483
rect 25188 25452 27721 25480
rect 25188 25440 25194 25452
rect 27709 25449 27721 25452
rect 27755 25480 27767 25483
rect 30006 25480 30012 25492
rect 27755 25452 30012 25480
rect 27755 25449 27767 25452
rect 27709 25443 27767 25449
rect 30006 25440 30012 25452
rect 30064 25440 30070 25492
rect 34238 25440 34244 25492
rect 34296 25480 34302 25492
rect 35342 25480 35348 25492
rect 34296 25452 35348 25480
rect 34296 25440 34302 25452
rect 35342 25440 35348 25452
rect 35400 25440 35406 25492
rect 37826 25440 37832 25492
rect 37884 25480 37890 25492
rect 37884 25452 39436 25480
rect 37884 25440 37890 25452
rect 10870 25372 10876 25424
rect 10928 25412 10934 25424
rect 14277 25415 14335 25421
rect 14277 25412 14289 25415
rect 10928 25384 14289 25412
rect 10928 25372 10934 25384
rect 14277 25381 14289 25384
rect 14323 25381 14335 25415
rect 14277 25375 14335 25381
rect 27246 25372 27252 25424
rect 27304 25412 27310 25424
rect 30745 25415 30803 25421
rect 27304 25384 28948 25412
rect 27304 25372 27310 25384
rect 12342 25344 12348 25356
rect 10796 25316 12348 25344
rect 2041 25307 2099 25313
rect 12342 25304 12348 25316
rect 12400 25304 12406 25356
rect 22925 25347 22983 25353
rect 22925 25313 22937 25347
rect 22971 25344 22983 25347
rect 24302 25344 24308 25356
rect 22971 25316 24308 25344
rect 22971 25313 22983 25316
rect 22925 25307 22983 25313
rect 24302 25304 24308 25316
rect 24360 25304 24366 25356
rect 25225 25347 25283 25353
rect 25225 25313 25237 25347
rect 25271 25344 25283 25347
rect 25682 25344 25688 25356
rect 25271 25316 25688 25344
rect 25271 25313 25283 25316
rect 25225 25307 25283 25313
rect 25682 25304 25688 25316
rect 25740 25304 25746 25356
rect 25961 25347 26019 25353
rect 25961 25313 25973 25347
rect 26007 25344 26019 25347
rect 27522 25344 27528 25356
rect 26007 25316 27528 25344
rect 26007 25313 26019 25316
rect 25961 25307 26019 25313
rect 27522 25304 27528 25316
rect 27580 25304 27586 25356
rect 28920 25353 28948 25384
rect 30745 25381 30757 25415
rect 30791 25412 30803 25415
rect 31662 25412 31668 25424
rect 30791 25384 31668 25412
rect 30791 25381 30803 25384
rect 30745 25375 30803 25381
rect 31662 25372 31668 25384
rect 31720 25372 31726 25424
rect 37366 25412 37372 25424
rect 33888 25384 37372 25412
rect 28905 25347 28963 25353
rect 28905 25313 28917 25347
rect 28951 25313 28963 25347
rect 28905 25307 28963 25313
rect 30006 25304 30012 25356
rect 30064 25344 30070 25356
rect 31297 25347 31355 25353
rect 31297 25344 31309 25347
rect 30064 25316 31309 25344
rect 30064 25304 30070 25316
rect 31297 25313 31309 25316
rect 31343 25313 31355 25347
rect 31297 25307 31355 25313
rect 31846 25304 31852 25356
rect 31904 25344 31910 25356
rect 32493 25347 32551 25353
rect 32493 25344 32505 25347
rect 31904 25316 32505 25344
rect 31904 25304 31910 25316
rect 32493 25313 32505 25316
rect 32539 25313 32551 25347
rect 32493 25307 32551 25313
rect 1765 25279 1823 25285
rect 1765 25245 1777 25279
rect 1811 25276 1823 25279
rect 4154 25276 4160 25288
rect 1811 25248 4160 25276
rect 1811 25245 1823 25248
rect 1765 25239 1823 25245
rect 4154 25236 4160 25248
rect 4212 25236 4218 25288
rect 5077 25279 5135 25285
rect 5077 25245 5089 25279
rect 5123 25276 5135 25279
rect 6270 25276 6276 25288
rect 5123 25248 6276 25276
rect 5123 25245 5135 25248
rect 5077 25239 5135 25245
rect 6270 25236 6276 25248
rect 6328 25236 6334 25288
rect 10594 25236 10600 25288
rect 10652 25236 10658 25288
rect 14461 25279 14519 25285
rect 14461 25245 14473 25279
rect 14507 25276 14519 25279
rect 16482 25276 16488 25288
rect 14507 25248 16488 25276
rect 14507 25245 14519 25248
rect 14461 25239 14519 25245
rect 16482 25236 16488 25248
rect 16540 25236 16546 25288
rect 22646 25236 22652 25288
rect 22704 25236 22710 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25276 24087 25279
rect 24949 25279 25007 25285
rect 24949 25276 24961 25279
rect 24075 25248 24961 25276
rect 24075 25245 24087 25248
rect 24029 25239 24087 25245
rect 24949 25245 24961 25248
rect 24995 25245 25007 25279
rect 24949 25239 25007 25245
rect 28258 25236 28264 25288
rect 28316 25276 28322 25288
rect 28721 25279 28779 25285
rect 28721 25276 28733 25279
rect 28316 25248 28733 25276
rect 28316 25236 28322 25248
rect 28721 25245 28733 25248
rect 28767 25245 28779 25279
rect 28721 25239 28779 25245
rect 28813 25279 28871 25285
rect 28813 25245 28825 25279
rect 28859 25276 28871 25279
rect 28994 25276 29000 25288
rect 28859 25248 29000 25276
rect 28859 25245 28871 25248
rect 28813 25239 28871 25245
rect 28994 25236 29000 25248
rect 29052 25236 29058 25288
rect 29086 25236 29092 25288
rect 29144 25276 29150 25288
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29144 25248 29929 25276
rect 29144 25236 29150 25248
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 31205 25279 31263 25285
rect 31205 25245 31217 25279
rect 31251 25276 31263 25279
rect 31754 25276 31760 25288
rect 31251 25248 31760 25276
rect 31251 25245 31263 25248
rect 31205 25239 31263 25245
rect 31754 25236 31760 25248
rect 31812 25236 31818 25288
rect 31938 25236 31944 25288
rect 31996 25276 32002 25288
rect 33888 25285 33916 25384
rect 37366 25372 37372 25384
rect 37424 25372 37430 25424
rect 39408 25412 39436 25452
rect 39482 25440 39488 25492
rect 39540 25440 39546 25492
rect 49142 25412 49148 25424
rect 39408 25384 49148 25412
rect 49142 25372 49148 25384
rect 49200 25372 49206 25424
rect 33962 25304 33968 25356
rect 34020 25304 34026 25356
rect 34054 25304 34060 25356
rect 34112 25304 34118 25356
rect 35618 25304 35624 25356
rect 35676 25344 35682 25356
rect 35713 25347 35771 25353
rect 35713 25344 35725 25347
rect 35676 25316 35725 25344
rect 35676 25304 35682 25316
rect 35713 25313 35725 25316
rect 35759 25313 35771 25347
rect 35713 25307 35771 25313
rect 35986 25304 35992 25356
rect 36044 25344 36050 25356
rect 37001 25347 37059 25353
rect 37001 25344 37013 25347
rect 36044 25316 37013 25344
rect 36044 25304 36050 25316
rect 37001 25313 37013 25316
rect 37047 25313 37059 25347
rect 37001 25307 37059 25313
rect 37185 25347 37243 25353
rect 37185 25313 37197 25347
rect 37231 25344 37243 25347
rect 38013 25347 38071 25353
rect 38013 25344 38025 25347
rect 37231 25316 38025 25344
rect 37231 25313 37243 25316
rect 37185 25307 37243 25313
rect 38013 25313 38025 25316
rect 38059 25344 38071 25347
rect 38562 25344 38568 25356
rect 38059 25316 38568 25344
rect 38059 25313 38071 25316
rect 38013 25307 38071 25313
rect 38562 25304 38568 25316
rect 38620 25304 38626 25356
rect 40494 25304 40500 25356
rect 40552 25304 40558 25356
rect 40678 25304 40684 25356
rect 40736 25304 40742 25356
rect 32401 25279 32459 25285
rect 32401 25276 32413 25279
rect 31996 25248 32413 25276
rect 31996 25236 32002 25248
rect 32401 25245 32413 25248
rect 32447 25245 32459 25279
rect 32401 25239 32459 25245
rect 33873 25279 33931 25285
rect 33873 25245 33885 25279
rect 33919 25245 33931 25279
rect 33873 25239 33931 25245
rect 34882 25236 34888 25288
rect 34940 25276 34946 25288
rect 37737 25279 37795 25285
rect 37737 25276 37749 25279
rect 34940 25248 37749 25276
rect 34940 25236 34946 25248
rect 37737 25245 37749 25248
rect 37783 25245 37795 25279
rect 37737 25239 37795 25245
rect 43438 25236 43444 25288
rect 43496 25276 43502 25288
rect 45281 25279 45339 25285
rect 45281 25276 45293 25279
rect 43496 25248 45293 25276
rect 43496 25236 43502 25248
rect 45281 25245 45293 25248
rect 45327 25245 45339 25279
rect 45281 25239 45339 25245
rect 45554 25236 45560 25288
rect 45612 25276 45618 25288
rect 46017 25279 46075 25285
rect 46017 25276 46029 25279
rect 45612 25248 46029 25276
rect 45612 25236 45618 25248
rect 46017 25245 46029 25248
rect 46063 25245 46075 25279
rect 46017 25239 46075 25245
rect 22741 25211 22799 25217
rect 22741 25177 22753 25211
rect 22787 25208 22799 25211
rect 25406 25208 25412 25220
rect 22787 25180 25412 25208
rect 22787 25177 22799 25180
rect 22741 25171 22799 25177
rect 25406 25168 25412 25180
rect 25464 25168 25470 25220
rect 26237 25211 26295 25217
rect 26237 25177 26249 25211
rect 26283 25177 26295 25211
rect 26237 25171 26295 25177
rect 22278 25100 22284 25152
rect 22336 25100 22342 25152
rect 23290 25100 23296 25152
rect 23348 25140 23354 25152
rect 24581 25143 24639 25149
rect 24581 25140 24593 25143
rect 23348 25112 24593 25140
rect 23348 25100 23354 25112
rect 24581 25109 24593 25112
rect 24627 25109 24639 25143
rect 24581 25103 24639 25109
rect 25041 25143 25099 25149
rect 25041 25109 25053 25143
rect 25087 25140 25099 25143
rect 26142 25140 26148 25152
rect 25087 25112 26148 25140
rect 25087 25109 25099 25112
rect 25041 25103 25099 25109
rect 26142 25100 26148 25112
rect 26200 25100 26206 25152
rect 26252 25140 26280 25171
rect 26694 25168 26700 25220
rect 26752 25168 26758 25220
rect 32214 25208 32220 25220
rect 28368 25180 32220 25208
rect 27614 25140 27620 25152
rect 26252 25112 27620 25140
rect 27614 25100 27620 25112
rect 27672 25100 27678 25152
rect 28368 25149 28396 25180
rect 32214 25168 32220 25180
rect 32272 25168 32278 25220
rect 32309 25211 32367 25217
rect 32309 25177 32321 25211
rect 32355 25208 32367 25211
rect 34514 25208 34520 25220
rect 32355 25180 34520 25208
rect 32355 25177 32367 25180
rect 32309 25171 32367 25177
rect 34514 25168 34520 25180
rect 34572 25168 34578 25220
rect 34790 25168 34796 25220
rect 34848 25208 34854 25220
rect 35621 25211 35679 25217
rect 35621 25208 35633 25211
rect 34848 25180 35633 25208
rect 34848 25168 34854 25180
rect 35621 25177 35633 25180
rect 35667 25177 35679 25211
rect 35621 25171 35679 25177
rect 36464 25180 36860 25208
rect 28353 25143 28411 25149
rect 28353 25109 28365 25143
rect 28399 25109 28411 25143
rect 28353 25103 28411 25109
rect 28994 25100 29000 25152
rect 29052 25140 29058 25152
rect 31113 25143 31171 25149
rect 31113 25140 31125 25143
rect 29052 25112 31125 25140
rect 29052 25100 29058 25112
rect 31113 25109 31125 25112
rect 31159 25109 31171 25143
rect 31113 25103 31171 25109
rect 31294 25100 31300 25152
rect 31352 25140 31358 25152
rect 31941 25143 31999 25149
rect 31941 25140 31953 25143
rect 31352 25112 31953 25140
rect 31352 25100 31358 25112
rect 31941 25109 31953 25112
rect 31987 25109 31999 25143
rect 31941 25103 31999 25109
rect 32766 25100 32772 25152
rect 32824 25140 32830 25152
rect 33505 25143 33563 25149
rect 33505 25140 33517 25143
rect 32824 25112 33517 25140
rect 32824 25100 32830 25112
rect 33505 25109 33517 25112
rect 33551 25109 33563 25143
rect 33505 25103 33563 25109
rect 35158 25100 35164 25152
rect 35216 25100 35222 25152
rect 35529 25143 35587 25149
rect 35529 25109 35541 25143
rect 35575 25140 35587 25143
rect 36464 25140 36492 25180
rect 35575 25112 36492 25140
rect 35575 25109 35587 25112
rect 35529 25103 35587 25109
rect 36538 25100 36544 25152
rect 36596 25100 36602 25152
rect 36832 25140 36860 25180
rect 36906 25168 36912 25220
rect 36964 25168 36970 25220
rect 39666 25208 39672 25220
rect 39238 25180 39672 25208
rect 39666 25168 39672 25180
rect 39724 25168 39730 25220
rect 44358 25168 44364 25220
rect 44416 25168 44422 25220
rect 45462 25168 45468 25220
rect 45520 25168 45526 25220
rect 46201 25211 46259 25217
rect 46201 25177 46213 25211
rect 46247 25208 46259 25211
rect 47486 25208 47492 25220
rect 46247 25180 47492 25208
rect 46247 25177 46259 25180
rect 46201 25171 46259 25177
rect 47486 25168 47492 25180
rect 47544 25168 47550 25220
rect 38746 25140 38752 25152
rect 36832 25112 38752 25140
rect 38746 25100 38752 25112
rect 38804 25100 38810 25152
rect 40034 25100 40040 25152
rect 40092 25100 40098 25152
rect 40402 25100 40408 25152
rect 40460 25100 40466 25152
rect 44450 25100 44456 25152
rect 44508 25100 44514 25152
rect 1104 25050 49864 25072
rect 1104 24998 7950 25050
rect 8002 24998 8014 25050
rect 8066 24998 8078 25050
rect 8130 24998 8142 25050
rect 8194 24998 8206 25050
rect 8258 24998 17950 25050
rect 18002 24998 18014 25050
rect 18066 24998 18078 25050
rect 18130 24998 18142 25050
rect 18194 24998 18206 25050
rect 18258 24998 27950 25050
rect 28002 24998 28014 25050
rect 28066 24998 28078 25050
rect 28130 24998 28142 25050
rect 28194 24998 28206 25050
rect 28258 24998 37950 25050
rect 38002 24998 38014 25050
rect 38066 24998 38078 25050
rect 38130 24998 38142 25050
rect 38194 24998 38206 25050
rect 38258 24998 47950 25050
rect 48002 24998 48014 25050
rect 48066 24998 48078 25050
rect 48130 24998 48142 25050
rect 48194 24998 48206 25050
rect 48258 24998 49864 25050
rect 1104 24976 49864 24998
rect 25774 24896 25780 24948
rect 25832 24896 25838 24948
rect 27430 24936 27436 24948
rect 27080 24908 27436 24936
rect 20990 24828 20996 24880
rect 21048 24828 21054 24880
rect 8440 24803 8498 24809
rect 8440 24769 8452 24803
rect 8486 24800 8498 24803
rect 9306 24800 9312 24812
rect 8486 24772 9312 24800
rect 8486 24769 8498 24772
rect 8440 24763 8498 24769
rect 9306 24760 9312 24772
rect 9364 24760 9370 24812
rect 8294 24692 8300 24744
rect 8352 24732 8358 24744
rect 8527 24735 8585 24741
rect 8527 24732 8539 24735
rect 8352 24704 8539 24732
rect 8352 24692 8358 24704
rect 8527 24701 8539 24704
rect 8573 24701 8585 24735
rect 8527 24695 8585 24701
rect 19702 24692 19708 24744
rect 19760 24692 19766 24744
rect 19981 24735 20039 24741
rect 19981 24701 19993 24735
rect 20027 24732 20039 24735
rect 21266 24732 21272 24744
rect 20027 24704 21272 24732
rect 20027 24701 20039 24704
rect 19981 24695 20039 24701
rect 21266 24692 21272 24704
rect 21324 24692 21330 24744
rect 25314 24692 25320 24744
rect 25372 24732 25378 24744
rect 25590 24732 25596 24744
rect 25372 24704 25596 24732
rect 25372 24692 25378 24704
rect 25590 24692 25596 24704
rect 25648 24732 25654 24744
rect 25869 24735 25927 24741
rect 25869 24732 25881 24735
rect 25648 24704 25881 24732
rect 25648 24692 25654 24704
rect 25869 24701 25881 24704
rect 25915 24701 25927 24735
rect 25869 24695 25927 24701
rect 26053 24735 26111 24741
rect 26053 24701 26065 24735
rect 26099 24732 26111 24735
rect 27080 24732 27108 24908
rect 27430 24896 27436 24908
rect 27488 24896 27494 24948
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 28902 24936 28908 24948
rect 27672 24908 28908 24936
rect 27672 24896 27678 24908
rect 28902 24896 28908 24908
rect 28960 24896 28966 24948
rect 30926 24896 30932 24948
rect 30984 24936 30990 24948
rect 32769 24939 32827 24945
rect 32769 24936 32781 24939
rect 30984 24908 32781 24936
rect 30984 24896 30990 24908
rect 32769 24905 32781 24908
rect 32815 24905 32827 24939
rect 35986 24936 35992 24948
rect 32769 24899 32827 24905
rect 32876 24908 35992 24936
rect 27522 24868 27528 24880
rect 27172 24840 27528 24868
rect 27172 24809 27200 24840
rect 27522 24828 27528 24840
rect 27580 24828 27586 24880
rect 27706 24828 27712 24880
rect 27764 24868 27770 24880
rect 29641 24871 29699 24877
rect 27764 24840 27922 24868
rect 27764 24828 27770 24840
rect 29641 24837 29653 24871
rect 29687 24868 29699 24871
rect 29914 24868 29920 24880
rect 29687 24840 29920 24868
rect 29687 24837 29699 24840
rect 29641 24831 29699 24837
rect 29914 24828 29920 24840
rect 29972 24828 29978 24880
rect 32214 24828 32220 24880
rect 32272 24868 32278 24880
rect 32876 24868 32904 24908
rect 35986 24896 35992 24908
rect 36044 24896 36050 24948
rect 36538 24896 36544 24948
rect 36596 24936 36602 24948
rect 37829 24939 37887 24945
rect 37829 24936 37841 24939
rect 36596 24908 37841 24936
rect 36596 24896 36602 24908
rect 37829 24905 37841 24908
rect 37875 24905 37887 24939
rect 37829 24899 37887 24905
rect 32272 24840 32904 24868
rect 32272 24828 32278 24840
rect 34238 24828 34244 24880
rect 34296 24828 34302 24880
rect 37458 24828 37464 24880
rect 37516 24868 37522 24880
rect 38470 24868 38476 24880
rect 37516 24840 38476 24868
rect 37516 24828 37522 24840
rect 38470 24828 38476 24840
rect 38528 24828 38534 24880
rect 27157 24803 27215 24809
rect 27157 24769 27169 24803
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 30742 24760 30748 24812
rect 30800 24760 30806 24812
rect 32858 24760 32864 24812
rect 32916 24760 32922 24812
rect 33870 24760 33876 24812
rect 33928 24800 33934 24812
rect 33965 24803 34023 24809
rect 33965 24800 33977 24803
rect 33928 24772 33977 24800
rect 33928 24760 33934 24772
rect 33965 24769 33977 24772
rect 34011 24769 34023 24803
rect 33965 24763 34023 24769
rect 35342 24760 35348 24812
rect 35400 24760 35406 24812
rect 37182 24760 37188 24812
rect 37240 24800 37246 24812
rect 37921 24803 37979 24809
rect 37921 24800 37933 24803
rect 37240 24772 37933 24800
rect 37240 24760 37246 24772
rect 37921 24769 37933 24772
rect 37967 24769 37979 24803
rect 37921 24763 37979 24769
rect 40221 24803 40279 24809
rect 40221 24769 40233 24803
rect 40267 24800 40279 24803
rect 40402 24800 40408 24812
rect 40267 24772 40408 24800
rect 40267 24769 40279 24772
rect 40221 24763 40279 24769
rect 40402 24760 40408 24772
rect 40460 24760 40466 24812
rect 47210 24760 47216 24812
rect 47268 24800 47274 24812
rect 47949 24803 48007 24809
rect 47949 24800 47961 24803
rect 47268 24772 47961 24800
rect 47268 24760 47274 24772
rect 47949 24769 47961 24772
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 26099 24704 27108 24732
rect 26099 24701 26111 24704
rect 26053 24695 26111 24701
rect 27430 24692 27436 24744
rect 27488 24692 27494 24744
rect 27522 24692 27528 24744
rect 27580 24732 27586 24744
rect 28166 24732 28172 24744
rect 27580 24704 28172 24732
rect 27580 24692 27586 24704
rect 28166 24692 28172 24704
rect 28224 24732 28230 24744
rect 29365 24735 29423 24741
rect 29365 24732 29377 24735
rect 28224 24704 29377 24732
rect 28224 24692 28230 24704
rect 29365 24701 29377 24704
rect 29411 24732 29423 24735
rect 30098 24732 30104 24744
rect 29411 24704 30104 24732
rect 29411 24701 29423 24704
rect 29365 24695 29423 24701
rect 30098 24692 30104 24704
rect 30156 24692 30162 24744
rect 21726 24624 21732 24676
rect 21784 24664 21790 24676
rect 21910 24664 21916 24676
rect 21784 24636 21916 24664
rect 21784 24624 21790 24636
rect 21910 24624 21916 24636
rect 21968 24664 21974 24676
rect 26878 24664 26884 24676
rect 21968 24636 26884 24664
rect 21968 24624 21974 24636
rect 26878 24624 26884 24636
rect 26936 24624 26942 24676
rect 30760 24664 30788 24760
rect 31110 24692 31116 24744
rect 31168 24692 31174 24744
rect 32582 24692 32588 24744
rect 32640 24732 32646 24744
rect 32953 24735 33011 24741
rect 32953 24732 32965 24735
rect 32640 24704 32965 24732
rect 32640 24692 32646 24704
rect 32953 24701 32965 24704
rect 32999 24701 33011 24735
rect 32953 24695 33011 24701
rect 33318 24692 33324 24744
rect 33376 24732 33382 24744
rect 35989 24735 36047 24741
rect 35989 24732 36001 24735
rect 33376 24704 36001 24732
rect 33376 24692 33382 24704
rect 35989 24701 36001 24704
rect 36035 24701 36047 24735
rect 35989 24695 36047 24701
rect 38105 24735 38163 24741
rect 38105 24701 38117 24735
rect 38151 24732 38163 24735
rect 39482 24732 39488 24744
rect 38151 24704 39488 24732
rect 38151 24701 38163 24704
rect 38105 24695 38163 24701
rect 39482 24692 39488 24704
rect 39540 24692 39546 24744
rect 49142 24692 49148 24744
rect 49200 24692 49206 24744
rect 31570 24664 31576 24676
rect 30760 24636 31576 24664
rect 31570 24624 31576 24636
rect 31628 24624 31634 24676
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 25409 24599 25467 24605
rect 25409 24565 25421 24599
rect 25455 24596 25467 24599
rect 28994 24596 29000 24608
rect 25455 24568 29000 24596
rect 25455 24565 25467 24568
rect 25409 24559 25467 24565
rect 28994 24556 29000 24568
rect 29052 24556 29058 24608
rect 32398 24556 32404 24608
rect 32456 24556 32462 24608
rect 33870 24556 33876 24608
rect 33928 24596 33934 24608
rect 34882 24596 34888 24608
rect 33928 24568 34888 24596
rect 33928 24556 33934 24568
rect 34882 24556 34888 24568
rect 34940 24556 34946 24608
rect 34974 24556 34980 24608
rect 35032 24596 35038 24608
rect 37461 24599 37519 24605
rect 37461 24596 37473 24599
rect 35032 24568 37473 24596
rect 35032 24556 35038 24568
rect 37461 24565 37473 24568
rect 37507 24565 37519 24599
rect 37461 24559 37519 24565
rect 1104 24506 49864 24528
rect 1104 24454 2950 24506
rect 3002 24454 3014 24506
rect 3066 24454 3078 24506
rect 3130 24454 3142 24506
rect 3194 24454 3206 24506
rect 3258 24454 12950 24506
rect 13002 24454 13014 24506
rect 13066 24454 13078 24506
rect 13130 24454 13142 24506
rect 13194 24454 13206 24506
rect 13258 24454 22950 24506
rect 23002 24454 23014 24506
rect 23066 24454 23078 24506
rect 23130 24454 23142 24506
rect 23194 24454 23206 24506
rect 23258 24454 32950 24506
rect 33002 24454 33014 24506
rect 33066 24454 33078 24506
rect 33130 24454 33142 24506
rect 33194 24454 33206 24506
rect 33258 24454 42950 24506
rect 43002 24454 43014 24506
rect 43066 24454 43078 24506
rect 43130 24454 43142 24506
rect 43194 24454 43206 24506
rect 43258 24454 49864 24506
rect 1104 24432 49864 24454
rect 10873 24395 10931 24401
rect 10873 24361 10885 24395
rect 10919 24361 10931 24395
rect 10873 24355 10931 24361
rect 10888 24324 10916 24355
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 16393 24395 16451 24401
rect 16393 24392 16405 24395
rect 12400 24364 16405 24392
rect 12400 24352 12406 24364
rect 16393 24361 16405 24364
rect 16439 24361 16451 24395
rect 25498 24392 25504 24404
rect 16393 24355 16451 24361
rect 17236 24364 25504 24392
rect 14550 24324 14556 24336
rect 10888 24296 14556 24324
rect 14550 24284 14556 24296
rect 14608 24284 14614 24336
rect 14645 24259 14703 24265
rect 14645 24225 14657 24259
rect 14691 24256 14703 24259
rect 15286 24256 15292 24268
rect 14691 24228 15292 24256
rect 14691 24225 14703 24228
rect 14645 24219 14703 24225
rect 15286 24216 15292 24228
rect 15344 24216 15350 24268
rect 10594 24148 10600 24200
rect 10652 24188 10658 24200
rect 12526 24188 12532 24200
rect 10652 24160 12532 24188
rect 10652 24148 10658 24160
rect 12526 24148 12532 24160
rect 12584 24148 12590 24200
rect 14921 24123 14979 24129
rect 14921 24089 14933 24123
rect 14967 24120 14979 24123
rect 15194 24120 15200 24132
rect 14967 24092 15200 24120
rect 14967 24089 14979 24092
rect 14921 24083 14979 24089
rect 15194 24080 15200 24092
rect 15252 24080 15258 24132
rect 15378 24080 15384 24132
rect 15436 24080 15442 24132
rect 7834 24012 7840 24064
rect 7892 24052 7898 24064
rect 11057 24055 11115 24061
rect 11057 24052 11069 24055
rect 7892 24024 11069 24052
rect 7892 24012 7898 24024
rect 11057 24021 11069 24024
rect 11103 24021 11115 24055
rect 11057 24015 11115 24021
rect 11146 24012 11152 24064
rect 11204 24052 11210 24064
rect 17236 24052 17264 24364
rect 25498 24352 25504 24364
rect 25556 24352 25562 24404
rect 27617 24395 27675 24401
rect 27617 24361 27629 24395
rect 27663 24392 27675 24395
rect 28442 24392 28448 24404
rect 27663 24364 28448 24392
rect 27663 24361 27675 24364
rect 27617 24355 27675 24361
rect 28442 24352 28448 24364
rect 28500 24352 28506 24404
rect 28902 24352 28908 24404
rect 28960 24392 28966 24404
rect 36630 24392 36636 24404
rect 28960 24364 30236 24392
rect 28960 24352 28966 24364
rect 29086 24324 29092 24336
rect 28184 24296 29092 24324
rect 19702 24216 19708 24268
rect 19760 24256 19766 24268
rect 20809 24259 20867 24265
rect 20809 24256 20821 24259
rect 19760 24228 20821 24256
rect 19760 24216 19766 24228
rect 20809 24225 20821 24228
rect 20855 24256 20867 24259
rect 21818 24256 21824 24268
rect 20855 24228 21824 24256
rect 20855 24225 20867 24228
rect 20809 24219 20867 24225
rect 21818 24216 21824 24228
rect 21876 24216 21882 24268
rect 22830 24216 22836 24268
rect 22888 24256 22894 24268
rect 25593 24259 25651 24265
rect 25593 24256 25605 24259
rect 22888 24228 25605 24256
rect 22888 24216 22894 24228
rect 25593 24225 25605 24228
rect 25639 24225 25651 24259
rect 25593 24219 25651 24225
rect 26878 24216 26884 24268
rect 26936 24216 26942 24268
rect 27065 24259 27123 24265
rect 27065 24225 27077 24259
rect 27111 24256 27123 24259
rect 27430 24256 27436 24268
rect 27111 24228 27436 24256
rect 27111 24225 27123 24228
rect 27065 24219 27123 24225
rect 27430 24216 27436 24228
rect 27488 24256 27494 24268
rect 28074 24256 28080 24268
rect 27488 24228 28080 24256
rect 27488 24216 27494 24228
rect 28074 24216 28080 24228
rect 28132 24216 28138 24268
rect 25498 24148 25504 24200
rect 25556 24188 25562 24200
rect 26237 24191 26295 24197
rect 26237 24188 26249 24191
rect 25556 24160 26249 24188
rect 25556 24148 25562 24160
rect 26237 24157 26249 24160
rect 26283 24157 26295 24191
rect 26237 24151 26295 24157
rect 27985 24191 28043 24197
rect 27985 24157 27997 24191
rect 28031 24188 28043 24191
rect 28184 24188 28212 24296
rect 29086 24284 29092 24296
rect 29144 24284 29150 24336
rect 29733 24327 29791 24333
rect 29733 24293 29745 24327
rect 29779 24293 29791 24327
rect 30208 24324 30236 24364
rect 33980 24364 36636 24392
rect 30208 24296 30328 24324
rect 29733 24287 29791 24293
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24225 28319 24259
rect 28261 24219 28319 24225
rect 28031 24160 28212 24188
rect 28276 24188 28304 24219
rect 28350 24216 28356 24268
rect 28408 24256 28414 24268
rect 28718 24256 28724 24268
rect 28408 24228 28724 24256
rect 28408 24216 28414 24228
rect 28718 24216 28724 24228
rect 28776 24216 28782 24268
rect 29546 24256 29552 24268
rect 28920 24228 29552 24256
rect 28276 24160 28396 24188
rect 28031 24157 28043 24160
rect 27985 24151 28043 24157
rect 21085 24123 21143 24129
rect 21085 24089 21097 24123
rect 21131 24120 21143 24123
rect 21358 24120 21364 24132
rect 21131 24092 21364 24120
rect 21131 24089 21143 24092
rect 21085 24083 21143 24089
rect 21358 24080 21364 24092
rect 21416 24080 21422 24132
rect 23474 24120 23480 24132
rect 22310 24092 23480 24120
rect 23474 24080 23480 24092
rect 23532 24080 23538 24132
rect 28368 24120 28396 24160
rect 28442 24148 28448 24200
rect 28500 24188 28506 24200
rect 28920 24188 28948 24228
rect 29546 24216 29552 24228
rect 29604 24216 29610 24268
rect 28500 24160 28948 24188
rect 29748 24188 29776 24287
rect 30190 24216 30196 24268
rect 30248 24216 30254 24268
rect 30300 24265 30328 24296
rect 32214 24284 32220 24336
rect 32272 24324 32278 24336
rect 33686 24324 33692 24336
rect 32272 24296 33692 24324
rect 32272 24284 32278 24296
rect 33686 24284 33692 24296
rect 33744 24284 33750 24336
rect 30285 24259 30343 24265
rect 30285 24225 30297 24259
rect 30331 24225 30343 24259
rect 33980 24256 34008 24364
rect 36630 24352 36636 24364
rect 36688 24352 36694 24404
rect 34057 24259 34115 24265
rect 34057 24256 34069 24259
rect 33980 24228 34069 24256
rect 30285 24219 30343 24225
rect 34057 24225 34069 24228
rect 34103 24225 34115 24259
rect 34057 24219 34115 24225
rect 34241 24259 34299 24265
rect 34241 24225 34253 24259
rect 34287 24256 34299 24259
rect 34514 24256 34520 24268
rect 34287 24228 34520 24256
rect 34287 24225 34299 24228
rect 34241 24219 34299 24225
rect 34514 24216 34520 24228
rect 34572 24256 34578 24268
rect 34572 24228 34836 24256
rect 34572 24216 34578 24228
rect 32858 24188 32864 24200
rect 29748 24160 32864 24188
rect 28500 24148 28506 24160
rect 32858 24148 32864 24160
rect 32916 24148 32922 24200
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 33965 24191 34023 24197
rect 33965 24188 33977 24191
rect 33836 24160 33977 24188
rect 33836 24148 33842 24160
rect 33965 24157 33977 24160
rect 34011 24188 34023 24191
rect 34330 24188 34336 24200
rect 34011 24160 34336 24188
rect 34011 24157 34023 24160
rect 33965 24151 34023 24157
rect 34330 24148 34336 24160
rect 34388 24148 34394 24200
rect 29822 24120 29828 24132
rect 26436 24092 28304 24120
rect 28368 24092 29828 24120
rect 11204 24024 17264 24052
rect 11204 24012 11210 24024
rect 21266 24012 21272 24064
rect 21324 24052 21330 24064
rect 22554 24052 22560 24064
rect 21324 24024 22560 24052
rect 21324 24012 21330 24024
rect 22554 24012 22560 24024
rect 22612 24012 22618 24064
rect 23842 24012 23848 24064
rect 23900 24052 23906 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 23900 24024 25053 24052
rect 23900 24012 23906 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25041 24015 25099 24021
rect 25409 24055 25467 24061
rect 25409 24021 25421 24055
rect 25455 24052 25467 24055
rect 26234 24052 26240 24064
rect 25455 24024 26240 24052
rect 25455 24021 25467 24024
rect 25409 24015 25467 24021
rect 26234 24012 26240 24024
rect 26292 24012 26298 24064
rect 26436 24061 26464 24092
rect 26421 24055 26479 24061
rect 26421 24021 26433 24055
rect 26467 24021 26479 24055
rect 26421 24015 26479 24021
rect 26786 24012 26792 24064
rect 26844 24012 26850 24064
rect 27798 24012 27804 24064
rect 27856 24052 27862 24064
rect 28077 24055 28135 24061
rect 28077 24052 28089 24055
rect 27856 24024 28089 24052
rect 27856 24012 27862 24024
rect 28077 24021 28089 24024
rect 28123 24021 28135 24055
rect 28276 24052 28304 24092
rect 29822 24080 29828 24092
rect 29880 24080 29886 24132
rect 30834 24080 30840 24132
rect 30892 24120 30898 24132
rect 34808 24120 34836 24228
rect 35342 24216 35348 24268
rect 35400 24256 35406 24268
rect 35400 24228 36308 24256
rect 35400 24216 35406 24228
rect 34882 24148 34888 24200
rect 34940 24188 34946 24200
rect 34977 24191 35035 24197
rect 34977 24188 34989 24191
rect 34940 24160 34989 24188
rect 34940 24148 34946 24160
rect 34977 24157 34989 24160
rect 35023 24157 35035 24191
rect 34977 24151 35035 24157
rect 36280 24132 36308 24228
rect 37274 24216 37280 24268
rect 37332 24256 37338 24268
rect 37737 24259 37795 24265
rect 37737 24256 37749 24259
rect 37332 24228 37749 24256
rect 37332 24216 37338 24228
rect 37737 24225 37749 24228
rect 37783 24225 37795 24259
rect 37737 24219 37795 24225
rect 40310 24216 40316 24268
rect 40368 24256 40374 24268
rect 40497 24259 40555 24265
rect 40497 24256 40509 24259
rect 40368 24228 40509 24256
rect 40368 24216 40374 24228
rect 40497 24225 40509 24228
rect 40543 24225 40555 24259
rect 40497 24219 40555 24225
rect 40681 24259 40739 24265
rect 40681 24225 40693 24259
rect 40727 24256 40739 24259
rect 40770 24256 40776 24268
rect 40727 24228 40776 24256
rect 40727 24225 40739 24228
rect 40681 24219 40739 24225
rect 40770 24216 40776 24228
rect 40828 24216 40834 24268
rect 37645 24191 37703 24197
rect 37645 24157 37657 24191
rect 37691 24188 37703 24191
rect 37826 24188 37832 24200
rect 37691 24160 37832 24188
rect 37691 24157 37703 24160
rect 37645 24151 37703 24157
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 40034 24148 40040 24200
rect 40092 24188 40098 24200
rect 40405 24191 40463 24197
rect 40405 24188 40417 24191
rect 40092 24160 40417 24188
rect 40092 24148 40098 24160
rect 40405 24157 40417 24160
rect 40451 24157 40463 24191
rect 40405 24151 40463 24157
rect 47854 24148 47860 24200
rect 47912 24188 47918 24200
rect 47949 24191 48007 24197
rect 47949 24188 47961 24191
rect 47912 24160 47961 24188
rect 47912 24148 47918 24160
rect 47949 24157 47961 24160
rect 47995 24157 48007 24191
rect 47949 24151 48007 24157
rect 35253 24123 35311 24129
rect 35253 24120 35265 24123
rect 30892 24092 34376 24120
rect 34808 24092 35265 24120
rect 30892 24080 30898 24092
rect 34348 24064 34376 24092
rect 35253 24089 35265 24092
rect 35299 24120 35311 24123
rect 35526 24120 35532 24132
rect 35299 24092 35532 24120
rect 35299 24089 35311 24092
rect 35253 24083 35311 24089
rect 35526 24080 35532 24092
rect 35584 24080 35590 24132
rect 36262 24080 36268 24132
rect 36320 24080 36326 24132
rect 49142 24080 49148 24132
rect 49200 24080 49206 24132
rect 30101 24055 30159 24061
rect 30101 24052 30113 24055
rect 28276 24024 30113 24052
rect 28077 24015 28135 24021
rect 30101 24021 30113 24024
rect 30147 24021 30159 24055
rect 30101 24015 30159 24021
rect 33597 24055 33655 24061
rect 33597 24021 33609 24055
rect 33643 24052 33655 24055
rect 33870 24052 33876 24064
rect 33643 24024 33876 24052
rect 33643 24021 33655 24024
rect 33597 24015 33655 24021
rect 33870 24012 33876 24024
rect 33928 24012 33934 24064
rect 34330 24012 34336 24064
rect 34388 24012 34394 24064
rect 35342 24012 35348 24064
rect 35400 24052 35406 24064
rect 35618 24052 35624 24064
rect 35400 24024 35624 24052
rect 35400 24012 35406 24024
rect 35618 24012 35624 24024
rect 35676 24052 35682 24064
rect 36725 24055 36783 24061
rect 36725 24052 36737 24055
rect 35676 24024 36737 24052
rect 35676 24012 35682 24024
rect 36725 24021 36737 24024
rect 36771 24021 36783 24055
rect 36725 24015 36783 24021
rect 37185 24055 37243 24061
rect 37185 24021 37197 24055
rect 37231 24052 37243 24055
rect 37366 24052 37372 24064
rect 37231 24024 37372 24052
rect 37231 24021 37243 24024
rect 37185 24015 37243 24021
rect 37366 24012 37372 24024
rect 37424 24012 37430 24064
rect 37553 24055 37611 24061
rect 37553 24021 37565 24055
rect 37599 24052 37611 24055
rect 37826 24052 37832 24064
rect 37599 24024 37832 24052
rect 37599 24021 37611 24024
rect 37553 24015 37611 24021
rect 37826 24012 37832 24024
rect 37884 24052 37890 24064
rect 39206 24052 39212 24064
rect 37884 24024 39212 24052
rect 37884 24012 37890 24024
rect 39206 24012 39212 24024
rect 39264 24012 39270 24064
rect 40034 24012 40040 24064
rect 40092 24012 40098 24064
rect 1104 23962 49864 23984
rect 1104 23910 7950 23962
rect 8002 23910 8014 23962
rect 8066 23910 8078 23962
rect 8130 23910 8142 23962
rect 8194 23910 8206 23962
rect 8258 23910 17950 23962
rect 18002 23910 18014 23962
rect 18066 23910 18078 23962
rect 18130 23910 18142 23962
rect 18194 23910 18206 23962
rect 18258 23910 27950 23962
rect 28002 23910 28014 23962
rect 28066 23910 28078 23962
rect 28130 23910 28142 23962
rect 28194 23910 28206 23962
rect 28258 23910 37950 23962
rect 38002 23910 38014 23962
rect 38066 23910 38078 23962
rect 38130 23910 38142 23962
rect 38194 23910 38206 23962
rect 38258 23910 47950 23962
rect 48002 23910 48014 23962
rect 48066 23910 48078 23962
rect 48130 23910 48142 23962
rect 48194 23910 48206 23962
rect 48258 23910 49864 23962
rect 1104 23888 49864 23910
rect 6270 23808 6276 23860
rect 6328 23848 6334 23860
rect 9401 23851 9459 23857
rect 9401 23848 9413 23851
rect 6328 23820 9413 23848
rect 6328 23808 6334 23820
rect 9401 23817 9413 23820
rect 9447 23817 9459 23851
rect 15286 23848 15292 23860
rect 9401 23811 9459 23817
rect 13004 23820 15292 23848
rect 13004 23780 13032 23820
rect 15286 23808 15292 23820
rect 15344 23808 15350 23860
rect 16482 23808 16488 23860
rect 16540 23848 16546 23860
rect 19337 23851 19395 23857
rect 19337 23848 19349 23851
rect 16540 23820 19349 23848
rect 16540 23808 16546 23820
rect 19337 23817 19349 23820
rect 19383 23817 19395 23851
rect 19337 23811 19395 23817
rect 19705 23851 19763 23857
rect 19705 23817 19717 23851
rect 19751 23848 19763 23851
rect 20717 23851 20775 23857
rect 20717 23848 20729 23851
rect 19751 23820 20729 23848
rect 19751 23817 19763 23820
rect 19705 23811 19763 23817
rect 20717 23817 20729 23820
rect 20763 23817 20775 23851
rect 20717 23811 20775 23817
rect 21085 23851 21143 23857
rect 21085 23817 21097 23851
rect 21131 23848 21143 23851
rect 23290 23848 23296 23860
rect 21131 23820 23296 23848
rect 21131 23817 21143 23820
rect 21085 23811 21143 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 26237 23851 26295 23857
rect 26237 23817 26249 23851
rect 26283 23848 26295 23851
rect 30834 23848 30840 23860
rect 26283 23820 30840 23848
rect 26283 23817 26295 23820
rect 26237 23811 26295 23817
rect 30834 23808 30840 23820
rect 30892 23808 30898 23860
rect 32582 23808 32588 23860
rect 32640 23848 32646 23860
rect 34514 23848 34520 23860
rect 32640 23820 34520 23848
rect 32640 23808 32646 23820
rect 34514 23808 34520 23820
rect 34572 23808 34578 23860
rect 38194 23808 38200 23860
rect 38252 23848 38258 23860
rect 38562 23848 38568 23860
rect 38252 23820 38568 23848
rect 38252 23808 38258 23820
rect 38562 23808 38568 23820
rect 38620 23808 38626 23860
rect 15378 23780 15384 23792
rect 12912 23752 13032 23780
rect 14398 23752 15384 23780
rect 8757 23715 8815 23721
rect 8757 23681 8769 23715
rect 8803 23712 8815 23715
rect 12250 23712 12256 23724
rect 8803 23684 12256 23712
rect 8803 23681 8815 23684
rect 8757 23675 8815 23681
rect 12250 23672 12256 23684
rect 12308 23672 12314 23724
rect 12912 23721 12940 23752
rect 15378 23740 15384 23752
rect 15436 23740 15442 23792
rect 21450 23780 21456 23792
rect 19996 23752 21456 23780
rect 12897 23715 12955 23721
rect 12897 23681 12909 23715
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 7834 23604 7840 23656
rect 7892 23644 7898 23656
rect 8941 23647 8999 23653
rect 8941 23644 8953 23647
rect 7892 23616 8953 23644
rect 7892 23604 7898 23616
rect 8941 23613 8953 23616
rect 8987 23613 8999 23647
rect 8941 23607 8999 23613
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 13173 23647 13231 23653
rect 13173 23644 13185 23647
rect 12400 23616 13185 23644
rect 12400 23604 12406 23616
rect 13173 23613 13185 23616
rect 13219 23613 13231 23647
rect 13173 23607 13231 23613
rect 14550 23604 14556 23656
rect 14608 23644 14614 23656
rect 19996 23653 20024 23752
rect 21450 23740 21456 23752
rect 21508 23780 21514 23792
rect 22281 23783 22339 23789
rect 22281 23780 22293 23783
rect 21508 23752 22293 23780
rect 21508 23740 21514 23752
rect 22281 23749 22293 23752
rect 22327 23749 22339 23783
rect 26786 23780 26792 23792
rect 22281 23743 22339 23749
rect 25424 23752 26792 23780
rect 22002 23672 22008 23724
rect 22060 23672 22066 23724
rect 25424 23721 25452 23752
rect 26786 23740 26792 23752
rect 26844 23740 26850 23792
rect 26896 23752 29040 23780
rect 25409 23715 25467 23721
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 14608 23616 14657 23644
rect 14608 23604 14614 23616
rect 14645 23613 14657 23616
rect 14691 23613 14703 23647
rect 14645 23607 14703 23613
rect 19797 23647 19855 23653
rect 19797 23613 19809 23647
rect 19843 23613 19855 23647
rect 19797 23607 19855 23613
rect 19981 23647 20039 23653
rect 19981 23613 19993 23647
rect 20027 23613 20039 23647
rect 19981 23607 20039 23613
rect 19812 23508 19840 23607
rect 21174 23604 21180 23656
rect 21232 23604 21238 23656
rect 21266 23604 21272 23656
rect 21324 23604 21330 23656
rect 23400 23644 23428 23698
rect 25409 23681 25421 23715
rect 25455 23681 25467 23715
rect 26896 23712 26924 23752
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 25409 23675 25467 23681
rect 25516 23684 26924 23712
rect 28460 23684 28641 23712
rect 23474 23644 23480 23656
rect 23400 23616 23480 23644
rect 23474 23604 23480 23616
rect 23532 23604 23538 23656
rect 23658 23604 23664 23656
rect 23716 23644 23722 23656
rect 24029 23647 24087 23653
rect 24029 23644 24041 23647
rect 23716 23616 24041 23644
rect 23716 23604 23722 23616
rect 24029 23613 24041 23616
rect 24075 23644 24087 23647
rect 24670 23644 24676 23656
rect 24075 23616 24676 23644
rect 24075 23613 24087 23616
rect 24029 23607 24087 23613
rect 24670 23604 24676 23616
rect 24728 23644 24734 23656
rect 25516 23644 25544 23684
rect 26329 23647 26387 23653
rect 26329 23644 26341 23647
rect 24728 23616 25544 23644
rect 25608 23616 26341 23644
rect 24728 23604 24734 23616
rect 23382 23536 23388 23588
rect 23440 23576 23446 23588
rect 25608 23576 25636 23616
rect 26329 23613 26341 23616
rect 26375 23613 26387 23647
rect 26329 23607 26387 23613
rect 26513 23647 26571 23653
rect 26513 23613 26525 23647
rect 26559 23644 26571 23647
rect 27062 23644 27068 23656
rect 26559 23616 27068 23644
rect 26559 23613 26571 23616
rect 26513 23607 26571 23613
rect 27062 23604 27068 23616
rect 27120 23604 27126 23656
rect 23440 23548 25636 23576
rect 23440 23536 23446 23548
rect 26694 23536 26700 23588
rect 26752 23576 26758 23588
rect 27890 23576 27896 23588
rect 26752 23548 27896 23576
rect 26752 23536 26758 23548
rect 27890 23536 27896 23548
rect 27948 23536 27954 23588
rect 28460 23576 28488 23684
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 28629 23675 28687 23681
rect 28721 23715 28779 23721
rect 28721 23681 28733 23715
rect 28767 23712 28779 23715
rect 28902 23712 28908 23724
rect 28767 23684 28908 23712
rect 28767 23681 28779 23684
rect 28721 23675 28779 23681
rect 28902 23672 28908 23684
rect 28960 23672 28966 23724
rect 28813 23647 28871 23653
rect 28813 23613 28825 23647
rect 28859 23644 28871 23647
rect 29012 23644 29040 23752
rect 29270 23740 29276 23792
rect 29328 23780 29334 23792
rect 31478 23780 31484 23792
rect 29328 23752 31484 23780
rect 29328 23740 29334 23752
rect 31478 23740 31484 23752
rect 31536 23740 31542 23792
rect 33870 23740 33876 23792
rect 33928 23780 33934 23792
rect 34977 23783 35035 23789
rect 34977 23780 34989 23783
rect 33928 23752 34989 23780
rect 33928 23740 33934 23752
rect 34977 23749 34989 23752
rect 35023 23749 35035 23783
rect 34977 23743 35035 23749
rect 37274 23740 37280 23792
rect 37332 23780 37338 23792
rect 39025 23783 39083 23789
rect 39025 23780 39037 23783
rect 37332 23752 39037 23780
rect 37332 23740 37338 23752
rect 39025 23749 39037 23752
rect 39071 23749 39083 23783
rect 39025 23743 39083 23749
rect 39666 23740 39672 23792
rect 39724 23740 39730 23792
rect 33686 23672 33692 23724
rect 33744 23672 33750 23724
rect 34885 23715 34943 23721
rect 34885 23681 34897 23715
rect 34931 23681 34943 23715
rect 34885 23675 34943 23681
rect 28859 23616 29040 23644
rect 28859 23613 28871 23616
rect 28813 23607 28871 23613
rect 30098 23604 30104 23656
rect 30156 23644 30162 23656
rect 32306 23644 32312 23656
rect 30156 23616 32312 23644
rect 30156 23604 30162 23616
rect 32306 23604 32312 23616
rect 32364 23604 32370 23656
rect 32674 23604 32680 23656
rect 32732 23644 32738 23656
rect 34900 23644 34928 23675
rect 38286 23672 38292 23724
rect 38344 23712 38350 23724
rect 38562 23712 38568 23724
rect 38344 23684 38568 23712
rect 38344 23672 38350 23684
rect 38562 23672 38568 23684
rect 38620 23712 38626 23724
rect 38749 23715 38807 23721
rect 38749 23712 38761 23715
rect 38620 23684 38761 23712
rect 38620 23672 38626 23684
rect 38749 23681 38761 23684
rect 38795 23681 38807 23715
rect 38749 23675 38807 23681
rect 46842 23672 46848 23724
rect 46900 23712 46906 23724
rect 47949 23715 48007 23721
rect 47949 23712 47961 23715
rect 46900 23684 47961 23712
rect 46900 23672 46906 23684
rect 47949 23681 47961 23684
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 32732 23616 34928 23644
rect 35161 23647 35219 23653
rect 32732 23604 32738 23616
rect 35161 23613 35173 23647
rect 35207 23644 35219 23647
rect 35250 23644 35256 23656
rect 35207 23616 35256 23644
rect 35207 23613 35219 23616
rect 35161 23607 35219 23613
rect 35250 23604 35256 23616
rect 35308 23604 35314 23656
rect 35526 23604 35532 23656
rect 35584 23644 35590 23656
rect 39482 23644 39488 23656
rect 35584 23616 39488 23644
rect 35584 23604 35590 23616
rect 39482 23604 39488 23616
rect 39540 23604 39546 23656
rect 47486 23604 47492 23656
rect 47544 23644 47550 23656
rect 47854 23644 47860 23656
rect 47544 23616 47860 23644
rect 47544 23604 47550 23616
rect 47854 23604 47860 23616
rect 47912 23604 47918 23656
rect 49142 23604 49148 23656
rect 49200 23604 49206 23656
rect 28460 23548 28672 23576
rect 22094 23508 22100 23520
rect 19812 23480 22100 23508
rect 22094 23468 22100 23480
rect 22152 23468 22158 23520
rect 24765 23511 24823 23517
rect 24765 23477 24777 23511
rect 24811 23508 24823 23511
rect 24946 23508 24952 23520
rect 24811 23480 24952 23508
rect 24811 23477 24823 23480
rect 24765 23471 24823 23477
rect 24946 23468 24952 23480
rect 25004 23468 25010 23520
rect 25866 23468 25872 23520
rect 25924 23468 25930 23520
rect 26142 23468 26148 23520
rect 26200 23508 26206 23520
rect 28261 23511 28319 23517
rect 28261 23508 28273 23511
rect 26200 23480 28273 23508
rect 26200 23468 26206 23480
rect 28261 23477 28273 23480
rect 28307 23477 28319 23511
rect 28644 23508 28672 23548
rect 28902 23536 28908 23588
rect 28960 23576 28966 23588
rect 31478 23576 31484 23588
rect 28960 23548 31484 23576
rect 28960 23536 28966 23548
rect 31478 23536 31484 23548
rect 31536 23576 31542 23588
rect 32030 23576 32036 23588
rect 31536 23548 32036 23576
rect 31536 23536 31542 23548
rect 32030 23536 32036 23548
rect 32088 23536 32094 23588
rect 34054 23536 34060 23588
rect 34112 23536 34118 23588
rect 32214 23508 32220 23520
rect 28644 23480 32220 23508
rect 28261 23471 28319 23477
rect 32214 23468 32220 23480
rect 32272 23468 32278 23520
rect 32572 23511 32630 23517
rect 32572 23477 32584 23511
rect 32618 23508 32630 23511
rect 34146 23508 34152 23520
rect 32618 23480 34152 23508
rect 32618 23477 32630 23480
rect 32572 23471 32630 23477
rect 34146 23468 34152 23480
rect 34204 23468 34210 23520
rect 34514 23468 34520 23520
rect 34572 23468 34578 23520
rect 38746 23468 38752 23520
rect 38804 23508 38810 23520
rect 39574 23508 39580 23520
rect 38804 23480 39580 23508
rect 38804 23468 38810 23480
rect 39574 23468 39580 23480
rect 39632 23508 39638 23520
rect 40497 23511 40555 23517
rect 40497 23508 40509 23511
rect 39632 23480 40509 23508
rect 39632 23468 39638 23480
rect 40497 23477 40509 23480
rect 40543 23477 40555 23511
rect 40497 23471 40555 23477
rect 1104 23418 49864 23440
rect 1104 23366 2950 23418
rect 3002 23366 3014 23418
rect 3066 23366 3078 23418
rect 3130 23366 3142 23418
rect 3194 23366 3206 23418
rect 3258 23366 12950 23418
rect 13002 23366 13014 23418
rect 13066 23366 13078 23418
rect 13130 23366 13142 23418
rect 13194 23366 13206 23418
rect 13258 23366 22950 23418
rect 23002 23366 23014 23418
rect 23066 23366 23078 23418
rect 23130 23366 23142 23418
rect 23194 23366 23206 23418
rect 23258 23366 32950 23418
rect 33002 23366 33014 23418
rect 33066 23366 33078 23418
rect 33130 23366 33142 23418
rect 33194 23366 33206 23418
rect 33258 23366 42950 23418
rect 43002 23366 43014 23418
rect 43066 23366 43078 23418
rect 43130 23366 43142 23418
rect 43194 23366 43206 23418
rect 43258 23366 49864 23418
rect 1104 23344 49864 23366
rect 4154 23264 4160 23316
rect 4212 23304 4218 23316
rect 5169 23307 5227 23313
rect 5169 23304 5181 23307
rect 4212 23276 5181 23304
rect 4212 23264 4218 23276
rect 5169 23273 5181 23276
rect 5215 23273 5227 23307
rect 5169 23267 5227 23273
rect 22186 23264 22192 23316
rect 22244 23304 22250 23316
rect 22557 23307 22615 23313
rect 22557 23304 22569 23307
rect 22244 23276 22569 23304
rect 22244 23264 22250 23276
rect 22557 23273 22569 23276
rect 22603 23304 22615 23307
rect 22738 23304 22744 23316
rect 22603 23276 22744 23304
rect 22603 23273 22615 23276
rect 22557 23267 22615 23273
rect 22738 23264 22744 23276
rect 22796 23264 22802 23316
rect 27430 23304 27436 23316
rect 27264 23276 27436 23304
rect 1302 23128 1308 23180
rect 1360 23168 1366 23180
rect 2041 23171 2099 23177
rect 2041 23168 2053 23171
rect 1360 23140 2053 23168
rect 1360 23128 1366 23140
rect 2041 23137 2053 23140
rect 2087 23137 2099 23171
rect 5534 23168 5540 23180
rect 2041 23131 2099 23137
rect 3528 23140 5540 23168
rect 1765 23103 1823 23109
rect 1765 23069 1777 23103
rect 1811 23100 1823 23103
rect 3528 23100 3556 23140
rect 5534 23128 5540 23140
rect 5592 23128 5598 23180
rect 9030 23128 9036 23180
rect 9088 23168 9094 23180
rect 9263 23171 9321 23177
rect 9263 23168 9275 23171
rect 9088 23140 9275 23168
rect 9088 23128 9094 23140
rect 9263 23137 9275 23140
rect 9309 23137 9321 23171
rect 9263 23131 9321 23137
rect 15286 23128 15292 23180
rect 15344 23168 15350 23180
rect 17129 23171 17187 23177
rect 17129 23168 17141 23171
rect 15344 23140 17141 23168
rect 15344 23128 15350 23140
rect 17129 23137 17141 23140
rect 17175 23168 17187 23171
rect 19429 23171 19487 23177
rect 19429 23168 19441 23171
rect 17175 23140 19441 23168
rect 17175 23137 17187 23140
rect 17129 23131 17187 23137
rect 19429 23137 19441 23140
rect 19475 23168 19487 23171
rect 19702 23168 19708 23180
rect 19475 23140 19708 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19702 23128 19708 23140
rect 19760 23128 19766 23180
rect 22756 23168 22784 23264
rect 27264 23236 27292 23276
rect 27430 23264 27436 23276
rect 27488 23304 27494 23316
rect 27488 23276 28488 23304
rect 27488 23264 27494 23276
rect 25240 23208 27292 23236
rect 28460 23236 28488 23276
rect 28718 23264 28724 23316
rect 28776 23304 28782 23316
rect 28905 23307 28963 23313
rect 28905 23304 28917 23307
rect 28776 23276 28917 23304
rect 28776 23264 28782 23276
rect 28905 23273 28917 23276
rect 28951 23273 28963 23307
rect 31110 23304 31116 23316
rect 28905 23267 28963 23273
rect 29012 23276 31116 23304
rect 29012 23236 29040 23276
rect 31110 23264 31116 23276
rect 31168 23264 31174 23316
rect 31846 23264 31852 23316
rect 31904 23264 31910 23316
rect 34057 23307 34115 23313
rect 34057 23273 34069 23307
rect 34103 23304 34115 23307
rect 34146 23304 34152 23316
rect 34103 23276 34152 23304
rect 34103 23273 34115 23276
rect 34057 23267 34115 23273
rect 34146 23264 34152 23276
rect 34204 23264 34210 23316
rect 34238 23264 34244 23316
rect 34296 23304 34302 23316
rect 36633 23307 36691 23313
rect 36633 23304 36645 23307
rect 34296 23276 36645 23304
rect 34296 23264 34302 23276
rect 36633 23273 36645 23276
rect 36679 23273 36691 23307
rect 36633 23267 36691 23273
rect 37461 23307 37519 23313
rect 37461 23273 37473 23307
rect 37507 23304 37519 23307
rect 41230 23304 41236 23316
rect 37507 23276 41236 23304
rect 37507 23273 37519 23276
rect 37461 23267 37519 23273
rect 41230 23264 41236 23276
rect 41288 23264 41294 23316
rect 32122 23236 32128 23248
rect 28460 23208 29040 23236
rect 31404 23208 32128 23236
rect 23477 23171 23535 23177
rect 23477 23168 23489 23171
rect 22756 23140 23489 23168
rect 23477 23137 23489 23140
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 23658 23128 23664 23180
rect 23716 23128 23722 23180
rect 25240 23177 25268 23208
rect 25225 23171 25283 23177
rect 25225 23137 25237 23171
rect 25271 23137 25283 23171
rect 25225 23131 25283 23137
rect 27157 23171 27215 23177
rect 27157 23137 27169 23171
rect 27203 23168 27215 23171
rect 27522 23168 27528 23180
rect 27203 23140 27528 23168
rect 27203 23137 27215 23140
rect 27157 23131 27215 23137
rect 27522 23128 27528 23140
rect 27580 23128 27586 23180
rect 27890 23128 27896 23180
rect 27948 23168 27954 23180
rect 27948 23140 28580 23168
rect 27948 23128 27954 23140
rect 28552 23112 28580 23140
rect 30098 23128 30104 23180
rect 30156 23128 30162 23180
rect 30377 23171 30435 23177
rect 30377 23137 30389 23171
rect 30423 23168 30435 23171
rect 31404 23168 31432 23208
rect 32122 23196 32128 23208
rect 32180 23196 32186 23248
rect 32232 23208 32444 23236
rect 30423 23140 31432 23168
rect 30423 23137 30435 23140
rect 30377 23131 30435 23137
rect 31570 23128 31576 23180
rect 31628 23128 31634 23180
rect 1811 23072 3556 23100
rect 4157 23103 4215 23109
rect 1811 23069 1823 23072
rect 1765 23063 1823 23069
rect 4157 23069 4169 23103
rect 4203 23100 4215 23103
rect 4982 23100 4988 23112
rect 4203 23072 4988 23100
rect 4203 23069 4215 23072
rect 4157 23063 4215 23069
rect 4982 23060 4988 23072
rect 5040 23060 5046 23112
rect 9176 23103 9234 23109
rect 9176 23069 9188 23103
rect 9222 23100 9234 23103
rect 9766 23100 9772 23112
rect 9222 23072 9772 23100
rect 9222 23069 9234 23072
rect 9176 23063 9234 23069
rect 9766 23060 9772 23072
rect 9824 23060 9830 23112
rect 23382 23060 23388 23112
rect 23440 23060 23446 23112
rect 24946 23060 24952 23112
rect 25004 23060 25010 23112
rect 28534 23060 28540 23112
rect 28592 23060 28598 23112
rect 31588 23100 31616 23128
rect 32232 23100 32260 23208
rect 32306 23128 32312 23180
rect 32364 23128 32370 23180
rect 32416 23168 32444 23208
rect 38378 23196 38384 23248
rect 38436 23236 38442 23248
rect 38436 23208 41414 23236
rect 38436 23196 38442 23208
rect 34885 23171 34943 23177
rect 32416 23140 33732 23168
rect 33704 23112 33732 23140
rect 34885 23137 34897 23171
rect 34931 23168 34943 23171
rect 37458 23168 37464 23180
rect 34931 23140 37464 23168
rect 34931 23137 34943 23140
rect 34885 23131 34943 23137
rect 37458 23128 37464 23140
rect 37516 23128 37522 23180
rect 38746 23128 38752 23180
rect 38804 23128 38810 23180
rect 31510 23072 32260 23100
rect 33686 23060 33692 23112
rect 33744 23100 33750 23112
rect 34422 23100 34428 23112
rect 33744 23072 34428 23100
rect 33744 23060 33750 23072
rect 34422 23060 34428 23072
rect 34480 23060 34486 23112
rect 37645 23103 37703 23109
rect 37645 23100 37657 23103
rect 36464 23072 37657 23100
rect 5077 23035 5135 23041
rect 5077 23001 5089 23035
rect 5123 23032 5135 23035
rect 9674 23032 9680 23044
rect 5123 23004 9680 23032
rect 5123 23001 5135 23004
rect 5077 22995 5135 23001
rect 9674 22992 9680 23004
rect 9732 22992 9738 23044
rect 17402 22992 17408 23044
rect 17460 22992 17466 23044
rect 19705 23035 19763 23041
rect 17788 23004 17894 23032
rect 18800 23004 19334 23032
rect 2774 22924 2780 22976
rect 2832 22964 2838 22976
rect 4249 22967 4307 22973
rect 4249 22964 4261 22967
rect 2832 22936 4261 22964
rect 2832 22924 2838 22936
rect 4249 22933 4261 22936
rect 4295 22933 4307 22967
rect 4249 22927 4307 22933
rect 15378 22924 15384 22976
rect 15436 22964 15442 22976
rect 17788 22964 17816 23004
rect 18800 22964 18828 23004
rect 15436 22936 18828 22964
rect 15436 22924 15442 22936
rect 18874 22924 18880 22976
rect 18932 22924 18938 22976
rect 19306 22964 19334 23004
rect 19705 23001 19717 23035
rect 19751 23032 19763 23035
rect 19978 23032 19984 23044
rect 19751 23004 19984 23032
rect 19751 23001 19763 23004
rect 19705 22995 19763 23001
rect 19978 22992 19984 23004
rect 20036 22992 20042 23044
rect 20990 23032 20996 23044
rect 20930 23004 20996 23032
rect 20990 22992 20996 23004
rect 21048 22992 21054 23044
rect 23658 22992 23664 23044
rect 23716 23032 23722 23044
rect 27433 23035 27491 23041
rect 23716 23004 27384 23032
rect 23716 22992 23722 23004
rect 21008 22964 21036 22992
rect 19306 22936 21036 22964
rect 21177 22967 21235 22973
rect 21177 22933 21189 22967
rect 21223 22964 21235 22967
rect 21266 22964 21272 22976
rect 21223 22936 21272 22964
rect 21223 22933 21235 22936
rect 21177 22927 21235 22933
rect 21266 22924 21272 22936
rect 21324 22924 21330 22976
rect 22646 22924 22652 22976
rect 22704 22964 22710 22976
rect 23017 22967 23075 22973
rect 23017 22964 23029 22967
rect 22704 22936 23029 22964
rect 22704 22924 22710 22936
rect 23017 22933 23029 22936
rect 23063 22933 23075 22967
rect 23017 22927 23075 22933
rect 24578 22924 24584 22976
rect 24636 22924 24642 22976
rect 25038 22924 25044 22976
rect 25096 22924 25102 22976
rect 27356 22964 27384 23004
rect 27433 23001 27445 23035
rect 27479 23032 27491 23035
rect 27522 23032 27528 23044
rect 27479 23004 27528 23032
rect 27479 23001 27491 23004
rect 27433 22995 27491 23001
rect 27522 22992 27528 23004
rect 27580 22992 27586 23044
rect 27890 22992 27896 23044
rect 27948 22992 27954 23044
rect 31754 22992 31760 23044
rect 31812 23032 31818 23044
rect 32585 23035 32643 23041
rect 32585 23032 32597 23035
rect 31812 23004 32597 23032
rect 31812 22992 31818 23004
rect 32585 23001 32597 23004
rect 32631 23001 32643 23035
rect 35161 23035 35219 23041
rect 32585 22995 32643 23001
rect 33980 23004 34192 23032
rect 29178 22964 29184 22976
rect 27356 22936 29184 22964
rect 29178 22924 29184 22936
rect 29236 22964 29242 22976
rect 29454 22964 29460 22976
rect 29236 22936 29460 22964
rect 29236 22924 29242 22936
rect 29454 22924 29460 22936
rect 29512 22924 29518 22976
rect 30650 22924 30656 22976
rect 30708 22964 30714 22976
rect 33980 22964 34008 23004
rect 30708 22936 34008 22964
rect 34164 22964 34192 23004
rect 35161 23001 35173 23035
rect 35207 23032 35219 23035
rect 35250 23032 35256 23044
rect 35207 23004 35256 23032
rect 35207 23001 35219 23004
rect 35161 22995 35219 23001
rect 35250 22992 35256 23004
rect 35308 22992 35314 23044
rect 36170 22992 36176 23044
rect 36228 22992 36234 23044
rect 36464 22964 36492 23072
rect 37645 23069 37657 23072
rect 37691 23069 37703 23103
rect 37645 23063 37703 23069
rect 38565 23103 38623 23109
rect 38565 23069 38577 23103
rect 38611 23100 38623 23103
rect 40221 23103 40279 23109
rect 40221 23100 40233 23103
rect 38611 23072 40233 23100
rect 38611 23069 38623 23072
rect 38565 23063 38623 23069
rect 40221 23069 40233 23072
rect 40267 23069 40279 23103
rect 41386 23100 41414 23208
rect 44177 23103 44235 23109
rect 44177 23100 44189 23103
rect 41386 23072 44189 23100
rect 40221 23063 40279 23069
rect 44177 23069 44189 23072
rect 44223 23069 44235 23103
rect 44177 23063 44235 23069
rect 47670 23060 47676 23112
rect 47728 23100 47734 23112
rect 47949 23103 48007 23109
rect 47949 23100 47961 23103
rect 47728 23072 47961 23100
rect 47728 23060 47734 23072
rect 47949 23069 47961 23072
rect 47995 23069 48007 23103
rect 47949 23063 48007 23069
rect 37366 22992 37372 23044
rect 37424 23032 37430 23044
rect 38657 23035 38715 23041
rect 38657 23032 38669 23035
rect 37424 23004 38669 23032
rect 37424 22992 37430 23004
rect 38657 23001 38669 23004
rect 38703 23001 38715 23035
rect 38657 22995 38715 23001
rect 44361 23035 44419 23041
rect 44361 23001 44373 23035
rect 44407 23032 44419 23035
rect 46658 23032 46664 23044
rect 44407 23004 46664 23032
rect 44407 23001 44419 23004
rect 44361 22995 44419 23001
rect 46658 22992 46664 23004
rect 46716 22992 46722 23044
rect 49142 22992 49148 23044
rect 49200 22992 49206 23044
rect 34164 22936 36492 22964
rect 30708 22924 30714 22936
rect 37182 22924 37188 22976
rect 37240 22964 37246 22976
rect 37826 22964 37832 22976
rect 37240 22936 37832 22964
rect 37240 22924 37246 22936
rect 37826 22924 37832 22936
rect 37884 22924 37890 22976
rect 38197 22967 38255 22973
rect 38197 22933 38209 22967
rect 38243 22964 38255 22967
rect 38286 22964 38292 22976
rect 38243 22936 38292 22964
rect 38243 22933 38255 22936
rect 38197 22927 38255 22933
rect 38286 22924 38292 22936
rect 38344 22924 38350 22976
rect 1104 22874 49864 22896
rect 1104 22822 7950 22874
rect 8002 22822 8014 22874
rect 8066 22822 8078 22874
rect 8130 22822 8142 22874
rect 8194 22822 8206 22874
rect 8258 22822 17950 22874
rect 18002 22822 18014 22874
rect 18066 22822 18078 22874
rect 18130 22822 18142 22874
rect 18194 22822 18206 22874
rect 18258 22822 27950 22874
rect 28002 22822 28014 22874
rect 28066 22822 28078 22874
rect 28130 22822 28142 22874
rect 28194 22822 28206 22874
rect 28258 22822 37950 22874
rect 38002 22822 38014 22874
rect 38066 22822 38078 22874
rect 38130 22822 38142 22874
rect 38194 22822 38206 22874
rect 38258 22822 47950 22874
rect 48002 22822 48014 22874
rect 48066 22822 48078 22874
rect 48130 22822 48142 22874
rect 48194 22822 48206 22874
rect 48258 22822 49864 22874
rect 1104 22800 49864 22822
rect 17773 22763 17831 22769
rect 17773 22729 17785 22763
rect 17819 22760 17831 22763
rect 19337 22763 19395 22769
rect 19337 22760 19349 22763
rect 17819 22732 19349 22760
rect 17819 22729 17831 22732
rect 17773 22723 17831 22729
rect 19337 22729 19349 22732
rect 19383 22729 19395 22763
rect 19337 22723 19395 22729
rect 19705 22763 19763 22769
rect 19705 22729 19717 22763
rect 19751 22760 19763 22763
rect 22278 22760 22284 22772
rect 19751 22732 22284 22760
rect 19751 22729 19763 22732
rect 19705 22723 19763 22729
rect 22278 22720 22284 22732
rect 22336 22720 22342 22772
rect 23658 22720 23664 22772
rect 23716 22720 23722 22772
rect 24578 22720 24584 22772
rect 24636 22760 24642 22772
rect 30009 22763 30067 22769
rect 30009 22760 30021 22763
rect 24636 22732 30021 22760
rect 24636 22720 24642 22732
rect 30009 22729 30021 22732
rect 30055 22729 30067 22763
rect 30009 22723 30067 22729
rect 30101 22763 30159 22769
rect 30101 22729 30113 22763
rect 30147 22760 30159 22763
rect 30466 22760 30472 22772
rect 30147 22732 30472 22760
rect 30147 22729 30159 22732
rect 30101 22723 30159 22729
rect 30466 22720 30472 22732
rect 30524 22720 30530 22772
rect 31021 22763 31079 22769
rect 31021 22729 31033 22763
rect 31067 22760 31079 22763
rect 32674 22760 32680 22772
rect 31067 22732 32680 22760
rect 31067 22729 31079 22732
rect 31021 22723 31079 22729
rect 32674 22720 32680 22732
rect 32732 22720 32738 22772
rect 34057 22763 34115 22769
rect 34057 22729 34069 22763
rect 34103 22760 34115 22763
rect 34514 22760 34520 22772
rect 34103 22732 34520 22760
rect 34103 22729 34115 22732
rect 34057 22723 34115 22729
rect 34514 22720 34520 22732
rect 34572 22720 34578 22772
rect 38562 22760 38568 22772
rect 37660 22732 38568 22760
rect 17402 22652 17408 22704
rect 17460 22692 17466 22704
rect 21177 22695 21235 22701
rect 17460 22664 19932 22692
rect 17460 22652 17466 22664
rect 15194 22584 15200 22636
rect 15252 22624 15258 22636
rect 18874 22624 18880 22636
rect 15252 22596 18880 22624
rect 15252 22584 15258 22596
rect 17972 22565 18000 22596
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 17865 22559 17923 22565
rect 17865 22525 17877 22559
rect 17911 22525 17923 22559
rect 17865 22519 17923 22525
rect 17957 22559 18015 22565
rect 17957 22525 17969 22559
rect 18003 22525 18015 22559
rect 17957 22519 18015 22525
rect 17880 22488 17908 22519
rect 19794 22516 19800 22568
rect 19852 22516 19858 22568
rect 19904 22565 19932 22664
rect 21177 22661 21189 22695
rect 21223 22692 21235 22695
rect 21910 22692 21916 22704
rect 21223 22664 21916 22692
rect 21223 22661 21235 22664
rect 21177 22655 21235 22661
rect 21910 22652 21916 22664
rect 21968 22652 21974 22704
rect 23750 22652 23756 22704
rect 23808 22692 23814 22704
rect 26326 22692 26332 22704
rect 23808 22664 26332 22692
rect 23808 22652 23814 22664
rect 26326 22652 26332 22664
rect 26384 22652 26390 22704
rect 27430 22652 27436 22704
rect 27488 22652 27494 22704
rect 30374 22652 30380 22704
rect 30432 22692 30438 22704
rect 31481 22695 31539 22701
rect 31481 22692 31493 22695
rect 30432 22664 31493 22692
rect 30432 22652 30438 22664
rect 31481 22661 31493 22664
rect 31527 22692 31539 22695
rect 34149 22695 34207 22701
rect 31527 22664 34100 22692
rect 31527 22661 31539 22664
rect 31481 22655 31539 22661
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22624 21143 22627
rect 23290 22624 23296 22636
rect 21131 22596 23296 22624
rect 21131 22593 21143 22596
rect 21085 22587 21143 22593
rect 23290 22584 23296 22596
rect 23348 22584 23354 22636
rect 24949 22627 25007 22633
rect 24949 22593 24961 22627
rect 24995 22624 25007 22627
rect 25961 22627 26019 22633
rect 25961 22624 25973 22627
rect 24995 22596 25973 22624
rect 24995 22593 25007 22596
rect 24949 22587 25007 22593
rect 25961 22593 25973 22596
rect 26007 22593 26019 22627
rect 25961 22587 26019 22593
rect 28534 22584 28540 22636
rect 28592 22584 28598 22636
rect 31389 22627 31447 22633
rect 31389 22593 31401 22627
rect 31435 22624 31447 22627
rect 32493 22627 32551 22633
rect 32493 22624 32505 22627
rect 31435 22596 32505 22624
rect 31435 22593 31447 22596
rect 31389 22587 31447 22593
rect 32493 22593 32505 22596
rect 32539 22593 32551 22627
rect 34072 22624 34100 22664
rect 34149 22661 34161 22695
rect 34195 22692 34207 22695
rect 35158 22692 35164 22704
rect 34195 22664 35164 22692
rect 34195 22661 34207 22664
rect 34149 22655 34207 22661
rect 35158 22652 35164 22664
rect 35216 22652 35222 22704
rect 37182 22624 37188 22636
rect 34072 22596 37188 22624
rect 32493 22587 32551 22593
rect 37182 22584 37188 22596
rect 37240 22584 37246 22636
rect 37458 22584 37464 22636
rect 37516 22624 37522 22636
rect 37660 22633 37688 22732
rect 38562 22720 38568 22732
rect 38620 22720 38626 22772
rect 39666 22760 39672 22772
rect 39040 22732 39672 22760
rect 37826 22652 37832 22704
rect 37884 22692 37890 22704
rect 37921 22695 37979 22701
rect 37921 22692 37933 22695
rect 37884 22664 37933 22692
rect 37884 22652 37890 22664
rect 37921 22661 37933 22664
rect 37967 22661 37979 22695
rect 37921 22655 37979 22661
rect 39040 22636 39068 22732
rect 39666 22720 39672 22732
rect 39724 22720 39730 22772
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 37516 22596 37657 22624
rect 37516 22584 37522 22596
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 39022 22584 39028 22636
rect 39080 22584 39086 22636
rect 19889 22559 19947 22565
rect 19889 22525 19901 22559
rect 19935 22556 19947 22559
rect 21266 22556 21272 22568
rect 19935 22528 21272 22556
rect 19935 22525 19947 22528
rect 19889 22519 19947 22525
rect 21266 22516 21272 22528
rect 21324 22516 21330 22568
rect 23937 22559 23995 22565
rect 23937 22525 23949 22559
rect 23983 22556 23995 22559
rect 25041 22559 25099 22565
rect 23983 22528 24992 22556
rect 23983 22525 23995 22528
rect 23937 22519 23995 22525
rect 20717 22491 20775 22497
rect 20717 22488 20729 22491
rect 17880 22460 20729 22488
rect 20717 22457 20729 22460
rect 20763 22457 20775 22491
rect 20717 22451 20775 22457
rect 17402 22380 17408 22432
rect 17460 22380 17466 22432
rect 21634 22380 21640 22432
rect 21692 22420 21698 22432
rect 23293 22423 23351 22429
rect 23293 22420 23305 22423
rect 21692 22392 23305 22420
rect 21692 22380 21698 22392
rect 23293 22389 23305 22392
rect 23339 22389 23351 22423
rect 23293 22383 23351 22389
rect 23382 22380 23388 22432
rect 23440 22420 23446 22432
rect 24581 22423 24639 22429
rect 24581 22420 24593 22423
rect 23440 22392 24593 22420
rect 23440 22380 23446 22392
rect 24581 22389 24593 22392
rect 24627 22389 24639 22423
rect 24964 22420 24992 22528
rect 25041 22525 25053 22559
rect 25087 22525 25099 22559
rect 25041 22519 25099 22525
rect 25056 22488 25084 22519
rect 25130 22516 25136 22568
rect 25188 22516 25194 22568
rect 27157 22559 27215 22565
rect 27157 22525 27169 22559
rect 27203 22525 27215 22559
rect 27157 22519 27215 22525
rect 26510 22488 26516 22500
rect 25056 22460 26516 22488
rect 26510 22448 26516 22460
rect 26568 22448 26574 22500
rect 25038 22420 25044 22432
rect 24964 22392 25044 22420
rect 24581 22383 24639 22389
rect 25038 22380 25044 22392
rect 25096 22420 25102 22432
rect 26602 22420 26608 22432
rect 25096 22392 26608 22420
rect 25096 22380 25102 22392
rect 26602 22380 26608 22392
rect 26660 22380 26666 22432
rect 27172 22420 27200 22519
rect 27522 22516 27528 22568
rect 27580 22556 27586 22568
rect 28905 22559 28963 22565
rect 28905 22556 28917 22559
rect 27580 22528 28917 22556
rect 27580 22516 27586 22528
rect 28905 22525 28917 22528
rect 28951 22556 28963 22559
rect 30193 22559 30251 22565
rect 30193 22556 30205 22559
rect 28951 22528 30205 22556
rect 28951 22525 28963 22528
rect 28905 22519 28963 22525
rect 30193 22525 30205 22528
rect 30239 22525 30251 22559
rect 30193 22519 30251 22525
rect 31665 22559 31723 22565
rect 31665 22525 31677 22559
rect 31711 22556 31723 22559
rect 32582 22556 32588 22568
rect 31711 22528 32588 22556
rect 31711 22525 31723 22528
rect 31665 22519 31723 22525
rect 32582 22516 32588 22528
rect 32640 22516 32646 22568
rect 34238 22516 34244 22568
rect 34296 22516 34302 22568
rect 39482 22516 39488 22568
rect 39540 22556 39546 22568
rect 39669 22559 39727 22565
rect 39669 22556 39681 22559
rect 39540 22528 39681 22556
rect 39540 22516 39546 22528
rect 39669 22525 39681 22528
rect 39715 22525 39727 22559
rect 39669 22519 39727 22525
rect 29641 22491 29699 22497
rect 29641 22457 29653 22491
rect 29687 22488 29699 22491
rect 34514 22488 34520 22500
rect 29687 22460 34520 22488
rect 29687 22457 29699 22460
rect 29641 22451 29699 22457
rect 34514 22448 34520 22460
rect 34572 22448 34578 22500
rect 27798 22420 27804 22432
rect 27172 22392 27804 22420
rect 27798 22380 27804 22392
rect 27856 22380 27862 22432
rect 32306 22380 32312 22432
rect 32364 22420 32370 22432
rect 33689 22423 33747 22429
rect 33689 22420 33701 22423
rect 32364 22392 33701 22420
rect 32364 22380 32370 22392
rect 33689 22389 33701 22392
rect 33735 22389 33747 22423
rect 33689 22383 33747 22389
rect 1104 22330 49864 22352
rect 1104 22278 2950 22330
rect 3002 22278 3014 22330
rect 3066 22278 3078 22330
rect 3130 22278 3142 22330
rect 3194 22278 3206 22330
rect 3258 22278 12950 22330
rect 13002 22278 13014 22330
rect 13066 22278 13078 22330
rect 13130 22278 13142 22330
rect 13194 22278 13206 22330
rect 13258 22278 22950 22330
rect 23002 22278 23014 22330
rect 23066 22278 23078 22330
rect 23130 22278 23142 22330
rect 23194 22278 23206 22330
rect 23258 22278 32950 22330
rect 33002 22278 33014 22330
rect 33066 22278 33078 22330
rect 33130 22278 33142 22330
rect 33194 22278 33206 22330
rect 33258 22278 42950 22330
rect 43002 22278 43014 22330
rect 43066 22278 43078 22330
rect 43130 22278 43142 22330
rect 43194 22278 43206 22330
rect 43258 22278 49864 22330
rect 1104 22256 49864 22278
rect 12805 22219 12863 22225
rect 12805 22185 12817 22219
rect 12851 22216 12863 22219
rect 14734 22216 14740 22228
rect 12851 22188 14740 22216
rect 12851 22185 12863 22188
rect 12805 22179 12863 22185
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 14994 22219 15052 22225
rect 14994 22216 15006 22219
rect 14844 22188 15006 22216
rect 5534 22108 5540 22160
rect 5592 22108 5598 22160
rect 14550 22108 14556 22160
rect 14608 22148 14614 22160
rect 14844 22148 14872 22188
rect 14994 22185 15006 22188
rect 15040 22185 15052 22219
rect 14994 22179 15052 22185
rect 15102 22176 15108 22228
rect 15160 22216 15166 22228
rect 16482 22216 16488 22228
rect 15160 22188 16488 22216
rect 15160 22176 15166 22188
rect 16482 22176 16488 22188
rect 16540 22176 16546 22228
rect 19692 22219 19750 22225
rect 19692 22185 19704 22219
rect 19738 22216 19750 22219
rect 19738 22188 23244 22216
rect 19738 22185 19750 22188
rect 19692 22179 19750 22185
rect 14608 22120 14872 22148
rect 14608 22108 14614 22120
rect 22554 22108 22560 22160
rect 22612 22148 22618 22160
rect 23216 22148 23244 22188
rect 23290 22176 23296 22228
rect 23348 22176 23354 22228
rect 32122 22216 32128 22228
rect 26252 22188 32128 22216
rect 23566 22148 23572 22160
rect 22612 22120 22692 22148
rect 23216 22120 23572 22148
rect 22612 22108 22618 22120
rect 14737 22083 14795 22089
rect 14737 22049 14749 22083
rect 14783 22080 14795 22083
rect 19426 22080 19432 22092
rect 14783 22052 19432 22080
rect 14783 22049 14795 22052
rect 14737 22043 14795 22049
rect 19426 22040 19432 22052
rect 19484 22040 19490 22092
rect 20162 22040 20168 22092
rect 20220 22080 20226 22092
rect 22664 22089 22692 22120
rect 23566 22108 23572 22120
rect 23624 22108 23630 22160
rect 23768 22120 24440 22148
rect 21177 22083 21235 22089
rect 21177 22080 21189 22083
rect 20220 22052 21189 22080
rect 20220 22040 20226 22052
rect 21177 22049 21189 22052
rect 21223 22049 21235 22083
rect 21177 22043 21235 22049
rect 22649 22083 22707 22089
rect 22649 22049 22661 22083
rect 22695 22049 22707 22083
rect 22649 22043 22707 22049
rect 23290 22040 23296 22092
rect 23348 22080 23354 22092
rect 23474 22080 23480 22092
rect 23348 22052 23480 22080
rect 23348 22040 23354 22052
rect 23474 22040 23480 22052
rect 23532 22040 23538 22092
rect 9122 21972 9128 22024
rect 9180 22012 9186 22024
rect 9180 21984 12434 22012
rect 9180 21972 9186 21984
rect 5353 21947 5411 21953
rect 5353 21913 5365 21947
rect 5399 21944 5411 21947
rect 10226 21944 10232 21956
rect 5399 21916 10232 21944
rect 5399 21913 5411 21916
rect 5353 21907 5411 21913
rect 10226 21904 10232 21916
rect 10284 21904 10290 21956
rect 12406 21944 12434 21984
rect 12526 21972 12532 22024
rect 12584 21972 12590 22024
rect 13630 21972 13636 22024
rect 13688 21972 13694 22024
rect 20990 22012 20996 22024
rect 20838 21984 20996 22012
rect 20990 21972 20996 21984
rect 21048 21972 21054 22024
rect 23768 22012 23796 22120
rect 23937 22083 23995 22089
rect 23937 22049 23949 22083
rect 23983 22080 23995 22083
rect 24302 22080 24308 22092
rect 23983 22052 24308 22080
rect 23983 22049 23995 22052
rect 23937 22043 23995 22049
rect 24302 22040 24308 22052
rect 24360 22040 24366 22092
rect 24412 22080 24440 22120
rect 26252 22089 26280 22188
rect 32122 22176 32128 22188
rect 32180 22176 32186 22228
rect 33410 22176 33416 22228
rect 33468 22176 33474 22228
rect 34238 22176 34244 22228
rect 34296 22216 34302 22228
rect 35602 22219 35660 22225
rect 35602 22216 35614 22219
rect 34296 22188 35614 22216
rect 34296 22176 34302 22188
rect 35602 22185 35614 22188
rect 35648 22185 35660 22219
rect 35602 22179 35660 22185
rect 26602 22108 26608 22160
rect 26660 22148 26666 22160
rect 33428 22148 33456 22176
rect 34330 22148 34336 22160
rect 26660 22120 29040 22148
rect 33428 22120 34336 22148
rect 26660 22108 26666 22120
rect 25133 22083 25191 22089
rect 25133 22080 25145 22083
rect 24412 22052 25145 22080
rect 25133 22049 25145 22052
rect 25179 22080 25191 22083
rect 26237 22083 26295 22089
rect 25179 22052 26096 22080
rect 25179 22049 25191 22052
rect 25133 22043 25191 22049
rect 22066 21984 23796 22012
rect 12406 21916 13584 21944
rect 9306 21836 9312 21888
rect 9364 21876 9370 21888
rect 12989 21879 13047 21885
rect 12989 21876 13001 21879
rect 9364 21848 13001 21876
rect 9364 21836 9370 21848
rect 12989 21845 13001 21848
rect 13035 21845 13047 21879
rect 12989 21839 13047 21845
rect 13446 21836 13452 21888
rect 13504 21836 13510 21888
rect 13556 21876 13584 21916
rect 15470 21904 15476 21956
rect 15528 21904 15534 21956
rect 22066 21944 22094 21984
rect 25958 21972 25964 22024
rect 26016 21972 26022 22024
rect 26068 22021 26096 22052
rect 26237 22049 26249 22083
rect 26283 22080 26295 22083
rect 26283 22052 26317 22080
rect 26283 22049 26295 22052
rect 26237 22043 26295 22049
rect 28534 22040 28540 22092
rect 28592 22080 28598 22092
rect 29012 22089 29040 22120
rect 34330 22108 34336 22120
rect 34388 22108 34394 22160
rect 28905 22083 28963 22089
rect 28905 22080 28917 22083
rect 28592 22052 28917 22080
rect 28592 22040 28598 22052
rect 28905 22049 28917 22052
rect 28951 22049 28963 22083
rect 28905 22043 28963 22049
rect 28997 22083 29055 22089
rect 28997 22049 29009 22083
rect 29043 22049 29055 22083
rect 33870 22080 33876 22092
rect 28997 22043 29055 22049
rect 31726 22052 33876 22080
rect 26053 22015 26111 22021
rect 26053 21981 26065 22015
rect 26099 22012 26111 22015
rect 26099 21984 28948 22012
rect 26099 21981 26111 21984
rect 26053 21975 26111 21981
rect 21008 21916 22094 21944
rect 23661 21947 23719 21953
rect 21008 21876 21036 21916
rect 23661 21913 23673 21947
rect 23707 21944 23719 21947
rect 23842 21944 23848 21956
rect 23707 21916 23848 21944
rect 23707 21913 23719 21916
rect 23661 21907 23719 21913
rect 23842 21904 23848 21916
rect 23900 21904 23906 21956
rect 26694 21944 26700 21956
rect 24964 21916 26700 21944
rect 13556 21848 21036 21876
rect 22094 21836 22100 21888
rect 22152 21836 22158 21888
rect 22462 21836 22468 21888
rect 22520 21836 22526 21888
rect 22557 21879 22615 21885
rect 22557 21845 22569 21879
rect 22603 21876 22615 21879
rect 23566 21876 23572 21888
rect 22603 21848 23572 21876
rect 22603 21845 22615 21848
rect 22557 21839 22615 21845
rect 23566 21836 23572 21848
rect 23624 21836 23630 21888
rect 23753 21879 23811 21885
rect 23753 21845 23765 21879
rect 23799 21876 23811 21879
rect 24964 21876 24992 21916
rect 26694 21904 26700 21916
rect 26752 21904 26758 21956
rect 23799 21848 24992 21876
rect 23799 21845 23811 21848
rect 23753 21839 23811 21845
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 27522 21836 27528 21888
rect 27580 21876 27586 21888
rect 28445 21879 28503 21885
rect 28445 21876 28457 21879
rect 27580 21848 28457 21876
rect 27580 21836 27586 21848
rect 28445 21845 28457 21848
rect 28491 21845 28503 21879
rect 28445 21839 28503 21845
rect 28810 21836 28816 21888
rect 28868 21836 28874 21888
rect 28920 21876 28948 21984
rect 29362 21972 29368 22024
rect 29420 22012 29426 22024
rect 29917 22015 29975 22021
rect 29917 22012 29929 22015
rect 29420 21984 29929 22012
rect 29420 21972 29426 21984
rect 29917 21981 29929 21984
rect 29963 21981 29975 22015
rect 31726 22012 31754 22052
rect 33870 22040 33876 22052
rect 33928 22040 33934 22092
rect 37093 22083 37151 22089
rect 37093 22049 37105 22083
rect 37139 22080 37151 22083
rect 37274 22080 37280 22092
rect 37139 22052 37280 22080
rect 37139 22049 37151 22052
rect 37093 22043 37151 22049
rect 37274 22040 37280 22052
rect 37332 22040 37338 22092
rect 29917 21975 29975 21981
rect 30852 21984 31754 22012
rect 30852 21876 30880 21984
rect 32490 21972 32496 22024
rect 32548 22012 32554 22024
rect 35345 22015 35403 22021
rect 35345 22012 35357 22015
rect 32548 21984 35357 22012
rect 32548 21972 32554 21984
rect 35345 21981 35357 21984
rect 35391 21981 35403 22015
rect 35345 21975 35403 21981
rect 37829 22015 37887 22021
rect 37829 21981 37841 22015
rect 37875 21981 37887 22015
rect 37829 21975 37887 21981
rect 36078 21904 36084 21956
rect 36136 21904 36142 21956
rect 37844 21944 37872 21975
rect 47578 21972 47584 22024
rect 47636 22012 47642 22024
rect 47949 22015 48007 22021
rect 47949 22012 47961 22015
rect 47636 21984 47961 22012
rect 47636 21972 47642 21984
rect 47949 21981 47961 21984
rect 47995 21981 48007 22015
rect 47949 21975 48007 21981
rect 49142 21972 49148 22024
rect 49200 21972 49206 22024
rect 36924 21916 37872 21944
rect 28920 21848 30880 21876
rect 31662 21836 31668 21888
rect 31720 21876 31726 21888
rect 36924 21876 36952 21916
rect 38470 21904 38476 21956
rect 38528 21944 38534 21956
rect 43806 21944 43812 21956
rect 38528 21916 43812 21944
rect 38528 21904 38534 21916
rect 43806 21904 43812 21916
rect 43864 21904 43870 21956
rect 31720 21848 36952 21876
rect 37645 21879 37703 21885
rect 31720 21836 31726 21848
rect 37645 21845 37657 21879
rect 37691 21876 37703 21879
rect 41322 21876 41328 21888
rect 37691 21848 41328 21876
rect 37691 21845 37703 21848
rect 37645 21839 37703 21845
rect 41322 21836 41328 21848
rect 41380 21836 41386 21888
rect 1104 21786 49864 21808
rect 1104 21734 7950 21786
rect 8002 21734 8014 21786
rect 8066 21734 8078 21786
rect 8130 21734 8142 21786
rect 8194 21734 8206 21786
rect 8258 21734 17950 21786
rect 18002 21734 18014 21786
rect 18066 21734 18078 21786
rect 18130 21734 18142 21786
rect 18194 21734 18206 21786
rect 18258 21734 27950 21786
rect 28002 21734 28014 21786
rect 28066 21734 28078 21786
rect 28130 21734 28142 21786
rect 28194 21734 28206 21786
rect 28258 21734 37950 21786
rect 38002 21734 38014 21786
rect 38066 21734 38078 21786
rect 38130 21734 38142 21786
rect 38194 21734 38206 21786
rect 38258 21734 47950 21786
rect 48002 21734 48014 21786
rect 48066 21734 48078 21786
rect 48130 21734 48142 21786
rect 48194 21734 48206 21786
rect 48258 21734 49864 21786
rect 1104 21712 49864 21734
rect 10226 21632 10232 21684
rect 10284 21632 10290 21684
rect 13630 21632 13636 21684
rect 13688 21672 13694 21684
rect 17402 21672 17408 21684
rect 13688 21644 17408 21672
rect 13688 21632 13694 21644
rect 17402 21632 17408 21644
rect 17460 21632 17466 21684
rect 19429 21675 19487 21681
rect 19429 21641 19441 21675
rect 19475 21672 19487 21675
rect 19794 21672 19800 21684
rect 19475 21644 19800 21672
rect 19475 21641 19487 21644
rect 19429 21635 19487 21641
rect 19794 21632 19800 21644
rect 19852 21632 19858 21684
rect 20717 21675 20775 21681
rect 20717 21641 20729 21675
rect 20763 21672 20775 21675
rect 21174 21672 21180 21684
rect 20763 21644 21180 21672
rect 20763 21641 20775 21644
rect 20717 21635 20775 21641
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 22462 21632 22468 21684
rect 22520 21672 22526 21684
rect 25133 21675 25191 21681
rect 25133 21672 25145 21675
rect 22520 21644 25145 21672
rect 22520 21632 22526 21644
rect 25133 21641 25145 21644
rect 25179 21641 25191 21675
rect 25133 21635 25191 21641
rect 25501 21675 25559 21681
rect 25501 21641 25513 21675
rect 25547 21672 25559 21675
rect 25866 21672 25872 21684
rect 25547 21644 25872 21672
rect 25547 21641 25559 21644
rect 25501 21635 25559 21641
rect 25866 21632 25872 21644
rect 25924 21632 25930 21684
rect 28997 21675 29055 21681
rect 28997 21641 29009 21675
rect 29043 21672 29055 21675
rect 29362 21672 29368 21684
rect 29043 21644 29368 21672
rect 29043 21641 29055 21644
rect 28997 21635 29055 21641
rect 29362 21632 29368 21644
rect 29420 21632 29426 21684
rect 32490 21672 32496 21684
rect 29840 21644 32496 21672
rect 21726 21604 21732 21616
rect 21100 21576 21732 21604
rect 21100 21548 21128 21576
rect 21726 21564 21732 21576
rect 21784 21564 21790 21616
rect 22094 21564 22100 21616
rect 22152 21604 22158 21616
rect 22741 21607 22799 21613
rect 22741 21604 22753 21607
rect 22152 21576 22753 21604
rect 22152 21564 22158 21576
rect 22741 21573 22753 21576
rect 22787 21604 22799 21607
rect 22830 21604 22836 21616
rect 22787 21576 22836 21604
rect 22787 21573 22799 21576
rect 22741 21567 22799 21573
rect 22830 21564 22836 21576
rect 22888 21564 22894 21616
rect 23290 21564 23296 21616
rect 23348 21564 23354 21616
rect 25590 21564 25596 21616
rect 25648 21604 25654 21616
rect 25648 21576 29132 21604
rect 25648 21564 25654 21576
rect 9585 21539 9643 21545
rect 9585 21505 9597 21539
rect 9631 21536 9643 21539
rect 13446 21536 13452 21548
rect 9631 21508 13452 21536
rect 9631 21505 9643 21508
rect 9585 21499 9643 21505
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 14461 21539 14519 21545
rect 14461 21505 14473 21539
rect 14507 21536 14519 21539
rect 16482 21536 16488 21548
rect 14507 21508 16488 21536
rect 14507 21505 14519 21508
rect 14461 21499 14519 21505
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 19518 21496 19524 21548
rect 19576 21536 19582 21548
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19576 21508 19809 21536
rect 19576 21496 19582 21508
rect 19797 21505 19809 21508
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 21082 21496 21088 21548
rect 21140 21496 21146 21548
rect 21177 21539 21235 21545
rect 21177 21505 21189 21539
rect 21223 21536 21235 21539
rect 22370 21536 22376 21548
rect 21223 21508 22376 21536
rect 21223 21505 21235 21508
rect 21177 21499 21235 21505
rect 22370 21496 22376 21508
rect 22428 21496 22434 21548
rect 28166 21496 28172 21548
rect 28224 21496 28230 21548
rect 29104 21545 29132 21576
rect 29840 21545 29868 21644
rect 32490 21632 32496 21644
rect 32548 21632 32554 21684
rect 34238 21632 34244 21684
rect 34296 21632 34302 21684
rect 37826 21632 37832 21684
rect 37884 21672 37890 21684
rect 40221 21675 40279 21681
rect 40221 21672 40233 21675
rect 37884 21644 40233 21672
rect 37884 21632 37890 21644
rect 40221 21641 40233 21644
rect 40267 21641 40279 21675
rect 40221 21635 40279 21641
rect 31570 21604 31576 21616
rect 31326 21576 31576 21604
rect 31570 21564 31576 21576
rect 31628 21564 31634 21616
rect 34422 21604 34428 21616
rect 33994 21576 34428 21604
rect 34422 21564 34428 21576
rect 34480 21604 34486 21616
rect 36078 21604 36084 21616
rect 34480 21576 36084 21604
rect 34480 21564 34486 21576
rect 36078 21564 36084 21576
rect 36136 21564 36142 21616
rect 38746 21564 38752 21616
rect 38804 21564 38810 21616
rect 39022 21564 39028 21616
rect 39080 21604 39086 21616
rect 39080 21576 39238 21604
rect 39080 21564 39086 21576
rect 43806 21564 43812 21616
rect 43864 21564 43870 21616
rect 29089 21539 29147 21545
rect 29089 21505 29101 21539
rect 29135 21505 29147 21539
rect 29825 21539 29883 21545
rect 29825 21536 29837 21539
rect 29089 21499 29147 21505
rect 29196 21508 29837 21536
rect 9766 21428 9772 21480
rect 9824 21428 9830 21480
rect 19886 21428 19892 21480
rect 19944 21428 19950 21480
rect 19978 21428 19984 21480
rect 20036 21468 20042 21480
rect 20073 21471 20131 21477
rect 20073 21468 20085 21471
rect 20036 21440 20085 21468
rect 20036 21428 20042 21440
rect 20073 21437 20085 21440
rect 20119 21437 20131 21471
rect 20073 21431 20131 21437
rect 12250 21360 12256 21412
rect 12308 21400 12314 21412
rect 14277 21403 14335 21409
rect 14277 21400 14289 21403
rect 12308 21372 14289 21400
rect 12308 21360 12314 21372
rect 14277 21369 14289 21372
rect 14323 21369 14335 21403
rect 20088 21400 20116 21431
rect 21358 21428 21364 21480
rect 21416 21428 21422 21480
rect 22462 21428 22468 21480
rect 22520 21428 22526 21480
rect 25593 21471 25651 21477
rect 25593 21437 25605 21471
rect 25639 21437 25651 21471
rect 25593 21431 25651 21437
rect 25608 21400 25636 21431
rect 25682 21428 25688 21480
rect 25740 21428 25746 21480
rect 27798 21428 27804 21480
rect 27856 21468 27862 21480
rect 29196 21468 29224 21508
rect 29825 21505 29837 21508
rect 29871 21505 29883 21539
rect 31846 21536 31852 21548
rect 29825 21499 29883 21505
rect 31312 21508 31852 21536
rect 27856 21440 29224 21468
rect 29273 21471 29331 21477
rect 27856 21428 27862 21440
rect 29273 21437 29285 21471
rect 29319 21468 29331 21471
rect 30101 21471 30159 21477
rect 30101 21468 30113 21471
rect 29319 21440 30113 21468
rect 29319 21437 29331 21440
rect 29273 21431 29331 21437
rect 30101 21437 30113 21440
rect 30147 21468 30159 21471
rect 31312 21468 31340 21508
rect 31846 21496 31852 21508
rect 31904 21496 31910 21548
rect 32490 21496 32496 21548
rect 32548 21496 32554 21548
rect 35342 21496 35348 21548
rect 35400 21496 35406 21548
rect 35986 21496 35992 21548
rect 36044 21496 36050 21548
rect 38470 21496 38476 21548
rect 38528 21496 38534 21548
rect 46198 21496 46204 21548
rect 46256 21536 46262 21548
rect 47949 21539 48007 21545
rect 47949 21536 47961 21539
rect 46256 21508 47961 21536
rect 46256 21496 46262 21508
rect 47949 21505 47961 21508
rect 47995 21505 48007 21539
rect 47949 21499 48007 21505
rect 30147 21440 31340 21468
rect 31573 21471 31631 21477
rect 30147 21437 30159 21440
rect 30101 21431 30159 21437
rect 31573 21437 31585 21471
rect 31619 21468 31631 21471
rect 31754 21468 31760 21480
rect 31619 21440 31760 21468
rect 31619 21437 31631 21440
rect 31573 21431 31631 21437
rect 31754 21428 31760 21440
rect 31812 21428 31818 21480
rect 32214 21428 32220 21480
rect 32272 21468 32278 21480
rect 32769 21471 32827 21477
rect 32769 21468 32781 21471
rect 32272 21440 32781 21468
rect 32272 21428 32278 21440
rect 32769 21437 32781 21440
rect 32815 21468 32827 21471
rect 34054 21468 34060 21480
rect 32815 21440 34060 21468
rect 32815 21437 32827 21440
rect 32769 21431 32827 21437
rect 34054 21428 34060 21440
rect 34112 21428 34118 21480
rect 49142 21428 49148 21480
rect 49200 21428 49206 21480
rect 27430 21400 27436 21412
rect 20088 21372 22094 21400
rect 25608 21372 27436 21400
rect 14277 21363 14335 21369
rect 22066 21332 22094 21372
rect 27430 21360 27436 21372
rect 27488 21360 27494 21412
rect 27985 21403 28043 21409
rect 27985 21369 27997 21403
rect 28031 21400 28043 21403
rect 28902 21400 28908 21412
rect 28031 21372 28908 21400
rect 28031 21369 28043 21372
rect 27985 21363 28043 21369
rect 28902 21360 28908 21372
rect 28960 21360 28966 21412
rect 35161 21403 35219 21409
rect 35161 21369 35173 21403
rect 35207 21400 35219 21403
rect 43993 21403 44051 21409
rect 35207 21372 38608 21400
rect 35207 21369 35219 21372
rect 35161 21363 35219 21369
rect 38580 21344 38608 21372
rect 43993 21369 44005 21403
rect 44039 21400 44051 21403
rect 45094 21400 45100 21412
rect 44039 21372 45100 21400
rect 44039 21369 44051 21372
rect 43993 21363 44051 21369
rect 45094 21360 45100 21372
rect 45152 21360 45158 21412
rect 24213 21335 24271 21341
rect 24213 21332 24225 21335
rect 22066 21304 24225 21332
rect 24213 21301 24225 21304
rect 24259 21332 24271 21335
rect 24302 21332 24308 21344
rect 24259 21304 24308 21332
rect 24259 21301 24271 21304
rect 24213 21295 24271 21301
rect 24302 21292 24308 21304
rect 24360 21292 24366 21344
rect 28629 21335 28687 21341
rect 28629 21301 28641 21335
rect 28675 21332 28687 21335
rect 30650 21332 30656 21344
rect 28675 21304 30656 21332
rect 28675 21301 28687 21304
rect 28629 21295 28687 21301
rect 30650 21292 30656 21304
rect 30708 21292 30714 21344
rect 33502 21292 33508 21344
rect 33560 21332 33566 21344
rect 35434 21332 35440 21344
rect 33560 21304 35440 21332
rect 33560 21292 33566 21304
rect 35434 21292 35440 21304
rect 35492 21292 35498 21344
rect 35805 21335 35863 21341
rect 35805 21301 35817 21335
rect 35851 21332 35863 21335
rect 37090 21332 37096 21344
rect 35851 21304 37096 21332
rect 35851 21301 35863 21304
rect 35805 21295 35863 21301
rect 37090 21292 37096 21304
rect 37148 21292 37154 21344
rect 38562 21292 38568 21344
rect 38620 21292 38626 21344
rect 1104 21242 49864 21264
rect 1104 21190 2950 21242
rect 3002 21190 3014 21242
rect 3066 21190 3078 21242
rect 3130 21190 3142 21242
rect 3194 21190 3206 21242
rect 3258 21190 12950 21242
rect 13002 21190 13014 21242
rect 13066 21190 13078 21242
rect 13130 21190 13142 21242
rect 13194 21190 13206 21242
rect 13258 21190 22950 21242
rect 23002 21190 23014 21242
rect 23066 21190 23078 21242
rect 23130 21190 23142 21242
rect 23194 21190 23206 21242
rect 23258 21190 32950 21242
rect 33002 21190 33014 21242
rect 33066 21190 33078 21242
rect 33130 21190 33142 21242
rect 33194 21190 33206 21242
rect 33258 21190 42950 21242
rect 43002 21190 43014 21242
rect 43066 21190 43078 21242
rect 43130 21190 43142 21242
rect 43194 21190 43206 21242
rect 43258 21190 49864 21242
rect 1104 21168 49864 21190
rect 9674 21088 9680 21140
rect 9732 21088 9738 21140
rect 28166 21088 28172 21140
rect 28224 21128 28230 21140
rect 30742 21128 30748 21140
rect 28224 21100 30748 21128
rect 28224 21088 28230 21100
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 27338 21020 27344 21072
rect 27396 21060 27402 21072
rect 35342 21060 35348 21072
rect 27396 21032 35348 21060
rect 27396 21020 27402 21032
rect 35342 21020 35348 21032
rect 35400 21020 35406 21072
rect 36633 21063 36691 21069
rect 36633 21029 36645 21063
rect 36679 21060 36691 21063
rect 43714 21060 43720 21072
rect 36679 21032 43720 21060
rect 36679 21029 36691 21032
rect 36633 21023 36691 21029
rect 43714 21020 43720 21032
rect 43772 21020 43778 21072
rect 9125 20995 9183 21001
rect 9125 20961 9137 20995
rect 9171 20992 9183 20995
rect 10962 20992 10968 21004
rect 9171 20964 10968 20992
rect 9171 20961 9183 20964
rect 9125 20955 9183 20961
rect 10962 20952 10968 20964
rect 11020 20952 11026 21004
rect 30929 20995 30987 21001
rect 30929 20961 30941 20995
rect 30975 20992 30987 20995
rect 31754 20992 31760 21004
rect 30975 20964 31760 20992
rect 30975 20961 30987 20964
rect 30929 20955 30987 20961
rect 31754 20952 31760 20964
rect 31812 20952 31818 21004
rect 32858 20952 32864 21004
rect 32916 20992 32922 21004
rect 32916 20964 36860 20992
rect 32916 20952 32922 20964
rect 4157 20927 4215 20933
rect 4157 20893 4169 20927
rect 4203 20924 4215 20927
rect 7834 20924 7840 20936
rect 4203 20896 7840 20924
rect 4203 20893 4215 20896
rect 4157 20887 4215 20893
rect 7834 20884 7840 20896
rect 7892 20884 7898 20936
rect 9306 20884 9312 20936
rect 9364 20884 9370 20936
rect 30650 20884 30656 20936
rect 30708 20884 30714 20936
rect 30742 20884 30748 20936
rect 30800 20924 30806 20936
rect 31665 20927 31723 20933
rect 31665 20924 31677 20927
rect 30800 20896 31677 20924
rect 30800 20884 30806 20896
rect 31665 20893 31677 20896
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 32309 20927 32367 20933
rect 32309 20893 32321 20927
rect 32355 20924 32367 20927
rect 35066 20924 35072 20936
rect 32355 20896 35072 20924
rect 32355 20893 32367 20896
rect 32309 20887 32367 20893
rect 35066 20884 35072 20896
rect 35124 20884 35130 20936
rect 36832 20933 36860 20964
rect 37826 20952 37832 21004
rect 37884 20992 37890 21004
rect 38381 20995 38439 21001
rect 38381 20992 38393 20995
rect 37884 20964 38393 20992
rect 37884 20952 37890 20964
rect 38381 20961 38393 20964
rect 38427 20961 38439 20995
rect 38381 20955 38439 20961
rect 36817 20927 36875 20933
rect 36817 20893 36829 20927
rect 36863 20893 36875 20927
rect 36817 20887 36875 20893
rect 38197 20927 38255 20933
rect 38197 20893 38209 20927
rect 38243 20924 38255 20927
rect 38286 20924 38292 20936
rect 38243 20896 38292 20924
rect 38243 20893 38255 20896
rect 38197 20887 38255 20893
rect 38286 20884 38292 20896
rect 38344 20884 38350 20936
rect 46934 20884 46940 20936
rect 46992 20924 46998 20936
rect 47949 20927 48007 20933
rect 47949 20924 47961 20927
rect 46992 20896 47961 20924
rect 46992 20884 46998 20896
rect 47949 20893 47961 20896
rect 47995 20893 48007 20927
rect 47949 20887 48007 20893
rect 28810 20816 28816 20868
rect 28868 20856 28874 20868
rect 36170 20856 36176 20868
rect 28868 20828 36176 20856
rect 28868 20816 28874 20828
rect 36170 20816 36176 20828
rect 36228 20816 36234 20868
rect 36354 20816 36360 20868
rect 36412 20856 36418 20868
rect 36412 20828 36768 20856
rect 36412 20816 36418 20828
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 4249 20791 4307 20797
rect 4249 20788 4261 20791
rect 2924 20760 4261 20788
rect 2924 20748 2930 20760
rect 4249 20757 4261 20760
rect 4295 20757 4307 20791
rect 4249 20751 4307 20757
rect 30282 20748 30288 20800
rect 30340 20748 30346 20800
rect 30745 20791 30803 20797
rect 30745 20757 30757 20791
rect 30791 20788 30803 20791
rect 31294 20788 31300 20800
rect 30791 20760 31300 20788
rect 30791 20757 30803 20760
rect 30745 20751 30803 20757
rect 31294 20748 31300 20760
rect 31352 20748 31358 20800
rect 31938 20748 31944 20800
rect 31996 20788 32002 20800
rect 32125 20791 32183 20797
rect 32125 20788 32137 20791
rect 31996 20760 32137 20788
rect 31996 20748 32002 20760
rect 32125 20757 32137 20760
rect 32171 20757 32183 20791
rect 36188 20788 36216 20816
rect 36538 20788 36544 20800
rect 36188 20760 36544 20788
rect 32125 20751 32183 20757
rect 36538 20748 36544 20760
rect 36596 20748 36602 20800
rect 36740 20788 36768 20828
rect 37642 20816 37648 20868
rect 37700 20856 37706 20868
rect 37700 20828 38332 20856
rect 37700 20816 37706 20828
rect 38304 20797 38332 20828
rect 49142 20816 49148 20868
rect 49200 20816 49206 20868
rect 37829 20791 37887 20797
rect 37829 20788 37841 20791
rect 36740 20760 37841 20788
rect 37829 20757 37841 20760
rect 37875 20757 37887 20791
rect 37829 20751 37887 20757
rect 38289 20791 38347 20797
rect 38289 20757 38301 20791
rect 38335 20757 38347 20791
rect 38289 20751 38347 20757
rect 1104 20698 49864 20720
rect 1104 20646 7950 20698
rect 8002 20646 8014 20698
rect 8066 20646 8078 20698
rect 8130 20646 8142 20698
rect 8194 20646 8206 20698
rect 8258 20646 17950 20698
rect 18002 20646 18014 20698
rect 18066 20646 18078 20698
rect 18130 20646 18142 20698
rect 18194 20646 18206 20698
rect 18258 20646 27950 20698
rect 28002 20646 28014 20698
rect 28066 20646 28078 20698
rect 28130 20646 28142 20698
rect 28194 20646 28206 20698
rect 28258 20646 37950 20698
rect 38002 20646 38014 20698
rect 38066 20646 38078 20698
rect 38130 20646 38142 20698
rect 38194 20646 38206 20698
rect 38258 20646 47950 20698
rect 48002 20646 48014 20698
rect 48066 20646 48078 20698
rect 48130 20646 48142 20698
rect 48194 20646 48206 20698
rect 48258 20646 49864 20698
rect 1104 20624 49864 20646
rect 21177 20587 21235 20593
rect 21177 20553 21189 20587
rect 21223 20584 21235 20587
rect 21634 20584 21640 20596
rect 21223 20556 21640 20584
rect 21223 20553 21235 20556
rect 21177 20547 21235 20553
rect 21634 20544 21640 20556
rect 21692 20544 21698 20596
rect 21818 20544 21824 20596
rect 21876 20584 21882 20596
rect 22462 20584 22468 20596
rect 21876 20556 22468 20584
rect 21876 20544 21882 20556
rect 22462 20544 22468 20556
rect 22520 20584 22526 20596
rect 24670 20584 24676 20596
rect 22520 20556 23060 20584
rect 22520 20544 22526 20556
rect 21358 20476 21364 20528
rect 21416 20516 21422 20528
rect 21416 20488 22968 20516
rect 21416 20476 21422 20488
rect 1765 20451 1823 20457
rect 1765 20417 1777 20451
rect 1811 20448 1823 20451
rect 2774 20448 2780 20460
rect 1811 20420 2780 20448
rect 1811 20417 1823 20420
rect 1765 20411 1823 20417
rect 2774 20408 2780 20420
rect 2832 20408 2838 20460
rect 20806 20408 20812 20460
rect 20864 20448 20870 20460
rect 21085 20451 21143 20457
rect 21085 20448 21097 20451
rect 20864 20420 21097 20448
rect 20864 20408 20870 20420
rect 21085 20417 21097 20420
rect 21131 20448 21143 20451
rect 22278 20448 22284 20460
rect 21131 20420 22284 20448
rect 21131 20417 21143 20420
rect 21085 20411 21143 20417
rect 22278 20408 22284 20420
rect 22336 20408 22342 20460
rect 1302 20340 1308 20392
rect 1360 20380 1366 20392
rect 2041 20383 2099 20389
rect 2041 20380 2053 20383
rect 1360 20352 2053 20380
rect 1360 20340 1366 20352
rect 2041 20349 2053 20352
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21726 20380 21732 20392
rect 21407 20352 21732 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 21726 20340 21732 20352
rect 21784 20340 21790 20392
rect 19794 20204 19800 20256
rect 19852 20244 19858 20256
rect 20717 20247 20775 20253
rect 20717 20244 20729 20247
rect 19852 20216 20729 20244
rect 19852 20204 19858 20216
rect 20717 20213 20729 20216
rect 20763 20213 20775 20247
rect 22940 20244 22968 20488
rect 23032 20457 23060 20556
rect 23676 20556 24676 20584
rect 23290 20476 23296 20528
rect 23348 20516 23354 20528
rect 23676 20516 23704 20556
rect 24670 20544 24676 20556
rect 24728 20544 24734 20596
rect 26142 20544 26148 20596
rect 26200 20584 26206 20596
rect 26237 20587 26295 20593
rect 26237 20584 26249 20587
rect 26200 20556 26249 20584
rect 26200 20544 26206 20556
rect 26237 20553 26249 20556
rect 26283 20553 26295 20587
rect 26237 20547 26295 20553
rect 30009 20587 30067 20593
rect 30009 20553 30021 20587
rect 30055 20553 30067 20587
rect 30009 20547 30067 20553
rect 23348 20488 23782 20516
rect 23348 20476 23354 20488
rect 23017 20451 23075 20457
rect 23017 20417 23029 20451
rect 23063 20417 23075 20451
rect 23017 20411 23075 20417
rect 26145 20451 26203 20457
rect 26145 20417 26157 20451
rect 26191 20448 26203 20451
rect 27154 20448 27160 20460
rect 26191 20420 27160 20448
rect 26191 20417 26203 20420
rect 26145 20411 26203 20417
rect 27154 20408 27160 20420
rect 27212 20408 27218 20460
rect 30024 20448 30052 20547
rect 30466 20544 30472 20596
rect 30524 20544 30530 20596
rect 32858 20544 32864 20596
rect 32916 20544 32922 20596
rect 30377 20519 30435 20525
rect 30377 20485 30389 20519
rect 30423 20516 30435 20519
rect 30742 20516 30748 20528
rect 30423 20488 30748 20516
rect 30423 20485 30435 20488
rect 30377 20479 30435 20485
rect 30742 20476 30748 20488
rect 30800 20476 30806 20528
rect 32769 20519 32827 20525
rect 32769 20516 32781 20519
rect 31726 20488 32781 20516
rect 31726 20448 31754 20488
rect 32769 20485 32781 20488
rect 32815 20485 32827 20519
rect 32769 20479 32827 20485
rect 30024 20420 31754 20448
rect 34514 20408 34520 20460
rect 34572 20448 34578 20460
rect 36909 20451 36967 20457
rect 36909 20448 36921 20451
rect 34572 20420 36921 20448
rect 34572 20408 34578 20420
rect 36909 20417 36921 20420
rect 36955 20417 36967 20451
rect 36909 20411 36967 20417
rect 47854 20408 47860 20460
rect 47912 20448 47918 20460
rect 47949 20451 48007 20457
rect 47949 20448 47961 20451
rect 47912 20420 47961 20448
rect 47912 20408 47918 20420
rect 47949 20417 47961 20420
rect 47995 20417 48007 20451
rect 47949 20411 48007 20417
rect 23290 20340 23296 20392
rect 23348 20340 23354 20392
rect 25130 20340 25136 20392
rect 25188 20380 25194 20392
rect 26421 20383 26479 20389
rect 26421 20380 26433 20383
rect 25188 20352 26433 20380
rect 25188 20340 25194 20352
rect 26421 20349 26433 20352
rect 26467 20380 26479 20383
rect 26602 20380 26608 20392
rect 26467 20352 26608 20380
rect 26467 20349 26479 20352
rect 26421 20343 26479 20349
rect 26602 20340 26608 20352
rect 26660 20340 26666 20392
rect 30653 20383 30711 20389
rect 30653 20349 30665 20383
rect 30699 20380 30711 20383
rect 32214 20380 32220 20392
rect 30699 20352 32220 20380
rect 30699 20349 30711 20352
rect 30653 20343 30711 20349
rect 32214 20340 32220 20352
rect 32272 20340 32278 20392
rect 33045 20383 33103 20389
rect 33045 20349 33057 20383
rect 33091 20380 33103 20383
rect 34238 20380 34244 20392
rect 33091 20352 34244 20380
rect 33091 20349 33103 20352
rect 33045 20343 33103 20349
rect 34238 20340 34244 20352
rect 34296 20340 34302 20392
rect 49142 20340 49148 20392
rect 49200 20340 49206 20392
rect 24765 20247 24823 20253
rect 24765 20244 24777 20247
rect 22940 20216 24777 20244
rect 20717 20207 20775 20213
rect 24765 20213 24777 20216
rect 24811 20244 24823 20247
rect 25682 20244 25688 20256
rect 24811 20216 25688 20244
rect 24811 20213 24823 20216
rect 24765 20207 24823 20213
rect 25682 20204 25688 20216
rect 25740 20204 25746 20256
rect 25774 20204 25780 20256
rect 25832 20204 25838 20256
rect 32401 20247 32459 20253
rect 32401 20213 32413 20247
rect 32447 20244 32459 20247
rect 32490 20244 32496 20256
rect 32447 20216 32496 20244
rect 32447 20213 32459 20216
rect 32401 20207 32459 20213
rect 32490 20204 32496 20216
rect 32548 20204 32554 20256
rect 36725 20247 36783 20253
rect 36725 20213 36737 20247
rect 36771 20244 36783 20247
rect 39942 20244 39948 20256
rect 36771 20216 39948 20244
rect 36771 20213 36783 20216
rect 36725 20207 36783 20213
rect 39942 20204 39948 20216
rect 40000 20204 40006 20256
rect 1104 20154 49864 20176
rect 1104 20102 2950 20154
rect 3002 20102 3014 20154
rect 3066 20102 3078 20154
rect 3130 20102 3142 20154
rect 3194 20102 3206 20154
rect 3258 20102 12950 20154
rect 13002 20102 13014 20154
rect 13066 20102 13078 20154
rect 13130 20102 13142 20154
rect 13194 20102 13206 20154
rect 13258 20102 22950 20154
rect 23002 20102 23014 20154
rect 23066 20102 23078 20154
rect 23130 20102 23142 20154
rect 23194 20102 23206 20154
rect 23258 20102 32950 20154
rect 33002 20102 33014 20154
rect 33066 20102 33078 20154
rect 33130 20102 33142 20154
rect 33194 20102 33206 20154
rect 33258 20102 42950 20154
rect 43002 20102 43014 20154
rect 43066 20102 43078 20154
rect 43130 20102 43142 20154
rect 43194 20102 43206 20154
rect 43258 20102 49864 20154
rect 1104 20080 49864 20102
rect 10962 20000 10968 20052
rect 11020 20040 11026 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 11020 20012 14289 20040
rect 11020 20000 11026 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 19876 20043 19934 20049
rect 19876 20009 19888 20043
rect 19922 20040 19934 20043
rect 19922 20012 23152 20040
rect 19922 20009 19934 20012
rect 19876 20003 19934 20009
rect 18141 19975 18199 19981
rect 18141 19941 18153 19975
rect 18187 19972 18199 19975
rect 19334 19972 19340 19984
rect 18187 19944 19340 19972
rect 18187 19941 18199 19944
rect 18141 19935 18199 19941
rect 19334 19932 19340 19944
rect 19392 19932 19398 19984
rect 21361 19975 21419 19981
rect 21361 19941 21373 19975
rect 21407 19972 21419 19975
rect 21542 19972 21548 19984
rect 21407 19944 21548 19972
rect 21407 19941 21419 19944
rect 21361 19935 21419 19941
rect 21542 19932 21548 19944
rect 21600 19932 21606 19984
rect 18785 19907 18843 19913
rect 18785 19873 18797 19907
rect 18831 19873 18843 19907
rect 18785 19867 18843 19873
rect 14461 19839 14519 19845
rect 14461 19805 14473 19839
rect 14507 19836 14519 19839
rect 17862 19836 17868 19848
rect 14507 19808 17868 19836
rect 14507 19805 14519 19808
rect 14461 19799 14519 19805
rect 17862 19796 17868 19808
rect 17920 19796 17926 19848
rect 18800 19768 18828 19867
rect 19426 19864 19432 19916
rect 19484 19904 19490 19916
rect 19613 19907 19671 19913
rect 19613 19904 19625 19907
rect 19484 19876 19625 19904
rect 19484 19864 19490 19876
rect 19613 19873 19625 19876
rect 19659 19904 19671 19907
rect 21818 19904 21824 19916
rect 19659 19876 21824 19904
rect 19659 19873 19671 19876
rect 19613 19867 19671 19873
rect 21818 19864 21824 19876
rect 21876 19864 21882 19916
rect 22097 19907 22155 19913
rect 22097 19873 22109 19907
rect 22143 19904 22155 19907
rect 22462 19904 22468 19916
rect 22143 19876 22468 19904
rect 22143 19873 22155 19876
rect 22097 19867 22155 19873
rect 22462 19864 22468 19876
rect 22520 19904 22526 19916
rect 22738 19904 22744 19916
rect 22520 19876 22744 19904
rect 22520 19864 22526 19876
rect 22738 19864 22744 19876
rect 22796 19864 22802 19916
rect 23124 19904 23152 20012
rect 23566 20000 23572 20052
rect 23624 20040 23630 20052
rect 25225 20043 25283 20049
rect 25225 20040 25237 20043
rect 23624 20012 25237 20040
rect 23624 20000 23630 20012
rect 25225 20009 25237 20012
rect 25271 20009 25283 20043
rect 25225 20003 25283 20009
rect 26694 20000 26700 20052
rect 26752 20000 26758 20052
rect 35158 20040 35164 20052
rect 31772 20012 35164 20040
rect 23198 19932 23204 19984
rect 23256 19972 23262 19984
rect 25130 19972 25136 19984
rect 23256 19944 25136 19972
rect 23256 19932 23262 19944
rect 25130 19932 25136 19944
rect 25188 19932 25194 19984
rect 23474 19904 23480 19916
rect 23124 19876 23480 19904
rect 23474 19864 23480 19876
rect 23532 19904 23538 19916
rect 23569 19907 23627 19913
rect 23569 19904 23581 19907
rect 23532 19876 23581 19904
rect 23532 19864 23538 19876
rect 23569 19873 23581 19876
rect 23615 19873 23627 19907
rect 23569 19867 23627 19873
rect 25682 19864 25688 19916
rect 25740 19904 25746 19916
rect 25777 19907 25835 19913
rect 25777 19904 25789 19907
rect 25740 19876 25789 19904
rect 25740 19864 25746 19876
rect 25777 19873 25789 19876
rect 25823 19873 25835 19907
rect 25777 19867 25835 19873
rect 27338 19864 27344 19916
rect 27396 19864 27402 19916
rect 20990 19796 20996 19848
rect 21048 19836 21054 19848
rect 21048 19808 21864 19836
rect 21048 19796 21054 19808
rect 19426 19768 19432 19780
rect 18800 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19768 19490 19780
rect 20162 19768 20168 19780
rect 19484 19740 20168 19768
rect 19484 19728 19490 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 21836 19768 21864 19808
rect 23842 19796 23848 19848
rect 23900 19836 23906 19848
rect 28902 19836 28908 19848
rect 23900 19808 28908 19836
rect 23900 19796 23906 19808
rect 28902 19796 28908 19808
rect 28960 19796 28966 19848
rect 22554 19768 22560 19780
rect 21284 19740 21496 19768
rect 21836 19740 22560 19768
rect 18414 19660 18420 19712
rect 18472 19700 18478 19712
rect 18509 19703 18567 19709
rect 18509 19700 18521 19703
rect 18472 19672 18521 19700
rect 18472 19660 18478 19672
rect 18509 19669 18521 19672
rect 18555 19669 18567 19703
rect 18509 19663 18567 19669
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19700 18659 19703
rect 21284 19700 21312 19740
rect 18647 19672 21312 19700
rect 21468 19700 21496 19740
rect 22554 19728 22560 19740
rect 22612 19728 22618 19780
rect 27065 19771 27123 19777
rect 27065 19737 27077 19771
rect 27111 19768 27123 19771
rect 31772 19768 31800 20012
rect 35158 20000 35164 20012
rect 35216 20040 35222 20052
rect 35216 20012 35894 20040
rect 35216 20000 35222 20012
rect 31846 19932 31852 19984
rect 31904 19972 31910 19984
rect 35621 19975 35679 19981
rect 35621 19972 35633 19975
rect 31904 19944 35633 19972
rect 31904 19932 31910 19944
rect 35621 19941 35633 19944
rect 35667 19941 35679 19975
rect 35621 19935 35679 19941
rect 32030 19864 32036 19916
rect 32088 19904 32094 19916
rect 35434 19904 35440 19916
rect 32088 19876 35440 19904
rect 32088 19864 32094 19876
rect 35434 19864 35440 19876
rect 35492 19864 35498 19916
rect 35866 19904 35894 20012
rect 36906 19904 36912 19916
rect 35866 19876 36912 19904
rect 36906 19864 36912 19876
rect 36964 19864 36970 19916
rect 32306 19796 32312 19848
rect 32364 19796 32370 19848
rect 33137 19839 33195 19845
rect 33137 19805 33149 19839
rect 33183 19836 33195 19839
rect 33318 19836 33324 19848
rect 33183 19808 33324 19836
rect 33183 19805 33195 19808
rect 33137 19799 33195 19805
rect 33318 19796 33324 19808
rect 33376 19796 33382 19848
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19836 33931 19839
rect 33962 19836 33968 19848
rect 33919 19808 33968 19836
rect 33919 19805 33931 19808
rect 33873 19799 33931 19805
rect 33962 19796 33968 19808
rect 34020 19796 34026 19848
rect 34974 19796 34980 19848
rect 35032 19796 35038 19848
rect 35805 19839 35863 19845
rect 35805 19805 35817 19839
rect 35851 19836 35863 19839
rect 36722 19836 36728 19848
rect 35851 19808 36728 19836
rect 35851 19805 35863 19808
rect 35805 19799 35863 19805
rect 36722 19796 36728 19808
rect 36780 19796 36786 19848
rect 41230 19796 41236 19848
rect 41288 19836 41294 19848
rect 44085 19839 44143 19845
rect 44085 19836 44097 19839
rect 41288 19808 44097 19836
rect 41288 19796 41294 19808
rect 44085 19805 44097 19808
rect 44131 19805 44143 19839
rect 44085 19799 44143 19805
rect 27111 19740 31800 19768
rect 27111 19737 27123 19740
rect 27065 19731 27123 19737
rect 32030 19728 32036 19780
rect 32088 19768 32094 19780
rect 34057 19771 34115 19777
rect 32088 19740 33272 19768
rect 32088 19728 32094 19740
rect 23934 19700 23940 19712
rect 21468 19672 23940 19700
rect 18647 19669 18659 19672
rect 18601 19663 18659 19669
rect 23934 19660 23940 19672
rect 23992 19660 23998 19712
rect 25590 19660 25596 19712
rect 25648 19660 25654 19712
rect 25685 19703 25743 19709
rect 25685 19669 25697 19703
rect 25731 19700 25743 19703
rect 26418 19700 26424 19712
rect 25731 19672 26424 19700
rect 25731 19669 25743 19672
rect 25685 19663 25743 19669
rect 26418 19660 26424 19672
rect 26476 19660 26482 19712
rect 26970 19660 26976 19712
rect 27028 19700 27034 19712
rect 27157 19703 27215 19709
rect 27157 19700 27169 19703
rect 27028 19672 27169 19700
rect 27028 19660 27034 19672
rect 27157 19669 27169 19672
rect 27203 19669 27215 19703
rect 27157 19663 27215 19669
rect 32306 19660 32312 19712
rect 32364 19700 32370 19712
rect 33244 19709 33272 19740
rect 34057 19737 34069 19771
rect 34103 19768 34115 19771
rect 34146 19768 34152 19780
rect 34103 19740 34152 19768
rect 34103 19737 34115 19740
rect 34057 19731 34115 19737
rect 34146 19728 34152 19740
rect 34204 19728 34210 19780
rect 44269 19771 44327 19777
rect 44269 19737 44281 19771
rect 44315 19768 44327 19771
rect 46198 19768 46204 19780
rect 44315 19740 46204 19768
rect 44315 19737 44327 19740
rect 44269 19731 44327 19737
rect 46198 19728 46204 19740
rect 46256 19728 46262 19780
rect 32401 19703 32459 19709
rect 32401 19700 32413 19703
rect 32364 19672 32413 19700
rect 32364 19660 32370 19672
rect 32401 19669 32413 19672
rect 32447 19669 32459 19703
rect 32401 19663 32459 19669
rect 33229 19703 33287 19709
rect 33229 19669 33241 19703
rect 33275 19669 33287 19703
rect 33229 19663 33287 19669
rect 34974 19660 34980 19712
rect 35032 19700 35038 19712
rect 35069 19703 35127 19709
rect 35069 19700 35081 19703
rect 35032 19672 35081 19700
rect 35032 19660 35038 19672
rect 35069 19669 35081 19672
rect 35115 19669 35127 19703
rect 35069 19663 35127 19669
rect 1104 19610 49864 19632
rect 1104 19558 7950 19610
rect 8002 19558 8014 19610
rect 8066 19558 8078 19610
rect 8130 19558 8142 19610
rect 8194 19558 8206 19610
rect 8258 19558 17950 19610
rect 18002 19558 18014 19610
rect 18066 19558 18078 19610
rect 18130 19558 18142 19610
rect 18194 19558 18206 19610
rect 18258 19558 27950 19610
rect 28002 19558 28014 19610
rect 28066 19558 28078 19610
rect 28130 19558 28142 19610
rect 28194 19558 28206 19610
rect 28258 19558 37950 19610
rect 38002 19558 38014 19610
rect 38066 19558 38078 19610
rect 38130 19558 38142 19610
rect 38194 19558 38206 19610
rect 38258 19558 47950 19610
rect 48002 19558 48014 19610
rect 48066 19558 48078 19610
rect 48130 19558 48142 19610
rect 48194 19558 48206 19610
rect 48258 19558 49864 19610
rect 1104 19536 49864 19558
rect 16482 19456 16488 19508
rect 16540 19496 16546 19508
rect 19889 19499 19947 19505
rect 19889 19496 19901 19499
rect 16540 19468 19901 19496
rect 16540 19456 16546 19468
rect 19889 19465 19901 19468
rect 19935 19465 19947 19499
rect 19889 19459 19947 19465
rect 22370 19456 22376 19508
rect 22428 19496 22434 19508
rect 23385 19499 23443 19505
rect 23385 19496 23397 19499
rect 22428 19468 23397 19496
rect 22428 19456 22434 19468
rect 23385 19465 23397 19468
rect 23431 19465 23443 19499
rect 23385 19459 23443 19465
rect 23753 19499 23811 19505
rect 23753 19465 23765 19499
rect 23799 19496 23811 19499
rect 23842 19496 23848 19508
rect 23799 19468 23848 19496
rect 23799 19465 23811 19468
rect 23753 19459 23811 19465
rect 23842 19456 23848 19468
rect 23900 19456 23906 19508
rect 27798 19496 27804 19508
rect 24596 19468 27804 19496
rect 20349 19431 20407 19437
rect 20349 19397 20361 19431
rect 20395 19428 20407 19431
rect 21174 19428 21180 19440
rect 20395 19400 21180 19428
rect 20395 19397 20407 19400
rect 20349 19391 20407 19397
rect 21174 19388 21180 19400
rect 21232 19388 21238 19440
rect 20257 19363 20315 19369
rect 20257 19329 20269 19363
rect 20303 19360 20315 19363
rect 22462 19360 22468 19372
rect 20303 19332 22468 19360
rect 20303 19329 20315 19332
rect 20257 19323 20315 19329
rect 22462 19320 22468 19332
rect 22520 19320 22526 19372
rect 23845 19363 23903 19369
rect 23845 19360 23857 19363
rect 23216 19332 23857 19360
rect 20533 19295 20591 19301
rect 20533 19261 20545 19295
rect 20579 19292 20591 19295
rect 21542 19292 21548 19304
rect 20579 19264 21548 19292
rect 20579 19261 20591 19264
rect 20533 19255 20591 19261
rect 21542 19252 21548 19264
rect 21600 19252 21606 19304
rect 23216 19292 23244 19332
rect 23845 19329 23857 19332
rect 23891 19360 23903 19363
rect 24486 19360 24492 19372
rect 23891 19332 24492 19360
rect 23891 19329 23903 19332
rect 23845 19323 23903 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24596 19369 24624 19468
rect 27798 19456 27804 19468
rect 27856 19496 27862 19508
rect 28810 19496 28816 19508
rect 27856 19468 28816 19496
rect 27856 19456 27862 19468
rect 28810 19456 28816 19468
rect 28868 19456 28874 19508
rect 33704 19468 35894 19496
rect 24762 19388 24768 19440
rect 24820 19428 24826 19440
rect 26605 19431 26663 19437
rect 24820 19400 25346 19428
rect 24820 19388 24826 19400
rect 26605 19397 26617 19431
rect 26651 19428 26663 19431
rect 26694 19428 26700 19440
rect 26651 19400 26700 19428
rect 26651 19397 26663 19400
rect 26605 19391 26663 19397
rect 26694 19388 26700 19400
rect 26752 19388 26758 19440
rect 26786 19388 26792 19440
rect 26844 19428 26850 19440
rect 27525 19431 27583 19437
rect 26844 19400 27292 19428
rect 26844 19388 26850 19400
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19329 24639 19363
rect 24581 19323 24639 19329
rect 22848 19264 23244 19292
rect 22848 19168 22876 19264
rect 23290 19252 23296 19304
rect 23348 19292 23354 19304
rect 23937 19295 23995 19301
rect 23937 19292 23949 19295
rect 23348 19264 23949 19292
rect 23348 19252 23354 19264
rect 23937 19261 23949 19264
rect 23983 19261 23995 19295
rect 24854 19292 24860 19304
rect 23937 19255 23995 19261
rect 24596 19264 24860 19292
rect 21910 19116 21916 19168
rect 21968 19156 21974 19168
rect 22738 19156 22744 19168
rect 21968 19128 22744 19156
rect 21968 19116 21974 19128
rect 22738 19116 22744 19128
rect 22796 19116 22802 19168
rect 22830 19116 22836 19168
rect 22888 19116 22894 19168
rect 23952 19156 23980 19255
rect 24596 19236 24624 19264
rect 24854 19252 24860 19264
rect 24912 19252 24918 19304
rect 27264 19292 27292 19400
rect 27525 19397 27537 19431
rect 27571 19428 27583 19431
rect 27571 19400 29224 19428
rect 27571 19397 27583 19400
rect 27525 19391 27583 19397
rect 27430 19320 27436 19372
rect 27488 19360 27494 19372
rect 28721 19363 28779 19369
rect 27488 19332 28396 19360
rect 27488 19320 27494 19332
rect 27617 19295 27675 19301
rect 27617 19292 27629 19295
rect 27264 19264 27629 19292
rect 27617 19261 27629 19264
rect 27663 19261 27675 19295
rect 27617 19255 27675 19261
rect 27798 19252 27804 19304
rect 27856 19252 27862 19304
rect 24578 19184 24584 19236
rect 24636 19184 24642 19236
rect 27062 19224 27068 19236
rect 26804 19196 27068 19224
rect 26804 19156 26832 19196
rect 27062 19184 27068 19196
rect 27120 19184 27126 19236
rect 27154 19184 27160 19236
rect 27212 19184 27218 19236
rect 28368 19233 28396 19332
rect 28721 19329 28733 19363
rect 28767 19360 28779 19363
rect 29086 19360 29092 19372
rect 28767 19332 29092 19360
rect 28767 19329 28779 19332
rect 28721 19323 28779 19329
rect 29086 19320 29092 19332
rect 29144 19320 29150 19372
rect 29196 19360 29224 19400
rect 33502 19360 33508 19372
rect 29196 19332 29408 19360
rect 28813 19295 28871 19301
rect 28813 19292 28825 19295
rect 28460 19264 28825 19292
rect 28353 19227 28411 19233
rect 28353 19193 28365 19227
rect 28399 19193 28411 19227
rect 28353 19187 28411 19193
rect 23952 19128 26832 19156
rect 26878 19116 26884 19168
rect 26936 19156 26942 19168
rect 27246 19156 27252 19168
rect 26936 19128 27252 19156
rect 26936 19116 26942 19128
rect 27246 19116 27252 19128
rect 27304 19156 27310 19168
rect 28460 19156 28488 19264
rect 28813 19261 28825 19264
rect 28859 19261 28871 19295
rect 28813 19255 28871 19261
rect 28905 19295 28963 19301
rect 28905 19261 28917 19295
rect 28951 19261 28963 19295
rect 29380 19292 29408 19332
rect 29564 19332 33508 19360
rect 29564 19292 29592 19332
rect 33502 19320 33508 19332
rect 33560 19320 33566 19372
rect 33704 19369 33732 19468
rect 35866 19428 35894 19468
rect 38470 19456 38476 19508
rect 38528 19496 38534 19508
rect 39209 19499 39267 19505
rect 39209 19496 39221 19499
rect 38528 19468 39221 19496
rect 38528 19456 38534 19468
rect 39209 19465 39221 19468
rect 39255 19465 39267 19499
rect 39209 19459 39267 19465
rect 39022 19428 39028 19440
rect 35866 19400 36032 19428
rect 38962 19400 39028 19428
rect 33689 19363 33747 19369
rect 33689 19329 33701 19363
rect 33735 19329 33747 19363
rect 35894 19360 35900 19372
rect 35098 19332 35900 19360
rect 33689 19323 33747 19329
rect 35894 19320 35900 19332
rect 35952 19320 35958 19372
rect 29380 19264 29592 19292
rect 33965 19295 34023 19301
rect 28905 19255 28963 19261
rect 33965 19261 33977 19295
rect 34011 19292 34023 19295
rect 36004 19292 36032 19400
rect 39022 19388 39028 19400
rect 39080 19388 39086 19440
rect 37458 19320 37464 19372
rect 37516 19320 37522 19372
rect 45462 19320 45468 19372
rect 45520 19360 45526 19372
rect 47949 19363 48007 19369
rect 47949 19360 47961 19363
rect 45520 19332 47961 19360
rect 45520 19320 45526 19332
rect 47949 19329 47961 19332
rect 47995 19329 48007 19363
rect 47949 19323 48007 19329
rect 49142 19320 49148 19372
rect 49200 19320 49206 19372
rect 37274 19292 37280 19304
rect 34011 19264 35894 19292
rect 36004 19264 37280 19292
rect 34011 19261 34023 19264
rect 33965 19255 34023 19261
rect 28534 19184 28540 19236
rect 28592 19224 28598 19236
rect 28920 19224 28948 19255
rect 35866 19224 35894 19264
rect 37274 19252 37280 19264
rect 37332 19292 37338 19304
rect 37476 19292 37504 19320
rect 37737 19295 37795 19301
rect 37737 19292 37749 19295
rect 37332 19264 37504 19292
rect 37568 19264 37749 19292
rect 37332 19252 37338 19264
rect 36630 19224 36636 19236
rect 28592 19196 28948 19224
rect 34992 19196 35572 19224
rect 35866 19196 36636 19224
rect 28592 19184 28598 19196
rect 27304 19128 28488 19156
rect 27304 19116 27310 19128
rect 34422 19116 34428 19168
rect 34480 19156 34486 19168
rect 34992 19156 35020 19196
rect 34480 19128 35020 19156
rect 34480 19116 34486 19128
rect 35434 19116 35440 19168
rect 35492 19116 35498 19168
rect 35544 19156 35572 19196
rect 36630 19184 36636 19196
rect 36688 19184 36694 19236
rect 37568 19168 37596 19264
rect 37737 19261 37749 19264
rect 37783 19261 37795 19295
rect 37737 19255 37795 19261
rect 36078 19156 36084 19168
rect 35544 19128 36084 19156
rect 36078 19116 36084 19128
rect 36136 19116 36142 19168
rect 37550 19116 37556 19168
rect 37608 19116 37614 19168
rect 1104 19066 49864 19088
rect 1104 19014 2950 19066
rect 3002 19014 3014 19066
rect 3066 19014 3078 19066
rect 3130 19014 3142 19066
rect 3194 19014 3206 19066
rect 3258 19014 12950 19066
rect 13002 19014 13014 19066
rect 13066 19014 13078 19066
rect 13130 19014 13142 19066
rect 13194 19014 13206 19066
rect 13258 19014 22950 19066
rect 23002 19014 23014 19066
rect 23066 19014 23078 19066
rect 23130 19014 23142 19066
rect 23194 19014 23206 19066
rect 23258 19014 32950 19066
rect 33002 19014 33014 19066
rect 33066 19014 33078 19066
rect 33130 19014 33142 19066
rect 33194 19014 33206 19066
rect 33258 19014 42950 19066
rect 43002 19014 43014 19066
rect 43066 19014 43078 19066
rect 43130 19014 43142 19066
rect 43194 19014 43206 19066
rect 43258 19014 49864 19066
rect 1104 18992 49864 19014
rect 18141 18955 18199 18961
rect 18141 18921 18153 18955
rect 18187 18952 18199 18955
rect 18782 18952 18788 18964
rect 18187 18924 18788 18952
rect 18187 18921 18199 18924
rect 18141 18915 18199 18921
rect 18782 18912 18788 18924
rect 18840 18912 18846 18964
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 19944 18924 20269 18952
rect 19944 18912 19950 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22370 18952 22376 18964
rect 22152 18924 22376 18952
rect 22152 18912 22158 18924
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 22462 18912 22468 18964
rect 22520 18912 22526 18964
rect 22738 18912 22744 18964
rect 22796 18952 22802 18964
rect 24581 18955 24639 18961
rect 24581 18952 24593 18955
rect 22796 18924 24593 18952
rect 22796 18912 22802 18924
rect 24581 18921 24593 18924
rect 24627 18921 24639 18955
rect 24581 18915 24639 18921
rect 24762 18912 24768 18964
rect 24820 18952 24826 18964
rect 27798 18952 27804 18964
rect 24820 18924 27804 18952
rect 24820 18912 24826 18924
rect 27798 18912 27804 18924
rect 27856 18952 27862 18964
rect 28534 18952 28540 18964
rect 27856 18924 28540 18952
rect 27856 18912 27862 18924
rect 28534 18912 28540 18924
rect 28592 18912 28598 18964
rect 37550 18912 37556 18964
rect 37608 18952 37614 18964
rect 38657 18955 38715 18961
rect 38657 18952 38669 18955
rect 37608 18924 38669 18952
rect 37608 18912 37614 18924
rect 38657 18921 38669 18924
rect 38703 18921 38715 18955
rect 38657 18915 38715 18921
rect 9766 18844 9772 18896
rect 9824 18884 9830 18896
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 9824 18856 18337 18884
rect 9824 18844 9830 18856
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 18325 18847 18383 18853
rect 21174 18844 21180 18896
rect 21232 18884 21238 18896
rect 23293 18887 23351 18893
rect 23293 18884 23305 18887
rect 21232 18856 23305 18884
rect 21232 18844 21238 18856
rect 23293 18853 23305 18856
rect 23339 18853 23351 18887
rect 23293 18847 23351 18853
rect 30929 18887 30987 18893
rect 30929 18853 30941 18887
rect 30975 18884 30987 18887
rect 32858 18884 32864 18896
rect 30975 18856 32864 18884
rect 30975 18853 30987 18856
rect 30929 18847 30987 18853
rect 32858 18844 32864 18856
rect 32916 18844 32922 18896
rect 20901 18819 20959 18825
rect 20901 18785 20913 18819
rect 20947 18816 20959 18819
rect 20947 18788 21404 18816
rect 20947 18785 20959 18788
rect 20901 18779 20959 18785
rect 4617 18751 4675 18757
rect 4617 18717 4629 18751
rect 4663 18748 4675 18751
rect 9306 18748 9312 18760
rect 4663 18720 9312 18748
rect 4663 18717 4675 18720
rect 4617 18711 4675 18717
rect 9306 18708 9312 18720
rect 9364 18708 9370 18760
rect 12526 18708 12532 18760
rect 12584 18748 12590 18760
rect 17865 18751 17923 18757
rect 17865 18748 17877 18751
rect 12584 18720 17877 18748
rect 12584 18708 12590 18720
rect 17865 18717 17877 18720
rect 17911 18717 17923 18751
rect 17865 18711 17923 18717
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 20588 18652 20729 18680
rect 20588 18640 20594 18652
rect 20717 18649 20729 18652
rect 20763 18649 20775 18683
rect 20717 18643 20775 18649
rect 2774 18572 2780 18624
rect 2832 18612 2838 18624
rect 4709 18615 4767 18621
rect 4709 18612 4721 18615
rect 2832 18584 4721 18612
rect 2832 18572 2838 18584
rect 4709 18581 4721 18584
rect 4755 18581 4767 18615
rect 4709 18575 4767 18581
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 21376 18612 21404 18788
rect 21818 18776 21824 18828
rect 21876 18816 21882 18828
rect 23109 18819 23167 18825
rect 21876 18788 22324 18816
rect 21876 18776 21882 18788
rect 22296 18692 22324 18788
rect 23109 18785 23121 18819
rect 23155 18816 23167 18819
rect 23474 18816 23480 18828
rect 23155 18788 23480 18816
rect 23155 18785 23167 18788
rect 23109 18779 23167 18785
rect 23474 18776 23480 18788
rect 23532 18816 23538 18828
rect 23845 18819 23903 18825
rect 23845 18816 23857 18819
rect 23532 18788 23857 18816
rect 23532 18776 23538 18788
rect 23845 18785 23857 18788
rect 23891 18785 23903 18819
rect 23845 18779 23903 18785
rect 24302 18776 24308 18828
rect 24360 18816 24366 18828
rect 25133 18819 25191 18825
rect 25133 18816 25145 18819
rect 24360 18788 25145 18816
rect 24360 18776 24366 18788
rect 25133 18785 25145 18788
rect 25179 18785 25191 18819
rect 25133 18779 25191 18785
rect 26602 18776 26608 18828
rect 26660 18776 26666 18828
rect 26970 18776 26976 18828
rect 27028 18816 27034 18828
rect 27028 18788 28488 18816
rect 27028 18776 27034 18788
rect 22462 18708 22468 18760
rect 22520 18748 22526 18760
rect 22925 18751 22983 18757
rect 22925 18748 22937 18751
rect 22520 18720 22937 18748
rect 22520 18708 22526 18720
rect 22925 18717 22937 18720
rect 22971 18717 22983 18751
rect 22925 18711 22983 18717
rect 23661 18751 23719 18757
rect 23661 18717 23673 18751
rect 23707 18748 23719 18751
rect 25774 18748 25780 18760
rect 23707 18720 25780 18748
rect 23707 18717 23719 18720
rect 23661 18711 23719 18717
rect 25774 18708 25780 18720
rect 25832 18708 25838 18760
rect 26421 18751 26479 18757
rect 26421 18717 26433 18751
rect 26467 18748 26479 18751
rect 27522 18748 27528 18760
rect 26467 18720 27528 18748
rect 26467 18717 26479 18720
rect 26421 18711 26479 18717
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 27614 18708 27620 18760
rect 27672 18748 27678 18760
rect 28350 18748 28356 18760
rect 27672 18720 28356 18748
rect 27672 18708 27678 18720
rect 28350 18708 28356 18720
rect 28408 18708 28414 18760
rect 28460 18748 28488 18788
rect 28810 18776 28816 18828
rect 28868 18816 28874 18828
rect 28997 18819 29055 18825
rect 28997 18816 29009 18819
rect 28868 18788 29009 18816
rect 28868 18776 28874 18788
rect 28997 18785 29009 18788
rect 29043 18785 29055 18819
rect 28997 18779 29055 18785
rect 31386 18776 31392 18828
rect 31444 18776 31450 18828
rect 31573 18819 31631 18825
rect 31573 18785 31585 18819
rect 31619 18816 31631 18819
rect 32582 18816 32588 18828
rect 31619 18788 32588 18816
rect 31619 18785 31631 18788
rect 31573 18779 31631 18785
rect 32582 18776 32588 18788
rect 32640 18776 32646 18828
rect 36909 18819 36967 18825
rect 36909 18785 36921 18819
rect 36955 18816 36967 18819
rect 37274 18816 37280 18828
rect 36955 18788 37280 18816
rect 36955 18785 36967 18788
rect 36909 18779 36967 18785
rect 37274 18776 37280 18788
rect 37332 18776 37338 18828
rect 31297 18751 31355 18757
rect 31297 18748 31309 18751
rect 28460 18720 31309 18748
rect 31297 18717 31309 18720
rect 31343 18717 31355 18751
rect 31297 18711 31355 18717
rect 41322 18708 41328 18760
rect 41380 18748 41386 18760
rect 44177 18751 44235 18757
rect 44177 18748 44189 18751
rect 41380 18720 44189 18748
rect 41380 18708 41386 18720
rect 44177 18717 44189 18720
rect 44223 18717 44235 18751
rect 44177 18711 44235 18717
rect 44450 18708 44456 18760
rect 44508 18748 44514 18760
rect 47949 18751 48007 18757
rect 47949 18748 47961 18751
rect 44508 18720 47961 18748
rect 44508 18708 44514 18720
rect 47949 18717 47961 18720
rect 47995 18717 48007 18751
rect 47949 18711 48007 18717
rect 21450 18640 21456 18692
rect 21508 18680 21514 18692
rect 21508 18652 22232 18680
rect 21508 18640 21514 18652
rect 22094 18612 22100 18624
rect 21376 18584 22100 18612
rect 22094 18572 22100 18584
rect 22152 18572 22158 18624
rect 22204 18612 22232 18652
rect 22278 18640 22284 18692
rect 22336 18640 22342 18692
rect 28261 18683 28319 18689
rect 28261 18680 28273 18683
rect 22388 18652 28273 18680
rect 22388 18612 22416 18652
rect 28261 18649 28273 18652
rect 28307 18680 28319 18683
rect 28442 18680 28448 18692
rect 28307 18652 28448 18680
rect 28307 18649 28319 18652
rect 28261 18643 28319 18649
rect 28442 18640 28448 18652
rect 28500 18640 28506 18692
rect 36265 18683 36323 18689
rect 36265 18649 36277 18683
rect 36311 18649 36323 18683
rect 36265 18643 36323 18649
rect 36449 18683 36507 18689
rect 36449 18649 36461 18683
rect 36495 18680 36507 18683
rect 36722 18680 36728 18692
rect 36495 18652 36728 18680
rect 36495 18649 36507 18652
rect 36449 18643 36507 18649
rect 22204 18584 22416 18612
rect 22833 18615 22891 18621
rect 22833 18581 22845 18615
rect 22879 18612 22891 18615
rect 23382 18612 23388 18624
rect 22879 18584 23388 18612
rect 22879 18581 22891 18584
rect 22833 18575 22891 18581
rect 23382 18572 23388 18584
rect 23440 18572 23446 18624
rect 23753 18615 23811 18621
rect 23753 18581 23765 18615
rect 23799 18612 23811 18615
rect 24854 18612 24860 18624
rect 23799 18584 24860 18612
rect 23799 18581 23811 18584
rect 23753 18575 23811 18581
rect 24854 18572 24860 18584
rect 24912 18572 24918 18624
rect 24946 18572 24952 18624
rect 25004 18572 25010 18624
rect 25041 18615 25099 18621
rect 25041 18581 25053 18615
rect 25087 18612 25099 18615
rect 25866 18612 25872 18624
rect 25087 18584 25872 18612
rect 25087 18581 25099 18584
rect 25041 18575 25099 18581
rect 25866 18572 25872 18584
rect 25924 18572 25930 18624
rect 25958 18572 25964 18624
rect 26016 18572 26022 18624
rect 26329 18615 26387 18621
rect 26329 18581 26341 18615
rect 26375 18612 26387 18615
rect 27246 18612 27252 18624
rect 26375 18584 27252 18612
rect 26375 18581 26387 18584
rect 26329 18575 26387 18581
rect 27246 18572 27252 18584
rect 27304 18572 27310 18624
rect 27338 18572 27344 18624
rect 27396 18612 27402 18624
rect 29270 18612 29276 18624
rect 27396 18584 29276 18612
rect 27396 18572 27402 18584
rect 29270 18572 29276 18584
rect 29328 18572 29334 18624
rect 36280 18612 36308 18643
rect 36722 18640 36728 18652
rect 36780 18640 36786 18692
rect 37182 18640 37188 18692
rect 37240 18640 37246 18692
rect 38654 18680 38660 18692
rect 38410 18652 38660 18680
rect 38654 18640 38660 18652
rect 38712 18640 38718 18692
rect 44361 18683 44419 18689
rect 44361 18649 44373 18683
rect 44407 18680 44419 18683
rect 47854 18680 47860 18692
rect 44407 18652 47860 18680
rect 44407 18649 44419 18652
rect 44361 18643 44419 18649
rect 47854 18640 47860 18652
rect 47912 18640 47918 18692
rect 49142 18640 49148 18692
rect 49200 18640 49206 18692
rect 36998 18612 37004 18624
rect 36280 18584 37004 18612
rect 36998 18572 37004 18584
rect 37056 18572 37062 18624
rect 1104 18522 49864 18544
rect 1104 18470 7950 18522
rect 8002 18470 8014 18522
rect 8066 18470 8078 18522
rect 8130 18470 8142 18522
rect 8194 18470 8206 18522
rect 8258 18470 17950 18522
rect 18002 18470 18014 18522
rect 18066 18470 18078 18522
rect 18130 18470 18142 18522
rect 18194 18470 18206 18522
rect 18258 18470 27950 18522
rect 28002 18470 28014 18522
rect 28066 18470 28078 18522
rect 28130 18470 28142 18522
rect 28194 18470 28206 18522
rect 28258 18470 37950 18522
rect 38002 18470 38014 18522
rect 38066 18470 38078 18522
rect 38130 18470 38142 18522
rect 38194 18470 38206 18522
rect 38258 18470 47950 18522
rect 48002 18470 48014 18522
rect 48066 18470 48078 18522
rect 48130 18470 48142 18522
rect 48194 18470 48206 18522
rect 48258 18470 49864 18522
rect 1104 18448 49864 18470
rect 19794 18368 19800 18420
rect 19852 18368 19858 18420
rect 20622 18368 20628 18420
rect 20680 18408 20686 18420
rect 20680 18380 24808 18408
rect 20680 18368 20686 18380
rect 20533 18343 20591 18349
rect 20533 18309 20545 18343
rect 20579 18340 20591 18343
rect 21450 18340 21456 18352
rect 20579 18312 21456 18340
rect 20579 18309 20591 18312
rect 20533 18303 20591 18309
rect 21450 18300 21456 18312
rect 21508 18300 21514 18352
rect 21542 18300 21548 18352
rect 21600 18340 21606 18352
rect 23293 18343 23351 18349
rect 23293 18340 23305 18343
rect 21600 18312 23305 18340
rect 21600 18300 21606 18312
rect 23293 18309 23305 18312
rect 23339 18309 23351 18343
rect 24578 18340 24584 18352
rect 24518 18312 24584 18340
rect 23293 18303 23351 18309
rect 24578 18300 24584 18312
rect 24636 18300 24642 18352
rect 1765 18275 1823 18281
rect 1765 18241 1777 18275
rect 1811 18272 1823 18275
rect 2866 18272 2872 18284
rect 1811 18244 2872 18272
rect 1811 18241 1823 18244
rect 1765 18235 1823 18241
rect 2866 18232 2872 18244
rect 2924 18232 2930 18284
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 22094 18272 22100 18284
rect 19751 18244 22100 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 22094 18232 22100 18244
rect 22152 18232 22158 18284
rect 22278 18232 22284 18284
rect 22336 18272 22342 18284
rect 23017 18275 23075 18281
rect 23017 18272 23029 18275
rect 22336 18244 23029 18272
rect 22336 18232 22342 18244
rect 23017 18241 23029 18244
rect 23063 18241 23075 18275
rect 24780 18272 24808 18380
rect 24946 18368 24952 18420
rect 25004 18408 25010 18420
rect 27249 18411 27307 18417
rect 27249 18408 27261 18411
rect 25004 18380 27261 18408
rect 25004 18368 25010 18380
rect 27249 18377 27261 18380
rect 27295 18377 27307 18411
rect 27249 18371 27307 18377
rect 27614 18368 27620 18420
rect 27672 18408 27678 18420
rect 34057 18411 34115 18417
rect 27672 18380 29040 18408
rect 27672 18368 27678 18380
rect 24854 18300 24860 18352
rect 24912 18340 24918 18352
rect 27154 18340 27160 18352
rect 24912 18312 27160 18340
rect 24912 18300 24918 18312
rect 27154 18300 27160 18312
rect 27212 18300 27218 18352
rect 28442 18300 28448 18352
rect 28500 18300 28506 18352
rect 29012 18340 29040 18380
rect 34057 18377 34069 18411
rect 34103 18408 34115 18411
rect 34790 18408 34796 18420
rect 34103 18380 34796 18408
rect 34103 18377 34115 18380
rect 34057 18371 34115 18377
rect 34790 18368 34796 18380
rect 34848 18368 34854 18420
rect 37734 18368 37740 18420
rect 37792 18408 37798 18420
rect 37921 18411 37979 18417
rect 37921 18408 37933 18411
rect 37792 18380 37933 18408
rect 37792 18368 37798 18380
rect 37921 18377 37933 18380
rect 37967 18377 37979 18411
rect 37921 18371 37979 18377
rect 32306 18340 32312 18352
rect 29012 18312 32312 18340
rect 32306 18300 32312 18312
rect 32364 18300 32370 18352
rect 32582 18300 32588 18352
rect 32640 18300 32646 18352
rect 34422 18340 34428 18352
rect 33810 18326 34428 18340
rect 33796 18312 34428 18326
rect 24780 18244 24900 18272
rect 23017 18235 23075 18241
rect 1302 18164 1308 18216
rect 1360 18204 1366 18216
rect 2041 18207 2099 18213
rect 2041 18204 2053 18207
rect 1360 18176 2053 18204
rect 1360 18164 1366 18176
rect 2041 18173 2053 18176
rect 2087 18173 2099 18207
rect 2041 18167 2099 18173
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18204 20039 18207
rect 20070 18204 20076 18216
rect 20027 18176 20076 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 20070 18164 20076 18176
rect 20128 18164 20134 18216
rect 20990 18164 20996 18216
rect 21048 18204 21054 18216
rect 21269 18207 21327 18213
rect 21269 18204 21281 18207
rect 21048 18176 21281 18204
rect 21048 18164 21054 18176
rect 21269 18173 21281 18176
rect 21315 18173 21327 18207
rect 21269 18167 21327 18173
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 18840 18108 20024 18136
rect 18840 18096 18846 18108
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19794 18068 19800 18080
rect 19383 18040 19800 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19794 18028 19800 18040
rect 19852 18028 19858 18080
rect 19996 18068 20024 18108
rect 21910 18096 21916 18148
rect 21968 18136 21974 18148
rect 22554 18136 22560 18148
rect 21968 18108 22560 18136
rect 21968 18096 21974 18108
rect 22554 18096 22560 18108
rect 22612 18096 22618 18148
rect 24762 18068 24768 18080
rect 19996 18040 24768 18068
rect 24762 18028 24768 18040
rect 24820 18028 24826 18080
rect 24872 18068 24900 18244
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 27338 18232 27344 18284
rect 27396 18272 27402 18284
rect 27709 18275 27767 18281
rect 27709 18272 27721 18275
rect 27396 18244 27721 18272
rect 27396 18232 27402 18244
rect 27709 18241 27721 18244
rect 27755 18241 27767 18275
rect 30193 18275 30251 18281
rect 30193 18272 30205 18275
rect 27709 18235 27767 18241
rect 28460 18244 30205 18272
rect 27430 18164 27436 18216
rect 27488 18204 27494 18216
rect 27801 18207 27859 18213
rect 27801 18204 27813 18207
rect 27488 18176 27813 18204
rect 27488 18164 27494 18176
rect 27801 18173 27813 18176
rect 27847 18173 27859 18207
rect 27801 18167 27859 18173
rect 26786 18096 26792 18148
rect 26844 18136 26850 18148
rect 28460 18136 28488 18244
rect 30193 18241 30205 18244
rect 30239 18241 30251 18275
rect 30193 18235 30251 18241
rect 30285 18275 30343 18281
rect 30285 18241 30297 18275
rect 30331 18272 30343 18275
rect 31202 18272 31208 18284
rect 30331 18244 31208 18272
rect 30331 18241 30343 18244
rect 30285 18235 30343 18241
rect 31202 18232 31208 18244
rect 31260 18232 31266 18284
rect 29273 18207 29331 18213
rect 29273 18173 29285 18207
rect 29319 18204 29331 18207
rect 30006 18204 30012 18216
rect 29319 18176 30012 18204
rect 29319 18173 29331 18176
rect 29273 18167 29331 18173
rect 30006 18164 30012 18176
rect 30064 18164 30070 18216
rect 30374 18164 30380 18216
rect 30432 18164 30438 18216
rect 32309 18207 32367 18213
rect 32309 18173 32321 18207
rect 32355 18173 32367 18207
rect 32309 18167 32367 18173
rect 26844 18108 28488 18136
rect 30024 18136 30052 18164
rect 32324 18136 32352 18167
rect 33318 18164 33324 18216
rect 33376 18204 33382 18216
rect 33796 18204 33824 18312
rect 34422 18300 34428 18312
rect 34480 18300 34486 18352
rect 36078 18340 36084 18352
rect 36018 18312 36084 18340
rect 36078 18300 36084 18312
rect 36136 18340 36142 18352
rect 36814 18340 36820 18352
rect 36136 18312 36820 18340
rect 36136 18300 36142 18312
rect 36814 18300 36820 18312
rect 36872 18300 36878 18352
rect 37366 18232 37372 18284
rect 37424 18272 37430 18284
rect 37829 18275 37887 18281
rect 37829 18272 37841 18275
rect 37424 18244 37841 18272
rect 37424 18232 37430 18244
rect 37829 18241 37841 18244
rect 37875 18241 37887 18275
rect 37829 18235 37887 18241
rect 46658 18232 46664 18284
rect 46716 18272 46722 18284
rect 47949 18275 48007 18281
rect 47949 18272 47961 18275
rect 46716 18244 47961 18272
rect 46716 18232 46722 18244
rect 47949 18241 47961 18244
rect 47995 18241 48007 18275
rect 47949 18235 48007 18241
rect 33376 18176 33824 18204
rect 34517 18207 34575 18213
rect 33376 18164 33382 18176
rect 34517 18173 34529 18207
rect 34563 18173 34575 18207
rect 34517 18167 34575 18173
rect 30024 18108 32352 18136
rect 26844 18096 26850 18108
rect 29086 18068 29092 18080
rect 24872 18040 29092 18068
rect 29086 18028 29092 18040
rect 29144 18028 29150 18080
rect 29825 18071 29883 18077
rect 29825 18037 29837 18071
rect 29871 18068 29883 18071
rect 33686 18068 33692 18080
rect 29871 18040 33692 18068
rect 29871 18037 29883 18040
rect 29825 18031 29883 18037
rect 33686 18028 33692 18040
rect 33744 18028 33750 18080
rect 34532 18068 34560 18167
rect 34790 18164 34796 18216
rect 34848 18204 34854 18216
rect 35250 18204 35256 18216
rect 34848 18176 35256 18204
rect 34848 18164 34854 18176
rect 35250 18164 35256 18176
rect 35308 18164 35314 18216
rect 38010 18164 38016 18216
rect 38068 18204 38074 18216
rect 38105 18207 38163 18213
rect 38105 18204 38117 18207
rect 38068 18176 38117 18204
rect 38068 18164 38074 18176
rect 38105 18173 38117 18176
rect 38151 18204 38163 18207
rect 38470 18204 38476 18216
rect 38151 18176 38476 18204
rect 38151 18173 38163 18176
rect 38105 18167 38163 18173
rect 38470 18164 38476 18176
rect 38528 18164 38534 18216
rect 49142 18164 49148 18216
rect 49200 18164 49206 18216
rect 34882 18068 34888 18080
rect 34532 18040 34888 18068
rect 34882 18028 34888 18040
rect 34940 18028 34946 18080
rect 36078 18028 36084 18080
rect 36136 18068 36142 18080
rect 36265 18071 36323 18077
rect 36265 18068 36277 18071
rect 36136 18040 36277 18068
rect 36136 18028 36142 18040
rect 36265 18037 36277 18040
rect 36311 18037 36323 18071
rect 36265 18031 36323 18037
rect 37461 18071 37519 18077
rect 37461 18037 37473 18071
rect 37507 18068 37519 18071
rect 41782 18068 41788 18080
rect 37507 18040 41788 18068
rect 37507 18037 37519 18040
rect 37461 18031 37519 18037
rect 41782 18028 41788 18040
rect 41840 18028 41846 18080
rect 1104 17978 49864 18000
rect 1104 17926 2950 17978
rect 3002 17926 3014 17978
rect 3066 17926 3078 17978
rect 3130 17926 3142 17978
rect 3194 17926 3206 17978
rect 3258 17926 12950 17978
rect 13002 17926 13014 17978
rect 13066 17926 13078 17978
rect 13130 17926 13142 17978
rect 13194 17926 13206 17978
rect 13258 17926 22950 17978
rect 23002 17926 23014 17978
rect 23066 17926 23078 17978
rect 23130 17926 23142 17978
rect 23194 17926 23206 17978
rect 23258 17926 32950 17978
rect 33002 17926 33014 17978
rect 33066 17926 33078 17978
rect 33130 17926 33142 17978
rect 33194 17926 33206 17978
rect 33258 17926 42950 17978
rect 43002 17926 43014 17978
rect 43066 17926 43078 17978
rect 43130 17926 43142 17978
rect 43194 17926 43206 17978
rect 43258 17926 49864 17978
rect 1104 17904 49864 17926
rect 17862 17824 17868 17876
rect 17920 17864 17926 17876
rect 19429 17867 19487 17873
rect 19429 17864 19441 17867
rect 17920 17836 19441 17864
rect 17920 17824 17926 17836
rect 19429 17833 19441 17836
rect 19475 17833 19487 17867
rect 21910 17864 21916 17876
rect 19429 17827 19487 17833
rect 19996 17836 21916 17864
rect 18141 17799 18199 17805
rect 18141 17765 18153 17799
rect 18187 17796 18199 17799
rect 19886 17796 19892 17808
rect 18187 17768 19892 17796
rect 18187 17765 18199 17768
rect 18141 17759 18199 17765
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 18785 17731 18843 17737
rect 18785 17697 18797 17731
rect 18831 17728 18843 17731
rect 19996 17728 20024 17836
rect 21910 17824 21916 17836
rect 21968 17824 21974 17876
rect 22002 17824 22008 17876
rect 22060 17864 22066 17876
rect 22462 17864 22468 17876
rect 22060 17836 22468 17864
rect 22060 17824 22066 17836
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 25590 17824 25596 17876
rect 25648 17864 25654 17876
rect 27341 17867 27399 17873
rect 27341 17864 27353 17867
rect 25648 17836 27353 17864
rect 25648 17824 25654 17836
rect 27341 17833 27353 17836
rect 27387 17833 27399 17867
rect 27341 17827 27399 17833
rect 32401 17867 32459 17873
rect 32401 17833 32413 17867
rect 32447 17864 32459 17867
rect 32582 17864 32588 17876
rect 32447 17836 32588 17864
rect 32447 17833 32459 17836
rect 32401 17827 32459 17833
rect 32582 17824 32588 17836
rect 32640 17824 32646 17876
rect 37182 17824 37188 17876
rect 37240 17864 37246 17876
rect 37277 17867 37335 17873
rect 37277 17864 37289 17867
rect 37240 17836 37289 17864
rect 37240 17824 37246 17836
rect 37277 17833 37289 17836
rect 37323 17833 37335 17867
rect 37277 17827 37335 17833
rect 37384 17836 39712 17864
rect 22370 17756 22376 17808
rect 22428 17796 22434 17808
rect 22428 17768 23060 17796
rect 22428 17756 22434 17768
rect 18831 17700 20024 17728
rect 20073 17731 20131 17737
rect 18831 17697 18843 17700
rect 18785 17691 18843 17697
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 21266 17728 21272 17740
rect 20119 17700 21272 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 21266 17688 21272 17700
rect 21324 17688 21330 17740
rect 21358 17688 21364 17740
rect 21416 17728 21422 17740
rect 22646 17728 22652 17740
rect 21416 17700 22652 17728
rect 21416 17688 21422 17700
rect 22646 17688 22652 17700
rect 22704 17688 22710 17740
rect 23032 17737 23060 17768
rect 27062 17756 27068 17808
rect 27120 17796 27126 17808
rect 34330 17796 34336 17808
rect 27120 17768 27936 17796
rect 27120 17756 27126 17768
rect 23017 17731 23075 17737
rect 23017 17697 23029 17731
rect 23063 17728 23075 17731
rect 27430 17728 27436 17740
rect 23063 17700 27436 17728
rect 23063 17697 23075 17700
rect 23017 17691 23075 17697
rect 27430 17688 27436 17700
rect 27488 17688 27494 17740
rect 27908 17737 27936 17768
rect 33704 17768 34336 17796
rect 27893 17731 27951 17737
rect 27893 17697 27905 17731
rect 27939 17697 27951 17731
rect 27893 17691 27951 17697
rect 30006 17688 30012 17740
rect 30064 17728 30070 17740
rect 33704 17737 33732 17768
rect 34330 17756 34336 17768
rect 34388 17756 34394 17808
rect 37090 17756 37096 17808
rect 37148 17796 37154 17808
rect 37384 17796 37412 17836
rect 37148 17768 37412 17796
rect 37148 17756 37154 17768
rect 30653 17731 30711 17737
rect 30653 17728 30665 17731
rect 30064 17700 30665 17728
rect 30064 17688 30070 17700
rect 30653 17697 30665 17700
rect 30699 17697 30711 17731
rect 30653 17691 30711 17697
rect 33689 17731 33747 17737
rect 33689 17697 33701 17731
rect 33735 17697 33747 17731
rect 33689 17691 33747 17697
rect 33873 17731 33931 17737
rect 33873 17697 33885 17731
rect 33919 17697 33931 17731
rect 33873 17691 33931 17697
rect 35529 17731 35587 17737
rect 35529 17697 35541 17731
rect 35575 17728 35587 17731
rect 35894 17728 35900 17740
rect 35575 17700 35900 17728
rect 35575 17697 35587 17700
rect 35529 17691 35587 17697
rect 19242 17620 19248 17672
rect 19300 17660 19306 17672
rect 20990 17660 20996 17672
rect 19300 17632 20996 17660
rect 19300 17620 19306 17632
rect 20990 17620 20996 17632
rect 21048 17620 21054 17672
rect 23290 17620 23296 17672
rect 23348 17660 23354 17672
rect 23661 17663 23719 17669
rect 23661 17660 23673 17663
rect 23348 17632 23673 17660
rect 23348 17620 23354 17632
rect 23661 17629 23673 17632
rect 23707 17629 23719 17663
rect 23661 17623 23719 17629
rect 27614 17620 27620 17672
rect 27672 17660 27678 17672
rect 27709 17663 27767 17669
rect 27709 17660 27721 17663
rect 27672 17632 27721 17660
rect 27672 17620 27678 17632
rect 27709 17629 27721 17632
rect 27755 17629 27767 17663
rect 33318 17660 33324 17672
rect 32062 17646 33324 17660
rect 27709 17623 27767 17629
rect 32048 17632 33324 17646
rect 18601 17595 18659 17601
rect 18601 17561 18613 17595
rect 18647 17592 18659 17595
rect 21358 17592 21364 17604
rect 18647 17564 21364 17592
rect 18647 17561 18659 17564
rect 18601 17555 18659 17561
rect 21358 17552 21364 17564
rect 21416 17552 21422 17604
rect 22278 17552 22284 17604
rect 22336 17552 22342 17604
rect 30009 17595 30067 17601
rect 30009 17561 30021 17595
rect 30055 17592 30067 17595
rect 30282 17592 30288 17604
rect 30055 17564 30288 17592
rect 30055 17561 30067 17564
rect 30009 17555 30067 17561
rect 30282 17552 30288 17564
rect 30340 17552 30346 17604
rect 30926 17552 30932 17604
rect 30984 17552 30990 17604
rect 18509 17527 18567 17533
rect 18509 17493 18521 17527
rect 18555 17524 18567 17527
rect 18782 17524 18788 17536
rect 18555 17496 18788 17524
rect 18555 17493 18567 17496
rect 18509 17487 18567 17493
rect 18782 17484 18788 17496
rect 18840 17484 18846 17536
rect 19794 17484 19800 17536
rect 19852 17484 19858 17536
rect 19886 17484 19892 17536
rect 19944 17484 19950 17536
rect 19978 17484 19984 17536
rect 20036 17524 20042 17536
rect 22002 17524 22008 17536
rect 20036 17496 22008 17524
rect 20036 17484 20042 17496
rect 22002 17484 22008 17496
rect 22060 17484 22066 17536
rect 24578 17484 24584 17536
rect 24636 17524 24642 17536
rect 26142 17524 26148 17536
rect 24636 17496 26148 17524
rect 24636 17484 24642 17496
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 27338 17484 27344 17536
rect 27396 17524 27402 17536
rect 27801 17527 27859 17533
rect 27801 17524 27813 17527
rect 27396 17496 27813 17524
rect 27396 17484 27402 17496
rect 27801 17493 27813 17496
rect 27847 17493 27859 17527
rect 27801 17487 27859 17493
rect 29730 17484 29736 17536
rect 29788 17524 29794 17536
rect 30101 17527 30159 17533
rect 30101 17524 30113 17527
rect 29788 17496 30113 17524
rect 29788 17484 29794 17496
rect 30101 17493 30113 17496
rect 30147 17493 30159 17527
rect 30101 17487 30159 17493
rect 30558 17484 30564 17536
rect 30616 17524 30622 17536
rect 32048 17524 32076 17632
rect 33318 17620 33324 17632
rect 33376 17620 33382 17672
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17660 33655 17663
rect 33778 17660 33784 17672
rect 33643 17632 33784 17660
rect 33643 17629 33655 17632
rect 33597 17623 33655 17629
rect 33778 17620 33784 17632
rect 33836 17620 33842 17672
rect 33888 17660 33916 17691
rect 35894 17688 35900 17700
rect 35952 17728 35958 17740
rect 37274 17728 37280 17740
rect 35952 17700 37280 17728
rect 35952 17688 35958 17700
rect 37274 17688 37280 17700
rect 37332 17728 37338 17740
rect 37737 17731 37795 17737
rect 37737 17728 37749 17731
rect 37332 17700 37749 17728
rect 37332 17688 37338 17700
rect 37737 17697 37749 17700
rect 37783 17697 37795 17731
rect 37737 17691 37795 17697
rect 38010 17688 38016 17740
rect 38068 17688 38074 17740
rect 38562 17688 38568 17740
rect 38620 17728 38626 17740
rect 39684 17728 39712 17836
rect 43165 17799 43223 17805
rect 43165 17765 43177 17799
rect 43211 17796 43223 17799
rect 44818 17796 44824 17808
rect 43211 17768 44824 17796
rect 43211 17765 43223 17768
rect 43165 17759 43223 17765
rect 44818 17756 44824 17768
rect 44876 17756 44882 17808
rect 44637 17731 44695 17737
rect 38620 17700 39528 17728
rect 39684 17700 43760 17728
rect 38620 17688 38626 17700
rect 33888 17632 35204 17660
rect 35176 17592 35204 17632
rect 35805 17595 35863 17601
rect 35805 17592 35817 17595
rect 33244 17564 34560 17592
rect 35176 17564 35817 17592
rect 33244 17533 33272 17564
rect 30616 17496 32076 17524
rect 33229 17527 33287 17533
rect 30616 17484 30622 17496
rect 33229 17493 33241 17527
rect 33275 17493 33287 17527
rect 34532 17524 34560 17564
rect 35805 17561 35817 17564
rect 35851 17592 35863 17595
rect 36078 17592 36084 17604
rect 35851 17564 36084 17592
rect 35851 17561 35863 17564
rect 35805 17555 35863 17561
rect 36078 17552 36084 17564
rect 36136 17552 36142 17604
rect 36814 17552 36820 17604
rect 36872 17552 36878 17604
rect 37090 17552 37096 17604
rect 37148 17592 37154 17604
rect 37148 17564 37964 17592
rect 37148 17552 37154 17564
rect 37826 17524 37832 17536
rect 34532 17496 37832 17524
rect 33229 17487 33287 17493
rect 37826 17484 37832 17496
rect 37884 17484 37890 17536
rect 37936 17524 37964 17564
rect 38654 17552 38660 17604
rect 38712 17552 38718 17604
rect 39500 17592 39528 17700
rect 43732 17601 43760 17700
rect 44637 17697 44649 17731
rect 44683 17728 44695 17731
rect 44683 17700 45048 17728
rect 44683 17697 44695 17700
rect 44637 17691 44695 17697
rect 43901 17663 43959 17669
rect 43901 17629 43913 17663
rect 43947 17660 43959 17663
rect 43947 17632 44680 17660
rect 43947 17629 43959 17632
rect 43901 17623 43959 17629
rect 42981 17595 43039 17601
rect 42981 17592 42993 17595
rect 39500 17564 42993 17592
rect 42981 17561 42993 17564
rect 43027 17561 43039 17595
rect 42981 17555 43039 17561
rect 43717 17595 43775 17601
rect 43717 17561 43729 17595
rect 43763 17561 43775 17595
rect 43717 17555 43775 17561
rect 44453 17595 44511 17601
rect 44453 17561 44465 17595
rect 44499 17561 44511 17595
rect 44453 17555 44511 17561
rect 39485 17527 39543 17533
rect 39485 17524 39497 17527
rect 37936 17496 39497 17524
rect 39485 17493 39497 17496
rect 39531 17493 39543 17527
rect 39485 17487 39543 17493
rect 39942 17484 39948 17536
rect 40000 17524 40006 17536
rect 44468 17524 44496 17555
rect 40000 17496 44496 17524
rect 44652 17524 44680 17632
rect 45020 17592 45048 17700
rect 45094 17620 45100 17672
rect 45152 17660 45158 17672
rect 47949 17663 48007 17669
rect 47949 17660 47961 17663
rect 45152 17632 47961 17660
rect 45152 17620 45158 17632
rect 47949 17629 47961 17632
rect 47995 17629 48007 17663
rect 47949 17623 48007 17629
rect 46842 17592 46848 17604
rect 45020 17564 46848 17592
rect 46842 17552 46848 17564
rect 46900 17552 46906 17604
rect 49142 17552 49148 17604
rect 49200 17552 49206 17604
rect 46658 17524 46664 17536
rect 44652 17496 46664 17524
rect 40000 17484 40006 17496
rect 46658 17484 46664 17496
rect 46716 17484 46722 17536
rect 1104 17434 49864 17456
rect 1104 17382 7950 17434
rect 8002 17382 8014 17434
rect 8066 17382 8078 17434
rect 8130 17382 8142 17434
rect 8194 17382 8206 17434
rect 8258 17382 17950 17434
rect 18002 17382 18014 17434
rect 18066 17382 18078 17434
rect 18130 17382 18142 17434
rect 18194 17382 18206 17434
rect 18258 17382 27950 17434
rect 28002 17382 28014 17434
rect 28066 17382 28078 17434
rect 28130 17382 28142 17434
rect 28194 17382 28206 17434
rect 28258 17382 37950 17434
rect 38002 17382 38014 17434
rect 38066 17382 38078 17434
rect 38130 17382 38142 17434
rect 38194 17382 38206 17434
rect 38258 17382 47950 17434
rect 48002 17382 48014 17434
rect 48066 17382 48078 17434
rect 48130 17382 48142 17434
rect 48194 17382 48206 17434
rect 48258 17382 49864 17434
rect 1104 17360 49864 17382
rect 21266 17280 21272 17332
rect 21324 17320 21330 17332
rect 21453 17323 21511 17329
rect 21453 17320 21465 17323
rect 21324 17292 21465 17320
rect 21324 17280 21330 17292
rect 21453 17289 21465 17292
rect 21499 17289 21511 17323
rect 21453 17283 21511 17289
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22925 17323 22983 17329
rect 22925 17320 22937 17323
rect 22152 17292 22937 17320
rect 22152 17280 22158 17292
rect 22925 17289 22937 17292
rect 22971 17289 22983 17323
rect 22925 17283 22983 17289
rect 23290 17280 23296 17332
rect 23348 17280 23354 17332
rect 23385 17323 23443 17329
rect 23385 17289 23397 17323
rect 23431 17320 23443 17323
rect 24210 17320 24216 17332
rect 23431 17292 24216 17320
rect 23431 17289 23443 17292
rect 23385 17283 23443 17289
rect 24210 17280 24216 17292
rect 24268 17280 24274 17332
rect 24688 17292 26372 17320
rect 20714 17212 20720 17264
rect 20772 17212 20778 17264
rect 22278 17252 22284 17264
rect 21206 17238 22284 17252
rect 21192 17224 22284 17238
rect 19242 17076 19248 17128
rect 19300 17116 19306 17128
rect 19705 17119 19763 17125
rect 19705 17116 19717 17119
rect 19300 17088 19717 17116
rect 19300 17076 19306 17088
rect 19705 17085 19717 17088
rect 19751 17085 19763 17119
rect 19705 17079 19763 17085
rect 19981 17119 20039 17125
rect 19981 17085 19993 17119
rect 20027 17116 20039 17119
rect 20070 17116 20076 17128
rect 20027 17088 20076 17116
rect 20027 17085 20039 17088
rect 19981 17079 20039 17085
rect 20070 17076 20076 17088
rect 20128 17076 20134 17128
rect 20714 17076 20720 17128
rect 20772 17116 20778 17128
rect 21192 17116 21220 17224
rect 22278 17212 22284 17224
rect 22336 17212 22342 17264
rect 20772 17088 21220 17116
rect 20772 17076 20778 17088
rect 21726 17076 21732 17128
rect 21784 17116 21790 17128
rect 21910 17116 21916 17128
rect 21784 17088 21916 17116
rect 21784 17076 21790 17088
rect 21910 17076 21916 17088
rect 21968 17116 21974 17128
rect 23569 17119 23627 17125
rect 23569 17116 23581 17119
rect 21968 17088 23581 17116
rect 21968 17076 21974 17088
rect 23569 17085 23581 17088
rect 23615 17116 23627 17119
rect 24688 17116 24716 17292
rect 25038 17212 25044 17264
rect 25096 17212 25102 17264
rect 26344 17252 26372 17292
rect 27246 17280 27252 17332
rect 27304 17280 27310 17332
rect 27706 17280 27712 17332
rect 27764 17280 27770 17332
rect 28810 17280 28816 17332
rect 28868 17280 28874 17332
rect 31938 17320 31944 17332
rect 29656 17292 31944 17320
rect 26602 17252 26608 17264
rect 26344 17224 26608 17252
rect 26602 17212 26608 17224
rect 26660 17212 26666 17264
rect 27617 17255 27675 17261
rect 27617 17221 27629 17255
rect 27663 17252 27675 17255
rect 29656 17252 29684 17292
rect 31938 17280 31944 17292
rect 31996 17280 32002 17332
rect 32858 17280 32864 17332
rect 32916 17320 32922 17332
rect 35161 17323 35219 17329
rect 35161 17320 35173 17323
rect 32916 17292 35173 17320
rect 32916 17280 32922 17292
rect 35161 17289 35173 17292
rect 35207 17289 35219 17323
rect 35161 17283 35219 17289
rect 36446 17280 36452 17332
rect 36504 17320 36510 17332
rect 36814 17320 36820 17332
rect 36504 17292 36820 17320
rect 36504 17280 36510 17292
rect 36814 17280 36820 17292
rect 36872 17320 36878 17332
rect 38654 17320 38660 17332
rect 36872 17292 38660 17320
rect 36872 17280 36878 17292
rect 38654 17280 38660 17292
rect 38712 17280 38718 17332
rect 27663 17224 29684 17252
rect 27663 17221 27675 17224
rect 27617 17215 27675 17221
rect 30558 17212 30564 17264
rect 30616 17252 30622 17264
rect 30616 17224 30774 17252
rect 30616 17212 30622 17224
rect 33318 17212 33324 17264
rect 33376 17252 33382 17264
rect 33962 17252 33968 17264
rect 33376 17224 33968 17252
rect 33376 17212 33382 17224
rect 33962 17212 33968 17224
rect 34020 17212 34026 17264
rect 43714 17212 43720 17264
rect 43772 17212 43778 17264
rect 26142 17144 26148 17196
rect 26200 17184 26206 17196
rect 26200 17156 28396 17184
rect 26200 17144 26206 17156
rect 23615 17088 24716 17116
rect 24765 17119 24823 17125
rect 23615 17085 23627 17088
rect 23569 17079 23627 17085
rect 24765 17085 24777 17119
rect 24811 17085 24823 17119
rect 24765 17079 24823 17085
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 22002 16980 22008 16992
rect 20036 16952 22008 16980
rect 20036 16940 20042 16952
rect 22002 16940 22008 16952
rect 22060 16940 22066 16992
rect 24780 16980 24808 17079
rect 25038 17076 25044 17128
rect 25096 17116 25102 17128
rect 27801 17119 27859 17125
rect 27801 17116 27813 17119
rect 25096 17088 27813 17116
rect 25096 17076 25102 17088
rect 27801 17085 27813 17088
rect 27847 17116 27859 17119
rect 28258 17116 28264 17128
rect 27847 17088 28264 17116
rect 27847 17085 27859 17088
rect 27801 17079 27859 17085
rect 28258 17076 28264 17088
rect 28316 17076 28322 17128
rect 28368 17048 28396 17156
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28500 17156 29132 17184
rect 28500 17144 28506 17156
rect 28534 17076 28540 17128
rect 28592 17116 28598 17128
rect 29104 17125 29132 17156
rect 32398 17144 32404 17196
rect 32456 17184 32462 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32456 17156 32505 17184
rect 32456 17144 32462 17156
rect 32493 17153 32505 17156
rect 32539 17153 32551 17187
rect 32493 17147 32551 17153
rect 33410 17144 33416 17196
rect 33468 17184 33474 17196
rect 33873 17187 33931 17193
rect 33873 17184 33885 17187
rect 33468 17156 33885 17184
rect 33468 17144 33474 17156
rect 33873 17153 33885 17156
rect 33919 17153 33931 17187
rect 33873 17147 33931 17153
rect 35069 17187 35127 17193
rect 35069 17153 35081 17187
rect 35115 17184 35127 17187
rect 36081 17187 36139 17193
rect 36081 17184 36093 17187
rect 35115 17156 36093 17184
rect 35115 17153 35127 17156
rect 35069 17147 35127 17153
rect 36081 17153 36093 17156
rect 36127 17153 36139 17187
rect 36081 17147 36139 17153
rect 28905 17119 28963 17125
rect 28905 17116 28917 17119
rect 28592 17088 28917 17116
rect 28592 17076 28598 17088
rect 28905 17085 28917 17088
rect 28951 17085 28963 17119
rect 28905 17079 28963 17085
rect 29089 17119 29147 17125
rect 29089 17085 29101 17119
rect 29135 17116 29147 17119
rect 29546 17116 29552 17128
rect 29135 17088 29552 17116
rect 29135 17085 29147 17088
rect 29089 17079 29147 17085
rect 29546 17076 29552 17088
rect 29604 17076 29610 17128
rect 30006 17076 30012 17128
rect 30064 17076 30070 17128
rect 30282 17076 30288 17128
rect 30340 17076 30346 17128
rect 30926 17076 30932 17128
rect 30984 17116 30990 17128
rect 31757 17119 31815 17125
rect 31757 17116 31769 17119
rect 30984 17088 31769 17116
rect 30984 17076 30990 17088
rect 31757 17085 31769 17088
rect 31803 17116 31815 17119
rect 33594 17116 33600 17128
rect 31803 17088 33600 17116
rect 31803 17085 31815 17088
rect 31757 17079 31815 17085
rect 33594 17076 33600 17088
rect 33652 17076 33658 17128
rect 34149 17119 34207 17125
rect 34149 17085 34161 17119
rect 34195 17116 34207 17119
rect 34606 17116 34612 17128
rect 34195 17088 34612 17116
rect 34195 17085 34207 17088
rect 34149 17079 34207 17085
rect 34606 17076 34612 17088
rect 34664 17076 34670 17128
rect 35250 17076 35256 17128
rect 35308 17076 35314 17128
rect 33505 17051 33563 17057
rect 28368 17020 28580 17048
rect 25682 16980 25688 16992
rect 24780 16952 25688 16980
rect 25682 16940 25688 16952
rect 25740 16940 25746 16992
rect 26513 16983 26571 16989
rect 26513 16949 26525 16983
rect 26559 16980 26571 16983
rect 26602 16980 26608 16992
rect 26559 16952 26608 16980
rect 26559 16949 26571 16952
rect 26513 16943 26571 16949
rect 26602 16940 26608 16952
rect 26660 16940 26666 16992
rect 28442 16940 28448 16992
rect 28500 16940 28506 16992
rect 28552 16980 28580 17020
rect 33505 17017 33517 17051
rect 33551 17017 33563 17051
rect 33505 17011 33563 17017
rect 34701 17051 34759 17057
rect 34701 17017 34713 17051
rect 34747 17048 34759 17051
rect 40218 17048 40224 17060
rect 34747 17020 40224 17048
rect 34747 17017 34759 17020
rect 34701 17011 34759 17017
rect 30466 16980 30472 16992
rect 28552 16952 30472 16980
rect 30466 16940 30472 16952
rect 30524 16940 30530 16992
rect 32306 16940 32312 16992
rect 32364 16940 32370 16992
rect 33520 16980 33548 17011
rect 40218 17008 40224 17020
rect 40276 17008 40282 17060
rect 43901 17051 43959 17057
rect 43901 17017 43913 17051
rect 43947 17048 43959 17051
rect 46750 17048 46756 17060
rect 43947 17020 46756 17048
rect 43947 17017 43959 17020
rect 43901 17011 43959 17017
rect 46750 17008 46756 17020
rect 46808 17008 46814 17060
rect 36814 16980 36820 16992
rect 33520 16952 36820 16980
rect 36814 16940 36820 16952
rect 36872 16940 36878 16992
rect 38102 16940 38108 16992
rect 38160 16940 38166 16992
rect 1104 16890 49864 16912
rect 1104 16838 2950 16890
rect 3002 16838 3014 16890
rect 3066 16838 3078 16890
rect 3130 16838 3142 16890
rect 3194 16838 3206 16890
rect 3258 16838 12950 16890
rect 13002 16838 13014 16890
rect 13066 16838 13078 16890
rect 13130 16838 13142 16890
rect 13194 16838 13206 16890
rect 13258 16838 22950 16890
rect 23002 16838 23014 16890
rect 23066 16838 23078 16890
rect 23130 16838 23142 16890
rect 23194 16838 23206 16890
rect 23258 16838 32950 16890
rect 33002 16838 33014 16890
rect 33066 16838 33078 16890
rect 33130 16838 33142 16890
rect 33194 16838 33206 16890
rect 33258 16838 42950 16890
rect 43002 16838 43014 16890
rect 43066 16838 43078 16890
rect 43130 16838 43142 16890
rect 43194 16838 43206 16890
rect 43258 16838 49864 16890
rect 1104 16816 49864 16838
rect 19426 16736 19432 16788
rect 19484 16776 19490 16788
rect 19702 16785 19708 16788
rect 19686 16779 19708 16785
rect 19686 16776 19698 16779
rect 19484 16748 19698 16776
rect 19484 16736 19490 16748
rect 19686 16745 19698 16748
rect 19686 16739 19708 16745
rect 19702 16736 19708 16739
rect 19760 16736 19766 16788
rect 20070 16736 20076 16788
rect 20128 16776 20134 16788
rect 20128 16748 23428 16776
rect 20128 16736 20134 16748
rect 23400 16717 23428 16748
rect 24670 16736 24676 16788
rect 24728 16776 24734 16788
rect 26237 16779 26295 16785
rect 26237 16776 26249 16779
rect 24728 16748 26249 16776
rect 24728 16736 24734 16748
rect 26237 16745 26249 16748
rect 26283 16745 26295 16779
rect 36170 16776 36176 16788
rect 26237 16739 26295 16745
rect 34256 16748 36176 16776
rect 23385 16711 23443 16717
rect 23385 16677 23397 16711
rect 23431 16708 23443 16711
rect 23431 16680 25176 16708
rect 23431 16677 23443 16680
rect 23385 16671 23443 16677
rect 18598 16600 18604 16652
rect 18656 16640 18662 16652
rect 19242 16640 19248 16652
rect 18656 16612 19248 16640
rect 18656 16600 18662 16612
rect 19242 16600 19248 16612
rect 19300 16640 19306 16652
rect 19429 16643 19487 16649
rect 19429 16640 19441 16643
rect 19300 16612 19441 16640
rect 19300 16600 19306 16612
rect 19429 16609 19441 16612
rect 19475 16640 19487 16643
rect 21637 16643 21695 16649
rect 21637 16640 21649 16643
rect 19475 16612 21649 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 21637 16609 21649 16612
rect 21683 16640 21695 16643
rect 22462 16640 22468 16652
rect 21683 16612 22468 16640
rect 21683 16609 21695 16612
rect 21637 16603 21695 16609
rect 22462 16600 22468 16612
rect 22520 16600 22526 16652
rect 25038 16600 25044 16652
rect 25096 16600 25102 16652
rect 25148 16649 25176 16680
rect 25133 16643 25191 16649
rect 25133 16609 25145 16643
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 26694 16600 26700 16652
rect 26752 16640 26758 16652
rect 27709 16643 27767 16649
rect 27709 16640 27721 16643
rect 26752 16612 27721 16640
rect 26752 16600 26758 16612
rect 27709 16609 27721 16612
rect 27755 16609 27767 16643
rect 27709 16603 27767 16609
rect 34054 16600 34060 16652
rect 34112 16600 34118 16652
rect 34256 16649 34284 16748
rect 36170 16736 36176 16748
rect 36228 16776 36234 16788
rect 37090 16776 37096 16788
rect 36228 16748 37096 16776
rect 36228 16736 36234 16748
rect 37090 16736 37096 16748
rect 37148 16736 37154 16788
rect 34606 16668 34612 16720
rect 34664 16708 34670 16720
rect 34664 16680 35020 16708
rect 34664 16668 34670 16680
rect 34241 16643 34299 16649
rect 34241 16609 34253 16643
rect 34287 16609 34299 16643
rect 34241 16603 34299 16609
rect 34882 16600 34888 16652
rect 34940 16600 34946 16652
rect 34992 16640 35020 16680
rect 35161 16643 35219 16649
rect 35161 16640 35173 16643
rect 34992 16612 35173 16640
rect 35161 16609 35173 16612
rect 35207 16640 35219 16643
rect 35526 16640 35532 16652
rect 35207 16612 35532 16640
rect 35207 16609 35219 16612
rect 35161 16603 35219 16609
rect 35526 16600 35532 16612
rect 35584 16600 35590 16652
rect 37182 16600 37188 16652
rect 37240 16640 37246 16652
rect 38013 16643 38071 16649
rect 38013 16640 38025 16643
rect 37240 16612 38025 16640
rect 37240 16600 37246 16612
rect 38013 16609 38025 16612
rect 38059 16609 38071 16643
rect 38013 16603 38071 16609
rect 24578 16572 24584 16584
rect 23046 16544 24584 16572
rect 24578 16532 24584 16544
rect 24636 16532 24642 16584
rect 24949 16575 25007 16581
rect 24949 16541 24961 16575
rect 24995 16572 25007 16575
rect 25958 16572 25964 16584
rect 24995 16544 25964 16572
rect 24995 16541 25007 16544
rect 24949 16535 25007 16541
rect 25958 16532 25964 16544
rect 26016 16532 26022 16584
rect 26050 16532 26056 16584
rect 26108 16572 26114 16584
rect 26145 16575 26203 16581
rect 26145 16572 26157 16575
rect 26108 16544 26157 16572
rect 26108 16532 26114 16544
rect 26145 16541 26157 16544
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 28442 16572 28448 16584
rect 27571 16544 28448 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 28442 16532 28448 16544
rect 28500 16532 28506 16584
rect 30558 16532 30564 16584
rect 30616 16572 30622 16584
rect 33965 16575 34023 16581
rect 33965 16572 33977 16575
rect 30616 16544 33977 16572
rect 30616 16532 30622 16544
rect 33965 16541 33977 16544
rect 34011 16541 34023 16575
rect 33965 16535 34023 16541
rect 37826 16532 37832 16584
rect 37884 16572 37890 16584
rect 37921 16575 37979 16581
rect 37921 16572 37933 16575
rect 37884 16544 37933 16572
rect 37884 16532 37890 16544
rect 37921 16541 37933 16544
rect 37967 16541 37979 16575
rect 37921 16535 37979 16541
rect 46198 16532 46204 16584
rect 46256 16572 46262 16584
rect 47949 16575 48007 16581
rect 47949 16572 47961 16575
rect 46256 16544 47961 16572
rect 46256 16532 46262 16544
rect 47949 16541 47961 16544
rect 47995 16541 48007 16575
rect 47949 16535 48007 16541
rect 5537 16507 5595 16513
rect 5537 16473 5549 16507
rect 5583 16504 5595 16507
rect 9766 16504 9772 16516
rect 5583 16476 9772 16504
rect 5583 16473 5595 16476
rect 5537 16467 5595 16473
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 20088 16476 20194 16504
rect 21008 16476 21864 16504
rect 5626 16396 5632 16448
rect 5684 16396 5690 16448
rect 19242 16396 19248 16448
rect 19300 16436 19306 16448
rect 20088 16436 20116 16476
rect 20714 16436 20720 16448
rect 19300 16408 20720 16436
rect 19300 16396 19306 16408
rect 20714 16396 20720 16408
rect 20772 16436 20778 16448
rect 21008 16436 21036 16476
rect 20772 16408 21036 16436
rect 20772 16396 20778 16408
rect 21174 16396 21180 16448
rect 21232 16396 21238 16448
rect 21836 16436 21864 16476
rect 21910 16464 21916 16516
rect 21968 16464 21974 16516
rect 22020 16476 22402 16504
rect 23308 16476 24624 16504
rect 22020 16436 22048 16476
rect 21836 16408 22048 16436
rect 22094 16396 22100 16448
rect 22152 16436 22158 16448
rect 23308 16436 23336 16476
rect 24596 16445 24624 16476
rect 25774 16464 25780 16516
rect 25832 16504 25838 16516
rect 29454 16504 29460 16516
rect 25832 16476 29460 16504
rect 25832 16464 25838 16476
rect 29454 16464 29460 16476
rect 29512 16504 29518 16516
rect 31570 16504 31576 16516
rect 29512 16476 31576 16504
rect 29512 16464 29518 16476
rect 31570 16464 31576 16476
rect 31628 16464 31634 16516
rect 34514 16504 34520 16516
rect 33612 16476 34520 16504
rect 22152 16408 23336 16436
rect 24581 16439 24639 16445
rect 22152 16396 22158 16408
rect 24581 16405 24593 16439
rect 24627 16405 24639 16439
rect 24581 16399 24639 16405
rect 27154 16396 27160 16448
rect 27212 16396 27218 16448
rect 27522 16396 27528 16448
rect 27580 16436 27586 16448
rect 27617 16439 27675 16445
rect 27617 16436 27629 16439
rect 27580 16408 27629 16436
rect 27580 16396 27586 16408
rect 27617 16405 27629 16408
rect 27663 16405 27675 16439
rect 27617 16399 27675 16405
rect 28258 16396 28264 16448
rect 28316 16436 28322 16448
rect 28442 16436 28448 16448
rect 28316 16408 28448 16436
rect 28316 16396 28322 16408
rect 28442 16396 28448 16408
rect 28500 16396 28506 16448
rect 28534 16396 28540 16448
rect 28592 16436 28598 16448
rect 33134 16436 33140 16448
rect 28592 16408 33140 16436
rect 28592 16396 28598 16408
rect 33134 16396 33140 16408
rect 33192 16396 33198 16448
rect 33612 16445 33640 16476
rect 34514 16464 34520 16476
rect 34572 16464 34578 16516
rect 36446 16504 36452 16516
rect 36386 16476 36452 16504
rect 36446 16464 36452 16476
rect 36504 16464 36510 16516
rect 40126 16504 40132 16516
rect 37476 16476 40132 16504
rect 33597 16439 33655 16445
rect 33597 16405 33609 16439
rect 33643 16405 33655 16439
rect 33597 16399 33655 16405
rect 36630 16396 36636 16448
rect 36688 16436 36694 16448
rect 36906 16436 36912 16448
rect 36688 16408 36912 16436
rect 36688 16396 36694 16408
rect 36906 16396 36912 16408
rect 36964 16396 36970 16448
rect 37476 16445 37504 16476
rect 40126 16464 40132 16476
rect 40184 16464 40190 16516
rect 49142 16464 49148 16516
rect 49200 16464 49206 16516
rect 37461 16439 37519 16445
rect 37461 16405 37473 16439
rect 37507 16405 37519 16439
rect 37461 16399 37519 16405
rect 37829 16439 37887 16445
rect 37829 16405 37841 16439
rect 37875 16436 37887 16439
rect 38102 16436 38108 16448
rect 37875 16408 38108 16436
rect 37875 16405 37887 16408
rect 37829 16399 37887 16405
rect 38102 16396 38108 16408
rect 38160 16396 38166 16448
rect 1104 16346 49864 16368
rect 1104 16294 7950 16346
rect 8002 16294 8014 16346
rect 8066 16294 8078 16346
rect 8130 16294 8142 16346
rect 8194 16294 8206 16346
rect 8258 16294 17950 16346
rect 18002 16294 18014 16346
rect 18066 16294 18078 16346
rect 18130 16294 18142 16346
rect 18194 16294 18206 16346
rect 18258 16294 27950 16346
rect 28002 16294 28014 16346
rect 28066 16294 28078 16346
rect 28130 16294 28142 16346
rect 28194 16294 28206 16346
rect 28258 16294 37950 16346
rect 38002 16294 38014 16346
rect 38066 16294 38078 16346
rect 38130 16294 38142 16346
rect 38194 16294 38206 16346
rect 38258 16294 47950 16346
rect 48002 16294 48014 16346
rect 48066 16294 48078 16346
rect 48130 16294 48142 16346
rect 48194 16294 48206 16346
rect 48258 16294 49864 16346
rect 1104 16272 49864 16294
rect 18782 16192 18788 16244
rect 18840 16232 18846 16244
rect 25685 16235 25743 16241
rect 25685 16232 25697 16235
rect 18840 16204 25697 16232
rect 18840 16192 18846 16204
rect 25685 16201 25697 16204
rect 25731 16201 25743 16235
rect 25685 16195 25743 16201
rect 25774 16192 25780 16244
rect 25832 16192 25838 16244
rect 25866 16192 25872 16244
rect 25924 16232 25930 16244
rect 27157 16235 27215 16241
rect 27157 16232 27169 16235
rect 25924 16204 27169 16232
rect 25924 16192 25930 16204
rect 27157 16201 27169 16204
rect 27203 16201 27215 16235
rect 27157 16195 27215 16201
rect 27246 16192 27252 16244
rect 27304 16232 27310 16244
rect 27525 16235 27583 16241
rect 27525 16232 27537 16235
rect 27304 16204 27537 16232
rect 27304 16192 27310 16204
rect 27525 16201 27537 16204
rect 27571 16232 27583 16235
rect 29730 16232 29736 16244
rect 27571 16204 29736 16232
rect 27571 16201 27583 16204
rect 27525 16195 27583 16201
rect 29730 16192 29736 16204
rect 29788 16192 29794 16244
rect 32953 16235 33011 16241
rect 32953 16201 32965 16235
rect 32999 16232 33011 16235
rect 32999 16204 35894 16232
rect 32999 16201 33011 16204
rect 32953 16195 33011 16201
rect 16390 16124 16396 16176
rect 16448 16164 16454 16176
rect 23017 16167 23075 16173
rect 23017 16164 23029 16167
rect 16448 16136 23029 16164
rect 16448 16124 16454 16136
rect 23017 16133 23029 16136
rect 23063 16133 23075 16167
rect 24578 16164 24584 16176
rect 24242 16136 24584 16164
rect 23017 16127 23075 16133
rect 24578 16124 24584 16136
rect 24636 16124 24642 16176
rect 24762 16124 24768 16176
rect 24820 16124 24826 16176
rect 29362 16164 29368 16176
rect 27632 16136 29368 16164
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16096 1823 16099
rect 2774 16096 2780 16108
rect 1811 16068 2780 16096
rect 1811 16065 1823 16068
rect 1765 16059 1823 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 22462 16056 22468 16108
rect 22520 16096 22526 16108
rect 22741 16099 22799 16105
rect 22741 16096 22753 16099
rect 22520 16068 22753 16096
rect 22520 16056 22526 16068
rect 22741 16065 22753 16068
rect 22787 16065 22799 16099
rect 22741 16059 22799 16065
rect 26050 16056 26056 16108
rect 26108 16096 26114 16108
rect 27632 16105 27660 16136
rect 29362 16124 29368 16136
rect 29420 16124 29426 16176
rect 30466 16164 30472 16176
rect 30314 16136 30472 16164
rect 30466 16124 30472 16136
rect 30524 16124 30530 16176
rect 33410 16164 33416 16176
rect 31726 16136 33416 16164
rect 27617 16099 27675 16105
rect 27617 16096 27629 16099
rect 26108 16068 27629 16096
rect 26108 16056 26114 16068
rect 27617 16065 27629 16068
rect 27663 16065 27675 16099
rect 28810 16096 28816 16108
rect 27617 16059 27675 16065
rect 27816 16068 28816 16096
rect 1302 15988 1308 16040
rect 1360 16028 1366 16040
rect 2041 16031 2099 16037
rect 2041 16028 2053 16031
rect 1360 16000 2053 16028
rect 1360 15988 1366 16000
rect 2041 15997 2053 16000
rect 2087 15997 2099 16031
rect 2041 15991 2099 15997
rect 25961 16031 26019 16037
rect 25961 15997 25973 16031
rect 26007 16028 26019 16031
rect 26142 16028 26148 16040
rect 26007 16000 26148 16028
rect 26007 15997 26019 16000
rect 25961 15991 26019 15997
rect 26142 15988 26148 16000
rect 26200 15988 26206 16040
rect 27430 15988 27436 16040
rect 27488 16028 27494 16040
rect 27709 16031 27767 16037
rect 27709 16028 27721 16031
rect 27488 16000 27721 16028
rect 27488 15988 27494 16000
rect 27709 15997 27721 16000
rect 27755 15997 27767 16031
rect 27709 15991 27767 15997
rect 27614 15920 27620 15972
rect 27672 15960 27678 15972
rect 27816 15960 27844 16068
rect 28810 16056 28816 16068
rect 28868 16056 28874 16108
rect 29089 16031 29147 16037
rect 29089 15997 29101 16031
rect 29135 16028 29147 16031
rect 29178 16028 29184 16040
rect 29135 16000 29184 16028
rect 29135 15997 29147 16000
rect 29089 15991 29147 15997
rect 29178 15988 29184 16000
rect 29236 15988 29242 16040
rect 29454 15988 29460 16040
rect 29512 16028 29518 16040
rect 31726 16028 31754 16136
rect 33410 16124 33416 16136
rect 33468 16124 33474 16176
rect 35866 16164 35894 16204
rect 37366 16164 37372 16176
rect 35866 16136 37372 16164
rect 37366 16124 37372 16136
rect 37424 16124 37430 16176
rect 33321 16099 33379 16105
rect 33321 16065 33333 16099
rect 33367 16096 33379 16099
rect 34333 16099 34391 16105
rect 34333 16096 34345 16099
rect 33367 16068 34345 16096
rect 33367 16065 33379 16068
rect 33321 16059 33379 16065
rect 34333 16065 34345 16068
rect 34379 16065 34391 16099
rect 34333 16059 34391 16065
rect 36265 16099 36323 16105
rect 36265 16065 36277 16099
rect 36311 16096 36323 16099
rect 36354 16096 36360 16108
rect 36311 16068 36360 16096
rect 36311 16065 36323 16068
rect 36265 16059 36323 16065
rect 36354 16056 36360 16068
rect 36412 16056 36418 16108
rect 38841 16099 38899 16105
rect 38841 16065 38853 16099
rect 38887 16096 38899 16099
rect 40034 16096 40040 16108
rect 38887 16068 40040 16096
rect 38887 16065 38899 16068
rect 38841 16059 38899 16065
rect 40034 16056 40040 16068
rect 40092 16056 40098 16108
rect 47854 16056 47860 16108
rect 47912 16096 47918 16108
rect 47949 16099 48007 16105
rect 47949 16096 47961 16099
rect 47912 16068 47961 16096
rect 47912 16056 47918 16068
rect 47949 16065 47961 16068
rect 47995 16065 48007 16099
rect 47949 16059 48007 16065
rect 29512 16000 31754 16028
rect 29512 15988 29518 16000
rect 33134 15988 33140 16040
rect 33192 16028 33198 16040
rect 33413 16031 33471 16037
rect 33413 16028 33425 16031
rect 33192 16000 33425 16028
rect 33192 15988 33198 16000
rect 33413 15997 33425 16000
rect 33459 15997 33471 16031
rect 33413 15991 33471 15997
rect 33597 16031 33655 16037
rect 33597 15997 33609 16031
rect 33643 16028 33655 16031
rect 37550 16028 37556 16040
rect 33643 16000 37556 16028
rect 33643 15997 33655 16000
rect 33597 15991 33655 15997
rect 37550 15988 37556 16000
rect 37608 15988 37614 16040
rect 49142 15988 49148 16040
rect 49200 15988 49206 16040
rect 27672 15932 27844 15960
rect 27672 15920 27678 15932
rect 30190 15920 30196 15972
rect 30248 15960 30254 15972
rect 33226 15960 33232 15972
rect 30248 15932 33232 15960
rect 30248 15920 30254 15932
rect 33226 15920 33232 15932
rect 33284 15920 33290 15972
rect 33318 15920 33324 15972
rect 33376 15960 33382 15972
rect 39114 15960 39120 15972
rect 33376 15932 39120 15960
rect 33376 15920 33382 15932
rect 39114 15920 39120 15932
rect 39172 15920 39178 15972
rect 25317 15895 25375 15901
rect 25317 15861 25329 15895
rect 25363 15892 25375 15895
rect 29822 15892 29828 15904
rect 25363 15864 29828 15892
rect 25363 15861 25375 15864
rect 25317 15855 25375 15861
rect 29822 15852 29828 15864
rect 29880 15852 29886 15904
rect 30098 15852 30104 15904
rect 30156 15892 30162 15904
rect 30561 15895 30619 15901
rect 30561 15892 30573 15895
rect 30156 15864 30573 15892
rect 30156 15852 30162 15864
rect 30561 15861 30573 15864
rect 30607 15892 30619 15895
rect 32858 15892 32864 15904
rect 30607 15864 32864 15892
rect 30607 15861 30619 15864
rect 30561 15855 30619 15861
rect 32858 15852 32864 15864
rect 32916 15852 32922 15904
rect 33410 15852 33416 15904
rect 33468 15892 33474 15904
rect 34977 15895 35035 15901
rect 34977 15892 34989 15895
rect 33468 15864 34989 15892
rect 33468 15852 33474 15864
rect 34977 15861 34989 15864
rect 35023 15861 35035 15895
rect 34977 15855 35035 15861
rect 36078 15852 36084 15904
rect 36136 15852 36142 15904
rect 37642 15852 37648 15904
rect 37700 15852 37706 15904
rect 37826 15852 37832 15904
rect 37884 15892 37890 15904
rect 38657 15895 38715 15901
rect 38657 15892 38669 15895
rect 37884 15864 38669 15892
rect 37884 15852 37890 15864
rect 38657 15861 38669 15864
rect 38703 15861 38715 15895
rect 38657 15855 38715 15861
rect 1104 15802 49864 15824
rect 1104 15750 2950 15802
rect 3002 15750 3014 15802
rect 3066 15750 3078 15802
rect 3130 15750 3142 15802
rect 3194 15750 3206 15802
rect 3258 15750 12950 15802
rect 13002 15750 13014 15802
rect 13066 15750 13078 15802
rect 13130 15750 13142 15802
rect 13194 15750 13206 15802
rect 13258 15750 22950 15802
rect 23002 15750 23014 15802
rect 23066 15750 23078 15802
rect 23130 15750 23142 15802
rect 23194 15750 23206 15802
rect 23258 15750 32950 15802
rect 33002 15750 33014 15802
rect 33066 15750 33078 15802
rect 33130 15750 33142 15802
rect 33194 15750 33206 15802
rect 33258 15750 42950 15802
rect 43002 15750 43014 15802
rect 43066 15750 43078 15802
rect 43130 15750 43142 15802
rect 43194 15750 43206 15802
rect 43258 15750 49864 15802
rect 1104 15728 49864 15750
rect 26418 15648 26424 15700
rect 26476 15648 26482 15700
rect 30190 15688 30196 15700
rect 28092 15660 30196 15688
rect 23382 15512 23388 15564
rect 23440 15552 23446 15564
rect 28092 15561 28120 15660
rect 30190 15648 30196 15660
rect 30248 15648 30254 15700
rect 33045 15691 33103 15697
rect 33045 15657 33057 15691
rect 33091 15688 33103 15691
rect 33318 15688 33324 15700
rect 33091 15660 33324 15688
rect 33091 15657 33103 15660
rect 33045 15651 33103 15657
rect 33318 15648 33324 15660
rect 33376 15648 33382 15700
rect 29181 15623 29239 15629
rect 29181 15589 29193 15623
rect 29227 15620 29239 15623
rect 29454 15620 29460 15632
rect 29227 15592 29460 15620
rect 29227 15589 29239 15592
rect 29181 15583 29239 15589
rect 29454 15580 29460 15592
rect 29512 15580 29518 15632
rect 32306 15580 32312 15632
rect 32364 15620 32370 15632
rect 32582 15620 32588 15632
rect 32364 15592 32588 15620
rect 32364 15580 32370 15592
rect 32582 15580 32588 15592
rect 32640 15580 32646 15632
rect 26973 15555 27031 15561
rect 26973 15552 26985 15555
rect 23440 15524 26985 15552
rect 23440 15512 23446 15524
rect 26973 15521 26985 15524
rect 27019 15521 27031 15555
rect 26973 15515 27031 15521
rect 28077 15555 28135 15561
rect 28077 15521 28089 15555
rect 28123 15521 28135 15555
rect 28077 15515 28135 15521
rect 28261 15555 28319 15561
rect 28261 15521 28273 15555
rect 28307 15552 28319 15555
rect 28307 15524 28764 15552
rect 28307 15521 28319 15524
rect 28261 15515 28319 15521
rect 19886 15444 19892 15496
rect 19944 15484 19950 15496
rect 20530 15484 20536 15496
rect 19944 15456 20536 15484
rect 19944 15444 19950 15456
rect 20530 15444 20536 15456
rect 20588 15484 20594 15496
rect 27985 15487 28043 15493
rect 27985 15484 27997 15487
rect 20588 15456 27997 15484
rect 20588 15444 20594 15456
rect 27985 15453 27997 15456
rect 28031 15453 28043 15487
rect 27985 15447 28043 15453
rect 24673 15419 24731 15425
rect 24673 15385 24685 15419
rect 24719 15416 24731 15419
rect 25222 15416 25228 15428
rect 24719 15388 25228 15416
rect 24719 15385 24731 15388
rect 24673 15379 24731 15385
rect 25222 15376 25228 15388
rect 25280 15376 25286 15428
rect 26789 15419 26847 15425
rect 26789 15385 26801 15419
rect 26835 15416 26847 15419
rect 27246 15416 27252 15428
rect 26835 15388 27252 15416
rect 26835 15385 26847 15388
rect 26789 15379 26847 15385
rect 27246 15376 27252 15388
rect 27304 15376 27310 15428
rect 28736 15416 28764 15524
rect 28810 15512 28816 15564
rect 28868 15552 28874 15564
rect 29733 15555 29791 15561
rect 29733 15552 29745 15555
rect 28868 15524 29745 15552
rect 28868 15512 28874 15524
rect 29733 15521 29745 15524
rect 29779 15552 29791 15555
rect 30006 15552 30012 15564
rect 29779 15524 30012 15552
rect 29779 15521 29791 15524
rect 29733 15515 29791 15521
rect 30006 15512 30012 15524
rect 30064 15512 30070 15564
rect 33594 15512 33600 15564
rect 33652 15512 33658 15564
rect 35894 15512 35900 15564
rect 35952 15512 35958 15564
rect 36170 15512 36176 15564
rect 36228 15512 36234 15564
rect 28994 15444 29000 15496
rect 29052 15444 29058 15496
rect 32490 15444 32496 15496
rect 32548 15484 32554 15496
rect 32585 15487 32643 15493
rect 32585 15484 32597 15487
rect 32548 15456 32597 15484
rect 32548 15444 32554 15456
rect 32585 15453 32597 15456
rect 32631 15453 32643 15487
rect 32585 15447 32643 15453
rect 33410 15444 33416 15496
rect 33468 15444 33474 15496
rect 33505 15487 33563 15493
rect 33505 15453 33517 15487
rect 33551 15484 33563 15487
rect 33686 15484 33692 15496
rect 33551 15456 33692 15484
rect 33551 15453 33563 15456
rect 33505 15447 33563 15453
rect 33686 15444 33692 15456
rect 33744 15444 33750 15496
rect 46842 15444 46848 15496
rect 46900 15484 46906 15496
rect 47949 15487 48007 15493
rect 47949 15484 47961 15487
rect 46900 15456 47961 15484
rect 46900 15444 46906 15456
rect 47949 15453 47961 15456
rect 47995 15453 48007 15487
rect 47949 15447 48007 15453
rect 29178 15416 29184 15428
rect 28736 15388 29184 15416
rect 29178 15376 29184 15388
rect 29236 15376 29242 15428
rect 29638 15416 29644 15428
rect 29380 15388 29644 15416
rect 22646 15308 22652 15360
rect 22704 15348 22710 15360
rect 24765 15351 24823 15357
rect 24765 15348 24777 15351
rect 22704 15320 24777 15348
rect 22704 15308 22710 15320
rect 24765 15317 24777 15320
rect 24811 15317 24823 15351
rect 24765 15311 24823 15317
rect 25590 15308 25596 15360
rect 25648 15348 25654 15360
rect 26050 15348 26056 15360
rect 25648 15320 26056 15348
rect 25648 15308 25654 15320
rect 26050 15308 26056 15320
rect 26108 15348 26114 15360
rect 26881 15351 26939 15357
rect 26881 15348 26893 15351
rect 26108 15320 26893 15348
rect 26108 15308 26114 15320
rect 26881 15317 26893 15320
rect 26927 15317 26939 15351
rect 26881 15311 26939 15317
rect 27617 15351 27675 15357
rect 27617 15317 27629 15351
rect 27663 15348 27675 15351
rect 29380 15348 29408 15388
rect 29638 15376 29644 15388
rect 29696 15376 29702 15428
rect 30009 15419 30067 15425
rect 30009 15385 30021 15419
rect 30055 15416 30067 15419
rect 30098 15416 30104 15428
rect 30055 15388 30104 15416
rect 30055 15385 30067 15388
rect 30009 15379 30067 15385
rect 30098 15376 30104 15388
rect 30156 15376 30162 15428
rect 30466 15416 30472 15428
rect 30208 15388 30472 15416
rect 27663 15320 29408 15348
rect 27663 15317 27675 15320
rect 27617 15311 27675 15317
rect 29454 15308 29460 15360
rect 29512 15348 29518 15360
rect 30208 15348 30236 15388
rect 30466 15376 30472 15388
rect 30524 15376 30530 15428
rect 36446 15376 36452 15428
rect 36504 15416 36510 15428
rect 36630 15416 36636 15428
rect 36504 15388 36636 15416
rect 36504 15376 36510 15388
rect 36630 15376 36636 15388
rect 36688 15376 36694 15428
rect 49142 15376 49148 15428
rect 49200 15376 49206 15428
rect 29512 15320 30236 15348
rect 29512 15308 29518 15320
rect 30282 15308 30288 15360
rect 30340 15348 30346 15360
rect 31481 15351 31539 15357
rect 31481 15348 31493 15351
rect 30340 15320 31493 15348
rect 30340 15308 30346 15320
rect 31481 15317 31493 15320
rect 31527 15317 31539 15351
rect 31481 15311 31539 15317
rect 31570 15308 31576 15360
rect 31628 15348 31634 15360
rect 31754 15348 31760 15360
rect 31628 15320 31760 15348
rect 31628 15308 31634 15320
rect 31754 15308 31760 15320
rect 31812 15308 31818 15360
rect 32398 15308 32404 15360
rect 32456 15308 32462 15360
rect 37645 15351 37703 15357
rect 37645 15317 37657 15351
rect 37691 15348 37703 15351
rect 37734 15348 37740 15360
rect 37691 15320 37740 15348
rect 37691 15317 37703 15320
rect 37645 15311 37703 15317
rect 37734 15308 37740 15320
rect 37792 15308 37798 15360
rect 1104 15258 49864 15280
rect 1104 15206 7950 15258
rect 8002 15206 8014 15258
rect 8066 15206 8078 15258
rect 8130 15206 8142 15258
rect 8194 15206 8206 15258
rect 8258 15206 17950 15258
rect 18002 15206 18014 15258
rect 18066 15206 18078 15258
rect 18130 15206 18142 15258
rect 18194 15206 18206 15258
rect 18258 15206 27950 15258
rect 28002 15206 28014 15258
rect 28066 15206 28078 15258
rect 28130 15206 28142 15258
rect 28194 15206 28206 15258
rect 28258 15206 37950 15258
rect 38002 15206 38014 15258
rect 38066 15206 38078 15258
rect 38130 15206 38142 15258
rect 38194 15206 38206 15258
rect 38258 15206 47950 15258
rect 48002 15206 48014 15258
rect 48066 15206 48078 15258
rect 48130 15206 48142 15258
rect 48194 15206 48206 15258
rect 48258 15206 49864 15258
rect 1104 15184 49864 15206
rect 19334 15104 19340 15156
rect 19392 15144 19398 15156
rect 20901 15147 20959 15153
rect 20901 15144 20913 15147
rect 19392 15116 20913 15144
rect 19392 15104 19398 15116
rect 20901 15113 20913 15116
rect 20947 15113 20959 15147
rect 20901 15107 20959 15113
rect 25038 15104 25044 15156
rect 25096 15144 25102 15156
rect 25869 15147 25927 15153
rect 25869 15144 25881 15147
rect 25096 15116 25881 15144
rect 25096 15104 25102 15116
rect 25869 15113 25881 15116
rect 25915 15113 25927 15147
rect 25869 15107 25927 15113
rect 29178 15104 29184 15156
rect 29236 15144 29242 15156
rect 29365 15147 29423 15153
rect 29365 15144 29377 15147
rect 29236 15116 29377 15144
rect 29236 15104 29242 15116
rect 29365 15113 29377 15116
rect 29411 15113 29423 15147
rect 29365 15107 29423 15113
rect 29638 15104 29644 15156
rect 29696 15144 29702 15156
rect 32769 15147 32827 15153
rect 32769 15144 32781 15147
rect 29696 15116 32781 15144
rect 29696 15104 29702 15116
rect 32769 15113 32781 15116
rect 32815 15113 32827 15147
rect 32769 15107 32827 15113
rect 37642 15104 37648 15156
rect 37700 15144 37706 15156
rect 37829 15147 37887 15153
rect 37829 15144 37841 15147
rect 37700 15116 37841 15144
rect 37700 15104 37706 15116
rect 37829 15113 37841 15116
rect 37875 15113 37887 15147
rect 37829 15107 37887 15113
rect 24578 15076 24584 15088
rect 23966 15048 24584 15076
rect 24578 15036 24584 15048
rect 24636 15036 24642 15088
rect 26237 15079 26295 15085
rect 26237 15045 26249 15079
rect 26283 15076 26295 15079
rect 27798 15076 27804 15088
rect 26283 15048 27804 15076
rect 26283 15045 26295 15048
rect 26237 15039 26295 15045
rect 27798 15036 27804 15048
rect 27856 15036 27862 15088
rect 29454 15076 29460 15088
rect 29118 15048 29460 15076
rect 29454 15036 29460 15048
rect 29512 15036 29518 15088
rect 29914 15036 29920 15088
rect 29972 15036 29978 15088
rect 31478 15036 31484 15088
rect 31536 15076 31542 15088
rect 31573 15079 31631 15085
rect 31573 15076 31585 15079
rect 31536 15048 31585 15076
rect 31536 15036 31542 15048
rect 31573 15045 31585 15048
rect 31619 15045 31631 15079
rect 31573 15039 31631 15045
rect 36814 15036 36820 15088
rect 36872 15076 36878 15088
rect 37921 15079 37979 15085
rect 37921 15076 37933 15079
rect 36872 15048 37933 15076
rect 36872 15036 36878 15048
rect 37921 15045 37933 15048
rect 37967 15045 37979 15079
rect 37921 15039 37979 15045
rect 17862 14968 17868 15020
rect 17920 15008 17926 15020
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 17920 14980 20821 15008
rect 17920 14968 17926 14980
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 22462 14968 22468 15020
rect 22520 14968 22526 15020
rect 25682 14968 25688 15020
rect 25740 15008 25746 15020
rect 27614 15008 27620 15020
rect 25740 14980 27620 15008
rect 25740 14968 25746 14980
rect 27614 14968 27620 14980
rect 27672 14968 27678 15020
rect 32214 14968 32220 15020
rect 32272 15008 32278 15020
rect 32677 15011 32735 15017
rect 32677 15008 32689 15011
rect 32272 14980 32689 15008
rect 32272 14968 32278 14980
rect 32677 14977 32689 14980
rect 32723 14977 32735 15011
rect 32677 14971 32735 14977
rect 41782 14968 41788 15020
rect 41840 14968 41846 15020
rect 46750 14968 46756 15020
rect 46808 15008 46814 15020
rect 47949 15011 48007 15017
rect 47949 15008 47961 15011
rect 46808 14980 47961 15008
rect 46808 14968 46814 14980
rect 47949 14977 47961 14980
rect 47995 14977 48007 15011
rect 47949 14971 48007 14977
rect 21085 14943 21143 14949
rect 21085 14909 21097 14943
rect 21131 14940 21143 14943
rect 21174 14940 21180 14952
rect 21131 14912 21180 14940
rect 21131 14909 21143 14912
rect 21085 14903 21143 14909
rect 21174 14900 21180 14912
rect 21232 14940 21238 14952
rect 22741 14943 22799 14949
rect 22741 14940 22753 14943
rect 21232 14912 22753 14940
rect 21232 14900 21238 14912
rect 22741 14909 22753 14912
rect 22787 14909 22799 14943
rect 22741 14903 22799 14909
rect 24213 14943 24271 14949
rect 24213 14909 24225 14943
rect 24259 14940 24271 14943
rect 26142 14940 26148 14952
rect 24259 14912 26148 14940
rect 24259 14909 24271 14912
rect 24213 14903 24271 14909
rect 26142 14900 26148 14912
rect 26200 14900 26206 14952
rect 26329 14943 26387 14949
rect 26329 14909 26341 14943
rect 26375 14909 26387 14943
rect 26329 14903 26387 14909
rect 26513 14943 26571 14949
rect 26513 14909 26525 14943
rect 26559 14940 26571 14943
rect 26602 14940 26608 14952
rect 26559 14912 26608 14940
rect 26559 14909 26571 14912
rect 26513 14903 26571 14909
rect 20438 14764 20444 14816
rect 20496 14764 20502 14816
rect 26344 14804 26372 14903
rect 26602 14900 26608 14912
rect 26660 14900 26666 14952
rect 27890 14900 27896 14952
rect 27948 14900 27954 14952
rect 30101 14943 30159 14949
rect 30101 14909 30113 14943
rect 30147 14940 30159 14943
rect 32122 14940 32128 14952
rect 30147 14912 32128 14940
rect 30147 14909 30159 14912
rect 30101 14903 30159 14909
rect 32122 14900 32128 14912
rect 32180 14900 32186 14952
rect 32858 14900 32864 14952
rect 32916 14900 32922 14952
rect 36906 14900 36912 14952
rect 36964 14940 36970 14952
rect 38013 14943 38071 14949
rect 38013 14940 38025 14943
rect 36964 14912 38025 14940
rect 36964 14900 36970 14912
rect 38013 14909 38025 14912
rect 38059 14909 38071 14943
rect 38013 14903 38071 14909
rect 49142 14900 49148 14952
rect 49200 14900 49206 14952
rect 31757 14875 31815 14881
rect 31757 14841 31769 14875
rect 31803 14841 31815 14875
rect 31757 14835 31815 14841
rect 32309 14875 32367 14881
rect 32309 14841 32321 14875
rect 32355 14872 32367 14875
rect 38286 14872 38292 14884
rect 32355 14844 38292 14872
rect 32355 14841 32367 14844
rect 32309 14835 32367 14841
rect 30006 14804 30012 14816
rect 26344 14776 30012 14804
rect 30006 14764 30012 14776
rect 30064 14764 30070 14816
rect 30190 14764 30196 14816
rect 30248 14804 30254 14816
rect 30745 14807 30803 14813
rect 30745 14804 30757 14807
rect 30248 14776 30757 14804
rect 30248 14764 30254 14776
rect 30745 14773 30757 14776
rect 30791 14773 30803 14807
rect 31772 14804 31800 14835
rect 38286 14832 38292 14844
rect 38344 14832 38350 14884
rect 33778 14804 33784 14816
rect 31772 14776 33784 14804
rect 30745 14767 30803 14773
rect 33778 14764 33784 14776
rect 33836 14764 33842 14816
rect 37461 14807 37519 14813
rect 37461 14773 37473 14807
rect 37507 14804 37519 14807
rect 41230 14804 41236 14816
rect 37507 14776 41236 14804
rect 37507 14773 37519 14776
rect 37461 14767 37519 14773
rect 41230 14764 41236 14776
rect 41288 14764 41294 14816
rect 41601 14807 41659 14813
rect 41601 14773 41613 14807
rect 41647 14804 41659 14807
rect 44174 14804 44180 14816
rect 41647 14776 44180 14804
rect 41647 14773 41659 14776
rect 41601 14767 41659 14773
rect 44174 14764 44180 14776
rect 44232 14764 44238 14816
rect 1104 14714 49864 14736
rect 1104 14662 2950 14714
rect 3002 14662 3014 14714
rect 3066 14662 3078 14714
rect 3130 14662 3142 14714
rect 3194 14662 3206 14714
rect 3258 14662 12950 14714
rect 13002 14662 13014 14714
rect 13066 14662 13078 14714
rect 13130 14662 13142 14714
rect 13194 14662 13206 14714
rect 13258 14662 22950 14714
rect 23002 14662 23014 14714
rect 23066 14662 23078 14714
rect 23130 14662 23142 14714
rect 23194 14662 23206 14714
rect 23258 14662 32950 14714
rect 33002 14662 33014 14714
rect 33066 14662 33078 14714
rect 33130 14662 33142 14714
rect 33194 14662 33206 14714
rect 33258 14662 42950 14714
rect 43002 14662 43014 14714
rect 43066 14662 43078 14714
rect 43130 14662 43142 14714
rect 43194 14662 43206 14714
rect 43258 14662 49864 14714
rect 1104 14640 49864 14662
rect 20438 14560 20444 14612
rect 20496 14600 20502 14612
rect 26326 14600 26332 14612
rect 20496 14572 26332 14600
rect 20496 14560 20502 14572
rect 26326 14560 26332 14572
rect 26384 14560 26390 14612
rect 27617 14603 27675 14609
rect 27617 14569 27629 14603
rect 27663 14600 27675 14603
rect 27890 14600 27896 14612
rect 27663 14572 27896 14600
rect 27663 14569 27675 14572
rect 27617 14563 27675 14569
rect 27890 14560 27896 14572
rect 27948 14600 27954 14612
rect 27948 14572 28488 14600
rect 27948 14560 27954 14572
rect 25682 14424 25688 14476
rect 25740 14464 25746 14476
rect 25869 14467 25927 14473
rect 25869 14464 25881 14467
rect 25740 14436 25881 14464
rect 25740 14424 25746 14436
rect 25869 14433 25881 14436
rect 25915 14433 25927 14467
rect 28460 14464 28488 14572
rect 32214 14560 32220 14612
rect 32272 14560 32278 14612
rect 32677 14535 32735 14541
rect 32677 14501 32689 14535
rect 32723 14532 32735 14535
rect 34330 14532 34336 14544
rect 32723 14504 34336 14532
rect 32723 14501 32735 14504
rect 32677 14495 32735 14501
rect 34330 14492 34336 14504
rect 34388 14492 34394 14544
rect 37185 14535 37243 14541
rect 37185 14501 37197 14535
rect 37231 14532 37243 14535
rect 41322 14532 41328 14544
rect 37231 14504 41328 14532
rect 37231 14501 37243 14504
rect 37185 14495 37243 14501
rect 41322 14492 41328 14504
rect 41380 14492 41386 14544
rect 30377 14467 30435 14473
rect 30377 14464 30389 14467
rect 28460 14436 30389 14464
rect 25869 14427 25927 14433
rect 30377 14433 30389 14436
rect 30423 14433 30435 14467
rect 30377 14427 30435 14433
rect 31754 14424 31760 14476
rect 31812 14464 31818 14476
rect 33137 14467 33195 14473
rect 33137 14464 33149 14467
rect 31812 14436 33149 14464
rect 31812 14424 31818 14436
rect 33137 14433 33149 14436
rect 33183 14433 33195 14467
rect 33137 14427 33195 14433
rect 33321 14467 33379 14473
rect 33321 14433 33333 14467
rect 33367 14464 33379 14467
rect 33962 14464 33968 14476
rect 33367 14436 33968 14464
rect 33367 14433 33379 14436
rect 33321 14427 33379 14433
rect 33962 14424 33968 14436
rect 34020 14424 34026 14476
rect 34514 14424 34520 14476
rect 34572 14464 34578 14476
rect 37645 14467 37703 14473
rect 37645 14464 37657 14467
rect 34572 14436 37657 14464
rect 34572 14424 34578 14436
rect 37645 14433 37657 14436
rect 37691 14433 37703 14467
rect 37645 14427 37703 14433
rect 37734 14424 37740 14476
rect 37792 14424 37798 14476
rect 30190 14356 30196 14408
rect 30248 14356 30254 14408
rect 30282 14356 30288 14408
rect 30340 14396 30346 14408
rect 33045 14399 33103 14405
rect 33045 14396 33057 14399
rect 30340 14368 33057 14396
rect 30340 14356 30346 14368
rect 33045 14365 33057 14368
rect 33091 14365 33103 14399
rect 33045 14359 33103 14365
rect 34238 14356 34244 14408
rect 34296 14396 34302 14408
rect 34977 14399 35035 14405
rect 34977 14396 34989 14399
rect 34296 14368 34989 14396
rect 34296 14356 34302 14368
rect 34977 14365 34989 14368
rect 35023 14365 35035 14399
rect 34977 14359 35035 14365
rect 37553 14399 37611 14405
rect 37553 14365 37565 14399
rect 37599 14396 37611 14399
rect 38565 14399 38623 14405
rect 38565 14396 38577 14399
rect 37599 14368 38577 14396
rect 37599 14365 37611 14368
rect 37553 14359 37611 14365
rect 38565 14365 38577 14368
rect 38611 14365 38623 14399
rect 38565 14359 38623 14365
rect 40034 14356 40040 14408
rect 40092 14356 40098 14408
rect 40218 14356 40224 14408
rect 40276 14356 40282 14408
rect 26142 14288 26148 14340
rect 26200 14288 26206 14340
rect 29454 14328 29460 14340
rect 27370 14300 29460 14328
rect 29454 14288 29460 14300
rect 29512 14288 29518 14340
rect 29840 14300 33272 14328
rect 29840 14269 29868 14300
rect 29825 14263 29883 14269
rect 29825 14229 29837 14263
rect 29871 14229 29883 14263
rect 29825 14223 29883 14229
rect 29914 14220 29920 14272
rect 29972 14260 29978 14272
rect 30285 14263 30343 14269
rect 30285 14260 30297 14263
rect 29972 14232 30297 14260
rect 29972 14220 29978 14232
rect 30285 14229 30297 14232
rect 30331 14229 30343 14263
rect 33244 14260 33272 14300
rect 35158 14288 35164 14340
rect 35216 14288 35222 14340
rect 37734 14288 37740 14340
rect 37792 14328 37798 14340
rect 40052 14328 40080 14356
rect 37792 14300 40080 14328
rect 37792 14288 37798 14300
rect 36906 14260 36912 14272
rect 33244 14232 36912 14260
rect 30285 14223 30343 14229
rect 36906 14220 36912 14232
rect 36964 14220 36970 14272
rect 40037 14263 40095 14269
rect 40037 14229 40049 14263
rect 40083 14260 40095 14263
rect 42794 14260 42800 14272
rect 40083 14232 42800 14260
rect 40083 14229 40095 14232
rect 40037 14223 40095 14229
rect 42794 14220 42800 14232
rect 42852 14220 42858 14272
rect 1104 14170 49864 14192
rect 1104 14118 7950 14170
rect 8002 14118 8014 14170
rect 8066 14118 8078 14170
rect 8130 14118 8142 14170
rect 8194 14118 8206 14170
rect 8258 14118 17950 14170
rect 18002 14118 18014 14170
rect 18066 14118 18078 14170
rect 18130 14118 18142 14170
rect 18194 14118 18206 14170
rect 18258 14118 27950 14170
rect 28002 14118 28014 14170
rect 28066 14118 28078 14170
rect 28130 14118 28142 14170
rect 28194 14118 28206 14170
rect 28258 14118 37950 14170
rect 38002 14118 38014 14170
rect 38066 14118 38078 14170
rect 38130 14118 38142 14170
rect 38194 14118 38206 14170
rect 38258 14118 47950 14170
rect 48002 14118 48014 14170
rect 48066 14118 48078 14170
rect 48130 14118 48142 14170
rect 48194 14118 48206 14170
rect 48258 14118 49864 14170
rect 1104 14096 49864 14118
rect 34882 14056 34888 14068
rect 33980 14028 34888 14056
rect 26326 13948 26332 14000
rect 26384 13988 26390 14000
rect 33980 13988 34008 14028
rect 34882 14016 34888 14028
rect 34940 14056 34946 14068
rect 35894 14056 35900 14068
rect 34940 14028 35900 14056
rect 34940 14016 34946 14028
rect 35894 14016 35900 14028
rect 35952 14016 35958 14068
rect 36725 14059 36783 14065
rect 36725 14025 36737 14059
rect 36771 14056 36783 14059
rect 43714 14056 43720 14068
rect 36771 14028 43720 14056
rect 36771 14025 36783 14028
rect 36725 14019 36783 14025
rect 43714 14016 43720 14028
rect 43772 14016 43778 14068
rect 26384 13960 30696 13988
rect 26384 13948 26390 13960
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13920 1823 13923
rect 5626 13920 5632 13932
rect 1811 13892 5632 13920
rect 1811 13889 1823 13892
rect 1765 13883 1823 13889
rect 5626 13880 5632 13892
rect 5684 13880 5690 13932
rect 28997 13923 29055 13929
rect 28997 13889 29009 13923
rect 29043 13920 29055 13923
rect 29270 13920 29276 13932
rect 29043 13892 29276 13920
rect 29043 13889 29055 13892
rect 28997 13883 29055 13889
rect 29270 13880 29276 13892
rect 29328 13880 29334 13932
rect 30668 13929 30696 13960
rect 33888 13960 34008 13988
rect 33888 13929 33916 13960
rect 34698 13948 34704 14000
rect 34756 13948 34762 14000
rect 36538 13948 36544 14000
rect 36596 13988 36602 14000
rect 37553 13991 37611 13997
rect 37553 13988 37565 13991
rect 36596 13960 37565 13988
rect 36596 13948 36602 13960
rect 37553 13957 37565 13960
rect 37599 13957 37611 13991
rect 37553 13951 37611 13957
rect 37734 13948 37740 14000
rect 37792 13948 37798 14000
rect 38289 13991 38347 13997
rect 38289 13957 38301 13991
rect 38335 13988 38347 13991
rect 38378 13988 38384 14000
rect 38335 13960 38384 13988
rect 38335 13957 38347 13960
rect 38289 13951 38347 13957
rect 38378 13948 38384 13960
rect 38436 13948 38442 14000
rect 38930 13948 38936 14000
rect 38988 13988 38994 14000
rect 42702 13988 42708 14000
rect 38988 13960 42708 13988
rect 38988 13948 38994 13960
rect 42702 13948 42708 13960
rect 42760 13948 42766 14000
rect 30653 13923 30711 13929
rect 30653 13889 30665 13923
rect 30699 13889 30711 13923
rect 30653 13883 30711 13889
rect 33873 13923 33931 13929
rect 33873 13889 33885 13923
rect 33919 13889 33931 13923
rect 33873 13883 33931 13889
rect 35452 13892 35894 13920
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 29181 13855 29239 13861
rect 29181 13821 29193 13855
rect 29227 13852 29239 13855
rect 29730 13852 29736 13864
rect 29227 13824 29736 13852
rect 29227 13821 29239 13824
rect 29181 13815 29239 13821
rect 29730 13812 29736 13824
rect 29788 13812 29794 13864
rect 35452 13852 35480 13892
rect 30484 13824 35480 13852
rect 30484 13793 30512 13824
rect 35526 13812 35532 13864
rect 35584 13852 35590 13864
rect 35621 13855 35679 13861
rect 35621 13852 35633 13855
rect 35584 13824 35633 13852
rect 35584 13812 35590 13824
rect 35621 13821 35633 13824
rect 35667 13821 35679 13855
rect 35866 13852 35894 13892
rect 36906 13880 36912 13932
rect 36964 13880 36970 13932
rect 38212 13892 38608 13920
rect 38212 13852 38240 13892
rect 35866 13824 38240 13852
rect 35621 13815 35679 13821
rect 38470 13812 38476 13864
rect 38528 13812 38534 13864
rect 38580 13852 38608 13892
rect 39114 13880 39120 13932
rect 39172 13880 39178 13932
rect 40126 13880 40132 13932
rect 40184 13920 40190 13932
rect 41785 13923 41843 13929
rect 41785 13920 41797 13923
rect 40184 13892 41797 13920
rect 40184 13880 40190 13892
rect 41785 13889 41797 13892
rect 41831 13889 41843 13923
rect 41785 13883 41843 13889
rect 46658 13880 46664 13932
rect 46716 13920 46722 13932
rect 47949 13923 48007 13929
rect 47949 13920 47961 13923
rect 46716 13892 47961 13920
rect 46716 13880 46722 13892
rect 47949 13889 47961 13892
rect 47995 13889 48007 13923
rect 47949 13883 48007 13889
rect 40586 13852 40592 13864
rect 38580 13824 40592 13852
rect 40586 13812 40592 13824
rect 40644 13812 40650 13864
rect 44358 13852 44364 13864
rect 41616 13824 44364 13852
rect 30469 13787 30527 13793
rect 30469 13753 30481 13787
rect 30515 13753 30527 13787
rect 30469 13747 30527 13753
rect 38930 13744 38936 13796
rect 38988 13744 38994 13796
rect 41616 13793 41644 13824
rect 44358 13812 44364 13824
rect 44416 13812 44422 13864
rect 49142 13812 49148 13864
rect 49200 13812 49206 13864
rect 41601 13787 41659 13793
rect 41601 13753 41613 13787
rect 41647 13753 41659 13787
rect 41601 13747 41659 13753
rect 34136 13719 34194 13725
rect 34136 13685 34148 13719
rect 34182 13716 34194 13719
rect 35434 13716 35440 13728
rect 34182 13688 35440 13716
rect 34182 13685 34194 13688
rect 34136 13679 34194 13685
rect 35434 13676 35440 13688
rect 35492 13676 35498 13728
rect 1104 13626 49864 13648
rect 1104 13574 2950 13626
rect 3002 13574 3014 13626
rect 3066 13574 3078 13626
rect 3130 13574 3142 13626
rect 3194 13574 3206 13626
rect 3258 13574 12950 13626
rect 13002 13574 13014 13626
rect 13066 13574 13078 13626
rect 13130 13574 13142 13626
rect 13194 13574 13206 13626
rect 13258 13574 22950 13626
rect 23002 13574 23014 13626
rect 23066 13574 23078 13626
rect 23130 13574 23142 13626
rect 23194 13574 23206 13626
rect 23258 13574 32950 13626
rect 33002 13574 33014 13626
rect 33066 13574 33078 13626
rect 33130 13574 33142 13626
rect 33194 13574 33206 13626
rect 33258 13574 42950 13626
rect 43002 13574 43014 13626
rect 43066 13574 43078 13626
rect 43130 13574 43142 13626
rect 43194 13574 43206 13626
rect 43258 13574 49864 13626
rect 1104 13552 49864 13574
rect 27798 13472 27804 13524
rect 27856 13512 27862 13524
rect 28261 13515 28319 13521
rect 28261 13512 28273 13515
rect 27856 13484 28273 13512
rect 27856 13472 27862 13484
rect 28261 13481 28273 13484
rect 28307 13481 28319 13515
rect 28261 13475 28319 13481
rect 33962 13472 33968 13524
rect 34020 13512 34026 13524
rect 36633 13515 36691 13521
rect 36633 13512 36645 13515
rect 34020 13484 36645 13512
rect 34020 13472 34026 13484
rect 36633 13481 36645 13484
rect 36679 13481 36691 13515
rect 36633 13475 36691 13481
rect 27338 13336 27344 13388
rect 27396 13376 27402 13388
rect 27798 13376 27804 13388
rect 27396 13348 27804 13376
rect 27396 13336 27402 13348
rect 27798 13336 27804 13348
rect 27856 13336 27862 13388
rect 28442 13336 28448 13388
rect 28500 13376 28506 13388
rect 28813 13379 28871 13385
rect 28813 13376 28825 13379
rect 28500 13348 28825 13376
rect 28500 13336 28506 13348
rect 28813 13345 28825 13348
rect 28859 13345 28871 13379
rect 28813 13339 28871 13345
rect 34882 13336 34888 13388
rect 34940 13336 34946 13388
rect 35161 13379 35219 13385
rect 35161 13345 35173 13379
rect 35207 13376 35219 13379
rect 37642 13376 37648 13388
rect 35207 13348 37648 13376
rect 35207 13345 35219 13348
rect 35161 13339 35219 13345
rect 37642 13336 37648 13348
rect 37700 13336 37706 13388
rect 25406 13268 25412 13320
rect 25464 13308 25470 13320
rect 25685 13311 25743 13317
rect 25685 13308 25697 13311
rect 25464 13280 25697 13308
rect 25464 13268 25470 13280
rect 25685 13277 25697 13280
rect 25731 13277 25743 13311
rect 25685 13271 25743 13277
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 28902 13308 28908 13320
rect 28767 13280 28908 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 28902 13268 28908 13280
rect 28960 13308 28966 13320
rect 28960 13280 31754 13308
rect 28960 13268 28966 13280
rect 28629 13243 28687 13249
rect 28629 13209 28641 13243
rect 28675 13240 28687 13243
rect 31726 13240 31754 13280
rect 33502 13268 33508 13320
rect 33560 13308 33566 13320
rect 34149 13311 34207 13317
rect 34149 13308 34161 13311
rect 33560 13280 34161 13308
rect 33560 13268 33566 13280
rect 34149 13277 34161 13280
rect 34195 13277 34207 13311
rect 34149 13271 34207 13277
rect 37090 13268 37096 13320
rect 37148 13308 37154 13320
rect 37185 13311 37243 13317
rect 37185 13308 37197 13311
rect 37148 13280 37197 13308
rect 37148 13268 37154 13280
rect 37185 13277 37197 13280
rect 37231 13277 37243 13311
rect 37185 13271 37243 13277
rect 37274 13268 37280 13320
rect 37332 13308 37338 13320
rect 38013 13311 38071 13317
rect 38013 13308 38025 13311
rect 37332 13280 38025 13308
rect 37332 13268 37338 13280
rect 38013 13277 38025 13280
rect 38059 13277 38071 13311
rect 38013 13271 38071 13277
rect 38286 13268 38292 13320
rect 38344 13308 38350 13320
rect 38657 13311 38715 13317
rect 38657 13308 38669 13311
rect 38344 13280 38669 13308
rect 38344 13268 38350 13280
rect 38657 13277 38669 13280
rect 38703 13277 38715 13311
rect 38657 13271 38715 13277
rect 40586 13268 40592 13320
rect 40644 13268 40650 13320
rect 44818 13268 44824 13320
rect 44876 13308 44882 13320
rect 47949 13311 48007 13317
rect 47949 13308 47961 13311
rect 44876 13280 47961 13308
rect 44876 13268 44882 13280
rect 47949 13277 47961 13280
rect 47995 13277 48007 13311
rect 47949 13271 48007 13277
rect 33686 13240 33692 13252
rect 28675 13212 30236 13240
rect 31726 13212 33692 13240
rect 28675 13209 28687 13212
rect 28629 13203 28687 13209
rect 25774 13132 25780 13184
rect 25832 13132 25838 13184
rect 30208 13172 30236 13212
rect 33686 13200 33692 13212
rect 33744 13200 33750 13252
rect 36538 13240 36544 13252
rect 36386 13212 36544 13240
rect 31754 13172 31760 13184
rect 30208 13144 31760 13172
rect 31754 13132 31760 13144
rect 31812 13172 31818 13184
rect 32582 13172 32588 13184
rect 31812 13144 32588 13172
rect 31812 13132 31818 13144
rect 32582 13132 32588 13144
rect 32640 13132 32646 13184
rect 34238 13132 34244 13184
rect 34296 13132 34302 13184
rect 34698 13132 34704 13184
rect 34756 13172 34762 13184
rect 36464 13172 36492 13212
rect 36538 13200 36544 13212
rect 36596 13200 36602 13252
rect 37366 13200 37372 13252
rect 37424 13200 37430 13252
rect 49142 13200 49148 13252
rect 49200 13200 49206 13252
rect 34756 13144 36492 13172
rect 38473 13175 38531 13181
rect 34756 13132 34762 13144
rect 38473 13141 38485 13175
rect 38519 13172 38531 13175
rect 39850 13172 39856 13184
rect 38519 13144 39856 13172
rect 38519 13141 38531 13144
rect 38473 13135 38531 13141
rect 39850 13132 39856 13144
rect 39908 13132 39914 13184
rect 40681 13175 40739 13181
rect 40681 13141 40693 13175
rect 40727 13172 40739 13175
rect 46750 13172 46756 13184
rect 40727 13144 46756 13172
rect 40727 13141 40739 13144
rect 40681 13135 40739 13141
rect 46750 13132 46756 13144
rect 46808 13132 46814 13184
rect 1104 13082 49864 13104
rect 1104 13030 7950 13082
rect 8002 13030 8014 13082
rect 8066 13030 8078 13082
rect 8130 13030 8142 13082
rect 8194 13030 8206 13082
rect 8258 13030 17950 13082
rect 18002 13030 18014 13082
rect 18066 13030 18078 13082
rect 18130 13030 18142 13082
rect 18194 13030 18206 13082
rect 18258 13030 27950 13082
rect 28002 13030 28014 13082
rect 28066 13030 28078 13082
rect 28130 13030 28142 13082
rect 28194 13030 28206 13082
rect 28258 13030 37950 13082
rect 38002 13030 38014 13082
rect 38066 13030 38078 13082
rect 38130 13030 38142 13082
rect 38194 13030 38206 13082
rect 38258 13030 47950 13082
rect 48002 13030 48014 13082
rect 48066 13030 48078 13082
rect 48130 13030 48142 13082
rect 48194 13030 48206 13082
rect 48258 13030 49864 13082
rect 1104 13008 49864 13030
rect 27522 12928 27528 12980
rect 27580 12968 27586 12980
rect 28813 12971 28871 12977
rect 28813 12968 28825 12971
rect 27580 12940 28825 12968
rect 27580 12928 27586 12940
rect 28813 12937 28825 12940
rect 28859 12937 28871 12971
rect 28813 12931 28871 12937
rect 29270 12928 29276 12980
rect 29328 12968 29334 12980
rect 30282 12968 30288 12980
rect 29328 12940 30288 12968
rect 29328 12928 29334 12940
rect 30282 12928 30288 12940
rect 30340 12928 30346 12980
rect 30469 12971 30527 12977
rect 30469 12937 30481 12971
rect 30515 12968 30527 12971
rect 30558 12968 30564 12980
rect 30515 12940 30564 12968
rect 30515 12937 30527 12940
rect 30469 12931 30527 12937
rect 30558 12928 30564 12940
rect 30616 12928 30622 12980
rect 34790 12968 34796 12980
rect 33704 12940 34796 12968
rect 26510 12860 26516 12912
rect 26568 12900 26574 12912
rect 27249 12903 27307 12909
rect 27249 12900 27261 12903
rect 26568 12872 27261 12900
rect 26568 12860 26574 12872
rect 27249 12869 27261 12872
rect 27295 12869 27307 12903
rect 27249 12863 27307 12869
rect 27985 12903 28043 12909
rect 27985 12869 27997 12903
rect 28031 12900 28043 12903
rect 28350 12900 28356 12912
rect 28031 12872 28356 12900
rect 28031 12869 28043 12872
rect 27985 12863 28043 12869
rect 28350 12860 28356 12872
rect 28408 12860 28414 12912
rect 29181 12903 29239 12909
rect 29181 12869 29193 12903
rect 29227 12900 29239 12903
rect 32398 12900 32404 12912
rect 29227 12872 32404 12900
rect 29227 12869 29239 12872
rect 29181 12863 29239 12869
rect 32398 12860 32404 12872
rect 32456 12860 32462 12912
rect 28442 12792 28448 12844
rect 28500 12832 28506 12844
rect 33704 12841 33732 12940
rect 34790 12928 34796 12940
rect 34848 12928 34854 12980
rect 35434 12928 35440 12980
rect 35492 12968 35498 12980
rect 36265 12971 36323 12977
rect 35492 12940 35894 12968
rect 35492 12928 35498 12940
rect 33962 12860 33968 12912
rect 34020 12860 34026 12912
rect 34698 12860 34704 12912
rect 34756 12860 34762 12912
rect 35866 12900 35894 12940
rect 36265 12937 36277 12971
rect 36311 12968 36323 12971
rect 37274 12968 37280 12980
rect 36311 12940 37280 12968
rect 36311 12937 36323 12940
rect 36265 12931 36323 12937
rect 37274 12928 37280 12940
rect 37332 12928 37338 12980
rect 35866 12872 36492 12900
rect 30377 12835 30435 12841
rect 28500 12804 29684 12832
rect 28500 12792 28506 12804
rect 29457 12767 29515 12773
rect 29457 12733 29469 12767
rect 29503 12764 29515 12767
rect 29546 12764 29552 12776
rect 29503 12736 29552 12764
rect 29503 12733 29515 12736
rect 29457 12727 29515 12733
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 29656 12764 29684 12804
rect 30377 12801 30389 12835
rect 30423 12832 30435 12835
rect 33689 12835 33747 12841
rect 30423 12804 31754 12832
rect 30423 12801 30435 12804
rect 30377 12795 30435 12801
rect 30561 12767 30619 12773
rect 30561 12764 30573 12767
rect 29656 12736 30573 12764
rect 30561 12733 30573 12736
rect 30607 12733 30619 12767
rect 30561 12727 30619 12733
rect 27154 12656 27160 12708
rect 27212 12696 27218 12708
rect 28169 12699 28227 12705
rect 28169 12696 28181 12699
rect 27212 12668 28181 12696
rect 27212 12656 27218 12668
rect 28169 12665 28181 12668
rect 28215 12665 28227 12699
rect 28169 12659 28227 12665
rect 30006 12656 30012 12708
rect 30064 12656 30070 12708
rect 25222 12588 25228 12640
rect 25280 12628 25286 12640
rect 27341 12631 27399 12637
rect 27341 12628 27353 12631
rect 25280 12600 27353 12628
rect 25280 12588 25286 12600
rect 27341 12597 27353 12600
rect 27387 12597 27399 12631
rect 31726 12628 31754 12804
rect 33689 12801 33701 12835
rect 33735 12801 33747 12835
rect 33689 12795 33747 12801
rect 34330 12724 34336 12776
rect 34388 12764 34394 12776
rect 36464 12773 36492 12872
rect 43714 12860 43720 12912
rect 43772 12860 43778 12912
rect 46750 12792 46756 12844
rect 46808 12832 46814 12844
rect 47949 12835 48007 12841
rect 47949 12832 47961 12835
rect 46808 12804 47961 12832
rect 46808 12792 46814 12804
rect 47949 12801 47961 12804
rect 47995 12801 48007 12835
rect 47949 12795 48007 12801
rect 36357 12767 36415 12773
rect 36357 12764 36369 12767
rect 34388 12736 36369 12764
rect 34388 12724 34394 12736
rect 36357 12733 36369 12736
rect 36403 12733 36415 12767
rect 36357 12727 36415 12733
rect 36449 12767 36507 12773
rect 36449 12733 36461 12767
rect 36495 12733 36507 12767
rect 36449 12727 36507 12733
rect 49142 12724 49148 12776
rect 49200 12724 49206 12776
rect 36078 12696 36084 12708
rect 34992 12668 36084 12696
rect 34992 12628 35020 12668
rect 36078 12656 36084 12668
rect 36136 12696 36142 12708
rect 36814 12696 36820 12708
rect 36136 12668 36820 12696
rect 36136 12656 36142 12668
rect 36814 12656 36820 12668
rect 36872 12656 36878 12708
rect 43901 12699 43959 12705
rect 43901 12665 43913 12699
rect 43947 12696 43959 12699
rect 44726 12696 44732 12708
rect 43947 12668 44732 12696
rect 43947 12665 43959 12668
rect 43901 12659 43959 12665
rect 44726 12656 44732 12668
rect 44784 12656 44790 12708
rect 31726 12600 35020 12628
rect 35897 12631 35955 12637
rect 27341 12591 27399 12597
rect 35897 12597 35909 12631
rect 35943 12628 35955 12631
rect 39942 12628 39948 12640
rect 35943 12600 39948 12628
rect 35943 12597 35955 12600
rect 35897 12591 35955 12597
rect 39942 12588 39948 12600
rect 40000 12588 40006 12640
rect 1104 12538 49864 12560
rect 1104 12486 2950 12538
rect 3002 12486 3014 12538
rect 3066 12486 3078 12538
rect 3130 12486 3142 12538
rect 3194 12486 3206 12538
rect 3258 12486 12950 12538
rect 13002 12486 13014 12538
rect 13066 12486 13078 12538
rect 13130 12486 13142 12538
rect 13194 12486 13206 12538
rect 13258 12486 22950 12538
rect 23002 12486 23014 12538
rect 23066 12486 23078 12538
rect 23130 12486 23142 12538
rect 23194 12486 23206 12538
rect 23258 12486 32950 12538
rect 33002 12486 33014 12538
rect 33066 12486 33078 12538
rect 33130 12486 33142 12538
rect 33194 12486 33206 12538
rect 33258 12486 42950 12538
rect 43002 12486 43014 12538
rect 43066 12486 43078 12538
rect 43130 12486 43142 12538
rect 43194 12486 43206 12538
rect 43258 12486 49864 12538
rect 1104 12464 49864 12486
rect 3326 12316 3332 12368
rect 3384 12356 3390 12368
rect 9490 12356 9496 12368
rect 3384 12328 9496 12356
rect 3384 12316 3390 12328
rect 9490 12316 9496 12328
rect 9548 12316 9554 12368
rect 39850 12248 39856 12300
rect 39908 12288 39914 12300
rect 39908 12260 44496 12288
rect 39908 12248 39914 12260
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12220 28871 12223
rect 28902 12220 28908 12232
rect 28859 12192 28908 12220
rect 28859 12189 28871 12192
rect 28813 12183 28871 12189
rect 28902 12180 28908 12192
rect 28960 12180 28966 12232
rect 38930 12180 38936 12232
rect 38988 12180 38994 12232
rect 41230 12180 41236 12232
rect 41288 12180 41294 12232
rect 44468 12229 44496 12260
rect 44453 12223 44511 12229
rect 44453 12189 44465 12223
rect 44499 12189 44511 12223
rect 44453 12183 44511 12189
rect 44726 12180 44732 12232
rect 44784 12220 44790 12232
rect 47949 12223 48007 12229
rect 47949 12220 47961 12223
rect 44784 12192 47961 12220
rect 44784 12180 44790 12192
rect 47949 12189 47961 12192
rect 47995 12189 48007 12223
rect 47949 12183 48007 12189
rect 28997 12155 29055 12161
rect 28997 12121 29009 12155
rect 29043 12152 29055 12155
rect 29178 12152 29184 12164
rect 29043 12124 29184 12152
rect 29043 12121 29055 12124
rect 28997 12115 29055 12121
rect 29178 12112 29184 12124
rect 29236 12112 29242 12164
rect 39117 12155 39175 12161
rect 39117 12121 39129 12155
rect 39163 12152 39175 12155
rect 41874 12152 41880 12164
rect 39163 12124 41880 12152
rect 39163 12121 39175 12124
rect 39117 12115 39175 12121
rect 41874 12112 41880 12124
rect 41932 12112 41938 12164
rect 49142 12112 49148 12164
rect 49200 12112 49206 12164
rect 41049 12087 41107 12093
rect 41049 12053 41061 12087
rect 41095 12084 41107 12087
rect 43346 12084 43352 12096
rect 41095 12056 43352 12084
rect 41095 12053 41107 12056
rect 41049 12047 41107 12053
rect 43346 12044 43352 12056
rect 43404 12044 43410 12096
rect 44266 12044 44272 12096
rect 44324 12044 44330 12096
rect 1104 11994 49864 12016
rect 1104 11942 7950 11994
rect 8002 11942 8014 11994
rect 8066 11942 8078 11994
rect 8130 11942 8142 11994
rect 8194 11942 8206 11994
rect 8258 11942 17950 11994
rect 18002 11942 18014 11994
rect 18066 11942 18078 11994
rect 18130 11942 18142 11994
rect 18194 11942 18206 11994
rect 18258 11942 27950 11994
rect 28002 11942 28014 11994
rect 28066 11942 28078 11994
rect 28130 11942 28142 11994
rect 28194 11942 28206 11994
rect 28258 11942 37950 11994
rect 38002 11942 38014 11994
rect 38066 11942 38078 11994
rect 38130 11942 38142 11994
rect 38194 11942 38206 11994
rect 38258 11942 47950 11994
rect 48002 11942 48014 11994
rect 48066 11942 48078 11994
rect 48130 11942 48142 11994
rect 48194 11942 48206 11994
rect 48258 11942 49864 11994
rect 1104 11920 49864 11942
rect 44174 11772 44180 11824
rect 44232 11812 44238 11824
rect 46293 11815 46351 11821
rect 46293 11812 46305 11815
rect 44232 11784 46305 11812
rect 44232 11772 44238 11784
rect 46293 11781 46305 11784
rect 46339 11781 46351 11815
rect 46293 11775 46351 11781
rect 41322 11704 41328 11756
rect 41380 11744 41386 11756
rect 41601 11747 41659 11753
rect 41601 11744 41613 11747
rect 41380 11716 41613 11744
rect 41380 11704 41386 11716
rect 41601 11713 41613 11716
rect 41647 11713 41659 11747
rect 41601 11707 41659 11713
rect 42702 11704 42708 11756
rect 42760 11744 42766 11756
rect 44821 11747 44879 11753
rect 45557 11748 45615 11753
rect 44821 11744 44833 11747
rect 42760 11716 44833 11744
rect 42760 11704 42766 11716
rect 44821 11713 44833 11716
rect 44867 11713 44879 11747
rect 44821 11707 44879 11713
rect 45480 11747 45615 11748
rect 45480 11720 45569 11747
rect 42794 11636 42800 11688
rect 42852 11676 42858 11688
rect 45480 11676 45508 11720
rect 45557 11713 45569 11720
rect 45603 11713 45615 11747
rect 45557 11707 45615 11713
rect 42852 11648 45508 11676
rect 42852 11636 42858 11648
rect 45005 11611 45063 11617
rect 45005 11577 45017 11611
rect 45051 11608 45063 11611
rect 45646 11608 45652 11620
rect 45051 11580 45652 11608
rect 45051 11577 45063 11580
rect 45005 11571 45063 11577
rect 45646 11568 45652 11580
rect 45704 11568 45710 11620
rect 45741 11611 45799 11617
rect 45741 11577 45753 11611
rect 45787 11608 45799 11611
rect 46842 11608 46848 11620
rect 45787 11580 46848 11608
rect 45787 11577 45799 11580
rect 45741 11571 45799 11577
rect 46842 11568 46848 11580
rect 46900 11568 46906 11620
rect 41417 11543 41475 11549
rect 41417 11509 41429 11543
rect 41463 11540 41475 11543
rect 44174 11540 44180 11552
rect 41463 11512 44180 11540
rect 41463 11509 41475 11512
rect 41417 11503 41475 11509
rect 44174 11500 44180 11512
rect 44232 11500 44238 11552
rect 46382 11500 46388 11552
rect 46440 11500 46446 11552
rect 1104 11450 49864 11472
rect 1104 11398 2950 11450
rect 3002 11398 3014 11450
rect 3066 11398 3078 11450
rect 3130 11398 3142 11450
rect 3194 11398 3206 11450
rect 3258 11398 12950 11450
rect 13002 11398 13014 11450
rect 13066 11398 13078 11450
rect 13130 11398 13142 11450
rect 13194 11398 13206 11450
rect 13258 11398 22950 11450
rect 23002 11398 23014 11450
rect 23066 11398 23078 11450
rect 23130 11398 23142 11450
rect 23194 11398 23206 11450
rect 23258 11398 32950 11450
rect 33002 11398 33014 11450
rect 33066 11398 33078 11450
rect 33130 11398 33142 11450
rect 33194 11398 33206 11450
rect 33258 11398 42950 11450
rect 43002 11398 43014 11450
rect 43066 11398 43078 11450
rect 43130 11398 43142 11450
rect 43194 11398 43206 11450
rect 43258 11398 49864 11450
rect 1104 11376 49864 11398
rect 12989 11339 13047 11345
rect 12989 11305 13001 11339
rect 13035 11336 13047 11339
rect 17862 11336 17868 11348
rect 13035 11308 17868 11336
rect 13035 11305 13047 11308
rect 12989 11299 13047 11305
rect 17862 11296 17868 11308
rect 17920 11296 17926 11348
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 19702 11200 19708 11212
rect 13679 11172 19708 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13403 11104 14473 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 44266 11092 44272 11144
rect 44324 11132 44330 11144
rect 47949 11135 48007 11141
rect 47949 11132 47961 11135
rect 44324 11104 47961 11132
rect 44324 11092 44330 11104
rect 47949 11101 47961 11104
rect 47995 11101 48007 11135
rect 47949 11095 48007 11101
rect 49142 11092 49148 11144
rect 49200 11092 49206 11144
rect 7558 11024 7564 11076
rect 7616 11064 7622 11076
rect 12437 11067 12495 11073
rect 12437 11064 12449 11067
rect 7616 11036 12449 11064
rect 7616 11024 7622 11036
rect 12437 11033 12449 11036
rect 12483 11064 12495 11067
rect 13449 11067 13507 11073
rect 13449 11064 13461 11067
rect 12483 11036 13461 11064
rect 12483 11033 12495 11036
rect 12437 11027 12495 11033
rect 13449 11033 13461 11036
rect 13495 11033 13507 11067
rect 13449 11027 13507 11033
rect 44358 11024 44364 11076
rect 44416 11064 44422 11076
rect 46293 11067 46351 11073
rect 46293 11064 46305 11067
rect 44416 11036 46305 11064
rect 44416 11024 44422 11036
rect 46293 11033 46305 11036
rect 46339 11033 46351 11067
rect 46293 11027 46351 11033
rect 46474 11024 46480 11076
rect 46532 11024 46538 11076
rect 1104 10906 49864 10928
rect 1104 10854 7950 10906
rect 8002 10854 8014 10906
rect 8066 10854 8078 10906
rect 8130 10854 8142 10906
rect 8194 10854 8206 10906
rect 8258 10854 17950 10906
rect 18002 10854 18014 10906
rect 18066 10854 18078 10906
rect 18130 10854 18142 10906
rect 18194 10854 18206 10906
rect 18258 10854 27950 10906
rect 28002 10854 28014 10906
rect 28066 10854 28078 10906
rect 28130 10854 28142 10906
rect 28194 10854 28206 10906
rect 28258 10854 37950 10906
rect 38002 10854 38014 10906
rect 38066 10854 38078 10906
rect 38130 10854 38142 10906
rect 38194 10854 38206 10906
rect 38258 10854 47950 10906
rect 48002 10854 48014 10906
rect 48066 10854 48078 10906
rect 48130 10854 48142 10906
rect 48194 10854 48206 10906
rect 48258 10854 49864 10906
rect 1104 10832 49864 10854
rect 24210 10684 24216 10736
rect 24268 10724 24274 10736
rect 24489 10727 24547 10733
rect 24489 10724 24501 10727
rect 24268 10696 24501 10724
rect 24268 10684 24274 10696
rect 24489 10693 24501 10696
rect 24535 10693 24547 10727
rect 24489 10687 24547 10693
rect 39942 10616 39948 10668
rect 40000 10656 40006 10668
rect 40773 10659 40831 10665
rect 40773 10656 40785 10659
rect 40000 10628 40785 10656
rect 40000 10616 40006 10628
rect 40773 10625 40785 10628
rect 40819 10625 40831 10659
rect 40773 10619 40831 10625
rect 47578 10616 47584 10668
rect 47636 10656 47642 10668
rect 47949 10659 48007 10665
rect 47949 10656 47961 10659
rect 47636 10628 47961 10656
rect 47636 10616 47642 10628
rect 47949 10625 47961 10628
rect 47995 10625 48007 10659
rect 47949 10619 48007 10625
rect 49142 10548 49148 10600
rect 49200 10548 49206 10600
rect 24673 10523 24731 10529
rect 24673 10489 24685 10523
rect 24719 10520 24731 10523
rect 25130 10520 25136 10532
rect 24719 10492 25136 10520
rect 24719 10489 24731 10492
rect 24673 10483 24731 10489
rect 25130 10480 25136 10492
rect 25188 10480 25194 10532
rect 40589 10455 40647 10461
rect 40589 10421 40601 10455
rect 40635 10452 40647 10455
rect 42702 10452 42708 10464
rect 40635 10424 42708 10452
rect 40635 10421 40647 10424
rect 40589 10415 40647 10421
rect 42702 10412 42708 10424
rect 42760 10412 42766 10464
rect 1104 10362 49864 10384
rect 1104 10310 2950 10362
rect 3002 10310 3014 10362
rect 3066 10310 3078 10362
rect 3130 10310 3142 10362
rect 3194 10310 3206 10362
rect 3258 10310 12950 10362
rect 13002 10310 13014 10362
rect 13066 10310 13078 10362
rect 13130 10310 13142 10362
rect 13194 10310 13206 10362
rect 13258 10310 22950 10362
rect 23002 10310 23014 10362
rect 23066 10310 23078 10362
rect 23130 10310 23142 10362
rect 23194 10310 23206 10362
rect 23258 10310 32950 10362
rect 33002 10310 33014 10362
rect 33066 10310 33078 10362
rect 33130 10310 33142 10362
rect 33194 10310 33206 10362
rect 33258 10310 42950 10362
rect 43002 10310 43014 10362
rect 43066 10310 43078 10362
rect 43130 10310 43142 10362
rect 43194 10310 43206 10362
rect 43258 10310 49864 10362
rect 1104 10288 49864 10310
rect 28534 10004 28540 10056
rect 28592 10044 28598 10056
rect 28721 10047 28779 10053
rect 28721 10044 28733 10047
rect 28592 10016 28733 10044
rect 28592 10004 28598 10016
rect 28721 10013 28733 10016
rect 28767 10013 28779 10047
rect 28721 10007 28779 10013
rect 31846 10004 31852 10056
rect 31904 10004 31910 10056
rect 45646 10004 45652 10056
rect 45704 10044 45710 10056
rect 47949 10047 48007 10053
rect 47949 10044 47961 10047
rect 45704 10016 47961 10044
rect 45704 10004 45710 10016
rect 47949 10013 47961 10016
rect 47995 10013 48007 10047
rect 47949 10007 48007 10013
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 30098 9976 30104 9988
rect 28951 9948 30104 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 30098 9936 30104 9948
rect 30156 9936 30162 9988
rect 49142 9936 49148 9988
rect 49200 9936 49206 9988
rect 29914 9868 29920 9920
rect 29972 9908 29978 9920
rect 31941 9911 31999 9917
rect 31941 9908 31953 9911
rect 29972 9880 31953 9908
rect 29972 9868 29978 9880
rect 31941 9877 31953 9880
rect 31987 9877 31999 9911
rect 31941 9871 31999 9877
rect 1104 9818 49864 9840
rect 1104 9766 7950 9818
rect 8002 9766 8014 9818
rect 8066 9766 8078 9818
rect 8130 9766 8142 9818
rect 8194 9766 8206 9818
rect 8258 9766 17950 9818
rect 18002 9766 18014 9818
rect 18066 9766 18078 9818
rect 18130 9766 18142 9818
rect 18194 9766 18206 9818
rect 18258 9766 27950 9818
rect 28002 9766 28014 9818
rect 28066 9766 28078 9818
rect 28130 9766 28142 9818
rect 28194 9766 28206 9818
rect 28258 9766 37950 9818
rect 38002 9766 38014 9818
rect 38066 9766 38078 9818
rect 38130 9766 38142 9818
rect 38194 9766 38206 9818
rect 38258 9766 47950 9818
rect 48002 9766 48014 9818
rect 48066 9766 48078 9818
rect 48130 9766 48142 9818
rect 48194 9766 48206 9818
rect 48258 9766 49864 9818
rect 1104 9744 49864 9766
rect 31938 9596 31944 9648
rect 31996 9636 32002 9648
rect 32401 9639 32459 9645
rect 32401 9636 32413 9639
rect 31996 9608 32413 9636
rect 31996 9596 32002 9608
rect 32401 9605 32413 9608
rect 32447 9605 32459 9639
rect 32401 9599 32459 9605
rect 34974 9596 34980 9648
rect 35032 9636 35038 9648
rect 35897 9639 35955 9645
rect 35897 9636 35909 9639
rect 35032 9608 35909 9636
rect 35032 9596 35038 9608
rect 35897 9605 35909 9608
rect 35943 9605 35955 9639
rect 35897 9599 35955 9605
rect 44174 9528 44180 9580
rect 44232 9568 44238 9580
rect 46293 9571 46351 9577
rect 46293 9568 46305 9571
rect 44232 9540 46305 9568
rect 44232 9528 44238 9540
rect 46293 9537 46305 9540
rect 46339 9537 46351 9571
rect 46293 9531 46351 9537
rect 46842 9528 46848 9580
rect 46900 9568 46906 9580
rect 47949 9571 48007 9577
rect 47949 9568 47961 9571
rect 46900 9540 47961 9568
rect 46900 9528 46906 9540
rect 47949 9537 47961 9540
rect 47995 9537 48007 9571
rect 47949 9531 48007 9537
rect 47762 9460 47768 9512
rect 47820 9500 47826 9512
rect 48682 9500 48688 9512
rect 47820 9472 48688 9500
rect 47820 9460 47826 9472
rect 48682 9460 48688 9472
rect 48740 9460 48746 9512
rect 49142 9460 49148 9512
rect 49200 9460 49206 9512
rect 32585 9435 32643 9441
rect 32585 9401 32597 9435
rect 32631 9432 32643 9435
rect 33962 9432 33968 9444
rect 32631 9404 33968 9432
rect 32631 9401 32643 9404
rect 32585 9395 32643 9401
rect 33962 9392 33968 9404
rect 34020 9392 34026 9444
rect 36081 9435 36139 9441
rect 36081 9401 36093 9435
rect 36127 9432 36139 9435
rect 37274 9432 37280 9444
rect 36127 9404 37280 9432
rect 36127 9401 36139 9404
rect 36081 9395 36139 9401
rect 37274 9392 37280 9404
rect 37332 9392 37338 9444
rect 46109 9367 46167 9373
rect 46109 9333 46121 9367
rect 46155 9364 46167 9367
rect 47762 9364 47768 9376
rect 46155 9336 47768 9364
rect 46155 9333 46167 9336
rect 46109 9327 46167 9333
rect 47762 9324 47768 9336
rect 47820 9324 47826 9376
rect 1104 9274 49864 9296
rect 1104 9222 2950 9274
rect 3002 9222 3014 9274
rect 3066 9222 3078 9274
rect 3130 9222 3142 9274
rect 3194 9222 3206 9274
rect 3258 9222 12950 9274
rect 13002 9222 13014 9274
rect 13066 9222 13078 9274
rect 13130 9222 13142 9274
rect 13194 9222 13206 9274
rect 13258 9222 22950 9274
rect 23002 9222 23014 9274
rect 23066 9222 23078 9274
rect 23130 9222 23142 9274
rect 23194 9222 23206 9274
rect 23258 9222 32950 9274
rect 33002 9222 33014 9274
rect 33066 9222 33078 9274
rect 33130 9222 33142 9274
rect 33194 9222 33206 9274
rect 33258 9222 42950 9274
rect 43002 9222 43014 9274
rect 43066 9222 43078 9274
rect 43130 9222 43142 9274
rect 43194 9222 43206 9274
rect 43258 9222 49864 9274
rect 1104 9200 49864 9222
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 9398 9092 9404 9104
rect 3384 9064 9404 9092
rect 3384 9052 3390 9064
rect 9398 9052 9404 9064
rect 9456 9052 9462 9104
rect 43346 8916 43352 8968
rect 43404 8956 43410 8968
rect 46017 8959 46075 8965
rect 46017 8956 46029 8959
rect 43404 8928 46029 8956
rect 43404 8916 43410 8928
rect 46017 8925 46029 8928
rect 46063 8925 46075 8959
rect 46017 8919 46075 8925
rect 47670 8916 47676 8968
rect 47728 8956 47734 8968
rect 48869 8959 48927 8965
rect 48869 8956 48881 8959
rect 47728 8928 48881 8956
rect 47728 8916 47734 8928
rect 48869 8925 48881 8928
rect 48915 8925 48927 8959
rect 48869 8919 48927 8925
rect 46198 8848 46204 8900
rect 46256 8848 46262 8900
rect 47118 8848 47124 8900
rect 47176 8888 47182 8900
rect 47949 8891 48007 8897
rect 47949 8888 47961 8891
rect 47176 8860 47961 8888
rect 47176 8848 47182 8860
rect 47949 8857 47961 8860
rect 47995 8888 48007 8891
rect 48406 8888 48412 8900
rect 47995 8860 48412 8888
rect 47995 8857 48007 8860
rect 47949 8851 48007 8857
rect 48406 8848 48412 8860
rect 48464 8848 48470 8900
rect 48682 8848 48688 8900
rect 48740 8848 48746 8900
rect 47854 8780 47860 8832
rect 47912 8820 47918 8832
rect 48041 8823 48099 8829
rect 48041 8820 48053 8823
rect 47912 8792 48053 8820
rect 47912 8780 47918 8792
rect 48041 8789 48053 8792
rect 48087 8789 48099 8823
rect 48041 8783 48099 8789
rect 1104 8730 49864 8752
rect 1104 8678 7950 8730
rect 8002 8678 8014 8730
rect 8066 8678 8078 8730
rect 8130 8678 8142 8730
rect 8194 8678 8206 8730
rect 8258 8678 17950 8730
rect 18002 8678 18014 8730
rect 18066 8678 18078 8730
rect 18130 8678 18142 8730
rect 18194 8678 18206 8730
rect 18258 8678 27950 8730
rect 28002 8678 28014 8730
rect 28066 8678 28078 8730
rect 28130 8678 28142 8730
rect 28194 8678 28206 8730
rect 28258 8678 37950 8730
rect 38002 8678 38014 8730
rect 38066 8678 38078 8730
rect 38130 8678 38142 8730
rect 38194 8678 38206 8730
rect 38258 8678 47950 8730
rect 48002 8678 48014 8730
rect 48066 8678 48078 8730
rect 48130 8678 48142 8730
rect 48194 8678 48206 8730
rect 48258 8678 49864 8730
rect 1104 8656 49864 8678
rect 9140 8588 13676 8616
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5592 8520 6914 8548
rect 5592 8508 5598 8520
rect 6886 8412 6914 8520
rect 9140 8489 9168 8588
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 13648 8480 13676 8588
rect 16482 8508 16488 8560
rect 16540 8548 16546 8560
rect 19242 8548 19248 8560
rect 16540 8520 19248 8548
rect 16540 8508 16546 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 32306 8508 32312 8560
rect 32364 8548 32370 8560
rect 36541 8551 36599 8557
rect 36541 8548 36553 8551
rect 32364 8520 36553 8548
rect 32364 8508 32370 8520
rect 36541 8517 36553 8520
rect 36587 8517 36599 8551
rect 36541 8511 36599 8517
rect 37826 8508 37832 8560
rect 37884 8508 37890 8560
rect 42702 8508 42708 8560
rect 42760 8548 42766 8560
rect 45741 8551 45799 8557
rect 45741 8548 45753 8551
rect 42760 8520 45753 8548
rect 42760 8508 42766 8520
rect 45741 8517 45753 8520
rect 45787 8517 45799 8551
rect 45741 8511 45799 8517
rect 18598 8480 18604 8492
rect 9125 8443 9183 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 6886 8384 9413 8412
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 10520 8344 10548 8466
rect 13648 8452 18604 8480
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 46474 8440 46480 8492
rect 46532 8480 46538 8492
rect 47949 8483 48007 8489
rect 47949 8480 47961 8483
rect 46532 8452 47961 8480
rect 46532 8440 46538 8452
rect 47949 8449 47961 8452
rect 47995 8449 48007 8483
rect 47949 8443 48007 8449
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8412 11207 8415
rect 23382 8412 23388 8424
rect 11195 8384 23388 8412
rect 11195 8381 11207 8384
rect 11149 8375 11207 8381
rect 23382 8372 23388 8384
rect 23440 8372 23446 8424
rect 36725 8415 36783 8421
rect 36725 8381 36737 8415
rect 36771 8412 36783 8415
rect 42610 8412 42616 8424
rect 36771 8384 42616 8412
rect 36771 8381 36783 8384
rect 36725 8375 36783 8381
rect 42610 8372 42616 8384
rect 42668 8372 42674 8424
rect 49142 8372 49148 8424
rect 49200 8372 49206 8424
rect 16482 8344 16488 8356
rect 10520 8316 16488 8344
rect 16482 8304 16488 8316
rect 16540 8304 16546 8356
rect 37642 8304 37648 8356
rect 37700 8344 37706 8356
rect 38013 8347 38071 8353
rect 38013 8344 38025 8347
rect 37700 8316 38025 8344
rect 37700 8304 37706 8316
rect 38013 8313 38025 8316
rect 38059 8313 38071 8347
rect 38013 8307 38071 8313
rect 45922 8304 45928 8356
rect 45980 8304 45986 8356
rect 1104 8186 49864 8208
rect 1104 8134 2950 8186
rect 3002 8134 3014 8186
rect 3066 8134 3078 8186
rect 3130 8134 3142 8186
rect 3194 8134 3206 8186
rect 3258 8134 12950 8186
rect 13002 8134 13014 8186
rect 13066 8134 13078 8186
rect 13130 8134 13142 8186
rect 13194 8134 13206 8186
rect 13258 8134 22950 8186
rect 23002 8134 23014 8186
rect 23066 8134 23078 8186
rect 23130 8134 23142 8186
rect 23194 8134 23206 8186
rect 23258 8134 32950 8186
rect 33002 8134 33014 8186
rect 33066 8134 33078 8186
rect 33130 8134 33142 8186
rect 33194 8134 33206 8186
rect 33258 8134 42950 8186
rect 43002 8134 43014 8186
rect 43066 8134 43078 8186
rect 43130 8134 43142 8186
rect 43194 8134 43206 8186
rect 43258 8134 49864 8186
rect 1104 8112 49864 8134
rect 46382 7828 46388 7880
rect 46440 7868 46446 7880
rect 47949 7871 48007 7877
rect 47949 7868 47961 7871
rect 46440 7840 47961 7868
rect 46440 7828 46446 7840
rect 47949 7837 47961 7840
rect 47995 7837 48007 7871
rect 47949 7831 48007 7837
rect 49142 7760 49148 7812
rect 49200 7760 49206 7812
rect 1104 7642 49864 7664
rect 1104 7590 7950 7642
rect 8002 7590 8014 7642
rect 8066 7590 8078 7642
rect 8130 7590 8142 7642
rect 8194 7590 8206 7642
rect 8258 7590 17950 7642
rect 18002 7590 18014 7642
rect 18066 7590 18078 7642
rect 18130 7590 18142 7642
rect 18194 7590 18206 7642
rect 18258 7590 27950 7642
rect 28002 7590 28014 7642
rect 28066 7590 28078 7642
rect 28130 7590 28142 7642
rect 28194 7590 28206 7642
rect 28258 7590 37950 7642
rect 38002 7590 38014 7642
rect 38066 7590 38078 7642
rect 38130 7590 38142 7642
rect 38194 7590 38206 7642
rect 38258 7590 47950 7642
rect 48002 7590 48014 7642
rect 48066 7590 48078 7642
rect 48130 7590 48142 7642
rect 48194 7590 48206 7642
rect 48258 7590 49864 7642
rect 1104 7568 49864 7590
rect 31754 7420 31760 7472
rect 31812 7460 31818 7472
rect 35713 7463 35771 7469
rect 35713 7460 35725 7463
rect 31812 7432 35725 7460
rect 31812 7420 31818 7432
rect 35713 7429 35725 7432
rect 35759 7429 35771 7463
rect 35713 7423 35771 7429
rect 29638 7352 29644 7404
rect 29696 7392 29702 7404
rect 37553 7395 37611 7401
rect 37553 7392 37565 7395
rect 29696 7364 37565 7392
rect 29696 7352 29702 7364
rect 37553 7361 37565 7364
rect 37599 7361 37611 7395
rect 37553 7355 37611 7361
rect 47762 7352 47768 7404
rect 47820 7392 47826 7404
rect 47949 7395 48007 7401
rect 47949 7392 47961 7395
rect 47820 7364 47961 7392
rect 47820 7352 47826 7364
rect 47949 7361 47961 7364
rect 47995 7361 48007 7395
rect 47949 7355 48007 7361
rect 35897 7327 35955 7333
rect 35897 7293 35909 7327
rect 35943 7324 35955 7327
rect 41414 7324 41420 7336
rect 35943 7296 41420 7324
rect 35943 7293 35955 7296
rect 35897 7287 35955 7293
rect 41414 7284 41420 7296
rect 41472 7284 41478 7336
rect 49142 7284 49148 7336
rect 49200 7284 49206 7336
rect 37737 7259 37795 7265
rect 37737 7225 37749 7259
rect 37783 7256 37795 7259
rect 45186 7256 45192 7268
rect 37783 7228 45192 7256
rect 37783 7225 37795 7228
rect 37737 7219 37795 7225
rect 45186 7216 45192 7228
rect 45244 7216 45250 7268
rect 47578 7216 47584 7268
rect 47636 7256 47642 7268
rect 47762 7256 47768 7268
rect 47636 7228 47768 7256
rect 47636 7216 47642 7228
rect 47762 7216 47768 7228
rect 47820 7216 47826 7268
rect 1104 7098 49864 7120
rect 1104 7046 2950 7098
rect 3002 7046 3014 7098
rect 3066 7046 3078 7098
rect 3130 7046 3142 7098
rect 3194 7046 3206 7098
rect 3258 7046 12950 7098
rect 13002 7046 13014 7098
rect 13066 7046 13078 7098
rect 13130 7046 13142 7098
rect 13194 7046 13206 7098
rect 13258 7046 22950 7098
rect 23002 7046 23014 7098
rect 23066 7046 23078 7098
rect 23130 7046 23142 7098
rect 23194 7046 23206 7098
rect 23258 7046 32950 7098
rect 33002 7046 33014 7098
rect 33066 7046 33078 7098
rect 33130 7046 33142 7098
rect 33194 7046 33206 7098
rect 33258 7046 42950 7098
rect 43002 7046 43014 7098
rect 43066 7046 43078 7098
rect 43130 7046 43142 7098
rect 43194 7046 43206 7098
rect 43258 7046 49864 7098
rect 1104 7024 49864 7046
rect 36814 6740 36820 6792
rect 36872 6780 36878 6792
rect 37737 6783 37795 6789
rect 36872 6752 37688 6780
rect 36872 6740 36878 6752
rect 32398 6672 32404 6724
rect 32456 6712 32462 6724
rect 37553 6715 37611 6721
rect 37553 6712 37565 6715
rect 32456 6684 37565 6712
rect 32456 6672 32462 6684
rect 37553 6681 37565 6684
rect 37599 6681 37611 6715
rect 37660 6712 37688 6752
rect 37737 6749 37749 6783
rect 37783 6780 37795 6783
rect 40126 6780 40132 6792
rect 37783 6752 40132 6780
rect 37783 6749 37795 6752
rect 37737 6743 37795 6749
rect 40126 6740 40132 6752
rect 40184 6740 40190 6792
rect 45922 6740 45928 6792
rect 45980 6780 45986 6792
rect 47949 6783 48007 6789
rect 47949 6780 47961 6783
rect 45980 6752 47961 6780
rect 45980 6740 45986 6752
rect 47949 6749 47961 6752
rect 47995 6749 48007 6783
rect 47949 6743 48007 6749
rect 38289 6715 38347 6721
rect 38289 6712 38301 6715
rect 37660 6684 38301 6712
rect 37553 6675 37611 6681
rect 38289 6681 38301 6684
rect 38335 6681 38347 6715
rect 38289 6675 38347 6681
rect 38473 6715 38531 6721
rect 38473 6681 38485 6715
rect 38519 6712 38531 6715
rect 44450 6712 44456 6724
rect 38519 6684 44456 6712
rect 38519 6681 38531 6684
rect 38473 6675 38531 6681
rect 44450 6672 44456 6684
rect 44508 6672 44514 6724
rect 49142 6672 49148 6724
rect 49200 6672 49206 6724
rect 3418 6604 3424 6656
rect 3476 6644 3482 6656
rect 8938 6644 8944 6656
rect 3476 6616 8944 6644
rect 3476 6604 3482 6616
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 1104 6554 49864 6576
rect 1104 6502 7950 6554
rect 8002 6502 8014 6554
rect 8066 6502 8078 6554
rect 8130 6502 8142 6554
rect 8194 6502 8206 6554
rect 8258 6502 17950 6554
rect 18002 6502 18014 6554
rect 18066 6502 18078 6554
rect 18130 6502 18142 6554
rect 18194 6502 18206 6554
rect 18258 6502 27950 6554
rect 28002 6502 28014 6554
rect 28066 6502 28078 6554
rect 28130 6502 28142 6554
rect 28194 6502 28206 6554
rect 28258 6502 37950 6554
rect 38002 6502 38014 6554
rect 38066 6502 38078 6554
rect 38130 6502 38142 6554
rect 38194 6502 38206 6554
rect 38258 6502 47950 6554
rect 48002 6502 48014 6554
rect 48066 6502 48078 6554
rect 48130 6502 48142 6554
rect 48194 6502 48206 6554
rect 48258 6502 49864 6554
rect 1104 6480 49864 6502
rect 1104 6010 49864 6032
rect 1104 5958 2950 6010
rect 3002 5958 3014 6010
rect 3066 5958 3078 6010
rect 3130 5958 3142 6010
rect 3194 5958 3206 6010
rect 3258 5958 12950 6010
rect 13002 5958 13014 6010
rect 13066 5958 13078 6010
rect 13130 5958 13142 6010
rect 13194 5958 13206 6010
rect 13258 5958 22950 6010
rect 23002 5958 23014 6010
rect 23066 5958 23078 6010
rect 23130 5958 23142 6010
rect 23194 5958 23206 6010
rect 23258 5958 32950 6010
rect 33002 5958 33014 6010
rect 33066 5958 33078 6010
rect 33130 5958 33142 6010
rect 33194 5958 33206 6010
rect 33258 5958 42950 6010
rect 43002 5958 43014 6010
rect 43066 5958 43078 6010
rect 43130 5958 43142 6010
rect 43194 5958 43206 6010
rect 43258 5958 49864 6010
rect 1104 5936 49864 5958
rect 46198 5652 46204 5704
rect 46256 5692 46262 5704
rect 47949 5695 48007 5701
rect 47949 5692 47961 5695
rect 46256 5664 47961 5692
rect 46256 5652 46262 5664
rect 47949 5661 47961 5664
rect 47995 5661 48007 5695
rect 47949 5655 48007 5661
rect 49142 5652 49148 5704
rect 49200 5652 49206 5704
rect 1104 5466 49864 5488
rect 1104 5414 7950 5466
rect 8002 5414 8014 5466
rect 8066 5414 8078 5466
rect 8130 5414 8142 5466
rect 8194 5414 8206 5466
rect 8258 5414 17950 5466
rect 18002 5414 18014 5466
rect 18066 5414 18078 5466
rect 18130 5414 18142 5466
rect 18194 5414 18206 5466
rect 18258 5414 27950 5466
rect 28002 5414 28014 5466
rect 28066 5414 28078 5466
rect 28130 5414 28142 5466
rect 28194 5414 28206 5466
rect 28258 5414 37950 5466
rect 38002 5414 38014 5466
rect 38066 5414 38078 5466
rect 38130 5414 38142 5466
rect 38194 5414 38206 5466
rect 38258 5414 47950 5466
rect 48002 5414 48014 5466
rect 48066 5414 48078 5466
rect 48130 5414 48142 5466
rect 48194 5414 48206 5466
rect 48258 5414 49864 5466
rect 1104 5392 49864 5414
rect 3418 5244 3424 5296
rect 3476 5284 3482 5296
rect 9030 5284 9036 5296
rect 3476 5256 9036 5284
rect 3476 5244 3482 5256
rect 9030 5244 9036 5256
rect 9088 5244 9094 5296
rect 30101 5219 30159 5225
rect 30101 5216 30113 5219
rect 29472 5188 30113 5216
rect 29472 5024 29500 5188
rect 30101 5185 30113 5188
rect 30147 5185 30159 5219
rect 30101 5179 30159 5185
rect 29454 4972 29460 5024
rect 29512 4972 29518 5024
rect 30193 5015 30251 5021
rect 30193 4981 30205 5015
rect 30239 5012 30251 5015
rect 47762 5012 47768 5024
rect 30239 4984 47768 5012
rect 30239 4981 30251 4984
rect 30193 4975 30251 4981
rect 47762 4972 47768 4984
rect 47820 4972 47826 5024
rect 49326 4972 49332 5024
rect 49384 4972 49390 5024
rect 1104 4922 49864 4944
rect 1104 4870 2950 4922
rect 3002 4870 3014 4922
rect 3066 4870 3078 4922
rect 3130 4870 3142 4922
rect 3194 4870 3206 4922
rect 3258 4870 12950 4922
rect 13002 4870 13014 4922
rect 13066 4870 13078 4922
rect 13130 4870 13142 4922
rect 13194 4870 13206 4922
rect 13258 4870 22950 4922
rect 23002 4870 23014 4922
rect 23066 4870 23078 4922
rect 23130 4870 23142 4922
rect 23194 4870 23206 4922
rect 23258 4870 32950 4922
rect 33002 4870 33014 4922
rect 33066 4870 33078 4922
rect 33130 4870 33142 4922
rect 33194 4870 33206 4922
rect 33258 4870 42950 4922
rect 43002 4870 43014 4922
rect 43066 4870 43078 4922
rect 43130 4870 43142 4922
rect 43194 4870 43206 4922
rect 43258 4870 49864 4922
rect 1104 4848 49864 4870
rect 10042 4768 10048 4820
rect 10100 4808 10106 4820
rect 29454 4808 29460 4820
rect 10100 4780 29460 4808
rect 10100 4768 10106 4780
rect 29454 4768 29460 4780
rect 29512 4768 29518 4820
rect 24762 4564 24768 4616
rect 24820 4604 24826 4616
rect 47949 4607 48007 4613
rect 47949 4604 47961 4607
rect 24820 4576 47961 4604
rect 24820 4564 24826 4576
rect 47949 4573 47961 4576
rect 47995 4573 48007 4607
rect 47949 4567 48007 4573
rect 49142 4496 49148 4548
rect 49200 4496 49206 4548
rect 1104 4378 49864 4400
rect 1104 4326 7950 4378
rect 8002 4326 8014 4378
rect 8066 4326 8078 4378
rect 8130 4326 8142 4378
rect 8194 4326 8206 4378
rect 8258 4326 17950 4378
rect 18002 4326 18014 4378
rect 18066 4326 18078 4378
rect 18130 4326 18142 4378
rect 18194 4326 18206 4378
rect 18258 4326 27950 4378
rect 28002 4326 28014 4378
rect 28066 4326 28078 4378
rect 28130 4326 28142 4378
rect 28194 4326 28206 4378
rect 28258 4326 37950 4378
rect 38002 4326 38014 4378
rect 38066 4326 38078 4378
rect 38130 4326 38142 4378
rect 38194 4326 38206 4378
rect 38258 4326 47950 4378
rect 48002 4326 48014 4378
rect 48066 4326 48078 4378
rect 48130 4326 48142 4378
rect 48194 4326 48206 4378
rect 48258 4326 49864 4378
rect 1104 4304 49864 4326
rect 33962 4088 33968 4140
rect 34020 4088 34026 4140
rect 38470 4088 38476 4140
rect 38528 4128 38534 4140
rect 39117 4131 39175 4137
rect 39117 4128 39129 4131
rect 38528 4100 39129 4128
rect 38528 4088 38534 4100
rect 39117 4097 39129 4100
rect 39163 4097 39175 4131
rect 39117 4091 39175 4097
rect 40126 4088 40132 4140
rect 40184 4128 40190 4140
rect 43533 4131 43591 4137
rect 43533 4128 43545 4131
rect 40184 4100 43545 4128
rect 40184 4088 40190 4100
rect 43533 4097 43545 4100
rect 43579 4097 43591 4131
rect 43533 4091 43591 4097
rect 46014 4088 46020 4140
rect 46072 4088 46078 4140
rect 48590 4088 48596 4140
rect 48648 4128 48654 4140
rect 48685 4131 48743 4137
rect 48685 4128 48697 4131
rect 48648 4100 48697 4128
rect 48648 4088 48654 4100
rect 48685 4097 48697 4100
rect 48731 4097 48743 4131
rect 48685 4091 48743 4097
rect 33870 4020 33876 4072
rect 33928 4060 33934 4072
rect 34425 4063 34483 4069
rect 34425 4060 34437 4063
rect 33928 4032 34437 4060
rect 33928 4020 33934 4032
rect 34425 4029 34437 4032
rect 34471 4029 34483 4063
rect 34425 4023 34483 4029
rect 39022 4020 39028 4072
rect 39080 4060 39086 4072
rect 39577 4063 39635 4069
rect 39577 4060 39589 4063
rect 39080 4032 39589 4060
rect 39080 4020 39086 4032
rect 39577 4029 39589 4032
rect 39623 4029 39635 4063
rect 39577 4023 39635 4029
rect 43438 4020 43444 4072
rect 43496 4060 43502 4072
rect 43993 4063 44051 4069
rect 43993 4060 44005 4063
rect 43496 4032 44005 4060
rect 43496 4020 43502 4032
rect 43993 4029 44005 4032
rect 44039 4029 44051 4063
rect 43993 4023 44051 4029
rect 36538 3952 36544 4004
rect 36596 3992 36602 4004
rect 46014 3992 46020 4004
rect 36596 3964 46020 3992
rect 36596 3952 36602 3964
rect 46014 3952 46020 3964
rect 46072 3952 46078 4004
rect 48866 3952 48872 4004
rect 48924 3952 48930 4004
rect 45833 3927 45891 3933
rect 45833 3893 45845 3927
rect 45879 3924 45891 3927
rect 47762 3924 47768 3936
rect 45879 3896 47768 3924
rect 45879 3893 45891 3896
rect 45833 3887 45891 3893
rect 47762 3884 47768 3896
rect 47820 3884 47826 3936
rect 1104 3834 49864 3856
rect 1104 3782 2950 3834
rect 3002 3782 3014 3834
rect 3066 3782 3078 3834
rect 3130 3782 3142 3834
rect 3194 3782 3206 3834
rect 3258 3782 12950 3834
rect 13002 3782 13014 3834
rect 13066 3782 13078 3834
rect 13130 3782 13142 3834
rect 13194 3782 13206 3834
rect 13258 3782 22950 3834
rect 23002 3782 23014 3834
rect 23066 3782 23078 3834
rect 23130 3782 23142 3834
rect 23194 3782 23206 3834
rect 23258 3782 32950 3834
rect 33002 3782 33014 3834
rect 33066 3782 33078 3834
rect 33130 3782 33142 3834
rect 33194 3782 33206 3834
rect 33258 3782 42950 3834
rect 43002 3782 43014 3834
rect 43066 3782 43078 3834
rect 43130 3782 43142 3834
rect 43194 3782 43206 3834
rect 43258 3782 49864 3834
rect 1104 3760 49864 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 5534 3720 5540 3732
rect 1627 3692 5540 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 18322 3612 18328 3664
rect 18380 3652 18386 3664
rect 26878 3652 26884 3664
rect 18380 3624 26884 3652
rect 18380 3612 18386 3624
rect 26878 3612 26884 3624
rect 26936 3612 26942 3664
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 25041 3587 25099 3593
rect 25041 3584 25053 3587
rect 24360 3556 25053 3584
rect 24360 3544 24366 3556
rect 25041 3553 25053 3556
rect 25087 3553 25099 3587
rect 25041 3547 25099 3553
rect 29454 3544 29460 3596
rect 29512 3584 29518 3596
rect 30193 3587 30251 3593
rect 30193 3584 30205 3587
rect 29512 3556 30205 3584
rect 29512 3544 29518 3556
rect 30193 3553 30205 3556
rect 30239 3553 30251 3587
rect 30193 3547 30251 3553
rect 30926 3544 30932 3596
rect 30984 3584 30990 3596
rect 32033 3587 32091 3593
rect 32033 3584 32045 3587
rect 30984 3556 32045 3584
rect 30984 3544 30990 3556
rect 32033 3553 32045 3556
rect 32079 3553 32091 3587
rect 32033 3547 32091 3553
rect 34606 3544 34612 3596
rect 34664 3584 34670 3596
rect 35345 3587 35403 3593
rect 35345 3584 35357 3587
rect 34664 3556 35357 3584
rect 34664 3544 34670 3556
rect 35345 3553 35357 3556
rect 35391 3553 35403 3587
rect 35345 3547 35403 3553
rect 36078 3544 36084 3596
rect 36136 3584 36142 3596
rect 37185 3587 37243 3593
rect 37185 3584 37197 3587
rect 36136 3556 37197 3584
rect 36136 3544 36142 3556
rect 37185 3553 37197 3556
rect 37231 3553 37243 3587
rect 37185 3547 37243 3553
rect 39758 3544 39764 3596
rect 39816 3584 39822 3596
rect 40497 3587 40555 3593
rect 40497 3584 40509 3587
rect 39816 3556 40509 3584
rect 39816 3544 39822 3556
rect 40497 3553 40509 3556
rect 40543 3553 40555 3587
rect 40497 3547 40555 3553
rect 41230 3544 41236 3596
rect 41288 3584 41294 3596
rect 42337 3587 42395 3593
rect 42337 3584 42349 3587
rect 41288 3556 42349 3584
rect 41288 3544 41294 3556
rect 42337 3553 42349 3556
rect 42383 3553 42395 3587
rect 42337 3547 42395 3553
rect 44174 3544 44180 3596
rect 44232 3584 44238 3596
rect 45649 3587 45707 3593
rect 45649 3584 45661 3587
rect 44232 3556 45661 3584
rect 44232 3544 44238 3556
rect 45649 3553 45661 3556
rect 45695 3553 45707 3587
rect 45649 3547 45707 3553
rect 1765 3519 1823 3525
rect 1765 3485 1777 3519
rect 1811 3516 1823 3519
rect 2774 3516 2780 3528
rect 1811 3488 2780 3516
rect 1811 3485 1823 3488
rect 1765 3479 1823 3485
rect 2774 3476 2780 3488
rect 2832 3476 2838 3528
rect 24765 3519 24823 3525
rect 24765 3485 24777 3519
rect 24811 3516 24823 3519
rect 25774 3516 25780 3528
rect 24811 3488 25780 3516
rect 24811 3485 24823 3488
rect 24765 3479 24823 3485
rect 25774 3476 25780 3488
rect 25832 3476 25838 3528
rect 29730 3476 29736 3528
rect 29788 3476 29794 3528
rect 30098 3476 30104 3528
rect 30156 3516 30162 3528
rect 31573 3519 31631 3525
rect 31573 3516 31585 3519
rect 30156 3488 31585 3516
rect 30156 3476 30162 3488
rect 31573 3485 31585 3488
rect 31619 3485 31631 3519
rect 31573 3479 31631 3485
rect 34238 3476 34244 3528
rect 34296 3516 34302 3528
rect 34885 3519 34943 3525
rect 34885 3516 34897 3519
rect 34296 3488 34897 3516
rect 34296 3476 34302 3488
rect 34885 3485 34897 3488
rect 34931 3485 34943 3519
rect 34885 3479 34943 3485
rect 36722 3476 36728 3528
rect 36780 3476 36786 3528
rect 37274 3476 37280 3528
rect 37332 3516 37338 3528
rect 40037 3519 40095 3525
rect 40037 3516 40049 3519
rect 37332 3488 40049 3516
rect 37332 3476 37338 3488
rect 40037 3485 40049 3488
rect 40083 3485 40095 3519
rect 40037 3479 40095 3485
rect 41874 3476 41880 3528
rect 41932 3476 41938 3528
rect 45186 3476 45192 3528
rect 45244 3476 45250 3528
rect 47670 3476 47676 3528
rect 47728 3516 47734 3528
rect 47949 3519 48007 3525
rect 47949 3516 47961 3519
rect 47728 3488 47961 3516
rect 47728 3476 47734 3488
rect 47949 3485 47961 3488
rect 47995 3485 48007 3519
rect 47949 3479 48007 3485
rect 49145 3451 49203 3457
rect 49145 3417 49157 3451
rect 49191 3448 49203 3451
rect 49326 3448 49332 3460
rect 49191 3420 49332 3448
rect 49191 3417 49203 3420
rect 49145 3411 49203 3417
rect 49326 3408 49332 3420
rect 49384 3408 49390 3460
rect 12894 3340 12900 3392
rect 12952 3380 12958 3392
rect 26786 3380 26792 3392
rect 12952 3352 26792 3380
rect 12952 3340 12958 3352
rect 26786 3340 26792 3352
rect 26844 3340 26850 3392
rect 1104 3290 49864 3312
rect 1104 3238 7950 3290
rect 8002 3238 8014 3290
rect 8066 3238 8078 3290
rect 8130 3238 8142 3290
rect 8194 3238 8206 3290
rect 8258 3238 17950 3290
rect 18002 3238 18014 3290
rect 18066 3238 18078 3290
rect 18130 3238 18142 3290
rect 18194 3238 18206 3290
rect 18258 3238 27950 3290
rect 28002 3238 28014 3290
rect 28066 3238 28078 3290
rect 28130 3238 28142 3290
rect 28194 3238 28206 3290
rect 28258 3238 37950 3290
rect 38002 3238 38014 3290
rect 38066 3238 38078 3290
rect 38130 3238 38142 3290
rect 38194 3238 38206 3290
rect 38258 3238 47950 3290
rect 48002 3238 48014 3290
rect 48066 3238 48078 3290
rect 48130 3238 48142 3290
rect 48194 3238 48206 3290
rect 48258 3238 49864 3290
rect 1104 3216 49864 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3145 2375 3179
rect 2317 3139 2375 3145
rect 10597 3179 10655 3185
rect 10597 3145 10609 3179
rect 10643 3176 10655 3179
rect 14458 3176 14464 3188
rect 10643 3148 14464 3176
rect 10643 3145 10655 3148
rect 10597 3139 10655 3145
rect 2332 3108 2360 3139
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 19978 3176 19984 3188
rect 14568 3148 19984 3176
rect 7558 3108 7564 3120
rect 2332 3080 7564 3108
rect 7558 3068 7564 3080
rect 7616 3068 7622 3120
rect 10244 3080 12848 3108
rect 1486 3000 1492 3052
rect 1544 3040 1550 3052
rect 1581 3043 1639 3049
rect 1581 3040 1593 3043
rect 1544 3012 1593 3040
rect 1544 3000 1550 3012
rect 1581 3009 1593 3012
rect 1627 3009 1639 3043
rect 2501 3043 2559 3049
rect 2501 3040 2513 3043
rect 1581 3003 1639 3009
rect 1688 3012 2513 3040
rect 750 2932 756 2984
rect 808 2972 814 2984
rect 1688 2972 1716 3012
rect 2501 3009 2513 3012
rect 2547 3009 2559 3043
rect 2501 3003 2559 3009
rect 3694 3000 3700 3052
rect 3752 3040 3758 3052
rect 3881 3043 3939 3049
rect 3881 3040 3893 3043
rect 3752 3012 3893 3040
rect 3752 3000 3758 3012
rect 3881 3009 3893 3012
rect 3927 3009 3939 3043
rect 3881 3003 3939 3009
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5224 3012 5365 3040
rect 5224 3000 5230 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 6638 3000 6644 3052
rect 6696 3040 6702 3052
rect 6825 3043 6883 3049
rect 6825 3040 6837 3043
rect 6696 3012 6837 3040
rect 6696 3000 6702 3012
rect 6825 3009 6837 3012
rect 6871 3009 6883 3043
rect 6825 3003 6883 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 10244 3040 10272 3080
rect 7055 3012 10272 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 10318 3000 10324 3052
rect 10376 3040 10382 3052
rect 10413 3043 10471 3049
rect 10413 3040 10425 3043
rect 10376 3012 10425 3040
rect 10376 3000 10382 3012
rect 10413 3009 10425 3012
rect 10459 3009 10471 3043
rect 10413 3003 10471 3009
rect 12526 3000 12532 3052
rect 12584 3040 12590 3052
rect 12713 3043 12771 3049
rect 12713 3040 12725 3043
rect 12584 3012 12725 3040
rect 12584 3000 12590 3012
rect 12713 3009 12725 3012
rect 12759 3009 12771 3043
rect 12820 3040 12848 3080
rect 12894 3068 12900 3120
rect 12952 3068 12958 3120
rect 14568 3108 14596 3148
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 30558 3176 30564 3188
rect 20916 3148 30564 3176
rect 18414 3108 18420 3120
rect 13004 3080 14596 3108
rect 16546 3080 18420 3108
rect 13004 3040 13032 3080
rect 12820 3012 13032 3040
rect 12713 3003 12771 3009
rect 13998 3000 14004 3052
rect 14056 3040 14062 3052
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 14056 3012 14105 3040
rect 14056 3000 14062 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 14093 3003 14151 3009
rect 16546 2972 16574 3080
rect 18414 3068 18420 3080
rect 18472 3068 18478 3120
rect 17678 3000 17684 3052
rect 17736 3040 17742 3052
rect 17865 3043 17923 3049
rect 17865 3040 17877 3043
rect 17736 3012 17877 3040
rect 17736 3000 17742 3012
rect 17865 3009 17877 3012
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3040 18291 3043
rect 18322 3040 18328 3052
rect 18279 3012 18328 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 20916 3049 20944 3148
rect 30558 3136 30564 3148
rect 30616 3136 30622 3188
rect 47118 3136 47124 3188
rect 47176 3136 47182 3188
rect 25590 3108 25596 3120
rect 22296 3080 25596 3108
rect 22296 3049 22324 3080
rect 25590 3068 25596 3080
rect 25648 3068 25654 3120
rect 37366 3068 37372 3120
rect 37424 3108 37430 3120
rect 37424 3080 39344 3108
rect 37424 3068 37430 3080
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 22281 3043 22339 3049
rect 22281 3009 22293 3043
rect 22327 3009 22339 3043
rect 22281 3003 22339 3009
rect 23385 3043 23443 3049
rect 23385 3009 23397 3043
rect 23431 3040 23443 3043
rect 24670 3040 24676 3052
rect 23431 3012 24676 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 24670 3000 24676 3012
rect 24728 3000 24734 3052
rect 25130 3000 25136 3052
rect 25188 3000 25194 3052
rect 27525 3043 27583 3049
rect 27525 3009 27537 3043
rect 27571 3040 27583 3043
rect 29086 3040 29092 3052
rect 27571 3012 29092 3040
rect 27571 3009 27583 3012
rect 27525 3003 27583 3009
rect 29086 3000 29092 3012
rect 29144 3000 29150 3052
rect 29178 3000 29184 3052
rect 29236 3000 29242 3052
rect 32030 3000 32036 3052
rect 32088 3040 32094 3052
rect 32309 3043 32367 3049
rect 32309 3040 32321 3043
rect 32088 3012 32321 3040
rect 32088 3000 32094 3012
rect 32309 3009 32321 3012
rect 32355 3009 32367 3043
rect 32309 3003 32367 3009
rect 34146 3000 34152 3052
rect 34204 3000 34210 3052
rect 37642 3000 37648 3052
rect 37700 3000 37706 3052
rect 39316 3049 39344 3080
rect 47854 3068 47860 3120
rect 47912 3068 47918 3120
rect 39301 3043 39359 3049
rect 39301 3009 39313 3043
rect 39347 3009 39359 3043
rect 39301 3003 39359 3009
rect 42610 3000 42616 3052
rect 42668 3000 42674 3052
rect 44450 3000 44456 3052
rect 44508 3000 44514 3052
rect 46937 3043 46995 3049
rect 46937 3009 46949 3043
rect 46983 3040 46995 3043
rect 47118 3040 47124 3052
rect 46983 3012 47124 3040
rect 46983 3009 46995 3012
rect 46937 3003 46995 3009
rect 47118 3000 47124 3012
rect 47176 3000 47182 3052
rect 47872 3040 47900 3068
rect 47949 3043 48007 3049
rect 47949 3040 47961 3043
rect 47872 3012 47961 3040
rect 47949 3009 47961 3012
rect 47995 3009 48007 3043
rect 47949 3003 48007 3009
rect 808 2944 1716 2972
rect 1780 2944 16574 2972
rect 808 2932 814 2944
rect 1780 2913 1808 2944
rect 19150 2932 19156 2984
rect 19208 2972 19214 2984
rect 19245 2975 19303 2981
rect 19245 2972 19257 2975
rect 19208 2944 19257 2972
rect 19208 2932 19214 2944
rect 19245 2941 19257 2944
rect 19291 2941 19303 2975
rect 19245 2935 19303 2941
rect 19521 2975 19579 2981
rect 19521 2941 19533 2975
rect 19567 2941 19579 2975
rect 19521 2935 19579 2941
rect 1765 2907 1823 2913
rect 1765 2873 1777 2907
rect 1811 2873 1823 2907
rect 1765 2867 1823 2873
rect 4065 2907 4123 2913
rect 4065 2873 4077 2907
rect 4111 2904 4123 2907
rect 14277 2907 14335 2913
rect 4111 2876 12940 2904
rect 4111 2873 4123 2876
rect 4065 2867 4123 2873
rect 12912 2836 12940 2876
rect 14277 2873 14289 2907
rect 14323 2904 14335 2907
rect 17218 2904 17224 2916
rect 14323 2876 17224 2904
rect 14323 2873 14335 2876
rect 14277 2867 14335 2873
rect 17218 2864 17224 2876
rect 17276 2864 17282 2916
rect 18782 2904 18788 2916
rect 17696 2876 18788 2904
rect 17696 2836 17724 2876
rect 18782 2864 18788 2876
rect 18840 2864 18846 2916
rect 19536 2904 19564 2935
rect 20622 2932 20628 2984
rect 20680 2932 20686 2984
rect 22005 2975 22063 2981
rect 22005 2941 22017 2975
rect 22051 2972 22063 2975
rect 22094 2972 22100 2984
rect 22051 2944 22100 2972
rect 22051 2941 22063 2944
rect 22005 2935 22063 2941
rect 22094 2932 22100 2944
rect 22152 2932 22158 2984
rect 23566 2932 23572 2984
rect 23624 2972 23630 2984
rect 23753 2975 23811 2981
rect 23753 2972 23765 2975
rect 23624 2944 23765 2972
rect 23624 2932 23630 2944
rect 23753 2941 23765 2944
rect 23799 2941 23811 2975
rect 23753 2935 23811 2941
rect 25038 2932 25044 2984
rect 25096 2972 25102 2984
rect 25593 2975 25651 2981
rect 25593 2972 25605 2975
rect 25096 2944 25605 2972
rect 25096 2932 25102 2944
rect 25593 2941 25605 2944
rect 25639 2941 25651 2975
rect 25593 2935 25651 2941
rect 27246 2932 27252 2984
rect 27304 2972 27310 2984
rect 27801 2975 27859 2981
rect 27801 2972 27813 2975
rect 27304 2944 27813 2972
rect 27304 2932 27310 2944
rect 27801 2941 27813 2944
rect 27847 2941 27859 2975
rect 27801 2935 27859 2941
rect 28718 2932 28724 2984
rect 28776 2972 28782 2984
rect 29641 2975 29699 2981
rect 29641 2972 29653 2975
rect 28776 2944 29653 2972
rect 28776 2932 28782 2944
rect 29641 2941 29653 2944
rect 29687 2941 29699 2975
rect 29641 2935 29699 2941
rect 31662 2932 31668 2984
rect 31720 2972 31726 2984
rect 32769 2975 32827 2981
rect 32769 2972 32781 2975
rect 31720 2944 32781 2972
rect 31720 2932 31726 2944
rect 32769 2941 32781 2944
rect 32815 2941 32827 2975
rect 32769 2935 32827 2941
rect 34609 2975 34667 2981
rect 34609 2941 34621 2975
rect 34655 2941 34667 2975
rect 34609 2935 34667 2941
rect 28350 2904 28356 2916
rect 19536 2876 28356 2904
rect 28350 2864 28356 2876
rect 28408 2864 28414 2916
rect 32398 2864 32404 2916
rect 32456 2904 32462 2916
rect 34624 2904 34652 2935
rect 36814 2932 36820 2984
rect 36872 2972 36878 2984
rect 37921 2975 37979 2981
rect 37921 2972 37933 2975
rect 36872 2944 37933 2972
rect 36872 2932 36878 2944
rect 37921 2941 37933 2944
rect 37967 2941 37979 2975
rect 37921 2935 37979 2941
rect 39761 2975 39819 2981
rect 39761 2941 39773 2975
rect 39807 2941 39819 2975
rect 39761 2935 39819 2941
rect 32456 2876 34652 2904
rect 32456 2864 32462 2876
rect 37550 2864 37556 2916
rect 37608 2904 37614 2916
rect 39776 2904 39804 2935
rect 41966 2932 41972 2984
rect 42024 2972 42030 2984
rect 43073 2975 43131 2981
rect 43073 2972 43085 2975
rect 42024 2944 43085 2972
rect 42024 2932 42030 2944
rect 43073 2941 43085 2944
rect 43119 2941 43131 2975
rect 43073 2935 43131 2941
rect 44913 2975 44971 2981
rect 44913 2941 44925 2975
rect 44959 2941 44971 2975
rect 44913 2935 44971 2941
rect 37608 2876 39804 2904
rect 37608 2864 37614 2876
rect 42702 2864 42708 2916
rect 42760 2904 42766 2916
rect 44928 2904 44956 2935
rect 47854 2932 47860 2984
rect 47912 2972 47918 2984
rect 48409 2975 48467 2981
rect 48409 2972 48421 2975
rect 47912 2944 48421 2972
rect 47912 2932 47918 2944
rect 48409 2941 48421 2944
rect 48455 2941 48467 2975
rect 48409 2935 48467 2941
rect 42760 2876 44956 2904
rect 42760 2864 42766 2876
rect 12912 2808 17724 2836
rect 46382 2796 46388 2848
rect 46440 2836 46446 2848
rect 48314 2836 48320 2848
rect 46440 2808 48320 2836
rect 46440 2796 46446 2808
rect 48314 2796 48320 2808
rect 48372 2796 48378 2848
rect 1104 2746 49864 2768
rect 1104 2694 2950 2746
rect 3002 2694 3014 2746
rect 3066 2694 3078 2746
rect 3130 2694 3142 2746
rect 3194 2694 3206 2746
rect 3258 2694 12950 2746
rect 13002 2694 13014 2746
rect 13066 2694 13078 2746
rect 13130 2694 13142 2746
rect 13194 2694 13206 2746
rect 13258 2694 22950 2746
rect 23002 2694 23014 2746
rect 23066 2694 23078 2746
rect 23130 2694 23142 2746
rect 23194 2694 23206 2746
rect 23258 2694 32950 2746
rect 33002 2694 33014 2746
rect 33066 2694 33078 2746
rect 33130 2694 33142 2746
rect 33194 2694 33206 2746
rect 33258 2694 42950 2746
rect 43002 2694 43014 2746
rect 43066 2694 43078 2746
rect 43130 2694 43142 2746
rect 43194 2694 43206 2746
rect 43258 2694 49864 2746
rect 1104 2672 49864 2694
rect 10042 2592 10048 2644
rect 10100 2592 10106 2644
rect 11057 2635 11115 2641
rect 11057 2601 11069 2635
rect 11103 2632 11115 2635
rect 11146 2632 11152 2644
rect 11103 2604 11152 2632
rect 11103 2601 11115 2604
rect 11057 2595 11115 2601
rect 11146 2592 11152 2604
rect 11204 2592 11210 2644
rect 13630 2592 13636 2644
rect 13688 2592 13694 2644
rect 14553 2635 14611 2641
rect 14553 2601 14565 2635
rect 14599 2632 14611 2635
rect 18690 2632 18696 2644
rect 14599 2604 18696 2632
rect 14599 2601 14611 2604
rect 14553 2595 14611 2601
rect 18690 2592 18696 2604
rect 18748 2592 18754 2644
rect 20073 2635 20131 2641
rect 20073 2601 20085 2635
rect 20119 2632 20131 2635
rect 27798 2632 27804 2644
rect 20119 2604 27804 2632
rect 20119 2601 20131 2604
rect 20073 2595 20131 2601
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 46014 2592 46020 2644
rect 46072 2632 46078 2644
rect 46753 2635 46811 2641
rect 46753 2632 46765 2635
rect 46072 2604 46765 2632
rect 46072 2592 46078 2604
rect 46753 2601 46765 2604
rect 46799 2601 46811 2635
rect 46753 2595 46811 2601
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 27706 2564 27712 2576
rect 12299 2536 27712 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 27706 2524 27712 2536
rect 27764 2524 27770 2576
rect 9490 2456 9496 2508
rect 9548 2456 9554 2508
rect 18049 2499 18107 2505
rect 18049 2465 18061 2499
rect 18095 2496 18107 2499
rect 18414 2496 18420 2508
rect 18095 2468 18420 2496
rect 18095 2465 18107 2468
rect 18049 2459 18107 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 20625 2499 20683 2505
rect 20625 2465 20637 2499
rect 20671 2496 20683 2499
rect 21358 2496 21364 2508
rect 20671 2468 21364 2496
rect 20671 2465 20683 2468
rect 20625 2459 20683 2465
rect 21358 2456 21364 2468
rect 21416 2456 21422 2508
rect 22830 2456 22836 2508
rect 22888 2496 22894 2508
rect 23109 2499 23167 2505
rect 23109 2496 23121 2499
rect 22888 2468 23121 2496
rect 22888 2456 22894 2468
rect 23109 2465 23121 2468
rect 23155 2465 23167 2499
rect 23109 2459 23167 2465
rect 25774 2456 25780 2508
rect 25832 2456 25838 2508
rect 26510 2456 26516 2508
rect 26568 2496 26574 2508
rect 27617 2499 27675 2505
rect 27617 2496 27629 2499
rect 26568 2468 27629 2496
rect 26568 2456 26574 2468
rect 27617 2465 27629 2468
rect 27663 2465 27675 2499
rect 27617 2459 27675 2465
rect 28350 2456 28356 2508
rect 28408 2496 28414 2508
rect 30193 2499 30251 2505
rect 30193 2496 30205 2499
rect 28408 2468 30205 2496
rect 28408 2456 28414 2468
rect 30193 2465 30205 2468
rect 30239 2465 30251 2499
rect 30193 2459 30251 2465
rect 30282 2456 30288 2508
rect 30340 2496 30346 2508
rect 32769 2499 32827 2505
rect 32769 2496 32781 2499
rect 30340 2468 32781 2496
rect 30340 2456 30346 2468
rect 32769 2465 32781 2468
rect 32815 2465 32827 2499
rect 32769 2459 32827 2465
rect 35342 2456 35348 2508
rect 35400 2496 35406 2508
rect 37921 2499 37979 2505
rect 37921 2496 37933 2499
rect 35400 2468 37933 2496
rect 35400 2456 35406 2468
rect 37921 2465 37933 2468
rect 37967 2465 37979 2499
rect 37921 2459 37979 2465
rect 38286 2456 38292 2508
rect 38344 2496 38350 2508
rect 40497 2499 40555 2505
rect 40497 2496 40509 2499
rect 38344 2468 40509 2496
rect 38344 2456 38350 2468
rect 40497 2465 40509 2468
rect 40543 2465 40555 2499
rect 40497 2459 40555 2465
rect 40586 2456 40592 2508
rect 40644 2496 40650 2508
rect 43073 2499 43131 2505
rect 43073 2496 43085 2499
rect 40644 2468 43085 2496
rect 40644 2456 40650 2468
rect 43073 2465 43085 2468
rect 43119 2465 43131 2499
rect 43073 2459 43131 2465
rect 48314 2456 48320 2508
rect 48372 2456 48378 2508
rect 2133 2431 2191 2437
rect 2133 2397 2145 2431
rect 2179 2428 2191 2431
rect 2222 2428 2228 2440
rect 2179 2400 2228 2428
rect 2179 2397 2191 2400
rect 2133 2391 2191 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 7285 2431 7343 2437
rect 7285 2397 7297 2431
rect 7331 2428 7343 2431
rect 7374 2428 7380 2440
rect 7331 2400 7380 2428
rect 7331 2397 7343 2400
rect 7285 2391 7343 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 9582 2388 9588 2440
rect 9640 2428 9646 2440
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9640 2400 10241 2428
rect 9640 2388 9646 2400
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14734 2428 14740 2440
rect 14415 2400 14740 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 19797 2431 19855 2437
rect 19797 2397 19809 2431
rect 19843 2428 19855 2431
rect 19886 2428 19892 2440
rect 19843 2400 19892 2428
rect 19843 2397 19855 2400
rect 19797 2391 19855 2397
rect 2958 2320 2964 2372
rect 3016 2360 3022 2372
rect 3053 2363 3111 2369
rect 3053 2360 3065 2363
rect 3016 2332 3065 2360
rect 3016 2320 3022 2332
rect 3053 2329 3065 2332
rect 3099 2329 3111 2363
rect 3053 2323 3111 2329
rect 4430 2320 4436 2372
rect 4488 2360 4494 2372
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 4488 2332 4629 2360
rect 4488 2320 4494 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 4982 2320 4988 2372
rect 5040 2320 5046 2372
rect 5629 2363 5687 2369
rect 5629 2329 5641 2363
rect 5675 2360 5687 2363
rect 5902 2360 5908 2372
rect 5675 2332 5908 2360
rect 5675 2329 5687 2332
rect 5629 2323 5687 2329
rect 5902 2320 5908 2332
rect 5960 2320 5966 2372
rect 5994 2320 6000 2372
rect 6052 2320 6058 2372
rect 7834 2320 7840 2372
rect 7892 2360 7898 2372
rect 8205 2363 8263 2369
rect 8205 2360 8217 2363
rect 7892 2332 8217 2360
rect 7892 2320 7898 2332
rect 8205 2329 8217 2332
rect 8251 2329 8263 2363
rect 8205 2323 8263 2329
rect 8846 2320 8852 2372
rect 8904 2360 8910 2372
rect 9217 2363 9275 2369
rect 9217 2360 9229 2363
rect 8904 2332 9229 2360
rect 8904 2320 8910 2332
rect 9217 2329 9229 2332
rect 9263 2329 9275 2363
rect 9217 2323 9275 2329
rect 10781 2363 10839 2369
rect 10781 2329 10793 2363
rect 10827 2360 10839 2363
rect 11054 2360 11060 2372
rect 10827 2332 11060 2360
rect 10827 2329 10839 2332
rect 10781 2323 10839 2329
rect 11054 2320 11060 2332
rect 11112 2320 11118 2372
rect 11790 2320 11796 2372
rect 11848 2360 11854 2372
rect 11977 2363 12035 2369
rect 11977 2360 11989 2363
rect 11848 2332 11989 2360
rect 11848 2320 11854 2332
rect 11977 2329 11989 2332
rect 12023 2329 12035 2363
rect 11977 2323 12035 2329
rect 13262 2320 13268 2372
rect 13320 2360 13326 2372
rect 13357 2363 13415 2369
rect 13357 2360 13369 2363
rect 13320 2332 13369 2360
rect 13320 2320 13326 2332
rect 13357 2329 13369 2332
rect 13403 2329 13415 2363
rect 13357 2323 13415 2329
rect 15197 2363 15255 2369
rect 15197 2329 15209 2363
rect 15243 2360 15255 2363
rect 15470 2360 15476 2372
rect 15243 2332 15476 2360
rect 15243 2329 15255 2332
rect 15197 2323 15255 2329
rect 15470 2320 15476 2332
rect 15528 2320 15534 2372
rect 15933 2363 15991 2369
rect 15933 2329 15945 2363
rect 15979 2360 15991 2363
rect 16206 2360 16212 2372
rect 15979 2332 16212 2360
rect 15979 2329 15991 2332
rect 15933 2323 15991 2329
rect 16206 2320 16212 2332
rect 16264 2320 16270 2372
rect 16298 2320 16304 2372
rect 16356 2320 16362 2372
rect 16942 2320 16948 2372
rect 17000 2360 17006 2372
rect 17129 2363 17187 2369
rect 17129 2360 17141 2363
rect 17000 2332 17141 2360
rect 17000 2320 17006 2332
rect 17129 2329 17141 2332
rect 17175 2329 17187 2363
rect 18340 2360 18368 2391
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2428 20959 2431
rect 20947 2400 22094 2428
rect 20947 2397 20959 2400
rect 20901 2391 20959 2397
rect 22066 2360 22094 2400
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 25222 2388 25228 2440
rect 25280 2388 25286 2440
rect 27154 2388 27160 2440
rect 27212 2388 27218 2440
rect 29914 2388 29920 2440
rect 29972 2388 29978 2440
rect 32214 2388 32220 2440
rect 32272 2428 32278 2440
rect 32309 2431 32367 2437
rect 32309 2428 32321 2431
rect 32272 2400 32321 2428
rect 32272 2388 32278 2400
rect 32309 2397 32321 2400
rect 32355 2397 32367 2431
rect 32309 2391 32367 2397
rect 33778 2388 33784 2440
rect 33836 2428 33842 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 33836 2400 34897 2428
rect 33836 2388 33842 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 35250 2388 35256 2440
rect 35308 2428 35314 2440
rect 37461 2431 37519 2437
rect 37461 2428 37473 2431
rect 35308 2400 37473 2428
rect 35308 2388 35314 2400
rect 37461 2397 37473 2400
rect 37507 2397 37519 2431
rect 37461 2391 37519 2397
rect 40034 2388 40040 2440
rect 40092 2388 40098 2440
rect 41414 2388 41420 2440
rect 41472 2428 41478 2440
rect 42613 2431 42671 2437
rect 42613 2428 42625 2431
rect 41472 2400 42625 2428
rect 41472 2388 41478 2400
rect 42613 2397 42625 2400
rect 42659 2397 42671 2431
rect 42613 2391 42671 2397
rect 47762 2388 47768 2440
rect 47820 2388 47826 2440
rect 29270 2360 29276 2372
rect 18340 2332 20208 2360
rect 22066 2332 29276 2360
rect 17129 2323 17187 2329
rect 2406 2252 2412 2304
rect 2464 2252 2470 2304
rect 3326 2252 3332 2304
rect 3384 2252 3390 2304
rect 7558 2252 7564 2304
rect 7616 2252 7622 2304
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 15289 2295 15347 2301
rect 15289 2261 15301 2295
rect 15335 2292 15347 2295
rect 17310 2292 17316 2304
rect 15335 2264 17316 2292
rect 15335 2261 15347 2264
rect 15289 2255 15347 2261
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 17402 2252 17408 2304
rect 17460 2252 17466 2304
rect 20180 2292 20208 2332
rect 29270 2320 29276 2332
rect 29328 2320 29334 2372
rect 35805 2363 35863 2369
rect 35805 2329 35817 2363
rect 35851 2329 35863 2363
rect 35805 2323 35863 2329
rect 45465 2363 45523 2369
rect 45465 2329 45477 2363
rect 45511 2360 45523 2363
rect 45646 2360 45652 2372
rect 45511 2332 45652 2360
rect 45511 2329 45523 2332
rect 45465 2323 45523 2329
rect 28810 2292 28816 2304
rect 20180 2264 28816 2292
rect 28810 2252 28816 2264
rect 28868 2252 28874 2304
rect 33134 2252 33140 2304
rect 33192 2292 33198 2304
rect 35820 2292 35848 2323
rect 45646 2320 45652 2332
rect 45704 2320 45710 2372
rect 33192 2264 35848 2292
rect 33192 2252 33198 2264
rect 1104 2202 49864 2224
rect 1104 2150 7950 2202
rect 8002 2150 8014 2202
rect 8066 2150 8078 2202
rect 8130 2150 8142 2202
rect 8194 2150 8206 2202
rect 8258 2150 17950 2202
rect 18002 2150 18014 2202
rect 18066 2150 18078 2202
rect 18130 2150 18142 2202
rect 18194 2150 18206 2202
rect 18258 2150 27950 2202
rect 28002 2150 28014 2202
rect 28066 2150 28078 2202
rect 28130 2150 28142 2202
rect 28194 2150 28206 2202
rect 28258 2150 37950 2202
rect 38002 2150 38014 2202
rect 38066 2150 38078 2202
rect 38130 2150 38142 2202
rect 38194 2150 38206 2202
rect 38258 2150 47950 2202
rect 48002 2150 48014 2202
rect 48066 2150 48078 2202
rect 48130 2150 48142 2202
rect 48194 2150 48206 2202
rect 48258 2150 49864 2202
rect 1104 2128 49864 2150
rect 16298 2048 16304 2100
rect 16356 2088 16362 2100
rect 28442 2088 28448 2100
rect 16356 2060 28448 2088
rect 16356 2048 16362 2060
rect 28442 2048 28448 2060
rect 28500 2048 28506 2100
rect 5994 1980 6000 2032
rect 6052 2020 6058 2032
rect 17126 2020 17132 2032
rect 6052 1992 17132 2020
rect 6052 1980 6058 1992
rect 17126 1980 17132 1992
rect 17184 1980 17190 2032
rect 23750 2020 23756 2032
rect 17236 1992 23756 2020
rect 7558 1912 7564 1964
rect 7616 1952 7622 1964
rect 17236 1952 17264 1992
rect 23750 1980 23756 1992
rect 23808 1980 23814 2032
rect 7616 1924 17264 1952
rect 7616 1912 7622 1924
rect 17310 1912 17316 1964
rect 17368 1952 17374 1964
rect 26786 1952 26792 1964
rect 17368 1924 26792 1952
rect 17368 1912 17374 1924
rect 26786 1912 26792 1924
rect 26844 1912 26850 1964
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 2464 1856 12572 1884
rect 2464 1844 2470 1856
rect 12544 1816 12572 1856
rect 17402 1844 17408 1896
rect 17460 1884 17466 1896
rect 28626 1884 28632 1896
rect 17460 1856 28632 1884
rect 17460 1844 17466 1856
rect 28626 1844 28632 1856
rect 28684 1844 28690 1896
rect 19518 1816 19524 1828
rect 12544 1788 19524 1816
rect 19518 1776 19524 1788
rect 19576 1776 19582 1828
rect 8478 1708 8484 1760
rect 8536 1748 8542 1760
rect 22278 1748 22284 1760
rect 8536 1720 22284 1748
rect 8536 1708 8542 1720
rect 22278 1708 22284 1720
rect 22336 1708 22342 1760
rect 3326 1640 3332 1692
rect 3384 1680 3390 1692
rect 20714 1680 20720 1692
rect 3384 1652 20720 1680
rect 3384 1640 3390 1652
rect 20714 1640 20720 1652
rect 20772 1640 20778 1692
rect 17126 1572 17132 1624
rect 17184 1612 17190 1624
rect 25314 1612 25320 1624
rect 17184 1584 25320 1612
rect 17184 1572 17190 1584
rect 25314 1572 25320 1584
rect 25372 1572 25378 1624
<< via1 >>
rect 388 55700 440 55752
rect 2872 55700 2924 55752
rect 46848 55700 46900 55752
rect 50436 55700 50488 55752
rect 7950 54374 8002 54426
rect 8014 54374 8066 54426
rect 8078 54374 8130 54426
rect 8142 54374 8194 54426
rect 8206 54374 8258 54426
rect 17950 54374 18002 54426
rect 18014 54374 18066 54426
rect 18078 54374 18130 54426
rect 18142 54374 18194 54426
rect 18206 54374 18258 54426
rect 27950 54374 28002 54426
rect 28014 54374 28066 54426
rect 28078 54374 28130 54426
rect 28142 54374 28194 54426
rect 28206 54374 28258 54426
rect 37950 54374 38002 54426
rect 38014 54374 38066 54426
rect 38078 54374 38130 54426
rect 38142 54374 38194 54426
rect 38206 54374 38258 54426
rect 47950 54374 48002 54426
rect 48014 54374 48066 54426
rect 48078 54374 48130 54426
rect 48142 54374 48194 54426
rect 48206 54374 48258 54426
rect 3332 54204 3384 54256
rect 2780 54136 2832 54188
rect 10048 54272 10100 54324
rect 41696 54272 41748 54324
rect 6276 54204 6328 54256
rect 8484 54204 8536 54256
rect 11428 54204 11480 54256
rect 13636 54204 13688 54256
rect 16580 54204 16632 54256
rect 18788 54204 18840 54256
rect 20996 54247 21048 54256
rect 20996 54213 21005 54247
rect 21005 54213 21039 54247
rect 21039 54213 21048 54247
rect 20996 54204 21048 54213
rect 28356 54204 28408 54256
rect 32772 54204 32824 54256
rect 33508 54204 33560 54256
rect 37188 54204 37240 54256
rect 42340 54204 42392 54256
rect 3976 53975 4028 53984
rect 3976 53941 3985 53975
rect 3985 53941 4019 53975
rect 4019 53941 4028 53975
rect 3976 53932 4028 53941
rect 11704 54136 11756 54188
rect 14556 54136 14608 54188
rect 17684 54179 17736 54188
rect 17684 54145 17693 54179
rect 17693 54145 17727 54179
rect 17727 54145 17736 54179
rect 17684 54136 17736 54145
rect 20352 54136 20404 54188
rect 22744 54179 22796 54188
rect 22744 54145 22753 54179
rect 22753 54145 22787 54179
rect 22787 54145 22796 54179
rect 22744 54136 22796 54145
rect 24676 54136 24728 54188
rect 25412 54136 25464 54188
rect 26240 54136 26292 54188
rect 26884 54136 26936 54188
rect 27620 54136 27672 54188
rect 29828 54136 29880 54188
rect 30564 54136 30616 54188
rect 31300 54136 31352 54188
rect 34244 54136 34296 54188
rect 35716 54136 35768 54188
rect 36452 54136 36504 54188
rect 38660 54136 38712 54188
rect 39396 54136 39448 54188
rect 40132 54136 40184 54188
rect 40868 54136 40920 54188
rect 43076 54136 43128 54188
rect 44088 54136 44140 54188
rect 44548 54136 44600 54188
rect 46848 54136 46900 54188
rect 47492 54136 47544 54188
rect 47860 54136 47912 54188
rect 20168 54068 20220 54120
rect 22468 54068 22520 54120
rect 48228 54068 48280 54120
rect 14648 54000 14700 54052
rect 29644 54000 29696 54052
rect 33324 54000 33376 54052
rect 33968 54000 34020 54052
rect 40316 54000 40368 54052
rect 12348 53932 12400 53984
rect 24952 53975 25004 53984
rect 24952 53941 24961 53975
rect 24961 53941 24995 53975
rect 24995 53941 25004 53975
rect 24952 53932 25004 53941
rect 25688 53975 25740 53984
rect 25688 53941 25697 53975
rect 25697 53941 25731 53975
rect 25731 53941 25740 53975
rect 25688 53932 25740 53941
rect 26240 53975 26292 53984
rect 26240 53941 26249 53975
rect 26249 53941 26283 53975
rect 26283 53941 26292 53975
rect 26240 53932 26292 53941
rect 27436 53932 27488 53984
rect 28540 53932 28592 53984
rect 30012 53932 30064 53984
rect 30748 53932 30800 53984
rect 31392 53932 31444 53984
rect 35072 53975 35124 53984
rect 35072 53941 35081 53975
rect 35081 53941 35115 53975
rect 35115 53941 35124 53975
rect 35072 53932 35124 53941
rect 36544 53932 36596 53984
rect 36728 53975 36780 53984
rect 36728 53941 36737 53975
rect 36737 53941 36771 53975
rect 36771 53941 36780 53975
rect 36728 53932 36780 53941
rect 37648 53975 37700 53984
rect 37648 53941 37657 53975
rect 37657 53941 37691 53975
rect 37691 53941 37700 53975
rect 37648 53932 37700 53941
rect 38936 53975 38988 53984
rect 38936 53941 38945 53975
rect 38945 53941 38979 53975
rect 38979 53941 38988 53975
rect 38936 53932 38988 53941
rect 40408 53932 40460 53984
rect 41328 53932 41380 53984
rect 41512 53975 41564 53984
rect 41512 53941 41521 53975
rect 41521 53941 41555 53975
rect 41555 53941 41564 53975
rect 41512 53932 41564 53941
rect 43628 54000 43680 54052
rect 44180 53975 44232 53984
rect 44180 53941 44189 53975
rect 44189 53941 44223 53975
rect 44223 53941 44232 53975
rect 44180 53932 44232 53941
rect 46388 53975 46440 53984
rect 46388 53941 46397 53975
rect 46397 53941 46431 53975
rect 46431 53941 46440 53975
rect 46388 53932 46440 53941
rect 47032 53975 47084 53984
rect 47032 53941 47041 53975
rect 47041 53941 47075 53975
rect 47075 53941 47084 53975
rect 47032 53932 47084 53941
rect 2950 53830 3002 53882
rect 3014 53830 3066 53882
rect 3078 53830 3130 53882
rect 3142 53830 3194 53882
rect 3206 53830 3258 53882
rect 12950 53830 13002 53882
rect 13014 53830 13066 53882
rect 13078 53830 13130 53882
rect 13142 53830 13194 53882
rect 13206 53830 13258 53882
rect 22950 53830 23002 53882
rect 23014 53830 23066 53882
rect 23078 53830 23130 53882
rect 23142 53830 23194 53882
rect 23206 53830 23258 53882
rect 32950 53830 33002 53882
rect 33014 53830 33066 53882
rect 33078 53830 33130 53882
rect 33142 53830 33194 53882
rect 33206 53830 33258 53882
rect 42950 53830 43002 53882
rect 43014 53830 43066 53882
rect 43078 53830 43130 53882
rect 43142 53830 43194 53882
rect 43206 53830 43258 53882
rect 15844 53660 15896 53712
rect 27068 53660 27120 53712
rect 1860 53592 1912 53644
rect 5540 53592 5592 53644
rect 7012 53592 7064 53644
rect 10692 53592 10744 53644
rect 12164 53592 12216 53644
rect 18328 53635 18380 53644
rect 18328 53601 18337 53635
rect 18337 53601 18371 53635
rect 18371 53601 18380 53635
rect 18328 53592 18380 53601
rect 20260 53592 20312 53644
rect 21732 53592 21784 53644
rect 46756 53592 46808 53644
rect 6368 53456 6420 53508
rect 8944 53524 8996 53576
rect 10416 53567 10468 53576
rect 10416 53533 10425 53567
rect 10425 53533 10459 53567
rect 10459 53533 10468 53567
rect 10416 53524 10468 53533
rect 14740 53524 14792 53576
rect 10784 53456 10836 53508
rect 18420 53524 18472 53576
rect 22836 53524 22888 53576
rect 23296 53524 23348 53576
rect 23940 53524 23992 53576
rect 29092 53524 29144 53576
rect 32036 53524 32088 53576
rect 34980 53524 35032 53576
rect 37832 53524 37884 53576
rect 41604 53524 41656 53576
rect 46112 53524 46164 53576
rect 48964 53524 49016 53576
rect 22192 53456 22244 53508
rect 24952 53456 25004 53508
rect 20444 53388 20496 53440
rect 29736 53431 29788 53440
rect 29736 53397 29745 53431
rect 29745 53397 29779 53431
rect 29779 53397 29788 53431
rect 29736 53388 29788 53397
rect 32128 53431 32180 53440
rect 32128 53397 32137 53431
rect 32137 53397 32171 53431
rect 32171 53397 32180 53431
rect 32128 53388 32180 53397
rect 35348 53388 35400 53440
rect 36636 53388 36688 53440
rect 40684 53388 40736 53440
rect 48780 53388 48832 53440
rect 7950 53286 8002 53338
rect 8014 53286 8066 53338
rect 8078 53286 8130 53338
rect 8142 53286 8194 53338
rect 8206 53286 8258 53338
rect 17950 53286 18002 53338
rect 18014 53286 18066 53338
rect 18078 53286 18130 53338
rect 18142 53286 18194 53338
rect 18206 53286 18258 53338
rect 27950 53286 28002 53338
rect 28014 53286 28066 53338
rect 28078 53286 28130 53338
rect 28142 53286 28194 53338
rect 28206 53286 28258 53338
rect 37950 53286 38002 53338
rect 38014 53286 38066 53338
rect 38078 53286 38130 53338
rect 38142 53286 38194 53338
rect 38206 53286 38258 53338
rect 47950 53286 48002 53338
rect 48014 53286 48066 53338
rect 48078 53286 48130 53338
rect 48142 53286 48194 53338
rect 48206 53286 48258 53338
rect 46112 53227 46164 53236
rect 46112 53193 46121 53227
rect 46121 53193 46155 53227
rect 46155 53193 46164 53227
rect 46112 53184 46164 53193
rect 47032 53184 47084 53236
rect 940 53048 992 53100
rect 6276 53116 6328 53168
rect 9864 53116 9916 53168
rect 2596 52980 2648 53032
rect 4896 52980 4948 53032
rect 7748 52980 7800 53032
rect 9772 53091 9824 53100
rect 9772 53057 9781 53091
rect 9781 53057 9815 53091
rect 9815 53057 9824 53091
rect 9772 53048 9824 53057
rect 16948 53116 17000 53168
rect 15200 53048 15252 53100
rect 21272 53116 21324 53168
rect 49700 53116 49752 53168
rect 19616 53091 19668 53100
rect 19616 53057 19625 53091
rect 19625 53057 19659 53091
rect 19659 53057 19668 53091
rect 19616 53048 19668 53057
rect 46940 53048 46992 53100
rect 48320 53048 48372 53100
rect 9956 52980 10008 53032
rect 12808 52980 12860 53032
rect 15108 52980 15160 53032
rect 17316 52980 17368 53032
rect 19524 52980 19576 53032
rect 12440 52912 12492 52964
rect 1676 52844 1728 52896
rect 2950 52742 3002 52794
rect 3014 52742 3066 52794
rect 3078 52742 3130 52794
rect 3142 52742 3194 52794
rect 3206 52742 3258 52794
rect 12950 52742 13002 52794
rect 13014 52742 13066 52794
rect 13078 52742 13130 52794
rect 13142 52742 13194 52794
rect 13206 52742 13258 52794
rect 22950 52742 23002 52794
rect 23014 52742 23066 52794
rect 23078 52742 23130 52794
rect 23142 52742 23194 52794
rect 23206 52742 23258 52794
rect 32950 52742 33002 52794
rect 33014 52742 33066 52794
rect 33078 52742 33130 52794
rect 33142 52742 33194 52794
rect 33206 52742 33258 52794
rect 42950 52742 43002 52794
rect 43014 52742 43066 52794
rect 43078 52742 43130 52794
rect 43142 52742 43194 52794
rect 43206 52742 43258 52794
rect 1124 52504 1176 52556
rect 5816 52572 5868 52624
rect 9220 52572 9272 52624
rect 4068 52504 4120 52556
rect 14372 52504 14424 52556
rect 9220 52436 9272 52488
rect 14464 52436 14516 52488
rect 19156 52436 19208 52488
rect 49332 52479 49384 52488
rect 49332 52445 49341 52479
rect 49341 52445 49375 52479
rect 49375 52445 49384 52479
rect 49332 52436 49384 52445
rect 49148 52343 49200 52352
rect 49148 52309 49157 52343
rect 49157 52309 49191 52343
rect 49191 52309 49200 52343
rect 49148 52300 49200 52309
rect 7950 52198 8002 52250
rect 8014 52198 8066 52250
rect 8078 52198 8130 52250
rect 8142 52198 8194 52250
rect 8206 52198 8258 52250
rect 17950 52198 18002 52250
rect 18014 52198 18066 52250
rect 18078 52198 18130 52250
rect 18142 52198 18194 52250
rect 18206 52198 18258 52250
rect 27950 52198 28002 52250
rect 28014 52198 28066 52250
rect 28078 52198 28130 52250
rect 28142 52198 28194 52250
rect 28206 52198 28258 52250
rect 37950 52198 38002 52250
rect 38014 52198 38066 52250
rect 38078 52198 38130 52250
rect 38142 52198 38194 52250
rect 38206 52198 38258 52250
rect 47950 52198 48002 52250
rect 48014 52198 48066 52250
rect 48078 52198 48130 52250
rect 48142 52198 48194 52250
rect 48206 52198 48258 52250
rect 22744 52096 22796 52148
rect 2872 52028 2924 52080
rect 1584 52003 1636 52012
rect 1584 51969 1593 52003
rect 1593 51969 1627 52003
rect 1627 51969 1636 52003
rect 1584 51960 1636 51969
rect 23756 52003 23808 52012
rect 23756 51969 23765 52003
rect 23765 51969 23799 52003
rect 23799 51969 23808 52003
rect 23756 51960 23808 51969
rect 49056 52003 49108 52012
rect 49056 51969 49065 52003
rect 49065 51969 49099 52003
rect 49099 51969 49108 52003
rect 49056 51960 49108 51969
rect 38384 51756 38436 51808
rect 2950 51654 3002 51706
rect 3014 51654 3066 51706
rect 3078 51654 3130 51706
rect 3142 51654 3194 51706
rect 3206 51654 3258 51706
rect 12950 51654 13002 51706
rect 13014 51654 13066 51706
rect 13078 51654 13130 51706
rect 13142 51654 13194 51706
rect 13206 51654 13258 51706
rect 22950 51654 23002 51706
rect 23014 51654 23066 51706
rect 23078 51654 23130 51706
rect 23142 51654 23194 51706
rect 23206 51654 23258 51706
rect 32950 51654 33002 51706
rect 33014 51654 33066 51706
rect 33078 51654 33130 51706
rect 33142 51654 33194 51706
rect 33206 51654 33258 51706
rect 42950 51654 43002 51706
rect 43014 51654 43066 51706
rect 43078 51654 43130 51706
rect 43142 51654 43194 51706
rect 43206 51654 43258 51706
rect 10048 51552 10100 51604
rect 14464 51595 14516 51604
rect 14464 51561 14473 51595
rect 14473 51561 14507 51595
rect 14507 51561 14516 51595
rect 14464 51552 14516 51561
rect 22836 51552 22888 51604
rect 26700 51348 26752 51400
rect 49056 51391 49108 51400
rect 49056 51357 49065 51391
rect 49065 51357 49099 51391
rect 49099 51357 49108 51391
rect 49056 51348 49108 51357
rect 14280 51280 14332 51332
rect 15936 51280 15988 51332
rect 49332 51212 49384 51264
rect 7950 51110 8002 51162
rect 8014 51110 8066 51162
rect 8078 51110 8130 51162
rect 8142 51110 8194 51162
rect 8206 51110 8258 51162
rect 17950 51110 18002 51162
rect 18014 51110 18066 51162
rect 18078 51110 18130 51162
rect 18142 51110 18194 51162
rect 18206 51110 18258 51162
rect 27950 51110 28002 51162
rect 28014 51110 28066 51162
rect 28078 51110 28130 51162
rect 28142 51110 28194 51162
rect 28206 51110 28258 51162
rect 37950 51110 38002 51162
rect 38014 51110 38066 51162
rect 38078 51110 38130 51162
rect 38142 51110 38194 51162
rect 38206 51110 38258 51162
rect 47950 51110 48002 51162
rect 48014 51110 48066 51162
rect 48078 51110 48130 51162
rect 48142 51110 48194 51162
rect 48206 51110 48258 51162
rect 22192 51051 22244 51060
rect 22192 51017 22201 51051
rect 22201 51017 22235 51051
rect 22235 51017 22244 51051
rect 22192 51008 22244 51017
rect 20352 50940 20404 50992
rect 940 50872 992 50924
rect 22744 50872 22796 50924
rect 24124 50872 24176 50924
rect 48964 50915 49016 50924
rect 48964 50881 48973 50915
rect 48973 50881 49007 50915
rect 49007 50881 49016 50915
rect 48964 50872 49016 50881
rect 1952 50736 2004 50788
rect 38844 50668 38896 50720
rect 2950 50566 3002 50618
rect 3014 50566 3066 50618
rect 3078 50566 3130 50618
rect 3142 50566 3194 50618
rect 3206 50566 3258 50618
rect 12950 50566 13002 50618
rect 13014 50566 13066 50618
rect 13078 50566 13130 50618
rect 13142 50566 13194 50618
rect 13206 50566 13258 50618
rect 22950 50566 23002 50618
rect 23014 50566 23066 50618
rect 23078 50566 23130 50618
rect 23142 50566 23194 50618
rect 23206 50566 23258 50618
rect 32950 50566 33002 50618
rect 33014 50566 33066 50618
rect 33078 50566 33130 50618
rect 33142 50566 33194 50618
rect 33206 50566 33258 50618
rect 42950 50566 43002 50618
rect 43014 50566 43066 50618
rect 43078 50566 43130 50618
rect 43142 50566 43194 50618
rect 43206 50566 43258 50618
rect 17684 50464 17736 50516
rect 49056 50303 49108 50312
rect 49056 50269 49065 50303
rect 49065 50269 49099 50303
rect 49099 50269 49108 50303
rect 49056 50260 49108 50269
rect 22284 50192 22336 50244
rect 48872 50124 48924 50176
rect 7950 50022 8002 50074
rect 8014 50022 8066 50074
rect 8078 50022 8130 50074
rect 8142 50022 8194 50074
rect 8206 50022 8258 50074
rect 17950 50022 18002 50074
rect 18014 50022 18066 50074
rect 18078 50022 18130 50074
rect 18142 50022 18194 50074
rect 18206 50022 18258 50074
rect 27950 50022 28002 50074
rect 28014 50022 28066 50074
rect 28078 50022 28130 50074
rect 28142 50022 28194 50074
rect 28206 50022 28258 50074
rect 37950 50022 38002 50074
rect 38014 50022 38066 50074
rect 38078 50022 38130 50074
rect 38142 50022 38194 50074
rect 38206 50022 38258 50074
rect 47950 50022 48002 50074
rect 48014 50022 48066 50074
rect 48078 50022 48130 50074
rect 48142 50022 48194 50074
rect 48206 50022 48258 50074
rect 12348 49963 12400 49972
rect 12348 49929 12357 49963
rect 12357 49929 12391 49963
rect 12391 49929 12400 49963
rect 12348 49920 12400 49929
rect 14740 49963 14792 49972
rect 14740 49929 14749 49963
rect 14749 49929 14783 49963
rect 14783 49929 14792 49963
rect 14740 49920 14792 49929
rect 46204 49920 46256 49972
rect 20904 49852 20956 49904
rect 16856 49784 16908 49836
rect 49148 49784 49200 49836
rect 2950 49478 3002 49530
rect 3014 49478 3066 49530
rect 3078 49478 3130 49530
rect 3142 49478 3194 49530
rect 3206 49478 3258 49530
rect 12950 49478 13002 49530
rect 13014 49478 13066 49530
rect 13078 49478 13130 49530
rect 13142 49478 13194 49530
rect 13206 49478 13258 49530
rect 22950 49478 23002 49530
rect 23014 49478 23066 49530
rect 23078 49478 23130 49530
rect 23142 49478 23194 49530
rect 23206 49478 23258 49530
rect 32950 49478 33002 49530
rect 33014 49478 33066 49530
rect 33078 49478 33130 49530
rect 33142 49478 33194 49530
rect 33206 49478 33258 49530
rect 42950 49478 43002 49530
rect 43014 49478 43066 49530
rect 43078 49478 43130 49530
rect 43142 49478 43194 49530
rect 43206 49478 43258 49530
rect 15200 49376 15252 49428
rect 18420 49376 18472 49428
rect 20628 49172 20680 49224
rect 49240 49172 49292 49224
rect 22192 49104 22244 49156
rect 38660 49036 38712 49088
rect 7950 48934 8002 48986
rect 8014 48934 8066 48986
rect 8078 48934 8130 48986
rect 8142 48934 8194 48986
rect 8206 48934 8258 48986
rect 17950 48934 18002 48986
rect 18014 48934 18066 48986
rect 18078 48934 18130 48986
rect 18142 48934 18194 48986
rect 18206 48934 18258 48986
rect 27950 48934 28002 48986
rect 28014 48934 28066 48986
rect 28078 48934 28130 48986
rect 28142 48934 28194 48986
rect 28206 48934 28258 48986
rect 37950 48934 38002 48986
rect 38014 48934 38066 48986
rect 38078 48934 38130 48986
rect 38142 48934 38194 48986
rect 38206 48934 38258 48986
rect 47950 48934 48002 48986
rect 48014 48934 48066 48986
rect 48078 48934 48130 48986
rect 48142 48934 48194 48986
rect 48206 48934 48258 48986
rect 49056 48739 49108 48748
rect 49056 48705 49065 48739
rect 49065 48705 49099 48739
rect 49099 48705 49108 48739
rect 49056 48696 49108 48705
rect 40776 48492 40828 48544
rect 2950 48390 3002 48442
rect 3014 48390 3066 48442
rect 3078 48390 3130 48442
rect 3142 48390 3194 48442
rect 3206 48390 3258 48442
rect 12950 48390 13002 48442
rect 13014 48390 13066 48442
rect 13078 48390 13130 48442
rect 13142 48390 13194 48442
rect 13206 48390 13258 48442
rect 22950 48390 23002 48442
rect 23014 48390 23066 48442
rect 23078 48390 23130 48442
rect 23142 48390 23194 48442
rect 23206 48390 23258 48442
rect 32950 48390 33002 48442
rect 33014 48390 33066 48442
rect 33078 48390 33130 48442
rect 33142 48390 33194 48442
rect 33206 48390 33258 48442
rect 42950 48390 43002 48442
rect 43014 48390 43066 48442
rect 43078 48390 43130 48442
rect 43142 48390 43194 48442
rect 43206 48390 43258 48442
rect 46388 48220 46440 48272
rect 48320 48220 48372 48272
rect 21088 48152 21140 48204
rect 47768 48084 47820 48136
rect 940 48016 992 48068
rect 1860 48059 1912 48068
rect 1860 48025 1869 48059
rect 1869 48025 1903 48059
rect 1903 48025 1912 48059
rect 1860 48016 1912 48025
rect 3976 48016 4028 48068
rect 11980 48016 12032 48068
rect 22100 48016 22152 48068
rect 7950 47846 8002 47898
rect 8014 47846 8066 47898
rect 8078 47846 8130 47898
rect 8142 47846 8194 47898
rect 8206 47846 8258 47898
rect 17950 47846 18002 47898
rect 18014 47846 18066 47898
rect 18078 47846 18130 47898
rect 18142 47846 18194 47898
rect 18206 47846 18258 47898
rect 27950 47846 28002 47898
rect 28014 47846 28066 47898
rect 28078 47846 28130 47898
rect 28142 47846 28194 47898
rect 28206 47846 28258 47898
rect 37950 47846 38002 47898
rect 38014 47846 38066 47898
rect 38078 47846 38130 47898
rect 38142 47846 38194 47898
rect 38206 47846 38258 47898
rect 47950 47846 48002 47898
rect 48014 47846 48066 47898
rect 48078 47846 48130 47898
rect 48142 47846 48194 47898
rect 48206 47846 48258 47898
rect 23756 47744 23808 47796
rect 24860 47651 24912 47660
rect 24860 47617 24869 47651
rect 24869 47617 24903 47651
rect 24903 47617 24912 47651
rect 24860 47608 24912 47617
rect 49056 47651 49108 47660
rect 49056 47617 49065 47651
rect 49065 47617 49099 47651
rect 49099 47617 49108 47651
rect 49056 47608 49108 47617
rect 41052 47404 41104 47456
rect 2950 47302 3002 47354
rect 3014 47302 3066 47354
rect 3078 47302 3130 47354
rect 3142 47302 3194 47354
rect 3206 47302 3258 47354
rect 12950 47302 13002 47354
rect 13014 47302 13066 47354
rect 13078 47302 13130 47354
rect 13142 47302 13194 47354
rect 13206 47302 13258 47354
rect 22950 47302 23002 47354
rect 23014 47302 23066 47354
rect 23078 47302 23130 47354
rect 23142 47302 23194 47354
rect 23206 47302 23258 47354
rect 32950 47302 33002 47354
rect 33014 47302 33066 47354
rect 33078 47302 33130 47354
rect 33142 47302 33194 47354
rect 33206 47302 33258 47354
rect 42950 47302 43002 47354
rect 43014 47302 43066 47354
rect 43078 47302 43130 47354
rect 43142 47302 43194 47354
rect 43206 47302 43258 47354
rect 47860 47200 47912 47252
rect 48780 47243 48832 47252
rect 48780 47209 48789 47243
rect 48789 47209 48823 47243
rect 48823 47209 48832 47243
rect 48780 47200 48832 47209
rect 48412 46928 48464 46980
rect 7950 46758 8002 46810
rect 8014 46758 8066 46810
rect 8078 46758 8130 46810
rect 8142 46758 8194 46810
rect 8206 46758 8258 46810
rect 17950 46758 18002 46810
rect 18014 46758 18066 46810
rect 18078 46758 18130 46810
rect 18142 46758 18194 46810
rect 18206 46758 18258 46810
rect 27950 46758 28002 46810
rect 28014 46758 28066 46810
rect 28078 46758 28130 46810
rect 28142 46758 28194 46810
rect 28206 46758 28258 46810
rect 37950 46758 38002 46810
rect 38014 46758 38066 46810
rect 38078 46758 38130 46810
rect 38142 46758 38194 46810
rect 38206 46758 38258 46810
rect 47950 46758 48002 46810
rect 48014 46758 48066 46810
rect 48078 46758 48130 46810
rect 48142 46758 48194 46810
rect 48206 46758 48258 46810
rect 49332 46563 49384 46572
rect 49332 46529 49341 46563
rect 49341 46529 49375 46563
rect 49375 46529 49384 46563
rect 49332 46520 49384 46529
rect 48688 46316 48740 46368
rect 2950 46214 3002 46266
rect 3014 46214 3066 46266
rect 3078 46214 3130 46266
rect 3142 46214 3194 46266
rect 3206 46214 3258 46266
rect 12950 46214 13002 46266
rect 13014 46214 13066 46266
rect 13078 46214 13130 46266
rect 13142 46214 13194 46266
rect 13206 46214 13258 46266
rect 22950 46214 23002 46266
rect 23014 46214 23066 46266
rect 23078 46214 23130 46266
rect 23142 46214 23194 46266
rect 23206 46214 23258 46266
rect 32950 46214 33002 46266
rect 33014 46214 33066 46266
rect 33078 46214 33130 46266
rect 33142 46214 33194 46266
rect 33206 46214 33258 46266
rect 42950 46214 43002 46266
rect 43014 46214 43066 46266
rect 43078 46214 43130 46266
rect 43142 46214 43194 46266
rect 43206 46214 43258 46266
rect 15936 46112 15988 46164
rect 26700 46155 26752 46164
rect 26700 46121 26709 46155
rect 26709 46121 26743 46155
rect 26743 46121 26752 46155
rect 26700 46112 26752 46121
rect 940 45840 992 45892
rect 14280 45840 14332 45892
rect 22008 45908 22060 45960
rect 27712 45908 27764 45960
rect 48596 45908 48648 45960
rect 1768 45815 1820 45824
rect 1768 45781 1777 45815
rect 1777 45781 1811 45815
rect 1811 45781 1820 45815
rect 1768 45772 1820 45781
rect 20536 45840 20588 45892
rect 49148 45883 49200 45892
rect 49148 45849 49157 45883
rect 49157 45849 49191 45883
rect 49191 45849 49200 45883
rect 49148 45840 49200 45849
rect 7950 45670 8002 45722
rect 8014 45670 8066 45722
rect 8078 45670 8130 45722
rect 8142 45670 8194 45722
rect 8206 45670 8258 45722
rect 17950 45670 18002 45722
rect 18014 45670 18066 45722
rect 18078 45670 18130 45722
rect 18142 45670 18194 45722
rect 18206 45670 18258 45722
rect 27950 45670 28002 45722
rect 28014 45670 28066 45722
rect 28078 45670 28130 45722
rect 28142 45670 28194 45722
rect 28206 45670 28258 45722
rect 37950 45670 38002 45722
rect 38014 45670 38066 45722
rect 38078 45670 38130 45722
rect 38142 45670 38194 45722
rect 38206 45670 38258 45722
rect 47950 45670 48002 45722
rect 48014 45670 48066 45722
rect 48078 45670 48130 45722
rect 48142 45670 48194 45722
rect 48206 45670 48258 45722
rect 1768 45568 1820 45620
rect 22468 45568 22520 45620
rect 48596 45611 48648 45620
rect 48596 45577 48605 45611
rect 48605 45577 48639 45611
rect 48639 45577 48648 45611
rect 48596 45568 48648 45577
rect 10416 45500 10468 45552
rect 32128 45500 32180 45552
rect 33968 45543 34020 45552
rect 33968 45509 33977 45543
rect 33977 45509 34011 45543
rect 34011 45509 34020 45543
rect 33968 45500 34020 45509
rect 46940 45500 46992 45552
rect 14924 45475 14976 45484
rect 14924 45441 14933 45475
rect 14933 45441 14967 45475
rect 14967 45441 14976 45475
rect 14924 45432 14976 45441
rect 29736 45432 29788 45484
rect 33324 45432 33376 45484
rect 47860 45432 47912 45484
rect 32864 45407 32916 45416
rect 32864 45373 32873 45407
rect 32873 45373 32907 45407
rect 32907 45373 32916 45407
rect 32864 45364 32916 45373
rect 34152 45407 34204 45416
rect 34152 45373 34161 45407
rect 34161 45373 34195 45407
rect 34195 45373 34204 45407
rect 34152 45364 34204 45373
rect 49056 45296 49108 45348
rect 32680 45228 32732 45280
rect 33508 45271 33560 45280
rect 33508 45237 33517 45271
rect 33517 45237 33551 45271
rect 33551 45237 33560 45271
rect 33508 45228 33560 45237
rect 2950 45126 3002 45178
rect 3014 45126 3066 45178
rect 3078 45126 3130 45178
rect 3142 45126 3194 45178
rect 3206 45126 3258 45178
rect 12950 45126 13002 45178
rect 13014 45126 13066 45178
rect 13078 45126 13130 45178
rect 13142 45126 13194 45178
rect 13206 45126 13258 45178
rect 22950 45126 23002 45178
rect 23014 45126 23066 45178
rect 23078 45126 23130 45178
rect 23142 45126 23194 45178
rect 23206 45126 23258 45178
rect 32950 45126 33002 45178
rect 33014 45126 33066 45178
rect 33078 45126 33130 45178
rect 33142 45126 33194 45178
rect 33206 45126 33258 45178
rect 42950 45126 43002 45178
rect 43014 45126 43066 45178
rect 43078 45126 43130 45178
rect 43142 45126 43194 45178
rect 43206 45126 43258 45178
rect 22744 45024 22796 45076
rect 24124 45024 24176 45076
rect 35348 44931 35400 44940
rect 35348 44897 35357 44931
rect 35357 44897 35391 44931
rect 35391 44897 35400 44931
rect 35348 44888 35400 44897
rect 35532 44931 35584 44940
rect 35532 44897 35541 44931
rect 35541 44897 35575 44931
rect 35575 44897 35584 44931
rect 35532 44888 35584 44897
rect 24492 44820 24544 44872
rect 27160 44820 27212 44872
rect 38568 44820 38620 44872
rect 48504 44863 48556 44872
rect 48504 44829 48513 44863
rect 48513 44829 48547 44863
rect 48547 44829 48556 44863
rect 48504 44820 48556 44829
rect 32404 44752 32456 44804
rect 35072 44752 35124 44804
rect 34888 44727 34940 44736
rect 34888 44693 34897 44727
rect 34897 44693 34931 44727
rect 34931 44693 34940 44727
rect 34888 44684 34940 44693
rect 7950 44582 8002 44634
rect 8014 44582 8066 44634
rect 8078 44582 8130 44634
rect 8142 44582 8194 44634
rect 8206 44582 8258 44634
rect 17950 44582 18002 44634
rect 18014 44582 18066 44634
rect 18078 44582 18130 44634
rect 18142 44582 18194 44634
rect 18206 44582 18258 44634
rect 27950 44582 28002 44634
rect 28014 44582 28066 44634
rect 28078 44582 28130 44634
rect 28142 44582 28194 44634
rect 28206 44582 28258 44634
rect 37950 44582 38002 44634
rect 38014 44582 38066 44634
rect 38078 44582 38130 44634
rect 38142 44582 38194 44634
rect 38206 44582 38258 44634
rect 47950 44582 48002 44634
rect 48014 44582 48066 44634
rect 48078 44582 48130 44634
rect 48142 44582 48194 44634
rect 48206 44582 48258 44634
rect 9772 44480 9824 44532
rect 35440 44480 35492 44532
rect 36544 44523 36596 44532
rect 36544 44489 36553 44523
rect 36553 44489 36587 44523
rect 36587 44489 36596 44523
rect 36544 44480 36596 44489
rect 36636 44523 36688 44532
rect 36636 44489 36645 44523
rect 36645 44489 36679 44523
rect 36679 44489 36688 44523
rect 36636 44480 36688 44489
rect 40684 44480 40736 44532
rect 14464 44344 14516 44396
rect 37648 44344 37700 44396
rect 49332 44387 49384 44396
rect 49332 44353 49341 44387
rect 49341 44353 49375 44387
rect 49375 44353 49384 44387
rect 49332 44344 49384 44353
rect 36912 44276 36964 44328
rect 39304 44319 39356 44328
rect 39304 44285 39313 44319
rect 39313 44285 39347 44319
rect 39347 44285 39356 44319
rect 39304 44276 39356 44285
rect 36176 44183 36228 44192
rect 36176 44149 36185 44183
rect 36185 44149 36219 44183
rect 36219 44149 36228 44183
rect 36176 44140 36228 44149
rect 36544 44140 36596 44192
rect 37648 44140 37700 44192
rect 38752 44183 38804 44192
rect 38752 44149 38761 44183
rect 38761 44149 38795 44183
rect 38795 44149 38804 44183
rect 38752 44140 38804 44149
rect 43444 44140 43496 44192
rect 2950 44038 3002 44090
rect 3014 44038 3066 44090
rect 3078 44038 3130 44090
rect 3142 44038 3194 44090
rect 3206 44038 3258 44090
rect 12950 44038 13002 44090
rect 13014 44038 13066 44090
rect 13078 44038 13130 44090
rect 13142 44038 13194 44090
rect 13206 44038 13258 44090
rect 22950 44038 23002 44090
rect 23014 44038 23066 44090
rect 23078 44038 23130 44090
rect 23142 44038 23194 44090
rect 23206 44038 23258 44090
rect 32950 44038 33002 44090
rect 33014 44038 33066 44090
rect 33078 44038 33130 44090
rect 33142 44038 33194 44090
rect 33206 44038 33258 44090
rect 42950 44038 43002 44090
rect 43014 44038 43066 44090
rect 43078 44038 43130 44090
rect 43142 44038 43194 44090
rect 43206 44038 43258 44090
rect 11704 43936 11756 43988
rect 14648 43936 14700 43988
rect 16948 43979 17000 43988
rect 16948 43945 16957 43979
rect 16957 43945 16991 43979
rect 16991 43945 17000 43979
rect 16948 43936 17000 43945
rect 20444 43979 20496 43988
rect 20444 43945 20453 43979
rect 20453 43945 20487 43979
rect 20487 43945 20496 43979
rect 20444 43936 20496 43945
rect 21272 43979 21324 43988
rect 21272 43945 21281 43979
rect 21281 43945 21315 43979
rect 21315 43945 21324 43979
rect 21272 43936 21324 43945
rect 22284 43979 22336 43988
rect 22284 43945 22293 43979
rect 22293 43945 22327 43979
rect 22327 43945 22336 43979
rect 22284 43936 22336 43945
rect 32036 43936 32088 43988
rect 12440 43911 12492 43920
rect 12440 43877 12449 43911
rect 12449 43877 12483 43911
rect 12483 43877 12492 43911
rect 12440 43868 12492 43877
rect 19616 43868 19668 43920
rect 28816 43868 28868 43920
rect 29000 43843 29052 43852
rect 29000 43809 29009 43843
rect 29009 43809 29043 43843
rect 29043 43809 29052 43843
rect 29000 43800 29052 43809
rect 32956 43800 33008 43852
rect 38292 43800 38344 43852
rect 940 43732 992 43784
rect 21916 43732 21968 43784
rect 23296 43732 23348 43784
rect 26240 43732 26292 43784
rect 13452 43707 13504 43716
rect 13452 43673 13461 43707
rect 13461 43673 13495 43707
rect 13495 43673 13504 43707
rect 13452 43664 13504 43673
rect 2044 43596 2096 43648
rect 19984 43664 20036 43716
rect 20444 43664 20496 43716
rect 28632 43732 28684 43784
rect 32312 43775 32364 43784
rect 32312 43741 32321 43775
rect 32321 43741 32355 43775
rect 32355 43741 32364 43775
rect 32312 43732 32364 43741
rect 41512 43732 41564 43784
rect 48504 43775 48556 43784
rect 48504 43741 48513 43775
rect 48513 43741 48547 43775
rect 48547 43741 48556 43775
rect 48504 43732 48556 43741
rect 20996 43596 21048 43648
rect 24216 43596 24268 43648
rect 31668 43664 31720 43716
rect 30656 43596 30708 43648
rect 31760 43596 31812 43648
rect 33600 43664 33652 43716
rect 33324 43596 33376 43648
rect 33416 43596 33468 43648
rect 36728 43664 36780 43716
rect 40960 43664 41012 43716
rect 37280 43639 37332 43648
rect 37280 43605 37289 43639
rect 37289 43605 37323 43639
rect 37323 43605 37332 43639
rect 37280 43596 37332 43605
rect 7950 43494 8002 43546
rect 8014 43494 8066 43546
rect 8078 43494 8130 43546
rect 8142 43494 8194 43546
rect 8206 43494 8258 43546
rect 17950 43494 18002 43546
rect 18014 43494 18066 43546
rect 18078 43494 18130 43546
rect 18142 43494 18194 43546
rect 18206 43494 18258 43546
rect 27950 43494 28002 43546
rect 28014 43494 28066 43546
rect 28078 43494 28130 43546
rect 28142 43494 28194 43546
rect 28206 43494 28258 43546
rect 37950 43494 38002 43546
rect 38014 43494 38066 43546
rect 38078 43494 38130 43546
rect 38142 43494 38194 43546
rect 38206 43494 38258 43546
rect 47950 43494 48002 43546
rect 48014 43494 48066 43546
rect 48078 43494 48130 43546
rect 48142 43494 48194 43546
rect 48206 43494 48258 43546
rect 2044 43435 2096 43444
rect 2044 43401 2053 43435
rect 2053 43401 2087 43435
rect 2087 43401 2096 43435
rect 2044 43392 2096 43401
rect 8944 43392 8996 43444
rect 16856 43435 16908 43444
rect 16856 43401 16865 43435
rect 16865 43401 16899 43435
rect 16899 43401 16908 43435
rect 16856 43392 16908 43401
rect 19156 43435 19208 43444
rect 19156 43401 19165 43435
rect 19165 43401 19199 43435
rect 19199 43401 19208 43435
rect 19156 43392 19208 43401
rect 20352 43435 20404 43444
rect 20352 43401 20361 43435
rect 20361 43401 20395 43435
rect 20395 43401 20404 43435
rect 20352 43392 20404 43401
rect 20904 43435 20956 43444
rect 20904 43401 20913 43435
rect 20913 43401 20947 43435
rect 20947 43401 20956 43435
rect 20904 43392 20956 43401
rect 20996 43392 21048 43444
rect 24400 43392 24452 43444
rect 24860 43392 24912 43444
rect 28816 43392 28868 43444
rect 31392 43392 31444 43444
rect 32312 43392 32364 43444
rect 31668 43324 31720 43376
rect 40316 43435 40368 43444
rect 40316 43401 40325 43435
rect 40325 43401 40359 43435
rect 40359 43401 40368 43435
rect 40316 43392 40368 43401
rect 34796 43367 34848 43376
rect 34796 43333 34805 43367
rect 34805 43333 34839 43367
rect 34839 43333 34848 43367
rect 34796 43324 34848 43333
rect 11980 43256 12032 43308
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 19064 43299 19116 43308
rect 19064 43265 19073 43299
rect 19073 43265 19107 43299
rect 19107 43265 19116 43299
rect 19064 43256 19116 43265
rect 20260 43299 20312 43308
rect 20260 43265 20269 43299
rect 20269 43265 20303 43299
rect 20303 43265 20312 43299
rect 20260 43256 20312 43265
rect 21732 43256 21784 43308
rect 25964 43256 26016 43308
rect 32312 43299 32364 43308
rect 32312 43265 32321 43299
rect 32321 43265 32355 43299
rect 32355 43265 32364 43299
rect 32312 43256 32364 43265
rect 33600 43256 33652 43308
rect 19432 43188 19484 43240
rect 26332 43231 26384 43240
rect 26332 43197 26341 43231
rect 26341 43197 26375 43231
rect 26375 43197 26384 43231
rect 26332 43188 26384 43197
rect 27344 43188 27396 43240
rect 28632 43188 28684 43240
rect 31852 43188 31904 43240
rect 34520 43299 34572 43308
rect 34520 43265 34529 43299
rect 34529 43265 34563 43299
rect 34563 43265 34572 43299
rect 34520 43256 34572 43265
rect 38936 43256 38988 43308
rect 39856 43256 39908 43308
rect 13452 43120 13504 43172
rect 24032 43120 24084 43172
rect 35992 43188 36044 43240
rect 40592 43188 40644 43240
rect 42064 43188 42116 43240
rect 48504 43231 48556 43240
rect 48504 43197 48513 43231
rect 48513 43197 48547 43231
rect 48547 43197 48556 43231
rect 48504 43188 48556 43197
rect 34152 43120 34204 43172
rect 28908 43052 28960 43104
rect 34060 43095 34112 43104
rect 34060 43061 34069 43095
rect 34069 43061 34103 43095
rect 34103 43061 34112 43095
rect 34060 43052 34112 43061
rect 41236 43052 41288 43104
rect 2950 42950 3002 43002
rect 3014 42950 3066 43002
rect 3078 42950 3130 43002
rect 3142 42950 3194 43002
rect 3206 42950 3258 43002
rect 12950 42950 13002 43002
rect 13014 42950 13066 43002
rect 13078 42950 13130 43002
rect 13142 42950 13194 43002
rect 13206 42950 13258 43002
rect 22950 42950 23002 43002
rect 23014 42950 23066 43002
rect 23078 42950 23130 43002
rect 23142 42950 23194 43002
rect 23206 42950 23258 43002
rect 32950 42950 33002 43002
rect 33014 42950 33066 43002
rect 33078 42950 33130 43002
rect 33142 42950 33194 43002
rect 33206 42950 33258 43002
rect 42950 42950 43002 43002
rect 43014 42950 43066 43002
rect 43078 42950 43130 43002
rect 43142 42950 43194 43002
rect 43206 42950 43258 43002
rect 12072 42848 12124 42900
rect 21548 42848 21600 42900
rect 27344 42891 27396 42900
rect 27344 42857 27353 42891
rect 27353 42857 27387 42891
rect 27387 42857 27396 42891
rect 27344 42848 27396 42857
rect 40040 42780 40092 42832
rect 36912 42712 36964 42764
rect 24124 42644 24176 42696
rect 34520 42644 34572 42696
rect 37004 42644 37056 42696
rect 44180 42644 44232 42696
rect 48504 42687 48556 42696
rect 48504 42653 48513 42687
rect 48513 42653 48547 42687
rect 48547 42653 48556 42687
rect 48504 42644 48556 42653
rect 25872 42619 25924 42628
rect 25872 42585 25881 42619
rect 25881 42585 25915 42619
rect 25915 42585 25924 42619
rect 25872 42576 25924 42585
rect 26148 42576 26200 42628
rect 27252 42508 27304 42560
rect 36820 42508 36872 42560
rect 40224 42508 40276 42560
rect 40408 42551 40460 42560
rect 40408 42517 40417 42551
rect 40417 42517 40451 42551
rect 40451 42517 40460 42551
rect 40408 42508 40460 42517
rect 40500 42508 40552 42560
rect 7950 42406 8002 42458
rect 8014 42406 8066 42458
rect 8078 42406 8130 42458
rect 8142 42406 8194 42458
rect 8206 42406 8258 42458
rect 17950 42406 18002 42458
rect 18014 42406 18066 42458
rect 18078 42406 18130 42458
rect 18142 42406 18194 42458
rect 18206 42406 18258 42458
rect 27950 42406 28002 42458
rect 28014 42406 28066 42458
rect 28078 42406 28130 42458
rect 28142 42406 28194 42458
rect 28206 42406 28258 42458
rect 37950 42406 38002 42458
rect 38014 42406 38066 42458
rect 38078 42406 38130 42458
rect 38142 42406 38194 42458
rect 38206 42406 38258 42458
rect 47950 42406 48002 42458
rect 48014 42406 48066 42458
rect 48078 42406 48130 42458
rect 48142 42406 48194 42458
rect 48206 42406 48258 42458
rect 6368 42304 6420 42356
rect 9220 42347 9272 42356
rect 9220 42313 9229 42347
rect 9229 42313 9263 42347
rect 9263 42313 9272 42347
rect 9220 42304 9272 42313
rect 14556 42304 14608 42356
rect 20628 42347 20680 42356
rect 20628 42313 20637 42347
rect 20637 42313 20671 42347
rect 20671 42313 20680 42347
rect 20628 42304 20680 42313
rect 22192 42347 22244 42356
rect 22192 42313 22201 42347
rect 22201 42313 22235 42347
rect 22235 42313 22244 42347
rect 22192 42304 22244 42313
rect 25872 42347 25924 42356
rect 25872 42313 25881 42347
rect 25881 42313 25915 42347
rect 25915 42313 25924 42347
rect 25872 42304 25924 42313
rect 6276 42236 6328 42288
rect 24308 42236 24360 42288
rect 24860 42236 24912 42288
rect 7196 42211 7248 42220
rect 7196 42177 7205 42211
rect 7205 42177 7239 42211
rect 7239 42177 7248 42211
rect 7196 42168 7248 42177
rect 9128 42211 9180 42220
rect 9128 42177 9137 42211
rect 9137 42177 9171 42211
rect 9171 42177 9180 42211
rect 9128 42168 9180 42177
rect 17408 42168 17460 42220
rect 20812 42211 20864 42220
rect 20812 42177 20821 42211
rect 20821 42177 20855 42211
rect 20855 42177 20864 42211
rect 20812 42168 20864 42177
rect 22376 42211 22428 42220
rect 22376 42177 22385 42211
rect 22385 42177 22419 42211
rect 22419 42177 22428 42211
rect 22376 42168 22428 42177
rect 27344 42236 27396 42288
rect 31760 42304 31812 42356
rect 32772 42304 32824 42356
rect 34520 42304 34572 42356
rect 38292 42304 38344 42356
rect 41604 42347 41656 42356
rect 41604 42313 41613 42347
rect 41613 42313 41647 42347
rect 41647 42313 41656 42347
rect 41604 42304 41656 42313
rect 31668 42236 31720 42288
rect 35992 42236 36044 42288
rect 37004 42236 37056 42288
rect 17316 42100 17368 42152
rect 24124 42143 24176 42152
rect 24124 42109 24133 42143
rect 24133 42109 24167 42143
rect 24167 42109 24176 42143
rect 24124 42100 24176 42109
rect 27344 42100 27396 42152
rect 1584 42032 1636 42084
rect 23756 42032 23808 42084
rect 25872 41964 25924 42016
rect 26516 41964 26568 42016
rect 27252 41964 27304 42016
rect 39672 42168 39724 42220
rect 41328 42168 41380 42220
rect 46296 42168 46348 42220
rect 29184 42100 29236 42152
rect 31300 42100 31352 42152
rect 35532 42100 35584 42152
rect 37832 42100 37884 42152
rect 40316 42100 40368 42152
rect 43904 42100 43956 42152
rect 48504 42143 48556 42152
rect 48504 42109 48513 42143
rect 48513 42109 48547 42143
rect 48547 42109 48556 42143
rect 48504 42100 48556 42109
rect 29092 42032 29144 42084
rect 28632 41964 28684 42016
rect 29184 41964 29236 42016
rect 29828 41964 29880 42016
rect 31392 42032 31444 42084
rect 32496 42032 32548 42084
rect 31668 41964 31720 42016
rect 31852 41964 31904 42016
rect 35624 42007 35676 42016
rect 35624 41973 35633 42007
rect 35633 41973 35667 42007
rect 35667 41973 35676 42007
rect 35624 41964 35676 41973
rect 43536 41964 43588 42016
rect 2950 41862 3002 41914
rect 3014 41862 3066 41914
rect 3078 41862 3130 41914
rect 3142 41862 3194 41914
rect 3206 41862 3258 41914
rect 12950 41862 13002 41914
rect 13014 41862 13066 41914
rect 13078 41862 13130 41914
rect 13142 41862 13194 41914
rect 13206 41862 13258 41914
rect 22950 41862 23002 41914
rect 23014 41862 23066 41914
rect 23078 41862 23130 41914
rect 23142 41862 23194 41914
rect 23206 41862 23258 41914
rect 32950 41862 33002 41914
rect 33014 41862 33066 41914
rect 33078 41862 33130 41914
rect 33142 41862 33194 41914
rect 33206 41862 33258 41914
rect 42950 41862 43002 41914
rect 43014 41862 43066 41914
rect 43078 41862 43130 41914
rect 43142 41862 43194 41914
rect 43206 41862 43258 41914
rect 26332 41760 26384 41812
rect 31668 41760 31720 41812
rect 33048 41760 33100 41812
rect 35532 41760 35584 41812
rect 36912 41760 36964 41812
rect 48688 41760 48740 41812
rect 31392 41692 31444 41744
rect 24124 41624 24176 41676
rect 26516 41624 26568 41676
rect 23756 41599 23808 41608
rect 23756 41565 23765 41599
rect 23765 41565 23799 41599
rect 23799 41565 23808 41599
rect 23756 41556 23808 41565
rect 26424 41556 26476 41608
rect 34152 41624 34204 41676
rect 34520 41624 34572 41676
rect 34704 41624 34756 41676
rect 37832 41624 37884 41676
rect 31300 41556 31352 41608
rect 33048 41556 33100 41608
rect 48412 41556 48464 41608
rect 1676 41531 1728 41540
rect 1676 41497 1685 41531
rect 1685 41497 1719 41531
rect 1719 41497 1728 41531
rect 1676 41488 1728 41497
rect 11980 41488 12032 41540
rect 22468 41488 22520 41540
rect 10600 41420 10652 41472
rect 22100 41420 22152 41472
rect 31208 41488 31260 41540
rect 35072 41488 35124 41540
rect 33324 41420 33376 41472
rect 34060 41420 34112 41472
rect 35808 41420 35860 41472
rect 36636 41488 36688 41540
rect 37004 41420 37056 41472
rect 39672 41488 39724 41540
rect 7950 41318 8002 41370
rect 8014 41318 8066 41370
rect 8078 41318 8130 41370
rect 8142 41318 8194 41370
rect 8206 41318 8258 41370
rect 17950 41318 18002 41370
rect 18014 41318 18066 41370
rect 18078 41318 18130 41370
rect 18142 41318 18194 41370
rect 18206 41318 18258 41370
rect 27950 41318 28002 41370
rect 28014 41318 28066 41370
rect 28078 41318 28130 41370
rect 28142 41318 28194 41370
rect 28206 41318 28258 41370
rect 37950 41318 38002 41370
rect 38014 41318 38066 41370
rect 38078 41318 38130 41370
rect 38142 41318 38194 41370
rect 38206 41318 38258 41370
rect 47950 41318 48002 41370
rect 48014 41318 48066 41370
rect 48078 41318 48130 41370
rect 48142 41318 48194 41370
rect 48206 41318 48258 41370
rect 5816 41259 5868 41268
rect 5816 41225 5825 41259
rect 5825 41225 5859 41259
rect 5859 41225 5868 41259
rect 5816 41216 5868 41225
rect 9864 41259 9916 41268
rect 9864 41225 9873 41259
rect 9873 41225 9907 41259
rect 9907 41225 9916 41259
rect 9864 41216 9916 41225
rect 10784 41259 10836 41268
rect 10784 41225 10793 41259
rect 10793 41225 10827 41259
rect 10827 41225 10836 41259
rect 10784 41216 10836 41225
rect 22100 41216 22152 41268
rect 22468 41216 22520 41268
rect 24860 41216 24912 41268
rect 22192 41148 22244 41200
rect 26056 41216 26108 41268
rect 27712 41216 27764 41268
rect 29552 41216 29604 41268
rect 31944 41216 31996 41268
rect 5724 41123 5776 41132
rect 5724 41089 5733 41123
rect 5733 41089 5767 41123
rect 5767 41089 5776 41123
rect 5724 41080 5776 41089
rect 9772 41123 9824 41132
rect 9772 41089 9781 41123
rect 9781 41089 9815 41123
rect 9815 41089 9824 41123
rect 9772 41080 9824 41089
rect 10692 41123 10744 41132
rect 10692 41089 10701 41123
rect 10701 41089 10735 41123
rect 10735 41089 10744 41123
rect 10692 41080 10744 41089
rect 1768 41012 1820 41064
rect 22376 41123 22428 41132
rect 22376 41089 22385 41123
rect 22385 41089 22419 41123
rect 22419 41089 22428 41123
rect 22376 41080 22428 41089
rect 27988 41148 28040 41200
rect 30840 41148 30892 41200
rect 32864 41148 32916 41200
rect 24124 41080 24176 41132
rect 24584 41080 24636 41132
rect 27252 41123 27304 41132
rect 27252 41089 27261 41123
rect 27261 41089 27295 41123
rect 27295 41089 27304 41123
rect 27252 41080 27304 41089
rect 32588 41080 32640 41132
rect 22744 41012 22796 41064
rect 25044 41055 25096 41064
rect 25044 41021 25053 41055
rect 25053 41021 25087 41055
rect 25087 41021 25096 41055
rect 25044 41012 25096 41021
rect 27528 41055 27580 41064
rect 27528 41021 27537 41055
rect 27537 41021 27571 41055
rect 27571 41021 27580 41055
rect 27528 41012 27580 41021
rect 27988 41012 28040 41064
rect 29092 41012 29144 41064
rect 29920 40944 29972 40996
rect 32312 41012 32364 41064
rect 22560 40876 22612 40928
rect 22836 40876 22888 40928
rect 29000 40919 29052 40928
rect 29000 40885 29009 40919
rect 29009 40885 29043 40919
rect 29043 40885 29052 40919
rect 29000 40876 29052 40885
rect 29828 40876 29880 40928
rect 33048 40876 33100 40928
rect 33600 40876 33652 40928
rect 37004 41148 37056 41200
rect 39856 41148 39908 41200
rect 37832 41080 37884 41132
rect 38936 41012 38988 41064
rect 39948 41012 40000 41064
rect 39488 40944 39540 40996
rect 48504 41055 48556 41064
rect 48504 41021 48513 41055
rect 48513 41021 48547 41055
rect 48547 41021 48556 41055
rect 48504 41012 48556 41021
rect 34796 40876 34848 40928
rect 35164 40876 35216 40928
rect 39212 40876 39264 40928
rect 39764 40876 39816 40928
rect 39948 40919 40000 40928
rect 39948 40885 39957 40919
rect 39957 40885 39991 40919
rect 39991 40885 40000 40919
rect 39948 40876 40000 40885
rect 2950 40774 3002 40826
rect 3014 40774 3066 40826
rect 3078 40774 3130 40826
rect 3142 40774 3194 40826
rect 3206 40774 3258 40826
rect 12950 40774 13002 40826
rect 13014 40774 13066 40826
rect 13078 40774 13130 40826
rect 13142 40774 13194 40826
rect 13206 40774 13258 40826
rect 22950 40774 23002 40826
rect 23014 40774 23066 40826
rect 23078 40774 23130 40826
rect 23142 40774 23194 40826
rect 23206 40774 23258 40826
rect 32950 40774 33002 40826
rect 33014 40774 33066 40826
rect 33078 40774 33130 40826
rect 33142 40774 33194 40826
rect 33206 40774 33258 40826
rect 42950 40774 43002 40826
rect 43014 40774 43066 40826
rect 43078 40774 43130 40826
rect 43142 40774 43194 40826
rect 43206 40774 43258 40826
rect 20536 40672 20588 40724
rect 22008 40604 22060 40656
rect 25044 40536 25096 40588
rect 29552 40672 29604 40724
rect 29000 40604 29052 40656
rect 27252 40579 27304 40588
rect 27252 40545 27261 40579
rect 27261 40545 27295 40579
rect 27295 40545 27304 40579
rect 27252 40536 27304 40545
rect 22744 40468 22796 40520
rect 24308 40468 24360 40520
rect 23388 40400 23440 40452
rect 27068 40511 27120 40520
rect 27068 40477 27077 40511
rect 27077 40477 27111 40511
rect 27111 40477 27120 40511
rect 27068 40468 27120 40477
rect 31024 40672 31076 40724
rect 35072 40672 35124 40724
rect 39580 40672 39632 40724
rect 31024 40536 31076 40588
rect 32680 40579 32732 40588
rect 32680 40545 32689 40579
rect 32689 40545 32723 40579
rect 32723 40545 32732 40579
rect 32680 40536 32732 40545
rect 32772 40579 32824 40588
rect 32772 40545 32781 40579
rect 32781 40545 32815 40579
rect 32815 40545 32824 40579
rect 32772 40536 32824 40545
rect 33508 40536 33560 40588
rect 34152 40579 34204 40588
rect 34152 40545 34161 40579
rect 34161 40545 34195 40579
rect 34195 40545 34204 40579
rect 34152 40536 34204 40545
rect 38752 40536 38804 40588
rect 39396 40579 39448 40588
rect 39396 40545 39405 40579
rect 39405 40545 39439 40579
rect 39439 40545 39448 40579
rect 39396 40536 39448 40545
rect 39948 40536 40000 40588
rect 48780 40579 48832 40588
rect 48780 40545 48789 40579
rect 48789 40545 48823 40579
rect 48823 40545 48832 40579
rect 48780 40536 48832 40545
rect 29736 40511 29788 40520
rect 29736 40477 29745 40511
rect 29745 40477 29779 40511
rect 29779 40477 29788 40511
rect 29736 40468 29788 40477
rect 31668 40400 31720 40452
rect 22100 40332 22152 40384
rect 26608 40332 26660 40384
rect 26700 40375 26752 40384
rect 26700 40341 26709 40375
rect 26709 40341 26743 40375
rect 26743 40341 26752 40375
rect 26700 40332 26752 40341
rect 27068 40332 27120 40384
rect 29920 40332 29972 40384
rect 33324 40400 33376 40452
rect 33968 40443 34020 40452
rect 33968 40409 33977 40443
rect 33977 40409 34011 40443
rect 34011 40409 34020 40443
rect 33968 40400 34020 40409
rect 33876 40332 33928 40384
rect 37740 40468 37792 40520
rect 38568 40468 38620 40520
rect 48504 40511 48556 40520
rect 48504 40477 48513 40511
rect 48513 40477 48547 40511
rect 48547 40477 48556 40511
rect 48504 40468 48556 40477
rect 39948 40400 40000 40452
rect 37372 40332 37424 40384
rect 39120 40375 39172 40384
rect 39120 40341 39129 40375
rect 39129 40341 39163 40375
rect 39163 40341 39172 40375
rect 39120 40332 39172 40341
rect 7950 40230 8002 40282
rect 8014 40230 8066 40282
rect 8078 40230 8130 40282
rect 8142 40230 8194 40282
rect 8206 40230 8258 40282
rect 17950 40230 18002 40282
rect 18014 40230 18066 40282
rect 18078 40230 18130 40282
rect 18142 40230 18194 40282
rect 18206 40230 18258 40282
rect 27950 40230 28002 40282
rect 28014 40230 28066 40282
rect 28078 40230 28130 40282
rect 28142 40230 28194 40282
rect 28206 40230 28258 40282
rect 37950 40230 38002 40282
rect 38014 40230 38066 40282
rect 38078 40230 38130 40282
rect 38142 40230 38194 40282
rect 38206 40230 38258 40282
rect 47950 40230 48002 40282
rect 48014 40230 48066 40282
rect 48078 40230 48130 40282
rect 48142 40230 48194 40282
rect 48206 40230 48258 40282
rect 25044 40171 25096 40180
rect 25044 40137 25053 40171
rect 25053 40137 25087 40171
rect 25087 40137 25096 40171
rect 25044 40128 25096 40137
rect 24860 40060 24912 40112
rect 31668 40128 31720 40180
rect 32772 40128 32824 40180
rect 35256 40128 35308 40180
rect 35624 40128 35676 40180
rect 35900 40128 35952 40180
rect 36820 40128 36872 40180
rect 39856 40128 39908 40180
rect 29736 40060 29788 40112
rect 33600 40060 33652 40112
rect 21088 39924 21140 39976
rect 23572 39967 23624 39976
rect 23572 39933 23581 39967
rect 23581 39933 23615 39967
rect 23615 39933 23624 39967
rect 23572 39924 23624 39933
rect 24676 39856 24728 39908
rect 27712 39856 27764 39908
rect 22468 39788 22520 39840
rect 26056 39788 26108 39840
rect 28908 39924 28960 39976
rect 31300 39992 31352 40044
rect 32312 40035 32364 40044
rect 32312 40001 32321 40035
rect 32321 40001 32355 40035
rect 32355 40001 32364 40035
rect 32312 39992 32364 40001
rect 34520 40060 34572 40112
rect 37004 40060 37056 40112
rect 34704 40035 34756 40044
rect 34704 40001 34713 40035
rect 34713 40001 34747 40035
rect 34747 40001 34756 40035
rect 34704 39992 34756 40001
rect 37832 39992 37884 40044
rect 38568 40035 38620 40044
rect 38568 40001 38577 40035
rect 38577 40001 38611 40035
rect 38611 40001 38620 40035
rect 38568 39992 38620 40001
rect 40316 40171 40368 40180
rect 40316 40137 40325 40171
rect 40325 40137 40359 40171
rect 40359 40137 40368 40171
rect 40316 40128 40368 40137
rect 42432 40128 42484 40180
rect 41144 40103 41196 40112
rect 41144 40069 41153 40103
rect 41153 40069 41187 40103
rect 41187 40069 41196 40103
rect 41144 40060 41196 40069
rect 29828 39856 29880 39908
rect 33784 39856 33836 39908
rect 36452 39924 36504 39976
rect 36728 39924 36780 39976
rect 39396 39924 39448 39976
rect 41236 40035 41288 40044
rect 41236 40001 41245 40035
rect 41245 40001 41279 40035
rect 41279 40001 41288 40035
rect 41236 39992 41288 40001
rect 41696 39924 41748 39976
rect 48504 39967 48556 39976
rect 48504 39933 48513 39967
rect 48513 39933 48547 39967
rect 48547 39933 48556 39967
rect 48504 39924 48556 39933
rect 48596 39924 48648 39976
rect 41880 39856 41932 39908
rect 30196 39788 30248 39840
rect 30288 39788 30340 39840
rect 31576 39788 31628 39840
rect 34796 39788 34848 39840
rect 40960 39788 41012 39840
rect 2950 39686 3002 39738
rect 3014 39686 3066 39738
rect 3078 39686 3130 39738
rect 3142 39686 3194 39738
rect 3206 39686 3258 39738
rect 12950 39686 13002 39738
rect 13014 39686 13066 39738
rect 13078 39686 13130 39738
rect 13142 39686 13194 39738
rect 13206 39686 13258 39738
rect 22950 39686 23002 39738
rect 23014 39686 23066 39738
rect 23078 39686 23130 39738
rect 23142 39686 23194 39738
rect 23206 39686 23258 39738
rect 32950 39686 33002 39738
rect 33014 39686 33066 39738
rect 33078 39686 33130 39738
rect 33142 39686 33194 39738
rect 33206 39686 33258 39738
rect 42950 39686 43002 39738
rect 43014 39686 43066 39738
rect 43078 39686 43130 39738
rect 43142 39686 43194 39738
rect 43206 39686 43258 39738
rect 25964 39584 26016 39636
rect 29184 39584 29236 39636
rect 29644 39584 29696 39636
rect 30288 39584 30340 39636
rect 31024 39584 31076 39636
rect 31484 39584 31536 39636
rect 26056 39516 26108 39568
rect 22468 39491 22520 39500
rect 1860 39244 1912 39296
rect 22468 39457 22477 39491
rect 22477 39457 22511 39491
rect 22511 39457 22520 39491
rect 22468 39448 22520 39457
rect 22192 39380 22244 39432
rect 24584 39491 24636 39500
rect 24584 39457 24593 39491
rect 24593 39457 24627 39491
rect 24627 39457 24636 39491
rect 24584 39448 24636 39457
rect 25228 39448 25280 39500
rect 28448 39448 28500 39500
rect 31576 39516 31628 39568
rect 31116 39448 31168 39500
rect 26148 39380 26200 39432
rect 28724 39380 28776 39432
rect 30104 39380 30156 39432
rect 31576 39380 31628 39432
rect 32588 39627 32640 39636
rect 32588 39593 32597 39627
rect 32597 39593 32631 39627
rect 32631 39593 32640 39627
rect 32588 39584 32640 39593
rect 34336 39584 34388 39636
rect 39212 39584 39264 39636
rect 39856 39584 39908 39636
rect 32220 39516 32272 39568
rect 35992 39516 36044 39568
rect 38476 39516 38528 39568
rect 38844 39516 38896 39568
rect 38292 39448 38344 39500
rect 42800 39448 42852 39500
rect 48964 39516 49016 39568
rect 34336 39380 34388 39432
rect 34704 39380 34756 39432
rect 38844 39380 38896 39432
rect 40868 39423 40920 39432
rect 40868 39389 40877 39423
rect 40877 39389 40911 39423
rect 40911 39389 40920 39423
rect 40868 39380 40920 39389
rect 24860 39312 24912 39364
rect 26976 39312 27028 39364
rect 22376 39287 22428 39296
rect 22376 39253 22385 39287
rect 22385 39253 22419 39287
rect 22419 39253 22428 39287
rect 22376 39244 22428 39253
rect 23572 39244 23624 39296
rect 28816 39244 28868 39296
rect 30748 39244 30800 39296
rect 33600 39244 33652 39296
rect 37004 39312 37056 39364
rect 37556 39312 37608 39364
rect 41420 39312 41472 39364
rect 42616 39312 42668 39364
rect 37648 39244 37700 39296
rect 37832 39244 37884 39296
rect 39672 39244 39724 39296
rect 48780 39491 48832 39500
rect 48780 39457 48789 39491
rect 48789 39457 48823 39491
rect 48823 39457 48832 39491
rect 48780 39448 48832 39457
rect 43996 39380 44048 39432
rect 46940 39380 46992 39432
rect 48504 39423 48556 39432
rect 48504 39389 48513 39423
rect 48513 39389 48547 39423
rect 48547 39389 48556 39423
rect 48504 39380 48556 39389
rect 7950 39142 8002 39194
rect 8014 39142 8066 39194
rect 8078 39142 8130 39194
rect 8142 39142 8194 39194
rect 8206 39142 8258 39194
rect 17950 39142 18002 39194
rect 18014 39142 18066 39194
rect 18078 39142 18130 39194
rect 18142 39142 18194 39194
rect 18206 39142 18258 39194
rect 27950 39142 28002 39194
rect 28014 39142 28066 39194
rect 28078 39142 28130 39194
rect 28142 39142 28194 39194
rect 28206 39142 28258 39194
rect 37950 39142 38002 39194
rect 38014 39142 38066 39194
rect 38078 39142 38130 39194
rect 38142 39142 38194 39194
rect 38206 39142 38258 39194
rect 47950 39142 48002 39194
rect 48014 39142 48066 39194
rect 48078 39142 48130 39194
rect 48142 39142 48194 39194
rect 48206 39142 48258 39194
rect 24492 39083 24544 39092
rect 24492 39049 24501 39083
rect 24501 39049 24535 39083
rect 24535 39049 24544 39083
rect 24492 39040 24544 39049
rect 24584 39040 24636 39092
rect 25044 39040 25096 39092
rect 25872 39083 25924 39092
rect 25872 39049 25881 39083
rect 25881 39049 25915 39083
rect 25915 39049 25924 39083
rect 25872 39040 25924 39049
rect 26976 39040 27028 39092
rect 27160 39040 27212 39092
rect 32220 39040 32272 39092
rect 32404 39083 32456 39092
rect 32404 39049 32413 39083
rect 32413 39049 32447 39083
rect 32447 39049 32456 39083
rect 32404 39040 32456 39049
rect 33600 39083 33652 39092
rect 33600 39049 33609 39083
rect 33609 39049 33643 39083
rect 33643 39049 33652 39083
rect 33600 39040 33652 39049
rect 34796 39083 34848 39092
rect 34796 39049 34805 39083
rect 34805 39049 34839 39083
rect 34839 39049 34848 39083
rect 34796 39040 34848 39049
rect 34888 39040 34940 39092
rect 36176 39040 36228 39092
rect 37280 39040 37332 39092
rect 38844 39083 38896 39092
rect 38844 39049 38853 39083
rect 38853 39049 38887 39083
rect 38887 39049 38896 39083
rect 38844 39040 38896 39049
rect 39120 39040 39172 39092
rect 40040 39040 40092 39092
rect 40776 39040 40828 39092
rect 41420 39040 41472 39092
rect 42064 39040 42116 39092
rect 22836 38972 22888 39024
rect 24676 38972 24728 39024
rect 24860 39015 24912 39024
rect 24860 38981 24869 39015
rect 24869 38981 24903 39015
rect 24903 38981 24912 39015
rect 24860 38972 24912 38981
rect 27068 38972 27120 39024
rect 29828 38972 29880 39024
rect 37556 38972 37608 39024
rect 38568 38972 38620 39024
rect 940 38904 992 38956
rect 1952 38904 2004 38956
rect 26148 38904 26200 38956
rect 26240 38947 26292 38956
rect 26240 38913 26249 38947
rect 26249 38913 26283 38947
rect 26283 38913 26292 38947
rect 26240 38904 26292 38913
rect 26792 38904 26844 38956
rect 28448 38904 28500 38956
rect 24584 38836 24636 38888
rect 24952 38836 25004 38888
rect 26516 38879 26568 38888
rect 26516 38845 26525 38879
rect 26525 38845 26559 38879
rect 26559 38845 26568 38879
rect 26516 38836 26568 38845
rect 27896 38879 27948 38888
rect 27896 38845 27905 38879
rect 27905 38845 27939 38879
rect 27939 38845 27948 38879
rect 27896 38836 27948 38845
rect 27988 38836 28040 38888
rect 32588 38904 32640 38956
rect 26056 38768 26108 38820
rect 26792 38768 26844 38820
rect 28724 38768 28776 38820
rect 31576 38768 31628 38820
rect 7380 38700 7432 38752
rect 26976 38700 27028 38752
rect 28540 38743 28592 38752
rect 28540 38709 28549 38743
rect 28549 38709 28583 38743
rect 28583 38709 28592 38743
rect 28540 38700 28592 38709
rect 31116 38700 31168 38752
rect 34336 38836 34388 38888
rect 35256 38836 35308 38888
rect 34980 38743 35032 38752
rect 34980 38709 34989 38743
rect 34989 38709 35023 38743
rect 35023 38709 35032 38743
rect 34980 38700 35032 38709
rect 36176 38743 36228 38752
rect 36176 38709 36185 38743
rect 36185 38709 36219 38743
rect 36219 38709 36228 38743
rect 36176 38700 36228 38709
rect 36912 38904 36964 38956
rect 37832 38947 37884 38956
rect 37832 38913 37841 38947
rect 37841 38913 37875 38947
rect 37875 38913 37884 38947
rect 37832 38904 37884 38913
rect 39672 38947 39724 38956
rect 39672 38913 39681 38947
rect 39681 38913 39715 38947
rect 39715 38913 39724 38947
rect 39672 38904 39724 38913
rect 40868 38972 40920 39024
rect 41880 38972 41932 39024
rect 42616 38972 42668 39024
rect 36452 38836 36504 38888
rect 37188 38836 37240 38888
rect 37924 38836 37976 38888
rect 38660 38836 38712 38888
rect 39396 38836 39448 38888
rect 39856 38879 39908 38888
rect 39856 38845 39865 38879
rect 39865 38845 39899 38879
rect 39899 38845 39908 38879
rect 39856 38836 39908 38845
rect 40592 38879 40644 38888
rect 40592 38845 40601 38879
rect 40601 38845 40635 38879
rect 40635 38845 40644 38879
rect 40592 38836 40644 38845
rect 40040 38768 40092 38820
rect 37464 38743 37516 38752
rect 37464 38709 37473 38743
rect 37473 38709 37507 38743
rect 37507 38709 37516 38743
rect 37464 38700 37516 38709
rect 41236 38700 41288 38752
rect 41696 38700 41748 38752
rect 2950 38598 3002 38650
rect 3014 38598 3066 38650
rect 3078 38598 3130 38650
rect 3142 38598 3194 38650
rect 3206 38598 3258 38650
rect 12950 38598 13002 38650
rect 13014 38598 13066 38650
rect 13078 38598 13130 38650
rect 13142 38598 13194 38650
rect 13206 38598 13258 38650
rect 22950 38598 23002 38650
rect 23014 38598 23066 38650
rect 23078 38598 23130 38650
rect 23142 38598 23194 38650
rect 23206 38598 23258 38650
rect 32950 38598 33002 38650
rect 33014 38598 33066 38650
rect 33078 38598 33130 38650
rect 33142 38598 33194 38650
rect 33206 38598 33258 38650
rect 42950 38598 43002 38650
rect 43014 38598 43066 38650
rect 43078 38598 43130 38650
rect 43142 38598 43194 38650
rect 43206 38598 43258 38650
rect 23296 38539 23348 38548
rect 23296 38505 23305 38539
rect 23305 38505 23339 38539
rect 23339 38505 23348 38539
rect 23296 38496 23348 38505
rect 27068 38539 27120 38548
rect 27068 38505 27077 38539
rect 27077 38505 27111 38539
rect 27111 38505 27120 38539
rect 27068 38496 27120 38505
rect 36268 38496 36320 38548
rect 36636 38539 36688 38548
rect 36636 38505 36645 38539
rect 36645 38505 36679 38539
rect 36679 38505 36688 38539
rect 36636 38496 36688 38505
rect 41144 38496 41196 38548
rect 42800 38496 42852 38548
rect 43352 38496 43404 38548
rect 25228 38428 25280 38480
rect 26608 38428 26660 38480
rect 28816 38428 28868 38480
rect 21088 38403 21140 38412
rect 21088 38369 21097 38403
rect 21097 38369 21131 38403
rect 21131 38369 21140 38403
rect 21088 38360 21140 38369
rect 23848 38403 23900 38412
rect 23848 38369 23857 38403
rect 23857 38369 23891 38403
rect 23891 38369 23900 38403
rect 23848 38360 23900 38369
rect 27068 38360 27120 38412
rect 28540 38360 28592 38412
rect 31852 38428 31904 38480
rect 27160 38292 27212 38344
rect 30104 38360 30156 38412
rect 31668 38292 31720 38344
rect 33324 38403 33376 38412
rect 33324 38369 33333 38403
rect 33333 38369 33367 38403
rect 33367 38369 33376 38403
rect 33324 38360 33376 38369
rect 34520 38428 34572 38480
rect 34704 38360 34756 38412
rect 35256 38360 35308 38412
rect 37372 38360 37424 38412
rect 40408 38360 40460 38412
rect 40592 38403 40644 38412
rect 40592 38369 40601 38403
rect 40601 38369 40635 38403
rect 40635 38369 40644 38403
rect 40592 38360 40644 38369
rect 43168 38360 43220 38412
rect 36912 38292 36964 38344
rect 37556 38292 37608 38344
rect 41052 38292 41104 38344
rect 41512 38335 41564 38344
rect 41512 38301 41521 38335
rect 41521 38301 41555 38335
rect 41555 38301 41564 38335
rect 41512 38292 41564 38301
rect 42800 38292 42852 38344
rect 43996 38292 44048 38344
rect 49332 38335 49384 38344
rect 49332 38301 49341 38335
rect 49341 38301 49375 38335
rect 49375 38301 49384 38335
rect 49332 38292 49384 38301
rect 21364 38267 21416 38276
rect 21364 38233 21373 38267
rect 21373 38233 21407 38267
rect 21407 38233 21416 38267
rect 21364 38224 21416 38233
rect 24676 38224 24728 38276
rect 23664 38199 23716 38208
rect 23664 38165 23673 38199
rect 23673 38165 23707 38199
rect 23707 38165 23716 38199
rect 23664 38156 23716 38165
rect 25504 38156 25556 38208
rect 26976 38156 27028 38208
rect 28816 38199 28868 38208
rect 28816 38165 28825 38199
rect 28825 38165 28859 38199
rect 28859 38165 28868 38199
rect 28816 38156 28868 38165
rect 29920 38224 29972 38276
rect 30472 38224 30524 38276
rect 31576 38224 31628 38276
rect 32220 38224 32272 38276
rect 33232 38199 33284 38208
rect 33232 38165 33241 38199
rect 33241 38165 33275 38199
rect 33275 38165 33284 38199
rect 33232 38156 33284 38165
rect 35440 38224 35492 38276
rect 36452 38224 36504 38276
rect 37004 38224 37056 38276
rect 37096 38267 37148 38276
rect 37096 38233 37105 38267
rect 37105 38233 37139 38267
rect 37139 38233 37148 38267
rect 37096 38224 37148 38233
rect 38660 38224 38712 38276
rect 37280 38156 37332 38208
rect 38568 38156 38620 38208
rect 40408 38199 40460 38208
rect 40408 38165 40417 38199
rect 40417 38165 40451 38199
rect 40451 38165 40460 38199
rect 40408 38156 40460 38165
rect 40684 38156 40736 38208
rect 41696 38224 41748 38276
rect 43260 38224 43312 38276
rect 46204 38224 46256 38276
rect 43720 38156 43772 38208
rect 49148 38199 49200 38208
rect 49148 38165 49157 38199
rect 49157 38165 49191 38199
rect 49191 38165 49200 38199
rect 49148 38156 49200 38165
rect 7950 38054 8002 38106
rect 8014 38054 8066 38106
rect 8078 38054 8130 38106
rect 8142 38054 8194 38106
rect 8206 38054 8258 38106
rect 17950 38054 18002 38106
rect 18014 38054 18066 38106
rect 18078 38054 18130 38106
rect 18142 38054 18194 38106
rect 18206 38054 18258 38106
rect 27950 38054 28002 38106
rect 28014 38054 28066 38106
rect 28078 38054 28130 38106
rect 28142 38054 28194 38106
rect 28206 38054 28258 38106
rect 37950 38054 38002 38106
rect 38014 38054 38066 38106
rect 38078 38054 38130 38106
rect 38142 38054 38194 38106
rect 38206 38054 38258 38106
rect 47950 38054 48002 38106
rect 48014 38054 48066 38106
rect 48078 38054 48130 38106
rect 48142 38054 48194 38106
rect 48206 38054 48258 38106
rect 27160 37952 27212 38004
rect 27528 37952 27580 38004
rect 32864 37952 32916 38004
rect 33876 37952 33928 38004
rect 35348 37952 35400 38004
rect 37188 37952 37240 38004
rect 37832 37952 37884 38004
rect 39580 37952 39632 38004
rect 24676 37884 24728 37936
rect 28172 37884 28224 37936
rect 31300 37927 31352 37936
rect 31300 37893 31309 37927
rect 31309 37893 31343 37927
rect 31343 37893 31352 37927
rect 31300 37884 31352 37893
rect 31668 37884 31720 37936
rect 37096 37884 37148 37936
rect 41236 37995 41288 38004
rect 41236 37961 41245 37995
rect 41245 37961 41279 37995
rect 41279 37961 41288 37995
rect 41236 37952 41288 37961
rect 42800 37952 42852 38004
rect 43444 37952 43496 38004
rect 43720 37952 43772 38004
rect 48596 37952 48648 38004
rect 27160 37859 27212 37868
rect 27160 37825 27169 37859
rect 27169 37825 27203 37859
rect 27203 37825 27212 37859
rect 27160 37816 27212 37825
rect 30380 37816 30432 37868
rect 33508 37816 33560 37868
rect 26332 37748 26384 37800
rect 27068 37748 27120 37800
rect 27804 37748 27856 37800
rect 22468 37612 22520 37664
rect 24952 37612 25004 37664
rect 25044 37612 25096 37664
rect 29460 37748 29512 37800
rect 28908 37680 28960 37732
rect 32956 37791 33008 37800
rect 32956 37757 32965 37791
rect 32965 37757 32999 37791
rect 32999 37757 33008 37791
rect 32956 37748 33008 37757
rect 29736 37680 29788 37732
rect 34704 37816 34756 37868
rect 37832 37859 37884 37868
rect 37832 37825 37841 37859
rect 37841 37825 37875 37859
rect 37875 37825 37884 37859
rect 37832 37816 37884 37825
rect 40408 37816 40460 37868
rect 40684 37816 40736 37868
rect 43260 37884 43312 37936
rect 42248 37816 42300 37868
rect 34060 37791 34112 37800
rect 34060 37757 34069 37791
rect 34069 37757 34103 37791
rect 34103 37757 34112 37791
rect 34060 37748 34112 37757
rect 37924 37791 37976 37800
rect 37924 37757 37933 37791
rect 37933 37757 37967 37791
rect 37967 37757 37976 37791
rect 37924 37748 37976 37757
rect 38292 37748 38344 37800
rect 38660 37791 38712 37800
rect 38660 37757 38669 37791
rect 38669 37757 38703 37791
rect 38703 37757 38712 37791
rect 38660 37748 38712 37757
rect 40132 37748 40184 37800
rect 40316 37748 40368 37800
rect 43168 37791 43220 37800
rect 43168 37757 43177 37791
rect 43177 37757 43211 37791
rect 43211 37757 43220 37791
rect 43168 37748 43220 37757
rect 31300 37612 31352 37664
rect 31392 37612 31444 37664
rect 32496 37612 32548 37664
rect 32680 37612 32732 37664
rect 32956 37612 33008 37664
rect 34336 37612 34388 37664
rect 40316 37612 40368 37664
rect 43812 37680 43864 37732
rect 49332 37859 49384 37868
rect 49332 37825 49341 37859
rect 49341 37825 49375 37859
rect 49375 37825 49384 37859
rect 49332 37816 49384 37825
rect 40960 37612 41012 37664
rect 41420 37612 41472 37664
rect 2950 37510 3002 37562
rect 3014 37510 3066 37562
rect 3078 37510 3130 37562
rect 3142 37510 3194 37562
rect 3206 37510 3258 37562
rect 12950 37510 13002 37562
rect 13014 37510 13066 37562
rect 13078 37510 13130 37562
rect 13142 37510 13194 37562
rect 13206 37510 13258 37562
rect 22950 37510 23002 37562
rect 23014 37510 23066 37562
rect 23078 37510 23130 37562
rect 23142 37510 23194 37562
rect 23206 37510 23258 37562
rect 32950 37510 33002 37562
rect 33014 37510 33066 37562
rect 33078 37510 33130 37562
rect 33142 37510 33194 37562
rect 33206 37510 33258 37562
rect 42950 37510 43002 37562
rect 43014 37510 43066 37562
rect 43078 37510 43130 37562
rect 43142 37510 43194 37562
rect 43206 37510 43258 37562
rect 22100 37451 22152 37460
rect 22100 37417 22109 37451
rect 22109 37417 22143 37451
rect 22143 37417 22152 37451
rect 22100 37408 22152 37417
rect 25504 37451 25556 37460
rect 25504 37417 25513 37451
rect 25513 37417 25547 37451
rect 25547 37417 25556 37451
rect 25504 37408 25556 37417
rect 27528 37408 27580 37460
rect 27804 37408 27856 37460
rect 28816 37408 28868 37460
rect 34152 37408 34204 37460
rect 14464 37136 14516 37188
rect 23572 37272 23624 37324
rect 23756 37315 23808 37324
rect 23756 37281 23765 37315
rect 23765 37281 23799 37315
rect 23799 37281 23808 37315
rect 23756 37272 23808 37281
rect 29736 37383 29788 37392
rect 29736 37349 29745 37383
rect 29745 37349 29779 37383
rect 29779 37349 29788 37383
rect 29736 37340 29788 37349
rect 30196 37340 30248 37392
rect 23940 37272 23992 37324
rect 27160 37272 27212 37324
rect 27620 37272 27672 37324
rect 29092 37272 29144 37324
rect 31208 37272 31260 37324
rect 31484 37315 31536 37324
rect 31484 37281 31493 37315
rect 31493 37281 31527 37315
rect 31527 37281 31536 37315
rect 31484 37272 31536 37281
rect 32864 37272 32916 37324
rect 22468 37247 22520 37256
rect 22468 37213 22477 37247
rect 22477 37213 22511 37247
rect 22511 37213 22520 37247
rect 22468 37204 22520 37213
rect 14924 37068 14976 37120
rect 23388 37068 23440 37120
rect 28172 37204 28224 37256
rect 31300 37247 31352 37256
rect 31300 37213 31309 37247
rect 31309 37213 31343 37247
rect 31343 37213 31352 37247
rect 31300 37204 31352 37213
rect 32036 37204 32088 37256
rect 25596 37068 25648 37120
rect 25872 37111 25924 37120
rect 25872 37077 25881 37111
rect 25881 37077 25915 37111
rect 25915 37077 25924 37111
rect 25872 37068 25924 37077
rect 25964 37111 26016 37120
rect 25964 37077 25973 37111
rect 25973 37077 26007 37111
rect 26007 37077 26016 37111
rect 25964 37068 26016 37077
rect 27068 37179 27120 37188
rect 27068 37145 27077 37179
rect 27077 37145 27111 37179
rect 27111 37145 27120 37179
rect 27068 37136 27120 37145
rect 29276 37136 29328 37188
rect 31944 37136 31996 37188
rect 30840 37068 30892 37120
rect 31484 37068 31536 37120
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 33508 37136 33560 37188
rect 49148 37408 49200 37460
rect 38660 37340 38712 37392
rect 40132 37272 40184 37324
rect 40316 37272 40368 37324
rect 40684 37272 40736 37324
rect 41512 37272 41564 37324
rect 42524 37272 42576 37324
rect 48504 37315 48556 37324
rect 48504 37281 48513 37315
rect 48513 37281 48547 37315
rect 48547 37281 48556 37315
rect 48504 37272 48556 37281
rect 37004 37204 37056 37256
rect 37832 37204 37884 37256
rect 38476 37204 38528 37256
rect 40224 37204 40276 37256
rect 48780 37247 48832 37256
rect 48780 37213 48789 37247
rect 48789 37213 48823 37247
rect 48823 37213 48832 37247
rect 48780 37204 48832 37213
rect 34520 37068 34572 37120
rect 35440 37068 35492 37120
rect 35716 37068 35768 37120
rect 36452 37068 36504 37120
rect 39120 37068 39172 37120
rect 39488 37068 39540 37120
rect 43996 37136 44048 37188
rect 43444 37068 43496 37120
rect 43720 37068 43772 37120
rect 7950 36966 8002 37018
rect 8014 36966 8066 37018
rect 8078 36966 8130 37018
rect 8142 36966 8194 37018
rect 8206 36966 8258 37018
rect 17950 36966 18002 37018
rect 18014 36966 18066 37018
rect 18078 36966 18130 37018
rect 18142 36966 18194 37018
rect 18206 36966 18258 37018
rect 27950 36966 28002 37018
rect 28014 36966 28066 37018
rect 28078 36966 28130 37018
rect 28142 36966 28194 37018
rect 28206 36966 28258 37018
rect 37950 36966 38002 37018
rect 38014 36966 38066 37018
rect 38078 36966 38130 37018
rect 38142 36966 38194 37018
rect 38206 36966 38258 37018
rect 47950 36966 48002 37018
rect 48014 36966 48066 37018
rect 48078 36966 48130 37018
rect 48142 36966 48194 37018
rect 48206 36966 48258 37018
rect 19432 36907 19484 36916
rect 19432 36873 19441 36907
rect 19441 36873 19475 36907
rect 19475 36873 19484 36907
rect 19432 36864 19484 36873
rect 23756 36864 23808 36916
rect 29828 36864 29880 36916
rect 32404 36864 32456 36916
rect 24676 36796 24728 36848
rect 940 36728 992 36780
rect 17224 36728 17276 36780
rect 21824 36728 21876 36780
rect 21364 36660 21416 36712
rect 22560 36660 22612 36712
rect 24952 36660 25004 36712
rect 25780 36660 25832 36712
rect 26424 36703 26476 36712
rect 26424 36669 26433 36703
rect 26433 36669 26467 36703
rect 26467 36669 26476 36703
rect 26424 36660 26476 36669
rect 27344 36728 27396 36780
rect 27436 36660 27488 36712
rect 27804 36728 27856 36780
rect 34244 36796 34296 36848
rect 29000 36728 29052 36780
rect 31392 36728 31444 36780
rect 31760 36771 31812 36780
rect 31760 36737 31769 36771
rect 31769 36737 31803 36771
rect 31803 36737 31812 36771
rect 31760 36728 31812 36737
rect 37740 36864 37792 36916
rect 40592 36864 40644 36916
rect 42432 36864 42484 36916
rect 39028 36796 39080 36848
rect 39580 36796 39632 36848
rect 40408 36796 40460 36848
rect 42340 36796 42392 36848
rect 48780 36796 48832 36848
rect 35716 36728 35768 36780
rect 41236 36728 41288 36780
rect 30840 36660 30892 36712
rect 32128 36592 32180 36644
rect 33968 36660 34020 36712
rect 35256 36660 35308 36712
rect 7564 36524 7616 36576
rect 22836 36524 22888 36576
rect 25504 36524 25556 36576
rect 29644 36524 29696 36576
rect 29920 36567 29972 36576
rect 29920 36533 29929 36567
rect 29929 36533 29963 36567
rect 29963 36533 29972 36567
rect 29920 36524 29972 36533
rect 34060 36524 34112 36576
rect 38476 36660 38528 36712
rect 38660 36660 38712 36712
rect 39948 36703 40000 36712
rect 39948 36669 39957 36703
rect 39957 36669 39991 36703
rect 39991 36669 40000 36703
rect 39948 36660 40000 36669
rect 40960 36660 41012 36712
rect 43720 36728 43772 36780
rect 49332 36771 49384 36780
rect 49332 36737 49341 36771
rect 49341 36737 49375 36771
rect 49375 36737 49384 36771
rect 49332 36728 49384 36737
rect 43352 36660 43404 36712
rect 35808 36592 35860 36644
rect 36084 36567 36136 36576
rect 36084 36533 36093 36567
rect 36093 36533 36127 36567
rect 36127 36533 36136 36567
rect 36084 36524 36136 36533
rect 36544 36524 36596 36576
rect 36912 36524 36964 36576
rect 40408 36524 40460 36576
rect 40592 36524 40644 36576
rect 44088 36524 44140 36576
rect 49148 36567 49200 36576
rect 49148 36533 49157 36567
rect 49157 36533 49191 36567
rect 49191 36533 49200 36567
rect 49148 36524 49200 36533
rect 2950 36422 3002 36474
rect 3014 36422 3066 36474
rect 3078 36422 3130 36474
rect 3142 36422 3194 36474
rect 3206 36422 3258 36474
rect 12950 36422 13002 36474
rect 13014 36422 13066 36474
rect 13078 36422 13130 36474
rect 13142 36422 13194 36474
rect 13206 36422 13258 36474
rect 22950 36422 23002 36474
rect 23014 36422 23066 36474
rect 23078 36422 23130 36474
rect 23142 36422 23194 36474
rect 23206 36422 23258 36474
rect 32950 36422 33002 36474
rect 33014 36422 33066 36474
rect 33078 36422 33130 36474
rect 33142 36422 33194 36474
rect 33206 36422 33258 36474
rect 42950 36422 43002 36474
rect 43014 36422 43066 36474
rect 43078 36422 43130 36474
rect 43142 36422 43194 36474
rect 43206 36422 43258 36474
rect 21916 36363 21968 36372
rect 21916 36329 21925 36363
rect 21925 36329 21959 36363
rect 21959 36329 21968 36363
rect 21916 36320 21968 36329
rect 26240 36320 26292 36372
rect 27344 36363 27396 36372
rect 27344 36329 27353 36363
rect 27353 36329 27387 36363
rect 27387 36329 27396 36363
rect 27344 36320 27396 36329
rect 27436 36320 27488 36372
rect 32128 36320 32180 36372
rect 33876 36320 33928 36372
rect 34428 36320 34480 36372
rect 36360 36320 36412 36372
rect 37280 36320 37332 36372
rect 41236 36320 41288 36372
rect 25872 36252 25924 36304
rect 22652 36184 22704 36236
rect 22744 36184 22796 36236
rect 28632 36184 28684 36236
rect 22836 36159 22888 36168
rect 22836 36125 22845 36159
rect 22845 36125 22879 36159
rect 22879 36125 22888 36159
rect 22836 36116 22888 36125
rect 28172 36159 28224 36168
rect 28172 36125 28181 36159
rect 28181 36125 28215 36159
rect 28215 36125 28224 36159
rect 28172 36116 28224 36125
rect 28724 36116 28776 36168
rect 31760 36116 31812 36168
rect 32680 36227 32732 36236
rect 32680 36193 32689 36227
rect 32689 36193 32723 36227
rect 32723 36193 32732 36227
rect 32680 36184 32732 36193
rect 34612 36184 34664 36236
rect 34980 36184 35032 36236
rect 35072 36116 35124 36168
rect 35164 36116 35216 36168
rect 40592 36252 40644 36304
rect 49148 36252 49200 36304
rect 36452 36184 36504 36236
rect 36820 36227 36872 36236
rect 36820 36193 36829 36227
rect 36829 36193 36863 36227
rect 36863 36193 36872 36227
rect 36820 36184 36872 36193
rect 38016 36227 38068 36236
rect 38016 36193 38025 36227
rect 38025 36193 38059 36227
rect 38059 36193 38068 36227
rect 38016 36184 38068 36193
rect 38108 36184 38160 36236
rect 40500 36184 40552 36236
rect 41696 36184 41748 36236
rect 41788 36227 41840 36236
rect 41788 36193 41797 36227
rect 41797 36193 41831 36227
rect 41831 36193 41840 36227
rect 41788 36184 41840 36193
rect 41880 36227 41932 36236
rect 41880 36193 41889 36227
rect 41889 36193 41923 36227
rect 41923 36193 41932 36227
rect 41880 36184 41932 36193
rect 43352 36184 43404 36236
rect 41604 36116 41656 36168
rect 21732 36048 21784 36100
rect 29920 36048 29972 36100
rect 33140 36048 33192 36100
rect 35624 36048 35676 36100
rect 35808 36048 35860 36100
rect 36360 36048 36412 36100
rect 40224 36048 40276 36100
rect 40684 36048 40736 36100
rect 42800 36116 42852 36168
rect 43536 36116 43588 36168
rect 22652 35980 22704 36032
rect 26240 35980 26292 36032
rect 34520 35980 34572 36032
rect 36820 35980 36872 36032
rect 38108 35980 38160 36032
rect 38752 35980 38804 36032
rect 41328 36023 41380 36032
rect 41328 35989 41337 36023
rect 41337 35989 41371 36023
rect 41371 35989 41380 36023
rect 41328 35980 41380 35989
rect 42800 35980 42852 36032
rect 42892 36023 42944 36032
rect 42892 35989 42901 36023
rect 42901 35989 42935 36023
rect 42935 35989 42944 36023
rect 42892 35980 42944 35989
rect 43260 35980 43312 36032
rect 43904 35980 43956 36032
rect 7950 35878 8002 35930
rect 8014 35878 8066 35930
rect 8078 35878 8130 35930
rect 8142 35878 8194 35930
rect 8206 35878 8258 35930
rect 17950 35878 18002 35930
rect 18014 35878 18066 35930
rect 18078 35878 18130 35930
rect 18142 35878 18194 35930
rect 18206 35878 18258 35930
rect 27950 35878 28002 35930
rect 28014 35878 28066 35930
rect 28078 35878 28130 35930
rect 28142 35878 28194 35930
rect 28206 35878 28258 35930
rect 37950 35878 38002 35930
rect 38014 35878 38066 35930
rect 38078 35878 38130 35930
rect 38142 35878 38194 35930
rect 38206 35878 38258 35930
rect 47950 35878 48002 35930
rect 48014 35878 48066 35930
rect 48078 35878 48130 35930
rect 48142 35878 48194 35930
rect 48206 35878 48258 35930
rect 21088 35776 21140 35828
rect 21364 35776 21416 35828
rect 23296 35640 23348 35692
rect 23848 35776 23900 35828
rect 27160 35776 27212 35828
rect 30840 35819 30892 35828
rect 25044 35708 25096 35760
rect 27068 35708 27120 35760
rect 30840 35785 30849 35819
rect 30849 35785 30883 35819
rect 30883 35785 30892 35819
rect 30840 35776 30892 35785
rect 33140 35776 33192 35828
rect 35072 35776 35124 35828
rect 39304 35776 39356 35828
rect 39948 35819 40000 35828
rect 39948 35785 39957 35819
rect 39957 35785 39991 35819
rect 39991 35785 40000 35819
rect 39948 35776 40000 35785
rect 33968 35708 34020 35760
rect 17868 35572 17920 35624
rect 21088 35572 21140 35624
rect 22008 35615 22060 35624
rect 22008 35581 22017 35615
rect 22017 35581 22051 35615
rect 22051 35581 22060 35615
rect 22008 35572 22060 35581
rect 23940 35572 23992 35624
rect 26332 35572 26384 35624
rect 27160 35640 27212 35692
rect 30472 35640 30524 35692
rect 34520 35640 34572 35692
rect 38568 35708 38620 35760
rect 27620 35572 27672 35624
rect 29460 35572 29512 35624
rect 31576 35572 31628 35624
rect 32772 35615 32824 35624
rect 32772 35581 32781 35615
rect 32781 35581 32815 35615
rect 32815 35581 32824 35615
rect 32772 35572 32824 35581
rect 32864 35615 32916 35624
rect 32864 35581 32873 35615
rect 32873 35581 32907 35615
rect 32907 35581 32916 35615
rect 32864 35572 32916 35581
rect 35808 35572 35860 35624
rect 24676 35504 24728 35556
rect 35900 35504 35952 35556
rect 36176 35615 36228 35624
rect 36176 35581 36185 35615
rect 36185 35581 36219 35615
rect 36219 35581 36228 35615
rect 36176 35572 36228 35581
rect 39580 35640 39632 35692
rect 39120 35572 39172 35624
rect 49056 35776 49108 35828
rect 40776 35751 40828 35760
rect 40776 35717 40785 35751
rect 40785 35717 40819 35751
rect 40819 35717 40828 35751
rect 40776 35708 40828 35717
rect 40684 35640 40736 35692
rect 40960 35615 41012 35624
rect 40960 35581 40969 35615
rect 40969 35581 41003 35615
rect 41003 35581 41012 35615
rect 43168 35708 43220 35760
rect 42524 35640 42576 35692
rect 43996 35640 44048 35692
rect 49332 35683 49384 35692
rect 49332 35649 49341 35683
rect 49341 35649 49375 35683
rect 49375 35649 49384 35683
rect 49332 35640 49384 35649
rect 40960 35572 41012 35581
rect 41972 35572 42024 35624
rect 38200 35504 38252 35556
rect 23388 35436 23440 35488
rect 26516 35436 26568 35488
rect 27712 35436 27764 35488
rect 30104 35436 30156 35488
rect 30472 35436 30524 35488
rect 33600 35436 33652 35488
rect 37280 35436 37332 35488
rect 40316 35436 40368 35488
rect 42892 35436 42944 35488
rect 43352 35436 43404 35488
rect 2950 35334 3002 35386
rect 3014 35334 3066 35386
rect 3078 35334 3130 35386
rect 3142 35334 3194 35386
rect 3206 35334 3258 35386
rect 12950 35334 13002 35386
rect 13014 35334 13066 35386
rect 13078 35334 13130 35386
rect 13142 35334 13194 35386
rect 13206 35334 13258 35386
rect 22950 35334 23002 35386
rect 23014 35334 23066 35386
rect 23078 35334 23130 35386
rect 23142 35334 23194 35386
rect 23206 35334 23258 35386
rect 32950 35334 33002 35386
rect 33014 35334 33066 35386
rect 33078 35334 33130 35386
rect 33142 35334 33194 35386
rect 33206 35334 33258 35386
rect 42950 35334 43002 35386
rect 43014 35334 43066 35386
rect 43078 35334 43130 35386
rect 43142 35334 43194 35386
rect 43206 35334 43258 35386
rect 21824 35232 21876 35284
rect 26056 35275 26108 35284
rect 26056 35241 26065 35275
rect 26065 35241 26099 35275
rect 26099 35241 26108 35275
rect 26056 35232 26108 35241
rect 26608 35232 26660 35284
rect 27252 35232 27304 35284
rect 30472 35232 30524 35284
rect 23940 35164 23992 35216
rect 24216 35164 24268 35216
rect 29460 35164 29512 35216
rect 33876 35232 33928 35284
rect 38016 35232 38068 35284
rect 22008 35096 22060 35148
rect 22560 35096 22612 35148
rect 23388 35096 23440 35148
rect 27068 35096 27120 35148
rect 27160 35096 27212 35148
rect 29920 35096 29972 35148
rect 30564 35096 30616 35148
rect 31116 35096 31168 35148
rect 31668 35139 31720 35148
rect 31668 35105 31677 35139
rect 31677 35105 31711 35139
rect 31711 35105 31720 35139
rect 31668 35096 31720 35105
rect 32220 35139 32272 35148
rect 32220 35105 32229 35139
rect 32229 35105 32263 35139
rect 32263 35105 32272 35139
rect 32220 35096 32272 35105
rect 36084 35096 36136 35148
rect 36636 35139 36688 35148
rect 36636 35105 36645 35139
rect 36645 35105 36679 35139
rect 36679 35105 36688 35139
rect 36636 35096 36688 35105
rect 26240 35028 26292 35080
rect 26516 35028 26568 35080
rect 33600 35028 33652 35080
rect 35716 35028 35768 35080
rect 37464 35028 37516 35080
rect 22100 34960 22152 35012
rect 23296 34960 23348 35012
rect 24584 34892 24636 34944
rect 28448 34892 28500 34944
rect 28540 34892 28592 34944
rect 29828 34892 29880 34944
rect 30196 34892 30248 34944
rect 34244 34960 34296 35012
rect 41420 35164 41472 35216
rect 37832 35139 37884 35148
rect 37832 35105 37841 35139
rect 37841 35105 37875 35139
rect 37875 35105 37884 35139
rect 37832 35096 37884 35105
rect 37924 35139 37976 35148
rect 37924 35105 37933 35139
rect 37933 35105 37967 35139
rect 37967 35105 37976 35139
rect 37924 35096 37976 35105
rect 39212 35139 39264 35148
rect 39212 35105 39221 35139
rect 39221 35105 39255 35139
rect 39255 35105 39264 35139
rect 39212 35096 39264 35105
rect 42524 35096 42576 35148
rect 43352 35096 43404 35148
rect 43536 35096 43588 35148
rect 39580 35028 39632 35080
rect 40224 35028 40276 35080
rect 40684 35028 40736 35080
rect 35900 34892 35952 34944
rect 35992 34935 36044 34944
rect 35992 34901 36001 34935
rect 36001 34901 36035 34935
rect 36035 34901 36044 34935
rect 35992 34892 36044 34901
rect 36360 34935 36412 34944
rect 36360 34901 36369 34935
rect 36369 34901 36403 34935
rect 36403 34901 36412 34935
rect 36360 34892 36412 34901
rect 38660 34960 38712 35012
rect 39212 34960 39264 35012
rect 40132 34960 40184 35012
rect 37648 34892 37700 34944
rect 40592 34892 40644 34944
rect 41420 34935 41472 34944
rect 41420 34901 41429 34935
rect 41429 34901 41463 34935
rect 41463 34901 41472 34935
rect 41420 34892 41472 34901
rect 41788 34935 41840 34944
rect 41788 34901 41797 34935
rect 41797 34901 41831 34935
rect 41831 34901 41840 34935
rect 41788 34892 41840 34901
rect 49332 35071 49384 35080
rect 49332 35037 49341 35071
rect 49341 35037 49375 35071
rect 49375 35037 49384 35071
rect 49332 35028 49384 35037
rect 43996 34960 44048 35012
rect 43628 34892 43680 34944
rect 49148 34935 49200 34944
rect 49148 34901 49157 34935
rect 49157 34901 49191 34935
rect 49191 34901 49200 34935
rect 49148 34892 49200 34901
rect 7950 34790 8002 34842
rect 8014 34790 8066 34842
rect 8078 34790 8130 34842
rect 8142 34790 8194 34842
rect 8206 34790 8258 34842
rect 17950 34790 18002 34842
rect 18014 34790 18066 34842
rect 18078 34790 18130 34842
rect 18142 34790 18194 34842
rect 18206 34790 18258 34842
rect 27950 34790 28002 34842
rect 28014 34790 28066 34842
rect 28078 34790 28130 34842
rect 28142 34790 28194 34842
rect 28206 34790 28258 34842
rect 37950 34790 38002 34842
rect 38014 34790 38066 34842
rect 38078 34790 38130 34842
rect 38142 34790 38194 34842
rect 38206 34790 38258 34842
rect 47950 34790 48002 34842
rect 48014 34790 48066 34842
rect 48078 34790 48130 34842
rect 48142 34790 48194 34842
rect 48206 34790 48258 34842
rect 7840 34688 7892 34740
rect 19984 34688 20036 34740
rect 22192 34688 22244 34740
rect 24676 34620 24728 34672
rect 24860 34688 24912 34740
rect 28724 34688 28776 34740
rect 30472 34731 30524 34740
rect 30472 34697 30481 34731
rect 30481 34697 30515 34731
rect 30515 34697 30524 34731
rect 30472 34688 30524 34697
rect 30656 34688 30708 34740
rect 31392 34731 31444 34740
rect 31392 34697 31401 34731
rect 31401 34697 31435 34731
rect 31435 34697 31444 34731
rect 31392 34688 31444 34697
rect 34428 34688 34480 34740
rect 34612 34688 34664 34740
rect 35900 34688 35952 34740
rect 38936 34688 38988 34740
rect 28540 34620 28592 34672
rect 30564 34620 30616 34672
rect 1768 34595 1820 34604
rect 1768 34561 1777 34595
rect 1777 34561 1811 34595
rect 1811 34561 1820 34595
rect 1768 34552 1820 34561
rect 24952 34552 25004 34604
rect 27160 34552 27212 34604
rect 29828 34552 29880 34604
rect 22560 34484 22612 34536
rect 23848 34484 23900 34536
rect 25136 34484 25188 34536
rect 25872 34527 25924 34536
rect 25872 34493 25881 34527
rect 25881 34493 25915 34527
rect 25915 34493 25924 34527
rect 25872 34484 25924 34493
rect 26332 34484 26384 34536
rect 28540 34527 28592 34536
rect 28540 34493 28549 34527
rect 28549 34493 28583 34527
rect 28583 34493 28592 34527
rect 28540 34484 28592 34493
rect 29092 34484 29144 34536
rect 29920 34484 29972 34536
rect 30288 34484 30340 34536
rect 20444 34348 20496 34400
rect 28172 34416 28224 34468
rect 30104 34416 30156 34468
rect 30748 34484 30800 34536
rect 32680 34595 32732 34604
rect 32680 34561 32689 34595
rect 32689 34561 32723 34595
rect 32723 34561 32732 34595
rect 32680 34552 32732 34561
rect 25136 34348 25188 34400
rect 30564 34348 30616 34400
rect 30932 34348 30984 34400
rect 33784 34416 33836 34468
rect 35716 34620 35768 34672
rect 39488 34731 39540 34740
rect 39488 34697 39497 34731
rect 39497 34697 39531 34731
rect 39531 34697 39540 34731
rect 39488 34688 39540 34697
rect 39580 34688 39632 34740
rect 35808 34552 35860 34604
rect 33968 34484 34020 34536
rect 37188 34484 37240 34536
rect 37832 34552 37884 34604
rect 39856 34552 39908 34604
rect 40592 34595 40644 34604
rect 40592 34561 40601 34595
rect 40601 34561 40635 34595
rect 40635 34561 40644 34595
rect 40592 34552 40644 34561
rect 40868 34552 40920 34604
rect 39948 34484 40000 34536
rect 36084 34416 36136 34468
rect 40408 34416 40460 34468
rect 39948 34348 40000 34400
rect 40224 34391 40276 34400
rect 40224 34357 40233 34391
rect 40233 34357 40267 34391
rect 40267 34357 40276 34391
rect 40224 34348 40276 34357
rect 40776 34348 40828 34400
rect 41420 34688 41472 34740
rect 41788 34552 41840 34604
rect 42800 34620 42852 34672
rect 43628 34620 43680 34672
rect 49148 34620 49200 34672
rect 49332 34595 49384 34604
rect 49332 34561 49341 34595
rect 49341 34561 49375 34595
rect 49375 34561 49384 34595
rect 49332 34552 49384 34561
rect 43352 34484 43404 34536
rect 43444 34484 43496 34536
rect 43536 34527 43588 34536
rect 43536 34493 43545 34527
rect 43545 34493 43579 34527
rect 43579 34493 43588 34527
rect 43536 34484 43588 34493
rect 44272 34484 44324 34536
rect 49056 34484 49108 34536
rect 2950 34246 3002 34298
rect 3014 34246 3066 34298
rect 3078 34246 3130 34298
rect 3142 34246 3194 34298
rect 3206 34246 3258 34298
rect 12950 34246 13002 34298
rect 13014 34246 13066 34298
rect 13078 34246 13130 34298
rect 13142 34246 13194 34298
rect 13206 34246 13258 34298
rect 22950 34246 23002 34298
rect 23014 34246 23066 34298
rect 23078 34246 23130 34298
rect 23142 34246 23194 34298
rect 23206 34246 23258 34298
rect 32950 34246 33002 34298
rect 33014 34246 33066 34298
rect 33078 34246 33130 34298
rect 33142 34246 33194 34298
rect 33206 34246 33258 34298
rect 42950 34246 43002 34298
rect 43014 34246 43066 34298
rect 43078 34246 43130 34298
rect 43142 34246 43194 34298
rect 43206 34246 43258 34298
rect 20812 34144 20864 34196
rect 28172 34144 28224 34196
rect 30656 34144 30708 34196
rect 32680 34144 32732 34196
rect 34612 34144 34664 34196
rect 35348 34144 35400 34196
rect 35440 34144 35492 34196
rect 23388 34076 23440 34128
rect 22008 34008 22060 34060
rect 22376 34008 22428 34060
rect 36360 34076 36412 34128
rect 23940 34051 23992 34060
rect 23940 34017 23949 34051
rect 23949 34017 23983 34051
rect 23983 34017 23992 34051
rect 23940 34008 23992 34017
rect 25228 34051 25280 34060
rect 25228 34017 25237 34051
rect 25237 34017 25271 34051
rect 25271 34017 25280 34051
rect 25228 34008 25280 34017
rect 27160 34008 27212 34060
rect 34612 34008 34664 34060
rect 36084 34008 36136 34060
rect 22836 33940 22888 33992
rect 23296 33940 23348 33992
rect 23848 33940 23900 33992
rect 27620 33940 27672 33992
rect 29092 33940 29144 33992
rect 30564 33940 30616 33992
rect 35808 33940 35860 33992
rect 38614 34144 38666 34196
rect 38936 34144 38988 34196
rect 36636 34076 36688 34128
rect 37188 34008 37240 34060
rect 37740 34051 37792 34060
rect 37740 34017 37749 34051
rect 37749 34017 37783 34051
rect 37783 34017 37792 34051
rect 37740 34008 37792 34017
rect 38476 34008 38528 34060
rect 38660 34008 38712 34060
rect 38752 34051 38804 34060
rect 38752 34017 38761 34051
rect 38761 34017 38795 34051
rect 38795 34017 38804 34051
rect 38752 34008 38804 34017
rect 39580 34076 39632 34128
rect 42156 34076 42208 34128
rect 38844 33940 38896 33992
rect 41328 33940 41380 33992
rect 23480 33872 23532 33924
rect 26608 33872 26660 33924
rect 36452 33915 36504 33924
rect 36452 33881 36461 33915
rect 36461 33881 36495 33915
rect 36495 33881 36504 33915
rect 36452 33872 36504 33881
rect 36544 33872 36596 33924
rect 39396 33872 39448 33924
rect 23388 33804 23440 33856
rect 23756 33847 23808 33856
rect 23756 33813 23765 33847
rect 23765 33813 23799 33847
rect 23799 33813 23808 33847
rect 23756 33804 23808 33813
rect 27804 33804 27856 33856
rect 27988 33847 28040 33856
rect 27988 33813 27997 33847
rect 27997 33813 28031 33847
rect 28031 33813 28040 33847
rect 27988 33804 28040 33813
rect 31116 33847 31168 33856
rect 31116 33813 31125 33847
rect 31125 33813 31159 33847
rect 31159 33813 31168 33847
rect 31116 33804 31168 33813
rect 31208 33847 31260 33856
rect 31208 33813 31217 33847
rect 31217 33813 31251 33847
rect 31251 33813 31260 33847
rect 31208 33804 31260 33813
rect 33784 33804 33836 33856
rect 37096 33804 37148 33856
rect 37740 33804 37792 33856
rect 38614 33804 38666 33856
rect 39764 33804 39816 33856
rect 42248 33940 42300 33992
rect 49332 33983 49384 33992
rect 49332 33949 49341 33983
rect 49341 33949 49375 33983
rect 49375 33949 49384 33983
rect 49332 33940 49384 33949
rect 48320 33872 48372 33924
rect 48596 33804 48648 33856
rect 7950 33702 8002 33754
rect 8014 33702 8066 33754
rect 8078 33702 8130 33754
rect 8142 33702 8194 33754
rect 8206 33702 8258 33754
rect 17950 33702 18002 33754
rect 18014 33702 18066 33754
rect 18078 33702 18130 33754
rect 18142 33702 18194 33754
rect 18206 33702 18258 33754
rect 27950 33702 28002 33754
rect 28014 33702 28066 33754
rect 28078 33702 28130 33754
rect 28142 33702 28194 33754
rect 28206 33702 28258 33754
rect 37950 33702 38002 33754
rect 38014 33702 38066 33754
rect 38078 33702 38130 33754
rect 38142 33702 38194 33754
rect 38206 33702 38258 33754
rect 47950 33702 48002 33754
rect 48014 33702 48066 33754
rect 48078 33702 48130 33754
rect 48142 33702 48194 33754
rect 48206 33702 48258 33754
rect 23664 33643 23716 33652
rect 23664 33609 23673 33643
rect 23673 33609 23707 33643
rect 23707 33609 23716 33643
rect 23664 33600 23716 33609
rect 29000 33600 29052 33652
rect 29092 33643 29144 33652
rect 29092 33609 29101 33643
rect 29101 33609 29135 33643
rect 29135 33609 29144 33643
rect 29092 33600 29144 33609
rect 21456 33464 21508 33516
rect 25780 33464 25832 33516
rect 26700 33464 26752 33516
rect 24216 33439 24268 33448
rect 24216 33405 24225 33439
rect 24225 33405 24259 33439
rect 24259 33405 24268 33439
rect 24216 33396 24268 33405
rect 27344 33396 27396 33448
rect 27252 33328 27304 33380
rect 29092 33396 29144 33448
rect 29460 33396 29512 33448
rect 29644 33464 29696 33516
rect 37004 33600 37056 33652
rect 33876 33532 33928 33584
rect 31116 33464 31168 33516
rect 33968 33507 34020 33516
rect 33968 33473 33977 33507
rect 33977 33473 34011 33507
rect 34011 33473 34020 33507
rect 33968 33464 34020 33473
rect 34704 33396 34756 33448
rect 35716 33532 35768 33584
rect 36636 33532 36688 33584
rect 37372 33532 37424 33584
rect 38292 33532 38344 33584
rect 40132 33600 40184 33652
rect 39304 33532 39356 33584
rect 37832 33507 37884 33516
rect 37832 33473 37841 33507
rect 37841 33473 37875 33507
rect 37875 33473 37884 33507
rect 37832 33464 37884 33473
rect 41972 33600 42024 33652
rect 42616 33532 42668 33584
rect 43996 33532 44048 33584
rect 35716 33396 35768 33448
rect 37280 33396 37332 33448
rect 28816 33260 28868 33312
rect 28954 33260 29006 33312
rect 29184 33260 29236 33312
rect 30104 33260 30156 33312
rect 30656 33260 30708 33312
rect 36452 33328 36504 33380
rect 39396 33439 39448 33448
rect 39396 33405 39405 33439
rect 39405 33405 39439 33439
rect 39439 33405 39448 33439
rect 39396 33396 39448 33405
rect 40316 33439 40368 33448
rect 40316 33405 40325 33439
rect 40325 33405 40359 33439
rect 40359 33405 40368 33439
rect 40316 33396 40368 33405
rect 40592 33439 40644 33448
rect 40592 33405 40601 33439
rect 40601 33405 40635 33439
rect 40635 33405 40644 33439
rect 40592 33396 40644 33405
rect 41880 33396 41932 33448
rect 38384 33260 38436 33312
rect 39028 33260 39080 33312
rect 40960 33260 41012 33312
rect 42156 33260 42208 33312
rect 2950 33158 3002 33210
rect 3014 33158 3066 33210
rect 3078 33158 3130 33210
rect 3142 33158 3194 33210
rect 3206 33158 3258 33210
rect 12950 33158 13002 33210
rect 13014 33158 13066 33210
rect 13078 33158 13130 33210
rect 13142 33158 13194 33210
rect 13206 33158 13258 33210
rect 22950 33158 23002 33210
rect 23014 33158 23066 33210
rect 23078 33158 23130 33210
rect 23142 33158 23194 33210
rect 23206 33158 23258 33210
rect 32950 33158 33002 33210
rect 33014 33158 33066 33210
rect 33078 33158 33130 33210
rect 33142 33158 33194 33210
rect 33206 33158 33258 33210
rect 42950 33158 43002 33210
rect 43014 33158 43066 33210
rect 43078 33158 43130 33210
rect 43142 33158 43194 33210
rect 43206 33158 43258 33210
rect 27804 33056 27856 33108
rect 30288 33056 30340 33108
rect 31484 33056 31536 33108
rect 34796 33056 34848 33108
rect 23756 32988 23808 33040
rect 23940 32920 23992 32972
rect 22284 32895 22336 32904
rect 22284 32861 22293 32895
rect 22293 32861 22327 32895
rect 22327 32861 22336 32895
rect 22284 32852 22336 32861
rect 23848 32852 23900 32904
rect 24308 32920 24360 32972
rect 26976 32920 27028 32972
rect 27252 32963 27304 32972
rect 27252 32929 27261 32963
rect 27261 32929 27295 32963
rect 27295 32929 27304 32963
rect 27252 32920 27304 32929
rect 28632 32920 28684 32972
rect 28724 32852 28776 32904
rect 30196 32963 30248 32972
rect 30196 32929 30205 32963
rect 30205 32929 30239 32963
rect 30239 32929 30248 32963
rect 30196 32920 30248 32929
rect 22836 32784 22888 32836
rect 21548 32716 21600 32768
rect 26424 32784 26476 32836
rect 28908 32827 28960 32836
rect 28908 32793 28917 32827
rect 28917 32793 28951 32827
rect 28951 32793 28960 32827
rect 28908 32784 28960 32793
rect 29000 32784 29052 32836
rect 31300 32920 31352 32972
rect 31484 32963 31536 32972
rect 31484 32929 31493 32963
rect 31493 32929 31527 32963
rect 31527 32929 31536 32963
rect 31484 32920 31536 32929
rect 40592 33056 40644 33108
rect 40868 33056 40920 33108
rect 48780 33056 48832 33108
rect 35440 32920 35492 32972
rect 35716 32920 35768 32972
rect 38568 32988 38620 33040
rect 37740 32920 37792 32972
rect 38752 32920 38804 32972
rect 38936 32963 38988 32972
rect 38936 32929 38945 32963
rect 38945 32929 38979 32963
rect 38979 32929 38988 32963
rect 38936 32920 38988 32929
rect 43720 32988 43772 33040
rect 24032 32716 24084 32768
rect 24492 32716 24544 32768
rect 26516 32716 26568 32768
rect 26608 32759 26660 32768
rect 26608 32725 26617 32759
rect 26617 32725 26651 32759
rect 26651 32725 26660 32759
rect 26608 32716 26660 32725
rect 28724 32716 28776 32768
rect 29276 32716 29328 32768
rect 31760 32852 31812 32904
rect 32312 32852 32364 32904
rect 35900 32895 35952 32904
rect 35900 32861 35909 32895
rect 35909 32861 35943 32895
rect 35943 32861 35952 32895
rect 35900 32852 35952 32861
rect 37832 32852 37884 32904
rect 40592 32852 40644 32904
rect 40684 32852 40736 32904
rect 31300 32759 31352 32768
rect 31300 32725 31309 32759
rect 31309 32725 31343 32759
rect 31343 32725 31352 32759
rect 31300 32716 31352 32725
rect 32220 32716 32272 32768
rect 35716 32784 35768 32836
rect 36636 32784 36688 32836
rect 42064 32963 42116 32972
rect 42064 32929 42073 32963
rect 42073 32929 42107 32963
rect 42107 32929 42116 32963
rect 42064 32920 42116 32929
rect 42248 32963 42300 32972
rect 42248 32929 42257 32963
rect 42257 32929 42291 32963
rect 42291 32929 42300 32963
rect 42248 32920 42300 32929
rect 41972 32895 42024 32904
rect 41972 32861 41981 32895
rect 41981 32861 42015 32895
rect 42015 32861 42024 32895
rect 41972 32852 42024 32861
rect 43812 32895 43864 32904
rect 43812 32861 43821 32895
rect 43821 32861 43855 32895
rect 43855 32861 43864 32895
rect 43812 32852 43864 32861
rect 49332 32895 49384 32904
rect 49332 32861 49341 32895
rect 49341 32861 49375 32895
rect 49375 32861 49384 32895
rect 49332 32852 49384 32861
rect 34612 32716 34664 32768
rect 35348 32759 35400 32768
rect 35348 32725 35357 32759
rect 35357 32725 35391 32759
rect 35391 32725 35400 32759
rect 35348 32716 35400 32725
rect 37188 32716 37240 32768
rect 41328 32784 41380 32836
rect 41420 32784 41472 32836
rect 39120 32716 39172 32768
rect 40132 32716 40184 32768
rect 40500 32716 40552 32768
rect 40960 32716 41012 32768
rect 46388 32716 46440 32768
rect 49148 32759 49200 32768
rect 49148 32725 49157 32759
rect 49157 32725 49191 32759
rect 49191 32725 49200 32759
rect 49148 32716 49200 32725
rect 7950 32614 8002 32666
rect 8014 32614 8066 32666
rect 8078 32614 8130 32666
rect 8142 32614 8194 32666
rect 8206 32614 8258 32666
rect 17950 32614 18002 32666
rect 18014 32614 18066 32666
rect 18078 32614 18130 32666
rect 18142 32614 18194 32666
rect 18206 32614 18258 32666
rect 27950 32614 28002 32666
rect 28014 32614 28066 32666
rect 28078 32614 28130 32666
rect 28142 32614 28194 32666
rect 28206 32614 28258 32666
rect 37950 32614 38002 32666
rect 38014 32614 38066 32666
rect 38078 32614 38130 32666
rect 38142 32614 38194 32666
rect 38206 32614 38258 32666
rect 47950 32614 48002 32666
rect 48014 32614 48066 32666
rect 48078 32614 48130 32666
rect 48142 32614 48194 32666
rect 48206 32614 48258 32666
rect 17224 32555 17276 32564
rect 17224 32521 17233 32555
rect 17233 32521 17267 32555
rect 17267 32521 17276 32555
rect 17224 32512 17276 32521
rect 25228 32512 25280 32564
rect 26056 32512 26108 32564
rect 31300 32512 31352 32564
rect 36544 32512 36596 32564
rect 39580 32512 39632 32564
rect 41328 32512 41380 32564
rect 41512 32512 41564 32564
rect 47124 32512 47176 32564
rect 22836 32444 22888 32496
rect 24676 32444 24728 32496
rect 26516 32444 26568 32496
rect 940 32376 992 32428
rect 29092 32444 29144 32496
rect 34704 32444 34756 32496
rect 35624 32444 35676 32496
rect 36636 32444 36688 32496
rect 40040 32444 40092 32496
rect 41420 32444 41472 32496
rect 42616 32444 42668 32496
rect 5724 32308 5776 32360
rect 7472 32172 7524 32224
rect 17868 32351 17920 32360
rect 17868 32317 17877 32351
rect 17877 32317 17911 32351
rect 17911 32317 17920 32351
rect 17868 32308 17920 32317
rect 18512 32215 18564 32224
rect 18512 32181 18521 32215
rect 18521 32181 18555 32215
rect 18555 32181 18564 32215
rect 18512 32172 18564 32181
rect 22560 32172 22612 32224
rect 24216 32351 24268 32360
rect 24216 32317 24225 32351
rect 24225 32317 24259 32351
rect 24259 32317 24268 32351
rect 24216 32308 24268 32317
rect 24676 32308 24728 32360
rect 26240 32308 26292 32360
rect 28540 32308 28592 32360
rect 34612 32376 34664 32428
rect 37464 32376 37516 32428
rect 44088 32376 44140 32428
rect 48780 32419 48832 32428
rect 48780 32385 48789 32419
rect 48789 32385 48823 32419
rect 48823 32385 48832 32419
rect 48780 32376 48832 32385
rect 31944 32308 31996 32360
rect 26608 32240 26660 32292
rect 28724 32240 28776 32292
rect 34244 32283 34296 32292
rect 34244 32249 34253 32283
rect 34253 32249 34287 32283
rect 34287 32249 34296 32283
rect 34244 32240 34296 32249
rect 34980 32240 35032 32292
rect 35164 32308 35216 32360
rect 39028 32308 39080 32360
rect 42156 32308 42208 32360
rect 48504 32351 48556 32360
rect 48504 32317 48513 32351
rect 48513 32317 48547 32351
rect 48547 32317 48556 32351
rect 48504 32308 48556 32317
rect 36084 32240 36136 32292
rect 38476 32240 38528 32292
rect 41328 32240 41380 32292
rect 49148 32240 49200 32292
rect 24860 32172 24912 32224
rect 32128 32172 32180 32224
rect 34888 32172 34940 32224
rect 35716 32172 35768 32224
rect 39948 32172 40000 32224
rect 42800 32215 42852 32224
rect 42800 32181 42809 32215
rect 42809 32181 42843 32215
rect 42843 32181 42852 32215
rect 42800 32172 42852 32181
rect 44640 32215 44692 32224
rect 44640 32181 44649 32215
rect 44649 32181 44683 32215
rect 44683 32181 44692 32215
rect 44640 32172 44692 32181
rect 2950 32070 3002 32122
rect 3014 32070 3066 32122
rect 3078 32070 3130 32122
rect 3142 32070 3194 32122
rect 3206 32070 3258 32122
rect 12950 32070 13002 32122
rect 13014 32070 13066 32122
rect 13078 32070 13130 32122
rect 13142 32070 13194 32122
rect 13206 32070 13258 32122
rect 22950 32070 23002 32122
rect 23014 32070 23066 32122
rect 23078 32070 23130 32122
rect 23142 32070 23194 32122
rect 23206 32070 23258 32122
rect 32950 32070 33002 32122
rect 33014 32070 33066 32122
rect 33078 32070 33130 32122
rect 33142 32070 33194 32122
rect 33206 32070 33258 32122
rect 42950 32070 43002 32122
rect 43014 32070 43066 32122
rect 43078 32070 43130 32122
rect 43142 32070 43194 32122
rect 43206 32070 43258 32122
rect 22560 31968 22612 32020
rect 23940 31968 23992 32020
rect 23848 31832 23900 31884
rect 27068 31968 27120 32020
rect 28448 32011 28500 32020
rect 28448 31977 28457 32011
rect 28457 31977 28491 32011
rect 28491 31977 28500 32011
rect 28448 31968 28500 31977
rect 34336 31968 34388 32020
rect 26056 31875 26108 31884
rect 26056 31841 26065 31875
rect 26065 31841 26099 31875
rect 26099 31841 26108 31875
rect 26056 31832 26108 31841
rect 27252 31832 27304 31884
rect 31668 31900 31720 31952
rect 32036 31900 32088 31952
rect 28632 31832 28684 31884
rect 31760 31832 31812 31884
rect 33692 31832 33744 31884
rect 35256 31900 35308 31952
rect 36268 31900 36320 31952
rect 36728 31900 36780 31952
rect 38660 31900 38712 31952
rect 36176 31832 36228 31884
rect 37280 31832 37332 31884
rect 37648 31832 37700 31884
rect 21824 31807 21876 31816
rect 21824 31773 21833 31807
rect 21833 31773 21867 31807
rect 21867 31773 21876 31807
rect 21824 31764 21876 31773
rect 24768 31807 24820 31816
rect 24768 31773 24777 31807
rect 24777 31773 24811 31807
rect 24811 31773 24820 31807
rect 24768 31764 24820 31773
rect 37832 31764 37884 31816
rect 38476 31875 38528 31884
rect 38476 31841 38485 31875
rect 38485 31841 38519 31875
rect 38519 31841 38528 31875
rect 38476 31832 38528 31841
rect 38568 31832 38620 31884
rect 43444 31968 43496 32020
rect 43904 31968 43956 32020
rect 39028 31832 39080 31884
rect 40316 31832 40368 31884
rect 42708 31832 42760 31884
rect 47124 31832 47176 31884
rect 40040 31764 40092 31816
rect 41512 31764 41564 31816
rect 48504 31807 48556 31816
rect 48504 31773 48513 31807
rect 48513 31773 48547 31807
rect 48547 31773 48556 31807
rect 48504 31764 48556 31773
rect 22836 31696 22888 31748
rect 27528 31696 27580 31748
rect 27804 31696 27856 31748
rect 27712 31628 27764 31680
rect 40224 31696 40276 31748
rect 42616 31696 42668 31748
rect 34152 31628 34204 31680
rect 35808 31628 35860 31680
rect 36636 31628 36688 31680
rect 38476 31628 38528 31680
rect 41512 31628 41564 31680
rect 7950 31526 8002 31578
rect 8014 31526 8066 31578
rect 8078 31526 8130 31578
rect 8142 31526 8194 31578
rect 8206 31526 8258 31578
rect 17950 31526 18002 31578
rect 18014 31526 18066 31578
rect 18078 31526 18130 31578
rect 18142 31526 18194 31578
rect 18206 31526 18258 31578
rect 27950 31526 28002 31578
rect 28014 31526 28066 31578
rect 28078 31526 28130 31578
rect 28142 31526 28194 31578
rect 28206 31526 28258 31578
rect 37950 31526 38002 31578
rect 38014 31526 38066 31578
rect 38078 31526 38130 31578
rect 38142 31526 38194 31578
rect 38206 31526 38258 31578
rect 47950 31526 48002 31578
rect 48014 31526 48066 31578
rect 48078 31526 48130 31578
rect 48142 31526 48194 31578
rect 48206 31526 48258 31578
rect 23480 31467 23532 31476
rect 23480 31433 23489 31467
rect 23489 31433 23523 31467
rect 23523 31433 23532 31467
rect 23480 31424 23532 31433
rect 24768 31424 24820 31476
rect 25412 31424 25464 31476
rect 22468 31263 22520 31272
rect 22468 31229 22477 31263
rect 22477 31229 22511 31263
rect 22511 31229 22520 31263
rect 22468 31220 22520 31229
rect 25044 31356 25096 31408
rect 24860 31331 24912 31340
rect 24860 31297 24869 31331
rect 24869 31297 24903 31331
rect 24903 31297 24912 31331
rect 24860 31288 24912 31297
rect 26240 31288 26292 31340
rect 26700 31424 26752 31476
rect 32036 31424 32088 31476
rect 27160 31356 27212 31408
rect 27804 31288 27856 31340
rect 34612 31356 34664 31408
rect 36084 31424 36136 31476
rect 36820 31424 36872 31476
rect 37924 31356 37976 31408
rect 38568 31467 38620 31476
rect 38568 31433 38577 31467
rect 38577 31433 38611 31467
rect 38611 31433 38620 31467
rect 38568 31424 38620 31433
rect 38660 31424 38712 31476
rect 40040 31424 40092 31476
rect 40224 31424 40276 31476
rect 41328 31424 41380 31476
rect 42800 31424 42852 31476
rect 33600 31288 33652 31340
rect 36544 31288 36596 31340
rect 38384 31288 38436 31340
rect 38568 31288 38620 31340
rect 43536 31356 43588 31408
rect 22836 31220 22888 31272
rect 24216 31220 24268 31272
rect 25136 31263 25188 31272
rect 25136 31229 25145 31263
rect 25145 31229 25179 31263
rect 25179 31229 25188 31263
rect 25136 31220 25188 31229
rect 24952 31084 25004 31136
rect 32036 31220 32088 31272
rect 32404 31220 32456 31272
rect 32680 31220 32732 31272
rect 34336 31220 34388 31272
rect 26884 31084 26936 31136
rect 27528 31084 27580 31136
rect 29276 31084 29328 31136
rect 32864 31084 32916 31136
rect 35164 31220 35216 31272
rect 38476 31220 38528 31272
rect 42156 31288 42208 31340
rect 44272 31288 44324 31340
rect 48320 31288 48372 31340
rect 48504 31263 48556 31272
rect 48504 31229 48513 31263
rect 48513 31229 48547 31263
rect 48547 31229 48556 31263
rect 48504 31220 48556 31229
rect 35900 31084 35952 31136
rect 40408 31084 40460 31136
rect 40500 31084 40552 31136
rect 44364 31152 44416 31204
rect 45560 31152 45612 31204
rect 47860 31084 47912 31136
rect 2950 30982 3002 31034
rect 3014 30982 3066 31034
rect 3078 30982 3130 31034
rect 3142 30982 3194 31034
rect 3206 30982 3258 31034
rect 12950 30982 13002 31034
rect 13014 30982 13066 31034
rect 13078 30982 13130 31034
rect 13142 30982 13194 31034
rect 13206 30982 13258 31034
rect 22950 30982 23002 31034
rect 23014 30982 23066 31034
rect 23078 30982 23130 31034
rect 23142 30982 23194 31034
rect 23206 30982 23258 31034
rect 32950 30982 33002 31034
rect 33014 30982 33066 31034
rect 33078 30982 33130 31034
rect 33142 30982 33194 31034
rect 33206 30982 33258 31034
rect 42950 30982 43002 31034
rect 43014 30982 43066 31034
rect 43078 30982 43130 31034
rect 43142 30982 43194 31034
rect 43206 30982 43258 31034
rect 21456 30923 21508 30932
rect 21456 30889 21465 30923
rect 21465 30889 21499 30923
rect 21499 30889 21508 30923
rect 21456 30880 21508 30889
rect 23388 30880 23440 30932
rect 27528 30880 27580 30932
rect 30196 30880 30248 30932
rect 22100 30787 22152 30796
rect 22100 30753 22109 30787
rect 22109 30753 22143 30787
rect 22143 30753 22152 30787
rect 22100 30744 22152 30753
rect 23848 30787 23900 30796
rect 23848 30753 23857 30787
rect 23857 30753 23891 30787
rect 23891 30753 23900 30787
rect 23848 30744 23900 30753
rect 27068 30787 27120 30796
rect 27068 30753 27077 30787
rect 27077 30753 27111 30787
rect 27111 30753 27120 30787
rect 27068 30744 27120 30753
rect 28908 30812 28960 30864
rect 32588 30812 32640 30864
rect 34888 30812 34940 30864
rect 21824 30719 21876 30728
rect 21824 30685 21833 30719
rect 21833 30685 21867 30719
rect 21867 30685 21876 30719
rect 21824 30676 21876 30685
rect 23388 30676 23440 30728
rect 9128 30608 9180 30660
rect 21916 30651 21968 30660
rect 21916 30617 21925 30651
rect 21925 30617 21959 30651
rect 21959 30617 21968 30651
rect 21916 30608 21968 30617
rect 23296 30608 23348 30660
rect 24860 30719 24912 30728
rect 24860 30685 24869 30719
rect 24869 30685 24903 30719
rect 24903 30685 24912 30719
rect 24860 30676 24912 30685
rect 29276 30744 29328 30796
rect 23572 30583 23624 30592
rect 23572 30549 23581 30583
rect 23581 30549 23615 30583
rect 23615 30549 23624 30583
rect 23572 30540 23624 30549
rect 26884 30608 26936 30660
rect 27344 30651 27396 30660
rect 27344 30617 27353 30651
rect 27353 30617 27387 30651
rect 27387 30617 27396 30651
rect 27344 30608 27396 30617
rect 27252 30540 27304 30592
rect 27436 30540 27488 30592
rect 30564 30676 30616 30728
rect 31944 30744 31996 30796
rect 32312 30744 32364 30796
rect 33324 30676 33376 30728
rect 35440 30880 35492 30932
rect 37464 30880 37516 30932
rect 37556 30880 37608 30932
rect 38476 30880 38528 30932
rect 39672 30880 39724 30932
rect 40500 30880 40552 30932
rect 28816 30583 28868 30592
rect 28816 30549 28825 30583
rect 28825 30549 28859 30583
rect 28859 30549 28868 30583
rect 28816 30540 28868 30549
rect 30196 30583 30248 30592
rect 30196 30549 30205 30583
rect 30205 30549 30239 30583
rect 30239 30549 30248 30583
rect 30196 30540 30248 30549
rect 31576 30651 31628 30660
rect 31576 30617 31585 30651
rect 31585 30617 31619 30651
rect 31619 30617 31628 30651
rect 31576 30608 31628 30617
rect 35716 30744 35768 30796
rect 40224 30812 40276 30864
rect 40316 30812 40368 30864
rect 37924 30787 37976 30796
rect 37924 30753 37933 30787
rect 37933 30753 37967 30787
rect 37967 30753 37976 30787
rect 37924 30744 37976 30753
rect 38660 30744 38712 30796
rect 40040 30744 40092 30796
rect 37556 30676 37608 30728
rect 39488 30676 39540 30728
rect 40408 30719 40460 30728
rect 40408 30685 40417 30719
rect 40417 30685 40451 30719
rect 40451 30685 40460 30719
rect 40408 30676 40460 30685
rect 48596 30744 48648 30796
rect 41512 30719 41564 30728
rect 41512 30685 41521 30719
rect 41521 30685 41555 30719
rect 41555 30685 41564 30719
rect 41512 30676 41564 30685
rect 41604 30676 41656 30728
rect 43352 30676 43404 30728
rect 34980 30583 35032 30592
rect 34980 30549 34989 30583
rect 34989 30549 35023 30583
rect 35023 30549 35032 30583
rect 34980 30540 35032 30549
rect 35532 30540 35584 30592
rect 36544 30583 36596 30592
rect 36544 30549 36553 30583
rect 36553 30549 36587 30583
rect 36587 30549 36596 30583
rect 36544 30540 36596 30549
rect 37740 30583 37792 30592
rect 37740 30549 37749 30583
rect 37749 30549 37783 30583
rect 37783 30549 37792 30583
rect 37740 30540 37792 30549
rect 38752 30540 38804 30592
rect 41236 30540 41288 30592
rect 46020 30608 46072 30660
rect 42800 30540 42852 30592
rect 45468 30540 45520 30592
rect 7950 30438 8002 30490
rect 8014 30438 8066 30490
rect 8078 30438 8130 30490
rect 8142 30438 8194 30490
rect 8206 30438 8258 30490
rect 17950 30438 18002 30490
rect 18014 30438 18066 30490
rect 18078 30438 18130 30490
rect 18142 30438 18194 30490
rect 18206 30438 18258 30490
rect 27950 30438 28002 30490
rect 28014 30438 28066 30490
rect 28078 30438 28130 30490
rect 28142 30438 28194 30490
rect 28206 30438 28258 30490
rect 37950 30438 38002 30490
rect 38014 30438 38066 30490
rect 38078 30438 38130 30490
rect 38142 30438 38194 30490
rect 38206 30438 38258 30490
rect 47950 30438 48002 30490
rect 48014 30438 48066 30490
rect 48078 30438 48130 30490
rect 48142 30438 48194 30490
rect 48206 30438 48258 30490
rect 20260 30336 20312 30388
rect 27620 30336 27672 30388
rect 28264 30336 28316 30388
rect 30288 30336 30340 30388
rect 31576 30336 31628 30388
rect 34244 30336 34296 30388
rect 34428 30336 34480 30388
rect 38936 30336 38988 30388
rect 10692 30268 10744 30320
rect 25596 30311 25648 30320
rect 25596 30277 25605 30311
rect 25605 30277 25639 30311
rect 25639 30277 25648 30311
rect 25596 30268 25648 30277
rect 27068 30268 27120 30320
rect 30564 30268 30616 30320
rect 30656 30268 30708 30320
rect 33416 30268 33468 30320
rect 34336 30268 34388 30320
rect 35808 30268 35860 30320
rect 36268 30268 36320 30320
rect 37832 30311 37884 30320
rect 37832 30277 37841 30311
rect 37841 30277 37875 30311
rect 37875 30277 37884 30311
rect 37832 30268 37884 30277
rect 37924 30311 37976 30320
rect 37924 30277 37933 30311
rect 37933 30277 37967 30311
rect 37967 30277 37976 30311
rect 37924 30268 37976 30277
rect 7380 30243 7432 30252
rect 7380 30209 7389 30243
rect 7389 30209 7423 30243
rect 7423 30209 7432 30243
rect 7380 30200 7432 30209
rect 23572 30200 23624 30252
rect 29000 30200 29052 30252
rect 30012 30200 30064 30252
rect 7656 30132 7708 30184
rect 9128 30175 9180 30184
rect 9128 30141 9137 30175
rect 9137 30141 9171 30175
rect 9171 30141 9180 30175
rect 9128 30132 9180 30141
rect 25044 30175 25096 30184
rect 25044 30141 25053 30175
rect 25053 30141 25087 30175
rect 25087 30141 25096 30175
rect 25044 30132 25096 30141
rect 25872 30132 25924 30184
rect 24584 30064 24636 30116
rect 18696 29996 18748 30048
rect 28264 30064 28316 30116
rect 25780 29996 25832 30048
rect 28908 30175 28960 30184
rect 28908 30141 28917 30175
rect 28917 30141 28951 30175
rect 28951 30141 28960 30175
rect 28908 30132 28960 30141
rect 29828 30132 29880 30184
rect 30748 30064 30800 30116
rect 31024 30175 31076 30184
rect 31024 30141 31033 30175
rect 31033 30141 31067 30175
rect 31067 30141 31076 30175
rect 31024 30132 31076 30141
rect 34704 30200 34756 30252
rect 30932 30064 30984 30116
rect 32772 30064 32824 30116
rect 35992 30132 36044 30184
rect 36084 30175 36136 30184
rect 36084 30141 36093 30175
rect 36093 30141 36127 30175
rect 36127 30141 36136 30175
rect 36084 30132 36136 30141
rect 38016 30175 38068 30184
rect 38016 30141 38025 30175
rect 38025 30141 38059 30175
rect 38059 30141 38068 30175
rect 38016 30132 38068 30141
rect 39028 30268 39080 30320
rect 39580 30268 39632 30320
rect 41144 30268 41196 30320
rect 40224 30200 40276 30252
rect 34520 29996 34572 30048
rect 35900 30064 35952 30116
rect 38384 30064 38436 30116
rect 37372 29996 37424 30048
rect 37464 30039 37516 30048
rect 37464 30005 37473 30039
rect 37473 30005 37507 30039
rect 37507 30005 37516 30039
rect 37464 29996 37516 30005
rect 38568 29996 38620 30048
rect 39028 30132 39080 30184
rect 49332 30243 49384 30252
rect 49332 30209 49341 30243
rect 49341 30209 49375 30243
rect 49375 30209 49384 30243
rect 49332 30200 49384 30209
rect 39948 30064 40000 30116
rect 43536 30064 43588 30116
rect 40316 29996 40368 30048
rect 2950 29894 3002 29946
rect 3014 29894 3066 29946
rect 3078 29894 3130 29946
rect 3142 29894 3194 29946
rect 3206 29894 3258 29946
rect 12950 29894 13002 29946
rect 13014 29894 13066 29946
rect 13078 29894 13130 29946
rect 13142 29894 13194 29946
rect 13206 29894 13258 29946
rect 22950 29894 23002 29946
rect 23014 29894 23066 29946
rect 23078 29894 23130 29946
rect 23142 29894 23194 29946
rect 23206 29894 23258 29946
rect 32950 29894 33002 29946
rect 33014 29894 33066 29946
rect 33078 29894 33130 29946
rect 33142 29894 33194 29946
rect 33206 29894 33258 29946
rect 42950 29894 43002 29946
rect 43014 29894 43066 29946
rect 43078 29894 43130 29946
rect 43142 29894 43194 29946
rect 43206 29894 43258 29946
rect 25044 29792 25096 29844
rect 29552 29792 29604 29844
rect 22652 29724 22704 29776
rect 1308 29656 1360 29708
rect 22560 29656 22612 29708
rect 25872 29724 25924 29776
rect 27344 29656 27396 29708
rect 4896 29588 4948 29640
rect 27620 29656 27672 29708
rect 28908 29656 28960 29708
rect 35348 29792 35400 29844
rect 30012 29724 30064 29776
rect 29828 29588 29880 29640
rect 30104 29656 30156 29708
rect 31944 29724 31996 29776
rect 32680 29724 32732 29776
rect 34060 29724 34112 29776
rect 38016 29792 38068 29844
rect 38292 29792 38344 29844
rect 39028 29792 39080 29844
rect 39120 29792 39172 29844
rect 30012 29588 30064 29640
rect 35900 29656 35952 29708
rect 37648 29656 37700 29708
rect 40316 29656 40368 29708
rect 42708 29835 42760 29844
rect 42708 29801 42717 29835
rect 42717 29801 42751 29835
rect 42751 29801 42760 29835
rect 42708 29792 42760 29801
rect 40040 29588 40092 29640
rect 48504 29631 48556 29640
rect 48504 29597 48513 29631
rect 48513 29597 48547 29631
rect 48547 29597 48556 29631
rect 48504 29588 48556 29597
rect 22468 29563 22520 29572
rect 22468 29529 22477 29563
rect 22477 29529 22511 29563
rect 22511 29529 22520 29563
rect 22468 29520 22520 29529
rect 30196 29520 30248 29572
rect 32220 29520 32272 29572
rect 32680 29520 32732 29572
rect 33692 29520 33744 29572
rect 36636 29563 36688 29572
rect 36636 29529 36645 29563
rect 36645 29529 36679 29563
rect 36679 29529 36688 29563
rect 36636 29520 36688 29529
rect 37096 29520 37148 29572
rect 42616 29520 42668 29572
rect 29368 29452 29420 29504
rect 31300 29452 31352 29504
rect 31760 29452 31812 29504
rect 32404 29495 32456 29504
rect 32404 29461 32413 29495
rect 32413 29461 32447 29495
rect 32447 29461 32456 29495
rect 32404 29452 32456 29461
rect 35900 29452 35952 29504
rect 36268 29452 36320 29504
rect 7950 29350 8002 29402
rect 8014 29350 8066 29402
rect 8078 29350 8130 29402
rect 8142 29350 8194 29402
rect 8206 29350 8258 29402
rect 17950 29350 18002 29402
rect 18014 29350 18066 29402
rect 18078 29350 18130 29402
rect 18142 29350 18194 29402
rect 18206 29350 18258 29402
rect 27950 29350 28002 29402
rect 28014 29350 28066 29402
rect 28078 29350 28130 29402
rect 28142 29350 28194 29402
rect 28206 29350 28258 29402
rect 37950 29350 38002 29402
rect 38014 29350 38066 29402
rect 38078 29350 38130 29402
rect 38142 29350 38194 29402
rect 38206 29350 38258 29402
rect 47950 29350 48002 29402
rect 48014 29350 48066 29402
rect 48078 29350 48130 29402
rect 48142 29350 48194 29402
rect 48206 29350 48258 29402
rect 17316 29248 17368 29300
rect 22836 29248 22888 29300
rect 22100 29180 22152 29232
rect 28816 29248 28868 29300
rect 17408 29112 17460 29164
rect 29276 29180 29328 29232
rect 25136 29044 25188 29096
rect 27068 29112 27120 29164
rect 31208 29248 31260 29300
rect 31300 29248 31352 29300
rect 32404 29248 32456 29300
rect 34612 29248 34664 29300
rect 35164 29248 35216 29300
rect 36728 29248 36780 29300
rect 39672 29291 39724 29300
rect 39672 29257 39681 29291
rect 39681 29257 39715 29291
rect 39715 29257 39724 29291
rect 39672 29248 39724 29257
rect 39764 29291 39816 29300
rect 39764 29257 39773 29291
rect 39773 29257 39807 29291
rect 39807 29257 39816 29291
rect 39764 29248 39816 29257
rect 41236 29291 41288 29300
rect 41236 29257 41245 29291
rect 41245 29257 41279 29291
rect 41279 29257 41288 29291
rect 41236 29248 41288 29257
rect 30012 29180 30064 29232
rect 33784 29180 33836 29232
rect 35992 29180 36044 29232
rect 37188 29180 37240 29232
rect 39212 29180 39264 29232
rect 29460 29087 29512 29096
rect 29460 29053 29469 29087
rect 29469 29053 29503 29087
rect 29503 29053 29512 29087
rect 29460 29044 29512 29053
rect 29828 29044 29880 29096
rect 29000 28976 29052 29028
rect 30012 28976 30064 29028
rect 36636 29112 36688 29164
rect 39672 29112 39724 29164
rect 40776 29112 40828 29164
rect 41144 29155 41196 29164
rect 41144 29121 41153 29155
rect 41153 29121 41187 29155
rect 41187 29121 41196 29155
rect 41144 29112 41196 29121
rect 49332 29155 49384 29164
rect 49332 29121 49341 29155
rect 49341 29121 49375 29155
rect 49375 29121 49384 29155
rect 49332 29112 49384 29121
rect 33968 29087 34020 29096
rect 33968 29053 33977 29087
rect 33977 29053 34011 29087
rect 34011 29053 34020 29087
rect 33968 29044 34020 29053
rect 34612 29044 34664 29096
rect 37096 29044 37148 29096
rect 37832 29044 37884 29096
rect 39856 29087 39908 29096
rect 39856 29053 39865 29087
rect 39865 29053 39899 29087
rect 39899 29053 39908 29087
rect 39856 29044 39908 29053
rect 42708 29044 42760 29096
rect 33416 28976 33468 29028
rect 33692 28976 33744 29028
rect 38384 28976 38436 29028
rect 40040 28976 40092 29028
rect 43996 28976 44048 29028
rect 32312 28908 32364 28960
rect 33968 28908 34020 28960
rect 36268 28908 36320 28960
rect 36360 28951 36412 28960
rect 36360 28917 36369 28951
rect 36369 28917 36403 28951
rect 36403 28917 36412 28951
rect 36360 28908 36412 28917
rect 38660 28951 38712 28960
rect 38660 28917 38669 28951
rect 38669 28917 38703 28951
rect 38703 28917 38712 28951
rect 38660 28908 38712 28917
rect 2950 28806 3002 28858
rect 3014 28806 3066 28858
rect 3078 28806 3130 28858
rect 3142 28806 3194 28858
rect 3206 28806 3258 28858
rect 12950 28806 13002 28858
rect 13014 28806 13066 28858
rect 13078 28806 13130 28858
rect 13142 28806 13194 28858
rect 13206 28806 13258 28858
rect 22950 28806 23002 28858
rect 23014 28806 23066 28858
rect 23078 28806 23130 28858
rect 23142 28806 23194 28858
rect 23206 28806 23258 28858
rect 32950 28806 33002 28858
rect 33014 28806 33066 28858
rect 33078 28806 33130 28858
rect 33142 28806 33194 28858
rect 33206 28806 33258 28858
rect 42950 28806 43002 28858
rect 43014 28806 43066 28858
rect 43078 28806 43130 28858
rect 43142 28806 43194 28858
rect 43206 28806 43258 28858
rect 23296 28704 23348 28756
rect 33324 28704 33376 28756
rect 34612 28704 34664 28756
rect 35624 28704 35676 28756
rect 38568 28704 38620 28756
rect 41144 28704 41196 28756
rect 22192 28636 22244 28688
rect 7196 28500 7248 28552
rect 19524 28568 19576 28620
rect 21640 28500 21692 28552
rect 22008 28568 22060 28620
rect 22284 28568 22336 28620
rect 23204 28636 23256 28688
rect 27620 28636 27672 28688
rect 30380 28636 30432 28688
rect 31944 28636 31996 28688
rect 32956 28636 33008 28688
rect 34980 28636 35032 28688
rect 23388 28568 23440 28620
rect 29460 28568 29512 28620
rect 32864 28568 32916 28620
rect 34152 28611 34204 28620
rect 34152 28577 34161 28611
rect 34161 28577 34195 28611
rect 34195 28577 34204 28611
rect 34152 28568 34204 28577
rect 35624 28568 35676 28620
rect 36268 28568 36320 28620
rect 37372 28611 37424 28620
rect 37372 28577 37381 28611
rect 37381 28577 37415 28611
rect 37415 28577 37424 28611
rect 37372 28568 37424 28577
rect 38568 28568 38620 28620
rect 40316 28568 40368 28620
rect 40684 28611 40736 28620
rect 40684 28577 40693 28611
rect 40693 28577 40727 28611
rect 40727 28577 40736 28611
rect 40684 28568 40736 28577
rect 22376 28500 22428 28552
rect 22560 28500 22612 28552
rect 21824 28432 21876 28484
rect 22468 28432 22520 28484
rect 23204 28432 23256 28484
rect 29920 28543 29972 28552
rect 29920 28509 29929 28543
rect 29929 28509 29963 28543
rect 29963 28509 29972 28543
rect 29920 28500 29972 28509
rect 33600 28500 33652 28552
rect 34796 28500 34848 28552
rect 36360 28500 36412 28552
rect 38660 28500 38712 28552
rect 40960 28500 41012 28552
rect 49332 28543 49384 28552
rect 49332 28509 49341 28543
rect 49341 28509 49375 28543
rect 49375 28509 49384 28543
rect 49332 28500 49384 28509
rect 22008 28364 22060 28416
rect 22376 28407 22428 28416
rect 22376 28373 22385 28407
rect 22385 28373 22419 28407
rect 22419 28373 22428 28407
rect 23296 28407 23348 28416
rect 22376 28364 22428 28373
rect 23296 28373 23305 28407
rect 23305 28373 23339 28407
rect 23339 28373 23348 28407
rect 23296 28364 23348 28373
rect 27068 28475 27120 28484
rect 27068 28441 27077 28475
rect 27077 28441 27111 28475
rect 27111 28441 27120 28475
rect 27068 28432 27120 28441
rect 29736 28432 29788 28484
rect 30656 28407 30708 28416
rect 30656 28373 30665 28407
rect 30665 28373 30699 28407
rect 30699 28373 30708 28407
rect 30656 28364 30708 28373
rect 32220 28432 32272 28484
rect 31300 28364 31352 28416
rect 32772 28364 32824 28416
rect 34796 28364 34848 28416
rect 34980 28364 35032 28416
rect 35348 28407 35400 28416
rect 35348 28373 35357 28407
rect 35357 28373 35391 28407
rect 35391 28373 35400 28407
rect 35348 28364 35400 28373
rect 35440 28364 35492 28416
rect 36544 28407 36596 28416
rect 36544 28373 36553 28407
rect 36553 28373 36587 28407
rect 36587 28373 36596 28407
rect 36544 28364 36596 28373
rect 37188 28364 37240 28416
rect 40132 28432 40184 28484
rect 40316 28364 40368 28416
rect 49148 28407 49200 28416
rect 49148 28373 49157 28407
rect 49157 28373 49191 28407
rect 49191 28373 49200 28407
rect 49148 28364 49200 28373
rect 7950 28262 8002 28314
rect 8014 28262 8066 28314
rect 8078 28262 8130 28314
rect 8142 28262 8194 28314
rect 8206 28262 8258 28314
rect 17950 28262 18002 28314
rect 18014 28262 18066 28314
rect 18078 28262 18130 28314
rect 18142 28262 18194 28314
rect 18206 28262 18258 28314
rect 27950 28262 28002 28314
rect 28014 28262 28066 28314
rect 28078 28262 28130 28314
rect 28142 28262 28194 28314
rect 28206 28262 28258 28314
rect 37950 28262 38002 28314
rect 38014 28262 38066 28314
rect 38078 28262 38130 28314
rect 38142 28262 38194 28314
rect 38206 28262 38258 28314
rect 47950 28262 48002 28314
rect 48014 28262 48066 28314
rect 48078 28262 48130 28314
rect 48142 28262 48194 28314
rect 48206 28262 48258 28314
rect 4896 28203 4948 28212
rect 4896 28169 4905 28203
rect 4905 28169 4939 28203
rect 4939 28169 4948 28203
rect 4896 28160 4948 28169
rect 23388 28160 23440 28212
rect 27436 28160 27488 28212
rect 24952 28092 25004 28144
rect 27712 28092 27764 28144
rect 29460 28160 29512 28212
rect 32128 28160 32180 28212
rect 32404 28160 32456 28212
rect 34152 28160 34204 28212
rect 35900 28160 35952 28212
rect 36452 28203 36504 28212
rect 36452 28169 36461 28203
rect 36461 28169 36495 28203
rect 36495 28169 36504 28203
rect 36452 28160 36504 28169
rect 36544 28160 36596 28212
rect 39212 28160 39264 28212
rect 35348 28092 35400 28144
rect 7564 28067 7616 28076
rect 7564 28033 7573 28067
rect 7573 28033 7607 28067
rect 7607 28033 7616 28067
rect 7564 28024 7616 28033
rect 22008 28024 22060 28076
rect 22284 28024 22336 28076
rect 23756 28024 23808 28076
rect 29276 28024 29328 28076
rect 29460 28024 29512 28076
rect 32312 28067 32364 28076
rect 32312 28033 32321 28067
rect 32321 28033 32355 28067
rect 32355 28033 32364 28067
rect 32312 28024 32364 28033
rect 34152 28024 34204 28076
rect 34612 28024 34664 28076
rect 37464 28024 37516 28076
rect 38384 28135 38436 28144
rect 38384 28101 38393 28135
rect 38393 28101 38427 28135
rect 38427 28101 38436 28135
rect 38384 28092 38436 28101
rect 39304 28092 39356 28144
rect 39580 28092 39632 28144
rect 49148 28092 49200 28144
rect 38844 28024 38896 28076
rect 39212 28024 39264 28076
rect 47860 28024 47912 28076
rect 7748 27999 7800 28008
rect 7748 27965 7757 27999
rect 7757 27965 7791 27999
rect 7791 27965 7800 27999
rect 7748 27956 7800 27965
rect 9588 27956 9640 28008
rect 9680 27888 9732 27940
rect 24400 27820 24452 27872
rect 26608 27956 26660 28008
rect 27804 27956 27856 28008
rect 30104 27956 30156 28008
rect 24860 27820 24912 27872
rect 29184 27820 29236 27872
rect 30840 27863 30892 27872
rect 30840 27829 30849 27863
rect 30849 27829 30883 27863
rect 30883 27829 30892 27863
rect 30840 27820 30892 27829
rect 32956 27956 33008 28008
rect 33324 27956 33376 28008
rect 37280 27956 37332 28008
rect 38292 27956 38344 28008
rect 39672 27999 39724 28008
rect 39672 27965 39681 27999
rect 39681 27965 39715 27999
rect 39715 27965 39724 27999
rect 39672 27956 39724 27965
rect 31576 27888 31628 27940
rect 32220 27888 32272 27940
rect 32588 27820 32640 27872
rect 39396 27820 39448 27872
rect 47860 27820 47912 27872
rect 2950 27718 3002 27770
rect 3014 27718 3066 27770
rect 3078 27718 3130 27770
rect 3142 27718 3194 27770
rect 3206 27718 3258 27770
rect 12950 27718 13002 27770
rect 13014 27718 13066 27770
rect 13078 27718 13130 27770
rect 13142 27718 13194 27770
rect 13206 27718 13258 27770
rect 22950 27718 23002 27770
rect 23014 27718 23066 27770
rect 23078 27718 23130 27770
rect 23142 27718 23194 27770
rect 23206 27718 23258 27770
rect 32950 27718 33002 27770
rect 33014 27718 33066 27770
rect 33078 27718 33130 27770
rect 33142 27718 33194 27770
rect 33206 27718 33258 27770
rect 42950 27718 43002 27770
rect 43014 27718 43066 27770
rect 43078 27718 43130 27770
rect 43142 27718 43194 27770
rect 43206 27718 43258 27770
rect 7656 27548 7708 27600
rect 29460 27548 29512 27600
rect 35164 27548 35216 27600
rect 1308 27480 1360 27532
rect 30288 27480 30340 27532
rect 4896 27412 4948 27464
rect 5448 27412 5500 27464
rect 23112 27412 23164 27464
rect 24860 27455 24912 27464
rect 24860 27421 24869 27455
rect 24869 27421 24903 27455
rect 24903 27421 24912 27455
rect 24860 27412 24912 27421
rect 29920 27412 29972 27464
rect 30380 27412 30432 27464
rect 25136 27387 25188 27396
rect 25136 27353 25145 27387
rect 25145 27353 25179 27387
rect 25179 27353 25188 27387
rect 25136 27344 25188 27353
rect 23480 27276 23532 27328
rect 23756 27276 23808 27328
rect 24952 27276 25004 27328
rect 26700 27344 26752 27396
rect 28724 27344 28776 27396
rect 32220 27523 32272 27532
rect 32220 27489 32229 27523
rect 32229 27489 32263 27523
rect 32263 27489 32272 27523
rect 32220 27480 32272 27489
rect 35256 27480 35308 27532
rect 36084 27548 36136 27600
rect 38568 27548 38620 27600
rect 39672 27548 39724 27600
rect 40040 27523 40092 27532
rect 40040 27489 40049 27523
rect 40049 27489 40083 27523
rect 40083 27489 40092 27523
rect 40040 27480 40092 27489
rect 31668 27412 31720 27464
rect 33968 27412 34020 27464
rect 43996 27455 44048 27464
rect 43996 27421 44005 27455
rect 44005 27421 44039 27455
rect 44039 27421 44048 27455
rect 43996 27412 44048 27421
rect 46388 27412 46440 27464
rect 48504 27455 48556 27464
rect 48504 27421 48513 27455
rect 48513 27421 48547 27455
rect 48547 27421 48556 27455
rect 48504 27412 48556 27421
rect 48596 27412 48648 27464
rect 30932 27344 30984 27396
rect 32956 27344 33008 27396
rect 26608 27319 26660 27328
rect 26608 27285 26617 27319
rect 26617 27285 26651 27319
rect 26651 27285 26660 27319
rect 26608 27276 26660 27285
rect 27252 27276 27304 27328
rect 28448 27276 28500 27328
rect 30196 27319 30248 27328
rect 30196 27285 30205 27319
rect 30205 27285 30239 27319
rect 30239 27285 30248 27319
rect 30196 27276 30248 27285
rect 30564 27319 30616 27328
rect 30564 27285 30573 27319
rect 30573 27285 30607 27319
rect 30607 27285 30616 27319
rect 30564 27276 30616 27285
rect 31944 27276 31996 27328
rect 34612 27276 34664 27328
rect 35072 27276 35124 27328
rect 35440 27344 35492 27396
rect 37096 27344 37148 27396
rect 37832 27344 37884 27396
rect 40408 27344 40460 27396
rect 41604 27344 41656 27396
rect 42616 27344 42668 27396
rect 47584 27344 47636 27396
rect 40960 27276 41012 27328
rect 41052 27276 41104 27328
rect 43720 27276 43772 27328
rect 43812 27319 43864 27328
rect 43812 27285 43821 27319
rect 43821 27285 43855 27319
rect 43855 27285 43864 27319
rect 43812 27276 43864 27285
rect 7950 27174 8002 27226
rect 8014 27174 8066 27226
rect 8078 27174 8130 27226
rect 8142 27174 8194 27226
rect 8206 27174 8258 27226
rect 17950 27174 18002 27226
rect 18014 27174 18066 27226
rect 18078 27174 18130 27226
rect 18142 27174 18194 27226
rect 18206 27174 18258 27226
rect 27950 27174 28002 27226
rect 28014 27174 28066 27226
rect 28078 27174 28130 27226
rect 28142 27174 28194 27226
rect 28206 27174 28258 27226
rect 37950 27174 38002 27226
rect 38014 27174 38066 27226
rect 38078 27174 38130 27226
rect 38142 27174 38194 27226
rect 38206 27174 38258 27226
rect 47950 27174 48002 27226
rect 48014 27174 48066 27226
rect 48078 27174 48130 27226
rect 48142 27174 48194 27226
rect 48206 27174 48258 27226
rect 23112 27115 23164 27124
rect 23112 27081 23121 27115
rect 23121 27081 23155 27115
rect 23155 27081 23164 27115
rect 23112 27072 23164 27081
rect 23296 27072 23348 27124
rect 30288 27115 30340 27124
rect 30288 27081 30297 27115
rect 30297 27081 30331 27115
rect 30331 27081 30340 27115
rect 30288 27072 30340 27081
rect 30564 27072 30616 27124
rect 31392 27072 31444 27124
rect 32496 27072 32548 27124
rect 32680 27072 32732 27124
rect 24860 27004 24912 27056
rect 27804 27004 27856 27056
rect 7840 26979 7892 26988
rect 7840 26945 7849 26979
rect 7849 26945 7883 26979
rect 7883 26945 7892 26979
rect 7840 26936 7892 26945
rect 25504 26936 25556 26988
rect 27620 26936 27672 26988
rect 30104 27004 30156 27056
rect 30748 27004 30800 27056
rect 31208 27004 31260 27056
rect 31300 27004 31352 27056
rect 34152 27004 34204 27056
rect 8300 26868 8352 26920
rect 8944 26911 8996 26920
rect 8944 26877 8953 26911
rect 8953 26877 8987 26911
rect 8987 26877 8996 26911
rect 8944 26868 8996 26877
rect 23388 26911 23440 26920
rect 23388 26877 23397 26911
rect 23397 26877 23431 26911
rect 23431 26877 23440 26911
rect 23388 26868 23440 26877
rect 29184 26868 29236 26920
rect 30564 26868 30616 26920
rect 31576 26936 31628 26988
rect 33692 26936 33744 26988
rect 35900 27115 35952 27124
rect 35900 27081 35909 27115
rect 35909 27081 35943 27115
rect 35943 27081 35952 27115
rect 35900 27072 35952 27081
rect 37096 27072 37148 27124
rect 40684 27072 40736 27124
rect 37556 27004 37608 27056
rect 37464 26979 37516 26988
rect 37464 26945 37473 26979
rect 37473 26945 37507 26979
rect 37507 26945 37516 26979
rect 37464 26936 37516 26945
rect 31116 26800 31168 26852
rect 34060 26868 34112 26920
rect 24124 26732 24176 26784
rect 24216 26775 24268 26784
rect 24216 26741 24225 26775
rect 24225 26741 24259 26775
rect 24259 26741 24268 26775
rect 24216 26732 24268 26741
rect 26516 26732 26568 26784
rect 27344 26732 27396 26784
rect 30380 26732 30432 26784
rect 30472 26732 30524 26784
rect 33968 26732 34020 26784
rect 34428 26911 34480 26920
rect 34428 26877 34437 26911
rect 34437 26877 34471 26911
rect 34471 26877 34480 26911
rect 34428 26868 34480 26877
rect 38292 26911 38344 26920
rect 38292 26877 38301 26911
rect 38301 26877 38335 26911
rect 38335 26877 38344 26911
rect 38292 26868 38344 26877
rect 41604 27004 41656 27056
rect 44640 27004 44692 27056
rect 40040 26936 40092 26988
rect 45468 26936 45520 26988
rect 41788 26868 41840 26920
rect 42248 26868 42300 26920
rect 48504 26911 48556 26920
rect 48504 26877 48513 26911
rect 48513 26877 48547 26911
rect 48547 26877 48556 26911
rect 48504 26868 48556 26877
rect 48780 26911 48832 26920
rect 48780 26877 48789 26911
rect 48789 26877 48823 26911
rect 48823 26877 48832 26911
rect 48780 26868 48832 26877
rect 36636 26800 36688 26852
rect 34888 26732 34940 26784
rect 38384 26732 38436 26784
rect 41052 26732 41104 26784
rect 46848 26775 46900 26784
rect 46848 26741 46857 26775
rect 46857 26741 46891 26775
rect 46891 26741 46900 26775
rect 46848 26732 46900 26741
rect 47676 26732 47728 26784
rect 2950 26630 3002 26682
rect 3014 26630 3066 26682
rect 3078 26630 3130 26682
rect 3142 26630 3194 26682
rect 3206 26630 3258 26682
rect 12950 26630 13002 26682
rect 13014 26630 13066 26682
rect 13078 26630 13130 26682
rect 13142 26630 13194 26682
rect 13206 26630 13258 26682
rect 22950 26630 23002 26682
rect 23014 26630 23066 26682
rect 23078 26630 23130 26682
rect 23142 26630 23194 26682
rect 23206 26630 23258 26682
rect 32950 26630 33002 26682
rect 33014 26630 33066 26682
rect 33078 26630 33130 26682
rect 33142 26630 33194 26682
rect 33206 26630 33258 26682
rect 42950 26630 43002 26682
rect 43014 26630 43066 26682
rect 43078 26630 43130 26682
rect 43142 26630 43194 26682
rect 43206 26630 43258 26682
rect 7748 26528 7800 26580
rect 9680 26571 9732 26580
rect 9680 26537 9689 26571
rect 9689 26537 9723 26571
rect 9723 26537 9732 26571
rect 9680 26528 9732 26537
rect 24400 26528 24452 26580
rect 25044 26528 25096 26580
rect 25228 26528 25280 26580
rect 29184 26528 29236 26580
rect 23572 26460 23624 26512
rect 23940 26460 23992 26512
rect 10876 26392 10928 26444
rect 24860 26392 24912 26444
rect 7748 26367 7800 26376
rect 7748 26333 7792 26367
rect 7792 26333 7800 26367
rect 7748 26324 7800 26333
rect 4988 26256 5040 26308
rect 5448 26256 5500 26308
rect 10968 26324 11020 26376
rect 23480 26324 23532 26376
rect 31024 26460 31076 26512
rect 25044 26435 25096 26444
rect 25044 26401 25053 26435
rect 25053 26401 25087 26435
rect 25087 26401 25096 26435
rect 25044 26392 25096 26401
rect 23664 26256 23716 26308
rect 26424 26392 26476 26444
rect 27712 26392 27764 26444
rect 28356 26392 28408 26444
rect 28816 26392 28868 26444
rect 30564 26392 30616 26444
rect 30656 26392 30708 26444
rect 32588 26528 32640 26580
rect 34428 26528 34480 26580
rect 33692 26460 33744 26512
rect 37096 26528 37148 26580
rect 40500 26528 40552 26580
rect 40960 26528 41012 26580
rect 48780 26528 48832 26580
rect 34704 26460 34756 26512
rect 31668 26392 31720 26444
rect 27620 26324 27672 26376
rect 28632 26324 28684 26376
rect 37464 26392 37516 26444
rect 37556 26392 37608 26444
rect 40040 26435 40092 26444
rect 40040 26401 40049 26435
rect 40049 26401 40083 26435
rect 40083 26401 40092 26435
rect 40040 26392 40092 26401
rect 48596 26460 48648 26512
rect 41788 26435 41840 26444
rect 41788 26401 41797 26435
rect 41797 26401 41831 26435
rect 41831 26401 41840 26435
rect 41788 26392 41840 26401
rect 43720 26392 43772 26444
rect 25412 26188 25464 26240
rect 25688 26188 25740 26240
rect 26424 26231 26476 26240
rect 26424 26197 26433 26231
rect 26433 26197 26467 26231
rect 26467 26197 26476 26231
rect 26424 26188 26476 26197
rect 28356 26256 28408 26308
rect 39580 26324 39632 26376
rect 43812 26324 43864 26376
rect 48504 26367 48556 26376
rect 48504 26333 48513 26367
rect 48513 26333 48547 26367
rect 48547 26333 48556 26367
rect 48504 26324 48556 26333
rect 32312 26256 32364 26308
rect 32404 26299 32456 26308
rect 32404 26265 32413 26299
rect 32413 26265 32447 26299
rect 32447 26265 32456 26299
rect 32404 26256 32456 26265
rect 34244 26256 34296 26308
rect 39488 26256 39540 26308
rect 41604 26256 41656 26308
rect 30656 26231 30708 26240
rect 30656 26197 30665 26231
rect 30665 26197 30699 26231
rect 30699 26197 30708 26231
rect 30656 26188 30708 26197
rect 34888 26188 34940 26240
rect 37740 26231 37792 26240
rect 37740 26197 37749 26231
rect 37749 26197 37783 26231
rect 37783 26197 37792 26231
rect 37740 26188 37792 26197
rect 47216 26231 47268 26240
rect 47216 26197 47225 26231
rect 47225 26197 47259 26231
rect 47259 26197 47268 26231
rect 47216 26188 47268 26197
rect 7950 26086 8002 26138
rect 8014 26086 8066 26138
rect 8078 26086 8130 26138
rect 8142 26086 8194 26138
rect 8206 26086 8258 26138
rect 17950 26086 18002 26138
rect 18014 26086 18066 26138
rect 18078 26086 18130 26138
rect 18142 26086 18194 26138
rect 18206 26086 18258 26138
rect 27950 26086 28002 26138
rect 28014 26086 28066 26138
rect 28078 26086 28130 26138
rect 28142 26086 28194 26138
rect 28206 26086 28258 26138
rect 37950 26086 38002 26138
rect 38014 26086 38066 26138
rect 38078 26086 38130 26138
rect 38142 26086 38194 26138
rect 38206 26086 38258 26138
rect 47950 26086 48002 26138
rect 48014 26086 48066 26138
rect 48078 26086 48130 26138
rect 48142 26086 48194 26138
rect 48206 26086 48258 26138
rect 24124 25984 24176 26036
rect 27804 25984 27856 26036
rect 28448 25984 28500 26036
rect 29552 25984 29604 26036
rect 32680 26027 32732 26036
rect 32680 25993 32689 26027
rect 32689 25993 32723 26027
rect 32723 25993 32732 26027
rect 32680 25984 32732 25993
rect 37740 25984 37792 26036
rect 7656 25891 7708 25900
rect 7656 25857 7665 25891
rect 7665 25857 7699 25891
rect 7699 25857 7708 25891
rect 7656 25848 7708 25857
rect 25688 25916 25740 25968
rect 30748 25916 30800 25968
rect 32956 25916 33008 25968
rect 33784 25916 33836 25968
rect 26424 25848 26476 25900
rect 27528 25848 27580 25900
rect 34336 25848 34388 25900
rect 37648 25916 37700 25968
rect 39948 25984 40000 26036
rect 40408 25984 40460 26036
rect 40776 25984 40828 26036
rect 38292 25916 38344 25968
rect 37556 25848 37608 25900
rect 9036 25780 9088 25832
rect 9496 25823 9548 25832
rect 9496 25789 9505 25823
rect 9505 25789 9539 25823
rect 9539 25789 9548 25823
rect 9496 25780 9548 25789
rect 22100 25780 22152 25832
rect 22376 25780 22428 25832
rect 24308 25823 24360 25832
rect 24308 25789 24317 25823
rect 24317 25789 24351 25823
rect 24351 25789 24360 25823
rect 24308 25780 24360 25789
rect 24400 25780 24452 25832
rect 28356 25823 28408 25832
rect 28356 25789 28365 25823
rect 28365 25789 28399 25823
rect 28399 25789 28408 25823
rect 28356 25780 28408 25789
rect 22652 25644 22704 25696
rect 28264 25712 28316 25764
rect 25688 25644 25740 25696
rect 25780 25644 25832 25696
rect 27344 25644 27396 25696
rect 27436 25644 27488 25696
rect 30288 25780 30340 25832
rect 32404 25780 32456 25832
rect 29828 25712 29880 25764
rect 33324 25780 33376 25832
rect 34704 25780 34756 25832
rect 35900 25780 35952 25832
rect 38476 25848 38528 25900
rect 39396 25848 39448 25900
rect 40684 25916 40736 25968
rect 41604 25916 41656 25968
rect 42800 25916 42852 25968
rect 37464 25712 37516 25764
rect 37556 25712 37608 25764
rect 39580 25823 39632 25832
rect 39580 25789 39589 25823
rect 39589 25789 39623 25823
rect 39623 25789 39632 25823
rect 39580 25780 39632 25789
rect 39672 25780 39724 25832
rect 46020 25891 46072 25900
rect 46020 25857 46029 25891
rect 46029 25857 46063 25891
rect 46063 25857 46072 25891
rect 46020 25848 46072 25857
rect 49332 25891 49384 25900
rect 49332 25857 49341 25891
rect 49341 25857 49375 25891
rect 49375 25857 49384 25891
rect 49332 25848 49384 25857
rect 46204 25755 46256 25764
rect 46204 25721 46213 25755
rect 46213 25721 46247 25755
rect 46247 25721 46256 25755
rect 46204 25712 46256 25721
rect 46940 25755 46992 25764
rect 46940 25721 46949 25755
rect 46949 25721 46983 25755
rect 46983 25721 46992 25755
rect 46940 25712 46992 25721
rect 29920 25644 29972 25696
rect 30932 25687 30984 25696
rect 30932 25653 30941 25687
rect 30941 25653 30975 25687
rect 30975 25653 30984 25687
rect 30932 25644 30984 25653
rect 35992 25644 36044 25696
rect 36912 25687 36964 25696
rect 36912 25653 36921 25687
rect 36921 25653 36955 25687
rect 36955 25653 36964 25687
rect 36912 25644 36964 25653
rect 37740 25644 37792 25696
rect 49148 25687 49200 25696
rect 49148 25653 49157 25687
rect 49157 25653 49191 25687
rect 49191 25653 49200 25687
rect 49148 25644 49200 25653
rect 2950 25542 3002 25594
rect 3014 25542 3066 25594
rect 3078 25542 3130 25594
rect 3142 25542 3194 25594
rect 3206 25542 3258 25594
rect 12950 25542 13002 25594
rect 13014 25542 13066 25594
rect 13078 25542 13130 25594
rect 13142 25542 13194 25594
rect 13206 25542 13258 25594
rect 22950 25542 23002 25594
rect 23014 25542 23066 25594
rect 23078 25542 23130 25594
rect 23142 25542 23194 25594
rect 23206 25542 23258 25594
rect 32950 25542 33002 25594
rect 33014 25542 33066 25594
rect 33078 25542 33130 25594
rect 33142 25542 33194 25594
rect 33206 25542 33258 25594
rect 42950 25542 43002 25594
rect 43014 25542 43066 25594
rect 43078 25542 43130 25594
rect 43142 25542 43194 25594
rect 43206 25542 43258 25594
rect 4896 25483 4948 25492
rect 4896 25449 4905 25483
rect 4905 25449 4939 25483
rect 4939 25449 4948 25483
rect 4896 25440 4948 25449
rect 1308 25304 1360 25356
rect 10968 25440 11020 25492
rect 24308 25440 24360 25492
rect 25136 25440 25188 25492
rect 30012 25440 30064 25492
rect 34244 25440 34296 25492
rect 35348 25440 35400 25492
rect 37832 25440 37884 25492
rect 10876 25372 10928 25424
rect 27252 25372 27304 25424
rect 12348 25304 12400 25356
rect 24308 25304 24360 25356
rect 25688 25304 25740 25356
rect 27528 25304 27580 25356
rect 31668 25372 31720 25424
rect 30012 25304 30064 25356
rect 31852 25304 31904 25356
rect 4160 25236 4212 25288
rect 6276 25236 6328 25288
rect 10600 25279 10652 25288
rect 10600 25245 10609 25279
rect 10609 25245 10643 25279
rect 10643 25245 10652 25279
rect 10600 25236 10652 25245
rect 16488 25236 16540 25288
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 28264 25236 28316 25288
rect 29000 25236 29052 25288
rect 29092 25236 29144 25288
rect 31760 25236 31812 25288
rect 31944 25236 31996 25288
rect 37372 25372 37424 25424
rect 39488 25483 39540 25492
rect 39488 25449 39497 25483
rect 39497 25449 39531 25483
rect 39531 25449 39540 25483
rect 39488 25440 39540 25449
rect 49148 25372 49200 25424
rect 33968 25347 34020 25356
rect 33968 25313 33977 25347
rect 33977 25313 34011 25347
rect 34011 25313 34020 25347
rect 33968 25304 34020 25313
rect 34060 25347 34112 25356
rect 34060 25313 34069 25347
rect 34069 25313 34103 25347
rect 34103 25313 34112 25347
rect 34060 25304 34112 25313
rect 35624 25304 35676 25356
rect 35992 25304 36044 25356
rect 38568 25304 38620 25356
rect 40500 25347 40552 25356
rect 40500 25313 40509 25347
rect 40509 25313 40543 25347
rect 40543 25313 40552 25347
rect 40500 25304 40552 25313
rect 40684 25347 40736 25356
rect 40684 25313 40693 25347
rect 40693 25313 40727 25347
rect 40727 25313 40736 25347
rect 40684 25304 40736 25313
rect 34888 25236 34940 25288
rect 43444 25236 43496 25288
rect 45560 25236 45612 25288
rect 25412 25168 25464 25220
rect 22284 25143 22336 25152
rect 22284 25109 22293 25143
rect 22293 25109 22327 25143
rect 22327 25109 22336 25143
rect 22284 25100 22336 25109
rect 23296 25100 23348 25152
rect 26148 25100 26200 25152
rect 26700 25168 26752 25220
rect 27620 25100 27672 25152
rect 32220 25168 32272 25220
rect 34520 25168 34572 25220
rect 34796 25168 34848 25220
rect 29000 25100 29052 25152
rect 31300 25100 31352 25152
rect 32772 25100 32824 25152
rect 35164 25143 35216 25152
rect 35164 25109 35173 25143
rect 35173 25109 35207 25143
rect 35207 25109 35216 25143
rect 35164 25100 35216 25109
rect 36544 25143 36596 25152
rect 36544 25109 36553 25143
rect 36553 25109 36587 25143
rect 36587 25109 36596 25143
rect 36544 25100 36596 25109
rect 36912 25211 36964 25220
rect 36912 25177 36921 25211
rect 36921 25177 36955 25211
rect 36955 25177 36964 25211
rect 36912 25168 36964 25177
rect 39672 25168 39724 25220
rect 44364 25211 44416 25220
rect 44364 25177 44373 25211
rect 44373 25177 44407 25211
rect 44407 25177 44416 25211
rect 44364 25168 44416 25177
rect 45468 25211 45520 25220
rect 45468 25177 45477 25211
rect 45477 25177 45511 25211
rect 45511 25177 45520 25211
rect 45468 25168 45520 25177
rect 47492 25168 47544 25220
rect 38752 25100 38804 25152
rect 40040 25143 40092 25152
rect 40040 25109 40049 25143
rect 40049 25109 40083 25143
rect 40083 25109 40092 25143
rect 40040 25100 40092 25109
rect 40408 25143 40460 25152
rect 40408 25109 40417 25143
rect 40417 25109 40451 25143
rect 40451 25109 40460 25143
rect 40408 25100 40460 25109
rect 44456 25143 44508 25152
rect 44456 25109 44465 25143
rect 44465 25109 44499 25143
rect 44499 25109 44508 25143
rect 44456 25100 44508 25109
rect 7950 24998 8002 25050
rect 8014 24998 8066 25050
rect 8078 24998 8130 25050
rect 8142 24998 8194 25050
rect 8206 24998 8258 25050
rect 17950 24998 18002 25050
rect 18014 24998 18066 25050
rect 18078 24998 18130 25050
rect 18142 24998 18194 25050
rect 18206 24998 18258 25050
rect 27950 24998 28002 25050
rect 28014 24998 28066 25050
rect 28078 24998 28130 25050
rect 28142 24998 28194 25050
rect 28206 24998 28258 25050
rect 37950 24998 38002 25050
rect 38014 24998 38066 25050
rect 38078 24998 38130 25050
rect 38142 24998 38194 25050
rect 38206 24998 38258 25050
rect 47950 24998 48002 25050
rect 48014 24998 48066 25050
rect 48078 24998 48130 25050
rect 48142 24998 48194 25050
rect 48206 24998 48258 25050
rect 25780 24939 25832 24948
rect 25780 24905 25789 24939
rect 25789 24905 25823 24939
rect 25823 24905 25832 24939
rect 25780 24896 25832 24905
rect 20996 24828 21048 24880
rect 9312 24760 9364 24812
rect 8300 24692 8352 24744
rect 19708 24735 19760 24744
rect 19708 24701 19717 24735
rect 19717 24701 19751 24735
rect 19751 24701 19760 24735
rect 19708 24692 19760 24701
rect 21272 24692 21324 24744
rect 25320 24692 25372 24744
rect 25596 24692 25648 24744
rect 27436 24896 27488 24948
rect 27620 24896 27672 24948
rect 28908 24939 28960 24948
rect 28908 24905 28917 24939
rect 28917 24905 28951 24939
rect 28951 24905 28960 24939
rect 28908 24896 28960 24905
rect 30932 24896 30984 24948
rect 27528 24828 27580 24880
rect 27712 24828 27764 24880
rect 29920 24828 29972 24880
rect 32220 24828 32272 24880
rect 35992 24896 36044 24948
rect 36544 24896 36596 24948
rect 34244 24871 34296 24880
rect 34244 24837 34253 24871
rect 34253 24837 34287 24871
rect 34287 24837 34296 24871
rect 34244 24828 34296 24837
rect 37464 24828 37516 24880
rect 38476 24828 38528 24880
rect 30748 24760 30800 24812
rect 32864 24803 32916 24812
rect 32864 24769 32873 24803
rect 32873 24769 32907 24803
rect 32907 24769 32916 24803
rect 32864 24760 32916 24769
rect 33876 24760 33928 24812
rect 35348 24760 35400 24812
rect 37188 24760 37240 24812
rect 40408 24760 40460 24812
rect 47216 24760 47268 24812
rect 27436 24735 27488 24744
rect 27436 24701 27445 24735
rect 27445 24701 27479 24735
rect 27479 24701 27488 24735
rect 27436 24692 27488 24701
rect 27528 24692 27580 24744
rect 28172 24692 28224 24744
rect 30104 24692 30156 24744
rect 21732 24624 21784 24676
rect 21916 24624 21968 24676
rect 26884 24624 26936 24676
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 32588 24692 32640 24744
rect 33324 24692 33376 24744
rect 39488 24692 39540 24744
rect 49148 24735 49200 24744
rect 49148 24701 49157 24735
rect 49157 24701 49191 24735
rect 49191 24701 49200 24735
rect 49148 24692 49200 24701
rect 31576 24624 31628 24676
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 29000 24556 29052 24608
rect 32404 24599 32456 24608
rect 32404 24565 32413 24599
rect 32413 24565 32447 24599
rect 32447 24565 32456 24599
rect 32404 24556 32456 24565
rect 33876 24556 33928 24608
rect 34888 24556 34940 24608
rect 34980 24556 35032 24608
rect 2950 24454 3002 24506
rect 3014 24454 3066 24506
rect 3078 24454 3130 24506
rect 3142 24454 3194 24506
rect 3206 24454 3258 24506
rect 12950 24454 13002 24506
rect 13014 24454 13066 24506
rect 13078 24454 13130 24506
rect 13142 24454 13194 24506
rect 13206 24454 13258 24506
rect 22950 24454 23002 24506
rect 23014 24454 23066 24506
rect 23078 24454 23130 24506
rect 23142 24454 23194 24506
rect 23206 24454 23258 24506
rect 32950 24454 33002 24506
rect 33014 24454 33066 24506
rect 33078 24454 33130 24506
rect 33142 24454 33194 24506
rect 33206 24454 33258 24506
rect 42950 24454 43002 24506
rect 43014 24454 43066 24506
rect 43078 24454 43130 24506
rect 43142 24454 43194 24506
rect 43206 24454 43258 24506
rect 12348 24352 12400 24404
rect 14556 24284 14608 24336
rect 15292 24216 15344 24268
rect 10600 24191 10652 24200
rect 10600 24157 10609 24191
rect 10609 24157 10643 24191
rect 10643 24157 10652 24191
rect 10600 24148 10652 24157
rect 12532 24148 12584 24200
rect 15200 24080 15252 24132
rect 15384 24080 15436 24132
rect 7840 24012 7892 24064
rect 11152 24012 11204 24064
rect 25504 24352 25556 24404
rect 28448 24352 28500 24404
rect 28908 24352 28960 24404
rect 19708 24216 19760 24268
rect 21824 24216 21876 24268
rect 22836 24216 22888 24268
rect 26884 24259 26936 24268
rect 26884 24225 26893 24259
rect 26893 24225 26927 24259
rect 26927 24225 26936 24259
rect 26884 24216 26936 24225
rect 27436 24216 27488 24268
rect 28080 24216 28132 24268
rect 25504 24191 25556 24200
rect 25504 24157 25513 24191
rect 25513 24157 25547 24191
rect 25547 24157 25556 24191
rect 25504 24148 25556 24157
rect 29092 24284 29144 24336
rect 28356 24216 28408 24268
rect 28724 24216 28776 24268
rect 21364 24080 21416 24132
rect 23480 24080 23532 24132
rect 28448 24148 28500 24200
rect 29552 24216 29604 24268
rect 30196 24259 30248 24268
rect 30196 24225 30205 24259
rect 30205 24225 30239 24259
rect 30239 24225 30248 24259
rect 30196 24216 30248 24225
rect 32220 24284 32272 24336
rect 33692 24284 33744 24336
rect 36636 24352 36688 24404
rect 34520 24216 34572 24268
rect 32864 24148 32916 24200
rect 33784 24148 33836 24200
rect 34336 24148 34388 24200
rect 21272 24012 21324 24064
rect 22560 24055 22612 24064
rect 22560 24021 22569 24055
rect 22569 24021 22603 24055
rect 22603 24021 22612 24055
rect 22560 24012 22612 24021
rect 23848 24012 23900 24064
rect 26240 24012 26292 24064
rect 26792 24055 26844 24064
rect 26792 24021 26801 24055
rect 26801 24021 26835 24055
rect 26835 24021 26844 24055
rect 26792 24012 26844 24021
rect 27804 24012 27856 24064
rect 29828 24080 29880 24132
rect 30840 24080 30892 24132
rect 35348 24216 35400 24268
rect 34888 24148 34940 24200
rect 37280 24216 37332 24268
rect 40316 24216 40368 24268
rect 40776 24216 40828 24268
rect 37832 24148 37884 24200
rect 40040 24148 40092 24200
rect 47860 24148 47912 24200
rect 35532 24080 35584 24132
rect 36268 24080 36320 24132
rect 49148 24123 49200 24132
rect 49148 24089 49157 24123
rect 49157 24089 49191 24123
rect 49191 24089 49200 24123
rect 49148 24080 49200 24089
rect 33876 24012 33928 24064
rect 34336 24012 34388 24064
rect 35348 24012 35400 24064
rect 35624 24012 35676 24064
rect 37372 24012 37424 24064
rect 37832 24012 37884 24064
rect 39212 24012 39264 24064
rect 40040 24055 40092 24064
rect 40040 24021 40049 24055
rect 40049 24021 40083 24055
rect 40083 24021 40092 24055
rect 40040 24012 40092 24021
rect 7950 23910 8002 23962
rect 8014 23910 8066 23962
rect 8078 23910 8130 23962
rect 8142 23910 8194 23962
rect 8206 23910 8258 23962
rect 17950 23910 18002 23962
rect 18014 23910 18066 23962
rect 18078 23910 18130 23962
rect 18142 23910 18194 23962
rect 18206 23910 18258 23962
rect 27950 23910 28002 23962
rect 28014 23910 28066 23962
rect 28078 23910 28130 23962
rect 28142 23910 28194 23962
rect 28206 23910 28258 23962
rect 37950 23910 38002 23962
rect 38014 23910 38066 23962
rect 38078 23910 38130 23962
rect 38142 23910 38194 23962
rect 38206 23910 38258 23962
rect 47950 23910 48002 23962
rect 48014 23910 48066 23962
rect 48078 23910 48130 23962
rect 48142 23910 48194 23962
rect 48206 23910 48258 23962
rect 6276 23808 6328 23860
rect 15292 23808 15344 23860
rect 16488 23808 16540 23860
rect 23296 23808 23348 23860
rect 30840 23808 30892 23860
rect 32588 23808 32640 23860
rect 34520 23808 34572 23860
rect 38200 23808 38252 23860
rect 38568 23808 38620 23860
rect 12256 23672 12308 23724
rect 15384 23740 15436 23792
rect 7840 23604 7892 23656
rect 12348 23604 12400 23656
rect 14556 23604 14608 23656
rect 21456 23740 21508 23792
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 26792 23740 26844 23792
rect 21180 23647 21232 23656
rect 21180 23613 21189 23647
rect 21189 23613 21223 23647
rect 21223 23613 21232 23647
rect 21180 23604 21232 23613
rect 21272 23647 21324 23656
rect 21272 23613 21281 23647
rect 21281 23613 21315 23647
rect 21315 23613 21324 23647
rect 21272 23604 21324 23613
rect 23480 23604 23532 23656
rect 23664 23604 23716 23656
rect 24676 23604 24728 23656
rect 23388 23536 23440 23588
rect 27068 23604 27120 23656
rect 26700 23536 26752 23588
rect 27896 23536 27948 23588
rect 28908 23672 28960 23724
rect 29276 23740 29328 23792
rect 31484 23740 31536 23792
rect 33876 23740 33928 23792
rect 37280 23740 37332 23792
rect 39672 23740 39724 23792
rect 33692 23672 33744 23724
rect 30104 23604 30156 23656
rect 32312 23647 32364 23656
rect 32312 23613 32321 23647
rect 32321 23613 32355 23647
rect 32355 23613 32364 23647
rect 32312 23604 32364 23613
rect 32680 23604 32732 23656
rect 38292 23672 38344 23724
rect 38568 23672 38620 23724
rect 46848 23672 46900 23724
rect 35256 23604 35308 23656
rect 35532 23604 35584 23656
rect 39488 23604 39540 23656
rect 47492 23604 47544 23656
rect 47860 23604 47912 23656
rect 49148 23647 49200 23656
rect 49148 23613 49157 23647
rect 49157 23613 49191 23647
rect 49191 23613 49200 23647
rect 49148 23604 49200 23613
rect 22100 23468 22152 23520
rect 24952 23468 25004 23520
rect 25872 23511 25924 23520
rect 25872 23477 25881 23511
rect 25881 23477 25915 23511
rect 25915 23477 25924 23511
rect 25872 23468 25924 23477
rect 26148 23468 26200 23520
rect 28908 23536 28960 23588
rect 31484 23536 31536 23588
rect 32036 23536 32088 23588
rect 34060 23579 34112 23588
rect 34060 23545 34069 23579
rect 34069 23545 34103 23579
rect 34103 23545 34112 23579
rect 34060 23536 34112 23545
rect 32220 23468 32272 23520
rect 34152 23468 34204 23520
rect 34520 23511 34572 23520
rect 34520 23477 34529 23511
rect 34529 23477 34563 23511
rect 34563 23477 34572 23511
rect 34520 23468 34572 23477
rect 38752 23468 38804 23520
rect 39580 23468 39632 23520
rect 2950 23366 3002 23418
rect 3014 23366 3066 23418
rect 3078 23366 3130 23418
rect 3142 23366 3194 23418
rect 3206 23366 3258 23418
rect 12950 23366 13002 23418
rect 13014 23366 13066 23418
rect 13078 23366 13130 23418
rect 13142 23366 13194 23418
rect 13206 23366 13258 23418
rect 22950 23366 23002 23418
rect 23014 23366 23066 23418
rect 23078 23366 23130 23418
rect 23142 23366 23194 23418
rect 23206 23366 23258 23418
rect 32950 23366 33002 23418
rect 33014 23366 33066 23418
rect 33078 23366 33130 23418
rect 33142 23366 33194 23418
rect 33206 23366 33258 23418
rect 42950 23366 43002 23418
rect 43014 23366 43066 23418
rect 43078 23366 43130 23418
rect 43142 23366 43194 23418
rect 43206 23366 43258 23418
rect 4160 23264 4212 23316
rect 22192 23264 22244 23316
rect 22744 23264 22796 23316
rect 1308 23128 1360 23180
rect 5540 23128 5592 23180
rect 9036 23128 9088 23180
rect 15292 23128 15344 23180
rect 19708 23128 19760 23180
rect 27436 23264 27488 23316
rect 28724 23264 28776 23316
rect 31116 23264 31168 23316
rect 31852 23307 31904 23316
rect 31852 23273 31861 23307
rect 31861 23273 31895 23307
rect 31895 23273 31904 23307
rect 31852 23264 31904 23273
rect 34152 23264 34204 23316
rect 34244 23264 34296 23316
rect 41236 23264 41288 23316
rect 23664 23171 23716 23180
rect 23664 23137 23673 23171
rect 23673 23137 23707 23171
rect 23707 23137 23716 23171
rect 23664 23128 23716 23137
rect 27528 23128 27580 23180
rect 27896 23128 27948 23180
rect 30104 23171 30156 23180
rect 30104 23137 30113 23171
rect 30113 23137 30147 23171
rect 30147 23137 30156 23171
rect 30104 23128 30156 23137
rect 32128 23196 32180 23248
rect 31576 23128 31628 23180
rect 4988 23060 5040 23112
rect 9772 23060 9824 23112
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 24952 23103 25004 23112
rect 24952 23069 24961 23103
rect 24961 23069 24995 23103
rect 24995 23069 25004 23103
rect 24952 23060 25004 23069
rect 28540 23060 28592 23112
rect 32312 23171 32364 23180
rect 32312 23137 32321 23171
rect 32321 23137 32355 23171
rect 32355 23137 32364 23171
rect 32312 23128 32364 23137
rect 38384 23196 38436 23248
rect 37464 23128 37516 23180
rect 38752 23171 38804 23180
rect 38752 23137 38761 23171
rect 38761 23137 38795 23171
rect 38795 23137 38804 23171
rect 38752 23128 38804 23137
rect 33692 23060 33744 23112
rect 34428 23060 34480 23112
rect 9680 22992 9732 23044
rect 17408 23035 17460 23044
rect 17408 23001 17417 23035
rect 17417 23001 17451 23035
rect 17451 23001 17460 23035
rect 17408 22992 17460 23001
rect 2780 22924 2832 22976
rect 15384 22924 15436 22976
rect 18880 22967 18932 22976
rect 18880 22933 18889 22967
rect 18889 22933 18923 22967
rect 18923 22933 18932 22967
rect 18880 22924 18932 22933
rect 19984 22992 20036 23044
rect 20996 22992 21048 23044
rect 23664 22992 23716 23044
rect 21272 22924 21324 22976
rect 22652 22924 22704 22976
rect 24584 22967 24636 22976
rect 24584 22933 24593 22967
rect 24593 22933 24627 22967
rect 24627 22933 24636 22967
rect 24584 22924 24636 22933
rect 25044 22967 25096 22976
rect 25044 22933 25053 22967
rect 25053 22933 25087 22967
rect 25087 22933 25096 22967
rect 25044 22924 25096 22933
rect 27528 22992 27580 23044
rect 27896 22992 27948 23044
rect 31760 22992 31812 23044
rect 29184 22924 29236 22976
rect 29460 22924 29512 22976
rect 30656 22924 30708 22976
rect 35256 22992 35308 23044
rect 36176 22992 36228 23044
rect 47676 23060 47728 23112
rect 37372 22992 37424 23044
rect 46664 22992 46716 23044
rect 49148 23035 49200 23044
rect 49148 23001 49157 23035
rect 49157 23001 49191 23035
rect 49191 23001 49200 23035
rect 49148 22992 49200 23001
rect 37188 22924 37240 22976
rect 37832 22924 37884 22976
rect 38292 22924 38344 22976
rect 7950 22822 8002 22874
rect 8014 22822 8066 22874
rect 8078 22822 8130 22874
rect 8142 22822 8194 22874
rect 8206 22822 8258 22874
rect 17950 22822 18002 22874
rect 18014 22822 18066 22874
rect 18078 22822 18130 22874
rect 18142 22822 18194 22874
rect 18206 22822 18258 22874
rect 27950 22822 28002 22874
rect 28014 22822 28066 22874
rect 28078 22822 28130 22874
rect 28142 22822 28194 22874
rect 28206 22822 28258 22874
rect 37950 22822 38002 22874
rect 38014 22822 38066 22874
rect 38078 22822 38130 22874
rect 38142 22822 38194 22874
rect 38206 22822 38258 22874
rect 47950 22822 48002 22874
rect 48014 22822 48066 22874
rect 48078 22822 48130 22874
rect 48142 22822 48194 22874
rect 48206 22822 48258 22874
rect 22284 22720 22336 22772
rect 23664 22763 23716 22772
rect 23664 22729 23673 22763
rect 23673 22729 23707 22763
rect 23707 22729 23716 22763
rect 23664 22720 23716 22729
rect 24584 22720 24636 22772
rect 30472 22720 30524 22772
rect 32680 22720 32732 22772
rect 34520 22720 34572 22772
rect 17408 22652 17460 22704
rect 15200 22584 15252 22636
rect 18880 22584 18932 22636
rect 19800 22559 19852 22568
rect 19800 22525 19809 22559
rect 19809 22525 19843 22559
rect 19843 22525 19852 22559
rect 19800 22516 19852 22525
rect 21916 22652 21968 22704
rect 23756 22695 23808 22704
rect 23756 22661 23765 22695
rect 23765 22661 23799 22695
rect 23799 22661 23808 22695
rect 23756 22652 23808 22661
rect 26332 22652 26384 22704
rect 27436 22695 27488 22704
rect 27436 22661 27445 22695
rect 27445 22661 27479 22695
rect 27479 22661 27488 22695
rect 27436 22652 27488 22661
rect 30380 22652 30432 22704
rect 23296 22584 23348 22636
rect 28540 22584 28592 22636
rect 35164 22652 35216 22704
rect 37188 22584 37240 22636
rect 37464 22584 37516 22636
rect 38568 22720 38620 22772
rect 37832 22652 37884 22704
rect 39672 22720 39724 22772
rect 39028 22584 39080 22636
rect 21272 22559 21324 22568
rect 21272 22525 21281 22559
rect 21281 22525 21315 22559
rect 21315 22525 21324 22559
rect 21272 22516 21324 22525
rect 17408 22423 17460 22432
rect 17408 22389 17417 22423
rect 17417 22389 17451 22423
rect 17451 22389 17460 22423
rect 17408 22380 17460 22389
rect 21640 22380 21692 22432
rect 23388 22380 23440 22432
rect 25136 22559 25188 22568
rect 25136 22525 25145 22559
rect 25145 22525 25179 22559
rect 25179 22525 25188 22559
rect 25136 22516 25188 22525
rect 26516 22448 26568 22500
rect 25044 22380 25096 22432
rect 26608 22380 26660 22432
rect 27528 22516 27580 22568
rect 32588 22516 32640 22568
rect 34244 22559 34296 22568
rect 34244 22525 34253 22559
rect 34253 22525 34287 22559
rect 34287 22525 34296 22559
rect 34244 22516 34296 22525
rect 39488 22516 39540 22568
rect 34520 22448 34572 22500
rect 27804 22380 27856 22432
rect 32312 22380 32364 22432
rect 2950 22278 3002 22330
rect 3014 22278 3066 22330
rect 3078 22278 3130 22330
rect 3142 22278 3194 22330
rect 3206 22278 3258 22330
rect 12950 22278 13002 22330
rect 13014 22278 13066 22330
rect 13078 22278 13130 22330
rect 13142 22278 13194 22330
rect 13206 22278 13258 22330
rect 22950 22278 23002 22330
rect 23014 22278 23066 22330
rect 23078 22278 23130 22330
rect 23142 22278 23194 22330
rect 23206 22278 23258 22330
rect 32950 22278 33002 22330
rect 33014 22278 33066 22330
rect 33078 22278 33130 22330
rect 33142 22278 33194 22330
rect 33206 22278 33258 22330
rect 42950 22278 43002 22330
rect 43014 22278 43066 22330
rect 43078 22278 43130 22330
rect 43142 22278 43194 22330
rect 43206 22278 43258 22330
rect 14740 22176 14792 22228
rect 5540 22151 5592 22160
rect 5540 22117 5549 22151
rect 5549 22117 5583 22151
rect 5583 22117 5592 22151
rect 5540 22108 5592 22117
rect 14556 22108 14608 22160
rect 15108 22176 15160 22228
rect 16488 22219 16540 22228
rect 16488 22185 16497 22219
rect 16497 22185 16531 22219
rect 16531 22185 16540 22219
rect 16488 22176 16540 22185
rect 22560 22108 22612 22160
rect 23296 22219 23348 22228
rect 23296 22185 23305 22219
rect 23305 22185 23339 22219
rect 23339 22185 23348 22219
rect 23296 22176 23348 22185
rect 19432 22083 19484 22092
rect 19432 22049 19441 22083
rect 19441 22049 19475 22083
rect 19475 22049 19484 22083
rect 19432 22040 19484 22049
rect 20168 22040 20220 22092
rect 23572 22108 23624 22160
rect 23296 22040 23348 22092
rect 23480 22040 23532 22092
rect 9128 21972 9180 22024
rect 10232 21904 10284 21956
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 13636 22015 13688 22024
rect 13636 21981 13645 22015
rect 13645 21981 13679 22015
rect 13679 21981 13688 22015
rect 13636 21972 13688 21981
rect 20996 21972 21048 22024
rect 24308 22040 24360 22092
rect 32128 22176 32180 22228
rect 33416 22176 33468 22228
rect 34244 22176 34296 22228
rect 26608 22108 26660 22160
rect 9312 21836 9364 21888
rect 13452 21879 13504 21888
rect 13452 21845 13461 21879
rect 13461 21845 13495 21879
rect 13495 21845 13504 21879
rect 13452 21836 13504 21845
rect 15476 21904 15528 21956
rect 25964 22015 26016 22024
rect 25964 21981 25973 22015
rect 25973 21981 26007 22015
rect 26007 21981 26016 22015
rect 25964 21972 26016 21981
rect 28540 22040 28592 22092
rect 34336 22108 34388 22160
rect 23848 21904 23900 21956
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 22100 21836 22152 21845
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 23572 21836 23624 21888
rect 26700 21904 26752 21956
rect 25596 21879 25648 21888
rect 25596 21845 25605 21879
rect 25605 21845 25639 21879
rect 25639 21845 25648 21879
rect 25596 21836 25648 21845
rect 27528 21836 27580 21888
rect 28816 21879 28868 21888
rect 28816 21845 28825 21879
rect 28825 21845 28859 21879
rect 28859 21845 28868 21879
rect 28816 21836 28868 21845
rect 29368 21972 29420 22024
rect 33876 22040 33928 22092
rect 37280 22040 37332 22092
rect 32496 21972 32548 22024
rect 36084 21904 36136 21956
rect 47584 21972 47636 22024
rect 49148 22015 49200 22024
rect 49148 21981 49157 22015
rect 49157 21981 49191 22015
rect 49191 21981 49200 22015
rect 49148 21972 49200 21981
rect 31668 21836 31720 21888
rect 38476 21904 38528 21956
rect 43812 21904 43864 21956
rect 41328 21836 41380 21888
rect 7950 21734 8002 21786
rect 8014 21734 8066 21786
rect 8078 21734 8130 21786
rect 8142 21734 8194 21786
rect 8206 21734 8258 21786
rect 17950 21734 18002 21786
rect 18014 21734 18066 21786
rect 18078 21734 18130 21786
rect 18142 21734 18194 21786
rect 18206 21734 18258 21786
rect 27950 21734 28002 21786
rect 28014 21734 28066 21786
rect 28078 21734 28130 21786
rect 28142 21734 28194 21786
rect 28206 21734 28258 21786
rect 37950 21734 38002 21786
rect 38014 21734 38066 21786
rect 38078 21734 38130 21786
rect 38142 21734 38194 21786
rect 38206 21734 38258 21786
rect 47950 21734 48002 21786
rect 48014 21734 48066 21786
rect 48078 21734 48130 21786
rect 48142 21734 48194 21786
rect 48206 21734 48258 21786
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 13636 21632 13688 21684
rect 17408 21632 17460 21684
rect 19800 21632 19852 21684
rect 21180 21632 21232 21684
rect 22468 21632 22520 21684
rect 25872 21632 25924 21684
rect 29368 21632 29420 21684
rect 21732 21564 21784 21616
rect 22100 21564 22152 21616
rect 22836 21564 22888 21616
rect 23296 21564 23348 21616
rect 25596 21564 25648 21616
rect 13452 21496 13504 21548
rect 16488 21496 16540 21548
rect 19524 21496 19576 21548
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 22376 21496 22428 21548
rect 28172 21539 28224 21548
rect 28172 21505 28181 21539
rect 28181 21505 28215 21539
rect 28215 21505 28224 21539
rect 28172 21496 28224 21505
rect 32496 21632 32548 21684
rect 34244 21675 34296 21684
rect 34244 21641 34253 21675
rect 34253 21641 34287 21675
rect 34287 21641 34296 21675
rect 34244 21632 34296 21641
rect 37832 21632 37884 21684
rect 31576 21564 31628 21616
rect 34428 21564 34480 21616
rect 36084 21564 36136 21616
rect 38752 21607 38804 21616
rect 38752 21573 38761 21607
rect 38761 21573 38795 21607
rect 38795 21573 38804 21607
rect 38752 21564 38804 21573
rect 39028 21564 39080 21616
rect 43812 21607 43864 21616
rect 43812 21573 43821 21607
rect 43821 21573 43855 21607
rect 43855 21573 43864 21607
rect 43812 21564 43864 21573
rect 9772 21471 9824 21480
rect 9772 21437 9781 21471
rect 9781 21437 9815 21471
rect 9815 21437 9824 21471
rect 9772 21428 9824 21437
rect 19892 21471 19944 21480
rect 19892 21437 19901 21471
rect 19901 21437 19935 21471
rect 19935 21437 19944 21471
rect 19892 21428 19944 21437
rect 19984 21428 20036 21480
rect 12256 21360 12308 21412
rect 21364 21471 21416 21480
rect 21364 21437 21373 21471
rect 21373 21437 21407 21471
rect 21407 21437 21416 21471
rect 21364 21428 21416 21437
rect 22468 21471 22520 21480
rect 22468 21437 22477 21471
rect 22477 21437 22511 21471
rect 22511 21437 22520 21471
rect 22468 21428 22520 21437
rect 25688 21471 25740 21480
rect 25688 21437 25697 21471
rect 25697 21437 25731 21471
rect 25731 21437 25740 21471
rect 25688 21428 25740 21437
rect 27804 21428 27856 21480
rect 31852 21496 31904 21548
rect 32496 21539 32548 21548
rect 32496 21505 32505 21539
rect 32505 21505 32539 21539
rect 32539 21505 32548 21539
rect 32496 21496 32548 21505
rect 35348 21539 35400 21548
rect 35348 21505 35357 21539
rect 35357 21505 35391 21539
rect 35391 21505 35400 21539
rect 35348 21496 35400 21505
rect 35992 21539 36044 21548
rect 35992 21505 36001 21539
rect 36001 21505 36035 21539
rect 36035 21505 36044 21539
rect 35992 21496 36044 21505
rect 38476 21539 38528 21548
rect 38476 21505 38485 21539
rect 38485 21505 38519 21539
rect 38519 21505 38528 21539
rect 38476 21496 38528 21505
rect 46204 21496 46256 21548
rect 31760 21428 31812 21480
rect 32220 21428 32272 21480
rect 34060 21428 34112 21480
rect 49148 21471 49200 21480
rect 49148 21437 49157 21471
rect 49157 21437 49191 21471
rect 49191 21437 49200 21471
rect 49148 21428 49200 21437
rect 27436 21360 27488 21412
rect 28908 21360 28960 21412
rect 45100 21360 45152 21412
rect 24308 21292 24360 21344
rect 30656 21292 30708 21344
rect 33508 21292 33560 21344
rect 35440 21292 35492 21344
rect 37096 21292 37148 21344
rect 38568 21292 38620 21344
rect 2950 21190 3002 21242
rect 3014 21190 3066 21242
rect 3078 21190 3130 21242
rect 3142 21190 3194 21242
rect 3206 21190 3258 21242
rect 12950 21190 13002 21242
rect 13014 21190 13066 21242
rect 13078 21190 13130 21242
rect 13142 21190 13194 21242
rect 13206 21190 13258 21242
rect 22950 21190 23002 21242
rect 23014 21190 23066 21242
rect 23078 21190 23130 21242
rect 23142 21190 23194 21242
rect 23206 21190 23258 21242
rect 32950 21190 33002 21242
rect 33014 21190 33066 21242
rect 33078 21190 33130 21242
rect 33142 21190 33194 21242
rect 33206 21190 33258 21242
rect 42950 21190 43002 21242
rect 43014 21190 43066 21242
rect 43078 21190 43130 21242
rect 43142 21190 43194 21242
rect 43206 21190 43258 21242
rect 9680 21131 9732 21140
rect 9680 21097 9689 21131
rect 9689 21097 9723 21131
rect 9723 21097 9732 21131
rect 9680 21088 9732 21097
rect 28172 21088 28224 21140
rect 30748 21088 30800 21140
rect 27344 21020 27396 21072
rect 35348 21020 35400 21072
rect 43720 21020 43772 21072
rect 10968 20952 11020 21004
rect 31760 20952 31812 21004
rect 32864 20952 32916 21004
rect 7840 20884 7892 20936
rect 9312 20927 9364 20936
rect 9312 20893 9321 20927
rect 9321 20893 9355 20927
rect 9355 20893 9364 20927
rect 9312 20884 9364 20893
rect 30656 20927 30708 20936
rect 30656 20893 30665 20927
rect 30665 20893 30699 20927
rect 30699 20893 30708 20927
rect 30656 20884 30708 20893
rect 30748 20884 30800 20936
rect 35072 20884 35124 20936
rect 37832 20952 37884 21004
rect 38292 20884 38344 20936
rect 46940 20884 46992 20936
rect 28816 20816 28868 20868
rect 36176 20816 36228 20868
rect 36360 20816 36412 20868
rect 2872 20748 2924 20800
rect 30288 20791 30340 20800
rect 30288 20757 30297 20791
rect 30297 20757 30331 20791
rect 30331 20757 30340 20791
rect 30288 20748 30340 20757
rect 31300 20748 31352 20800
rect 31944 20748 31996 20800
rect 36544 20748 36596 20800
rect 37648 20816 37700 20868
rect 49148 20859 49200 20868
rect 49148 20825 49157 20859
rect 49157 20825 49191 20859
rect 49191 20825 49200 20859
rect 49148 20816 49200 20825
rect 7950 20646 8002 20698
rect 8014 20646 8066 20698
rect 8078 20646 8130 20698
rect 8142 20646 8194 20698
rect 8206 20646 8258 20698
rect 17950 20646 18002 20698
rect 18014 20646 18066 20698
rect 18078 20646 18130 20698
rect 18142 20646 18194 20698
rect 18206 20646 18258 20698
rect 27950 20646 28002 20698
rect 28014 20646 28066 20698
rect 28078 20646 28130 20698
rect 28142 20646 28194 20698
rect 28206 20646 28258 20698
rect 37950 20646 38002 20698
rect 38014 20646 38066 20698
rect 38078 20646 38130 20698
rect 38142 20646 38194 20698
rect 38206 20646 38258 20698
rect 47950 20646 48002 20698
rect 48014 20646 48066 20698
rect 48078 20646 48130 20698
rect 48142 20646 48194 20698
rect 48206 20646 48258 20698
rect 21640 20544 21692 20596
rect 21824 20544 21876 20596
rect 22468 20544 22520 20596
rect 21364 20476 21416 20528
rect 2780 20408 2832 20460
rect 20812 20408 20864 20460
rect 22284 20408 22336 20460
rect 1308 20340 1360 20392
rect 21732 20340 21784 20392
rect 19800 20204 19852 20256
rect 23296 20476 23348 20528
rect 24676 20544 24728 20596
rect 26148 20544 26200 20596
rect 27160 20408 27212 20460
rect 30472 20587 30524 20596
rect 30472 20553 30481 20587
rect 30481 20553 30515 20587
rect 30515 20553 30524 20587
rect 30472 20544 30524 20553
rect 32864 20587 32916 20596
rect 32864 20553 32873 20587
rect 32873 20553 32907 20587
rect 32907 20553 32916 20587
rect 32864 20544 32916 20553
rect 30748 20476 30800 20528
rect 34520 20408 34572 20460
rect 47860 20408 47912 20460
rect 23296 20383 23348 20392
rect 23296 20349 23305 20383
rect 23305 20349 23339 20383
rect 23339 20349 23348 20383
rect 23296 20340 23348 20349
rect 25136 20340 25188 20392
rect 26608 20340 26660 20392
rect 32220 20340 32272 20392
rect 34244 20340 34296 20392
rect 49148 20383 49200 20392
rect 49148 20349 49157 20383
rect 49157 20349 49191 20383
rect 49191 20349 49200 20383
rect 49148 20340 49200 20349
rect 25688 20204 25740 20256
rect 25780 20247 25832 20256
rect 25780 20213 25789 20247
rect 25789 20213 25823 20247
rect 25823 20213 25832 20247
rect 25780 20204 25832 20213
rect 32496 20204 32548 20256
rect 39948 20204 40000 20256
rect 2950 20102 3002 20154
rect 3014 20102 3066 20154
rect 3078 20102 3130 20154
rect 3142 20102 3194 20154
rect 3206 20102 3258 20154
rect 12950 20102 13002 20154
rect 13014 20102 13066 20154
rect 13078 20102 13130 20154
rect 13142 20102 13194 20154
rect 13206 20102 13258 20154
rect 22950 20102 23002 20154
rect 23014 20102 23066 20154
rect 23078 20102 23130 20154
rect 23142 20102 23194 20154
rect 23206 20102 23258 20154
rect 32950 20102 33002 20154
rect 33014 20102 33066 20154
rect 33078 20102 33130 20154
rect 33142 20102 33194 20154
rect 33206 20102 33258 20154
rect 42950 20102 43002 20154
rect 43014 20102 43066 20154
rect 43078 20102 43130 20154
rect 43142 20102 43194 20154
rect 43206 20102 43258 20154
rect 10968 20000 11020 20052
rect 19340 19932 19392 19984
rect 21548 19932 21600 19984
rect 17868 19796 17920 19848
rect 19432 19864 19484 19916
rect 21824 19907 21876 19916
rect 21824 19873 21833 19907
rect 21833 19873 21867 19907
rect 21867 19873 21876 19907
rect 21824 19864 21876 19873
rect 22468 19864 22520 19916
rect 22744 19864 22796 19916
rect 23572 20000 23624 20052
rect 26700 20043 26752 20052
rect 26700 20009 26709 20043
rect 26709 20009 26743 20043
rect 26743 20009 26752 20043
rect 26700 20000 26752 20009
rect 23204 19932 23256 19984
rect 25136 19932 25188 19984
rect 23480 19864 23532 19916
rect 25688 19864 25740 19916
rect 27344 19907 27396 19916
rect 27344 19873 27353 19907
rect 27353 19873 27387 19907
rect 27387 19873 27396 19907
rect 27344 19864 27396 19873
rect 20996 19796 21048 19848
rect 19432 19728 19484 19780
rect 20168 19728 20220 19780
rect 23848 19796 23900 19848
rect 28908 19796 28960 19848
rect 18420 19660 18472 19712
rect 22560 19728 22612 19780
rect 35164 20000 35216 20052
rect 31852 19932 31904 19984
rect 32036 19864 32088 19916
rect 35440 19864 35492 19916
rect 36912 19864 36964 19916
rect 32312 19839 32364 19848
rect 32312 19805 32321 19839
rect 32321 19805 32355 19839
rect 32355 19805 32364 19839
rect 32312 19796 32364 19805
rect 33324 19796 33376 19848
rect 33968 19796 34020 19848
rect 34980 19839 35032 19848
rect 34980 19805 34989 19839
rect 34989 19805 35023 19839
rect 35023 19805 35032 19839
rect 34980 19796 35032 19805
rect 36728 19796 36780 19848
rect 41236 19796 41288 19848
rect 32036 19728 32088 19780
rect 23940 19660 23992 19712
rect 25596 19703 25648 19712
rect 25596 19669 25605 19703
rect 25605 19669 25639 19703
rect 25639 19669 25648 19703
rect 25596 19660 25648 19669
rect 26424 19660 26476 19712
rect 26976 19660 27028 19712
rect 32312 19660 32364 19712
rect 34152 19728 34204 19780
rect 46204 19728 46256 19780
rect 34980 19660 35032 19712
rect 7950 19558 8002 19610
rect 8014 19558 8066 19610
rect 8078 19558 8130 19610
rect 8142 19558 8194 19610
rect 8206 19558 8258 19610
rect 17950 19558 18002 19610
rect 18014 19558 18066 19610
rect 18078 19558 18130 19610
rect 18142 19558 18194 19610
rect 18206 19558 18258 19610
rect 27950 19558 28002 19610
rect 28014 19558 28066 19610
rect 28078 19558 28130 19610
rect 28142 19558 28194 19610
rect 28206 19558 28258 19610
rect 37950 19558 38002 19610
rect 38014 19558 38066 19610
rect 38078 19558 38130 19610
rect 38142 19558 38194 19610
rect 38206 19558 38258 19610
rect 47950 19558 48002 19610
rect 48014 19558 48066 19610
rect 48078 19558 48130 19610
rect 48142 19558 48194 19610
rect 48206 19558 48258 19610
rect 16488 19456 16540 19508
rect 22376 19456 22428 19508
rect 23848 19456 23900 19508
rect 21180 19388 21232 19440
rect 22468 19320 22520 19372
rect 21548 19252 21600 19304
rect 24492 19320 24544 19372
rect 27804 19456 27856 19508
rect 28816 19456 28868 19508
rect 24768 19388 24820 19440
rect 26700 19388 26752 19440
rect 26792 19388 26844 19440
rect 23296 19252 23348 19304
rect 24860 19295 24912 19304
rect 21916 19116 21968 19168
rect 22744 19116 22796 19168
rect 22836 19159 22888 19168
rect 22836 19125 22845 19159
rect 22845 19125 22879 19159
rect 22879 19125 22888 19159
rect 22836 19116 22888 19125
rect 24860 19261 24869 19295
rect 24869 19261 24903 19295
rect 24903 19261 24912 19295
rect 24860 19252 24912 19261
rect 27436 19320 27488 19372
rect 27804 19295 27856 19304
rect 27804 19261 27813 19295
rect 27813 19261 27847 19295
rect 27847 19261 27856 19295
rect 27804 19252 27856 19261
rect 24584 19184 24636 19236
rect 27068 19184 27120 19236
rect 27160 19227 27212 19236
rect 27160 19193 27169 19227
rect 27169 19193 27203 19227
rect 27203 19193 27212 19227
rect 27160 19184 27212 19193
rect 29092 19320 29144 19372
rect 26884 19116 26936 19168
rect 27252 19116 27304 19168
rect 33508 19320 33560 19372
rect 38476 19456 38528 19508
rect 35900 19320 35952 19372
rect 39028 19388 39080 19440
rect 37464 19363 37516 19372
rect 37464 19329 37473 19363
rect 37473 19329 37507 19363
rect 37507 19329 37516 19363
rect 37464 19320 37516 19329
rect 45468 19320 45520 19372
rect 49148 19363 49200 19372
rect 49148 19329 49157 19363
rect 49157 19329 49191 19363
rect 49191 19329 49200 19363
rect 49148 19320 49200 19329
rect 28540 19184 28592 19236
rect 37280 19252 37332 19304
rect 34428 19116 34480 19168
rect 35440 19159 35492 19168
rect 35440 19125 35449 19159
rect 35449 19125 35483 19159
rect 35483 19125 35492 19159
rect 35440 19116 35492 19125
rect 36636 19184 36688 19236
rect 36084 19116 36136 19168
rect 37556 19116 37608 19168
rect 2950 19014 3002 19066
rect 3014 19014 3066 19066
rect 3078 19014 3130 19066
rect 3142 19014 3194 19066
rect 3206 19014 3258 19066
rect 12950 19014 13002 19066
rect 13014 19014 13066 19066
rect 13078 19014 13130 19066
rect 13142 19014 13194 19066
rect 13206 19014 13258 19066
rect 22950 19014 23002 19066
rect 23014 19014 23066 19066
rect 23078 19014 23130 19066
rect 23142 19014 23194 19066
rect 23206 19014 23258 19066
rect 32950 19014 33002 19066
rect 33014 19014 33066 19066
rect 33078 19014 33130 19066
rect 33142 19014 33194 19066
rect 33206 19014 33258 19066
rect 42950 19014 43002 19066
rect 43014 19014 43066 19066
rect 43078 19014 43130 19066
rect 43142 19014 43194 19066
rect 43206 19014 43258 19066
rect 18788 18912 18840 18964
rect 19892 18912 19944 18964
rect 22100 18912 22152 18964
rect 22376 18912 22428 18964
rect 22468 18955 22520 18964
rect 22468 18921 22477 18955
rect 22477 18921 22511 18955
rect 22511 18921 22520 18955
rect 22468 18912 22520 18921
rect 22744 18912 22796 18964
rect 24768 18912 24820 18964
rect 27804 18912 27856 18964
rect 28540 18912 28592 18964
rect 37556 18912 37608 18964
rect 9772 18844 9824 18896
rect 21180 18844 21232 18896
rect 32864 18844 32916 18896
rect 9312 18708 9364 18760
rect 12532 18708 12584 18760
rect 20536 18640 20588 18692
rect 2780 18572 2832 18624
rect 20628 18615 20680 18624
rect 20628 18581 20637 18615
rect 20637 18581 20671 18615
rect 20671 18581 20680 18615
rect 20628 18572 20680 18581
rect 21824 18776 21876 18828
rect 23480 18776 23532 18828
rect 24308 18776 24360 18828
rect 26608 18819 26660 18828
rect 26608 18785 26617 18819
rect 26617 18785 26651 18819
rect 26651 18785 26660 18819
rect 26608 18776 26660 18785
rect 26976 18776 27028 18828
rect 22468 18708 22520 18760
rect 25780 18708 25832 18760
rect 27528 18708 27580 18760
rect 27620 18708 27672 18760
rect 28356 18708 28408 18760
rect 28816 18776 28868 18828
rect 31392 18819 31444 18828
rect 31392 18785 31401 18819
rect 31401 18785 31435 18819
rect 31435 18785 31444 18819
rect 31392 18776 31444 18785
rect 32588 18776 32640 18828
rect 37280 18776 37332 18828
rect 41328 18708 41380 18760
rect 44456 18708 44508 18760
rect 21456 18683 21508 18692
rect 21456 18649 21465 18683
rect 21465 18649 21499 18683
rect 21499 18649 21508 18683
rect 21456 18640 21508 18649
rect 22100 18572 22152 18624
rect 22284 18683 22336 18692
rect 22284 18649 22293 18683
rect 22293 18649 22327 18683
rect 22327 18649 22336 18683
rect 22284 18640 22336 18649
rect 28448 18640 28500 18692
rect 23388 18572 23440 18624
rect 24860 18572 24912 18624
rect 24952 18615 25004 18624
rect 24952 18581 24961 18615
rect 24961 18581 24995 18615
rect 24995 18581 25004 18615
rect 24952 18572 25004 18581
rect 25872 18572 25924 18624
rect 25964 18615 26016 18624
rect 25964 18581 25973 18615
rect 25973 18581 26007 18615
rect 26007 18581 26016 18615
rect 25964 18572 26016 18581
rect 27252 18572 27304 18624
rect 27344 18572 27396 18624
rect 29276 18572 29328 18624
rect 36728 18640 36780 18692
rect 37188 18683 37240 18692
rect 37188 18649 37197 18683
rect 37197 18649 37231 18683
rect 37231 18649 37240 18683
rect 37188 18640 37240 18649
rect 38660 18640 38712 18692
rect 47860 18640 47912 18692
rect 49148 18683 49200 18692
rect 49148 18649 49157 18683
rect 49157 18649 49191 18683
rect 49191 18649 49200 18683
rect 49148 18640 49200 18649
rect 37004 18572 37056 18624
rect 7950 18470 8002 18522
rect 8014 18470 8066 18522
rect 8078 18470 8130 18522
rect 8142 18470 8194 18522
rect 8206 18470 8258 18522
rect 17950 18470 18002 18522
rect 18014 18470 18066 18522
rect 18078 18470 18130 18522
rect 18142 18470 18194 18522
rect 18206 18470 18258 18522
rect 27950 18470 28002 18522
rect 28014 18470 28066 18522
rect 28078 18470 28130 18522
rect 28142 18470 28194 18522
rect 28206 18470 28258 18522
rect 37950 18470 38002 18522
rect 38014 18470 38066 18522
rect 38078 18470 38130 18522
rect 38142 18470 38194 18522
rect 38206 18470 38258 18522
rect 47950 18470 48002 18522
rect 48014 18470 48066 18522
rect 48078 18470 48130 18522
rect 48142 18470 48194 18522
rect 48206 18470 48258 18522
rect 19800 18411 19852 18420
rect 19800 18377 19809 18411
rect 19809 18377 19843 18411
rect 19843 18377 19852 18411
rect 19800 18368 19852 18377
rect 20628 18368 20680 18420
rect 21456 18300 21508 18352
rect 21548 18300 21600 18352
rect 24584 18300 24636 18352
rect 2872 18232 2924 18284
rect 22100 18232 22152 18284
rect 22284 18232 22336 18284
rect 24952 18368 25004 18420
rect 27620 18411 27672 18420
rect 27620 18377 27629 18411
rect 27629 18377 27663 18411
rect 27663 18377 27672 18411
rect 27620 18368 27672 18377
rect 24860 18300 24912 18352
rect 27160 18300 27212 18352
rect 28448 18343 28500 18352
rect 28448 18309 28457 18343
rect 28457 18309 28491 18343
rect 28491 18309 28500 18343
rect 28448 18300 28500 18309
rect 34796 18368 34848 18420
rect 37740 18368 37792 18420
rect 32312 18300 32364 18352
rect 32588 18343 32640 18352
rect 32588 18309 32597 18343
rect 32597 18309 32631 18343
rect 32631 18309 32640 18343
rect 32588 18300 32640 18309
rect 1308 18164 1360 18216
rect 20076 18164 20128 18216
rect 20996 18164 21048 18216
rect 18788 18096 18840 18148
rect 19800 18028 19852 18080
rect 21916 18096 21968 18148
rect 22560 18096 22612 18148
rect 24768 18028 24820 18080
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 27344 18232 27396 18284
rect 27436 18164 27488 18216
rect 26792 18096 26844 18148
rect 31208 18232 31260 18284
rect 30012 18164 30064 18216
rect 30380 18207 30432 18216
rect 30380 18173 30389 18207
rect 30389 18173 30423 18207
rect 30423 18173 30432 18207
rect 30380 18164 30432 18173
rect 33324 18164 33376 18216
rect 34428 18300 34480 18352
rect 36084 18300 36136 18352
rect 36820 18300 36872 18352
rect 37372 18232 37424 18284
rect 46664 18232 46716 18284
rect 29092 18028 29144 18080
rect 33692 18028 33744 18080
rect 34796 18207 34848 18216
rect 34796 18173 34805 18207
rect 34805 18173 34839 18207
rect 34839 18173 34848 18207
rect 34796 18164 34848 18173
rect 35256 18164 35308 18216
rect 38016 18164 38068 18216
rect 38476 18164 38528 18216
rect 49148 18207 49200 18216
rect 49148 18173 49157 18207
rect 49157 18173 49191 18207
rect 49191 18173 49200 18207
rect 49148 18164 49200 18173
rect 34888 18028 34940 18080
rect 36084 18028 36136 18080
rect 41788 18028 41840 18080
rect 2950 17926 3002 17978
rect 3014 17926 3066 17978
rect 3078 17926 3130 17978
rect 3142 17926 3194 17978
rect 3206 17926 3258 17978
rect 12950 17926 13002 17978
rect 13014 17926 13066 17978
rect 13078 17926 13130 17978
rect 13142 17926 13194 17978
rect 13206 17926 13258 17978
rect 22950 17926 23002 17978
rect 23014 17926 23066 17978
rect 23078 17926 23130 17978
rect 23142 17926 23194 17978
rect 23206 17926 23258 17978
rect 32950 17926 33002 17978
rect 33014 17926 33066 17978
rect 33078 17926 33130 17978
rect 33142 17926 33194 17978
rect 33206 17926 33258 17978
rect 42950 17926 43002 17978
rect 43014 17926 43066 17978
rect 43078 17926 43130 17978
rect 43142 17926 43194 17978
rect 43206 17926 43258 17978
rect 17868 17824 17920 17876
rect 19892 17756 19944 17808
rect 21916 17824 21968 17876
rect 22008 17824 22060 17876
rect 22468 17824 22520 17876
rect 25596 17824 25648 17876
rect 32588 17824 32640 17876
rect 37188 17824 37240 17876
rect 22376 17756 22428 17808
rect 21272 17731 21324 17740
rect 21272 17697 21281 17731
rect 21281 17697 21315 17731
rect 21315 17697 21324 17731
rect 21272 17688 21324 17697
rect 21364 17688 21416 17740
rect 22652 17688 22704 17740
rect 27068 17756 27120 17808
rect 27436 17688 27488 17740
rect 30012 17688 30064 17740
rect 34336 17756 34388 17808
rect 37096 17756 37148 17808
rect 19248 17620 19300 17672
rect 20996 17663 21048 17672
rect 20996 17629 21005 17663
rect 21005 17629 21039 17663
rect 21039 17629 21048 17663
rect 20996 17620 21048 17629
rect 23296 17620 23348 17672
rect 27620 17620 27672 17672
rect 21364 17552 21416 17604
rect 22284 17552 22336 17604
rect 30288 17552 30340 17604
rect 30932 17595 30984 17604
rect 30932 17561 30941 17595
rect 30941 17561 30975 17595
rect 30975 17561 30984 17595
rect 30932 17552 30984 17561
rect 18788 17484 18840 17536
rect 19800 17527 19852 17536
rect 19800 17493 19809 17527
rect 19809 17493 19843 17527
rect 19843 17493 19852 17527
rect 19800 17484 19852 17493
rect 19892 17527 19944 17536
rect 19892 17493 19901 17527
rect 19901 17493 19935 17527
rect 19935 17493 19944 17527
rect 19892 17484 19944 17493
rect 19984 17484 20036 17536
rect 22008 17484 22060 17536
rect 24584 17484 24636 17536
rect 26148 17484 26200 17536
rect 27344 17484 27396 17536
rect 29736 17484 29788 17536
rect 30564 17484 30616 17536
rect 33324 17620 33376 17672
rect 33784 17620 33836 17672
rect 35900 17688 35952 17740
rect 37280 17688 37332 17740
rect 38016 17731 38068 17740
rect 38016 17697 38025 17731
rect 38025 17697 38059 17731
rect 38059 17697 38068 17731
rect 38016 17688 38068 17697
rect 38568 17688 38620 17740
rect 44824 17756 44876 17808
rect 36084 17552 36136 17604
rect 36820 17552 36872 17604
rect 37096 17552 37148 17604
rect 37832 17484 37884 17536
rect 38660 17552 38712 17604
rect 39948 17484 40000 17536
rect 45100 17620 45152 17672
rect 46848 17552 46900 17604
rect 49148 17595 49200 17604
rect 49148 17561 49157 17595
rect 49157 17561 49191 17595
rect 49191 17561 49200 17595
rect 49148 17552 49200 17561
rect 46664 17484 46716 17536
rect 7950 17382 8002 17434
rect 8014 17382 8066 17434
rect 8078 17382 8130 17434
rect 8142 17382 8194 17434
rect 8206 17382 8258 17434
rect 17950 17382 18002 17434
rect 18014 17382 18066 17434
rect 18078 17382 18130 17434
rect 18142 17382 18194 17434
rect 18206 17382 18258 17434
rect 27950 17382 28002 17434
rect 28014 17382 28066 17434
rect 28078 17382 28130 17434
rect 28142 17382 28194 17434
rect 28206 17382 28258 17434
rect 37950 17382 38002 17434
rect 38014 17382 38066 17434
rect 38078 17382 38130 17434
rect 38142 17382 38194 17434
rect 38206 17382 38258 17434
rect 47950 17382 48002 17434
rect 48014 17382 48066 17434
rect 48078 17382 48130 17434
rect 48142 17382 48194 17434
rect 48206 17382 48258 17434
rect 21272 17280 21324 17332
rect 22100 17280 22152 17332
rect 23296 17323 23348 17332
rect 23296 17289 23305 17323
rect 23305 17289 23339 17323
rect 23339 17289 23348 17323
rect 23296 17280 23348 17289
rect 24216 17280 24268 17332
rect 20720 17212 20772 17264
rect 19248 17076 19300 17128
rect 20076 17076 20128 17128
rect 20720 17076 20772 17128
rect 22284 17212 22336 17264
rect 21732 17076 21784 17128
rect 21916 17076 21968 17128
rect 25044 17255 25096 17264
rect 25044 17221 25053 17255
rect 25053 17221 25087 17255
rect 25087 17221 25096 17255
rect 25044 17212 25096 17221
rect 27252 17323 27304 17332
rect 27252 17289 27261 17323
rect 27261 17289 27295 17323
rect 27295 17289 27304 17323
rect 27252 17280 27304 17289
rect 27712 17323 27764 17332
rect 27712 17289 27721 17323
rect 27721 17289 27755 17323
rect 27755 17289 27764 17323
rect 27712 17280 27764 17289
rect 28816 17323 28868 17332
rect 28816 17289 28825 17323
rect 28825 17289 28859 17323
rect 28859 17289 28868 17323
rect 28816 17280 28868 17289
rect 26608 17212 26660 17264
rect 31944 17280 31996 17332
rect 32864 17280 32916 17332
rect 36452 17280 36504 17332
rect 36820 17280 36872 17332
rect 38660 17280 38712 17332
rect 30564 17212 30616 17264
rect 33324 17212 33376 17264
rect 33968 17255 34020 17264
rect 33968 17221 33977 17255
rect 33977 17221 34011 17255
rect 34011 17221 34020 17255
rect 33968 17212 34020 17221
rect 43720 17255 43772 17264
rect 43720 17221 43729 17255
rect 43729 17221 43763 17255
rect 43763 17221 43772 17255
rect 43720 17212 43772 17221
rect 26148 17144 26200 17196
rect 19984 16940 20036 16992
rect 22008 16940 22060 16992
rect 25044 17076 25096 17128
rect 28264 17076 28316 17128
rect 28448 17144 28500 17196
rect 28540 17076 28592 17128
rect 32404 17144 32456 17196
rect 33416 17144 33468 17196
rect 29552 17076 29604 17128
rect 30012 17119 30064 17128
rect 30012 17085 30021 17119
rect 30021 17085 30055 17119
rect 30055 17085 30064 17119
rect 30012 17076 30064 17085
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 30932 17076 30984 17128
rect 33600 17076 33652 17128
rect 34612 17076 34664 17128
rect 35256 17119 35308 17128
rect 35256 17085 35265 17119
rect 35265 17085 35299 17119
rect 35299 17085 35308 17119
rect 35256 17076 35308 17085
rect 25688 16940 25740 16992
rect 26608 16940 26660 16992
rect 28448 16983 28500 16992
rect 28448 16949 28457 16983
rect 28457 16949 28491 16983
rect 28491 16949 28500 16983
rect 28448 16940 28500 16949
rect 30472 16940 30524 16992
rect 32312 16983 32364 16992
rect 32312 16949 32321 16983
rect 32321 16949 32355 16983
rect 32355 16949 32364 16983
rect 32312 16940 32364 16949
rect 40224 17008 40276 17060
rect 46756 17008 46808 17060
rect 36820 16940 36872 16992
rect 38108 16983 38160 16992
rect 38108 16949 38117 16983
rect 38117 16949 38151 16983
rect 38151 16949 38160 16983
rect 38108 16940 38160 16949
rect 2950 16838 3002 16890
rect 3014 16838 3066 16890
rect 3078 16838 3130 16890
rect 3142 16838 3194 16890
rect 3206 16838 3258 16890
rect 12950 16838 13002 16890
rect 13014 16838 13066 16890
rect 13078 16838 13130 16890
rect 13142 16838 13194 16890
rect 13206 16838 13258 16890
rect 22950 16838 23002 16890
rect 23014 16838 23066 16890
rect 23078 16838 23130 16890
rect 23142 16838 23194 16890
rect 23206 16838 23258 16890
rect 32950 16838 33002 16890
rect 33014 16838 33066 16890
rect 33078 16838 33130 16890
rect 33142 16838 33194 16890
rect 33206 16838 33258 16890
rect 42950 16838 43002 16890
rect 43014 16838 43066 16890
rect 43078 16838 43130 16890
rect 43142 16838 43194 16890
rect 43206 16838 43258 16890
rect 19432 16736 19484 16788
rect 19708 16779 19760 16788
rect 19708 16745 19732 16779
rect 19732 16745 19760 16779
rect 19708 16736 19760 16745
rect 20076 16736 20128 16788
rect 24676 16736 24728 16788
rect 18604 16600 18656 16652
rect 19248 16600 19300 16652
rect 22468 16600 22520 16652
rect 25044 16643 25096 16652
rect 25044 16609 25053 16643
rect 25053 16609 25087 16643
rect 25087 16609 25096 16643
rect 25044 16600 25096 16609
rect 26700 16600 26752 16652
rect 34060 16643 34112 16652
rect 34060 16609 34069 16643
rect 34069 16609 34103 16643
rect 34103 16609 34112 16643
rect 34060 16600 34112 16609
rect 36176 16736 36228 16788
rect 37096 16736 37148 16788
rect 34612 16668 34664 16720
rect 34888 16643 34940 16652
rect 34888 16609 34897 16643
rect 34897 16609 34931 16643
rect 34931 16609 34940 16643
rect 34888 16600 34940 16609
rect 35532 16600 35584 16652
rect 37188 16600 37240 16652
rect 24584 16532 24636 16584
rect 25964 16532 26016 16584
rect 26056 16532 26108 16584
rect 28448 16532 28500 16584
rect 30564 16532 30616 16584
rect 37832 16532 37884 16584
rect 46204 16532 46256 16584
rect 9772 16464 9824 16516
rect 5632 16439 5684 16448
rect 5632 16405 5641 16439
rect 5641 16405 5675 16439
rect 5675 16405 5684 16439
rect 5632 16396 5684 16405
rect 19248 16396 19300 16448
rect 20720 16396 20772 16448
rect 21180 16439 21232 16448
rect 21180 16405 21189 16439
rect 21189 16405 21223 16439
rect 21223 16405 21232 16439
rect 21180 16396 21232 16405
rect 21916 16507 21968 16516
rect 21916 16473 21925 16507
rect 21925 16473 21959 16507
rect 21959 16473 21968 16507
rect 21916 16464 21968 16473
rect 22100 16396 22152 16448
rect 25780 16464 25832 16516
rect 29460 16464 29512 16516
rect 31576 16464 31628 16516
rect 27160 16439 27212 16448
rect 27160 16405 27169 16439
rect 27169 16405 27203 16439
rect 27203 16405 27212 16439
rect 27160 16396 27212 16405
rect 27528 16396 27580 16448
rect 28264 16396 28316 16448
rect 28448 16396 28500 16448
rect 28540 16396 28592 16448
rect 33140 16396 33192 16448
rect 34520 16464 34572 16516
rect 36452 16464 36504 16516
rect 36636 16439 36688 16448
rect 36636 16405 36645 16439
rect 36645 16405 36679 16439
rect 36679 16405 36688 16439
rect 36636 16396 36688 16405
rect 36912 16396 36964 16448
rect 40132 16464 40184 16516
rect 49148 16507 49200 16516
rect 49148 16473 49157 16507
rect 49157 16473 49191 16507
rect 49191 16473 49200 16507
rect 49148 16464 49200 16473
rect 38108 16396 38160 16448
rect 7950 16294 8002 16346
rect 8014 16294 8066 16346
rect 8078 16294 8130 16346
rect 8142 16294 8194 16346
rect 8206 16294 8258 16346
rect 17950 16294 18002 16346
rect 18014 16294 18066 16346
rect 18078 16294 18130 16346
rect 18142 16294 18194 16346
rect 18206 16294 18258 16346
rect 27950 16294 28002 16346
rect 28014 16294 28066 16346
rect 28078 16294 28130 16346
rect 28142 16294 28194 16346
rect 28206 16294 28258 16346
rect 37950 16294 38002 16346
rect 38014 16294 38066 16346
rect 38078 16294 38130 16346
rect 38142 16294 38194 16346
rect 38206 16294 38258 16346
rect 47950 16294 48002 16346
rect 48014 16294 48066 16346
rect 48078 16294 48130 16346
rect 48142 16294 48194 16346
rect 48206 16294 48258 16346
rect 18788 16192 18840 16244
rect 25780 16235 25832 16244
rect 25780 16201 25789 16235
rect 25789 16201 25823 16235
rect 25823 16201 25832 16235
rect 25780 16192 25832 16201
rect 25872 16192 25924 16244
rect 27252 16192 27304 16244
rect 29736 16192 29788 16244
rect 16396 16124 16448 16176
rect 24584 16124 24636 16176
rect 24768 16167 24820 16176
rect 24768 16133 24777 16167
rect 24777 16133 24811 16167
rect 24811 16133 24820 16167
rect 24768 16124 24820 16133
rect 2780 16056 2832 16108
rect 22468 16056 22520 16108
rect 26056 16056 26108 16108
rect 29368 16124 29420 16176
rect 30472 16124 30524 16176
rect 28816 16099 28868 16108
rect 1308 15988 1360 16040
rect 26148 15988 26200 16040
rect 27436 15988 27488 16040
rect 27620 15920 27672 15972
rect 28816 16065 28825 16099
rect 28825 16065 28859 16099
rect 28859 16065 28868 16099
rect 28816 16056 28868 16065
rect 29184 15988 29236 16040
rect 29460 15988 29512 16040
rect 33416 16124 33468 16176
rect 37372 16124 37424 16176
rect 36360 16056 36412 16108
rect 40040 16056 40092 16108
rect 47860 16056 47912 16108
rect 33140 15988 33192 16040
rect 37556 15988 37608 16040
rect 49148 16031 49200 16040
rect 49148 15997 49157 16031
rect 49157 15997 49191 16031
rect 49191 15997 49200 16031
rect 49148 15988 49200 15997
rect 30196 15920 30248 15972
rect 33232 15920 33284 15972
rect 33324 15920 33376 15972
rect 39120 15920 39172 15972
rect 29828 15852 29880 15904
rect 30104 15852 30156 15904
rect 32864 15852 32916 15904
rect 33416 15852 33468 15904
rect 36084 15895 36136 15904
rect 36084 15861 36093 15895
rect 36093 15861 36127 15895
rect 36127 15861 36136 15895
rect 36084 15852 36136 15861
rect 37648 15895 37700 15904
rect 37648 15861 37657 15895
rect 37657 15861 37691 15895
rect 37691 15861 37700 15895
rect 37648 15852 37700 15861
rect 37832 15852 37884 15904
rect 2950 15750 3002 15802
rect 3014 15750 3066 15802
rect 3078 15750 3130 15802
rect 3142 15750 3194 15802
rect 3206 15750 3258 15802
rect 12950 15750 13002 15802
rect 13014 15750 13066 15802
rect 13078 15750 13130 15802
rect 13142 15750 13194 15802
rect 13206 15750 13258 15802
rect 22950 15750 23002 15802
rect 23014 15750 23066 15802
rect 23078 15750 23130 15802
rect 23142 15750 23194 15802
rect 23206 15750 23258 15802
rect 32950 15750 33002 15802
rect 33014 15750 33066 15802
rect 33078 15750 33130 15802
rect 33142 15750 33194 15802
rect 33206 15750 33258 15802
rect 42950 15750 43002 15802
rect 43014 15750 43066 15802
rect 43078 15750 43130 15802
rect 43142 15750 43194 15802
rect 43206 15750 43258 15802
rect 26424 15691 26476 15700
rect 26424 15657 26433 15691
rect 26433 15657 26467 15691
rect 26467 15657 26476 15691
rect 26424 15648 26476 15657
rect 23388 15512 23440 15564
rect 30196 15648 30248 15700
rect 33324 15648 33376 15700
rect 29460 15580 29512 15632
rect 32312 15580 32364 15632
rect 32588 15580 32640 15632
rect 19892 15444 19944 15496
rect 20536 15444 20588 15496
rect 25228 15376 25280 15428
rect 27252 15376 27304 15428
rect 28816 15512 28868 15564
rect 30012 15512 30064 15564
rect 33600 15555 33652 15564
rect 33600 15521 33609 15555
rect 33609 15521 33643 15555
rect 33643 15521 33652 15555
rect 33600 15512 33652 15521
rect 35900 15555 35952 15564
rect 35900 15521 35909 15555
rect 35909 15521 35943 15555
rect 35943 15521 35952 15555
rect 35900 15512 35952 15521
rect 36176 15555 36228 15564
rect 36176 15521 36185 15555
rect 36185 15521 36219 15555
rect 36219 15521 36228 15555
rect 36176 15512 36228 15521
rect 29000 15487 29052 15496
rect 29000 15453 29009 15487
rect 29009 15453 29043 15487
rect 29043 15453 29052 15487
rect 29000 15444 29052 15453
rect 32496 15444 32548 15496
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 33692 15444 33744 15496
rect 46848 15444 46900 15496
rect 29184 15376 29236 15428
rect 22652 15308 22704 15360
rect 25596 15308 25648 15360
rect 26056 15308 26108 15360
rect 29644 15376 29696 15428
rect 30104 15376 30156 15428
rect 29460 15308 29512 15360
rect 30472 15376 30524 15428
rect 36452 15376 36504 15428
rect 36636 15376 36688 15428
rect 49148 15419 49200 15428
rect 49148 15385 49157 15419
rect 49157 15385 49191 15419
rect 49191 15385 49200 15419
rect 49148 15376 49200 15385
rect 30288 15308 30340 15360
rect 31576 15308 31628 15360
rect 31760 15308 31812 15360
rect 32404 15351 32456 15360
rect 32404 15317 32413 15351
rect 32413 15317 32447 15351
rect 32447 15317 32456 15351
rect 32404 15308 32456 15317
rect 37740 15308 37792 15360
rect 7950 15206 8002 15258
rect 8014 15206 8066 15258
rect 8078 15206 8130 15258
rect 8142 15206 8194 15258
rect 8206 15206 8258 15258
rect 17950 15206 18002 15258
rect 18014 15206 18066 15258
rect 18078 15206 18130 15258
rect 18142 15206 18194 15258
rect 18206 15206 18258 15258
rect 27950 15206 28002 15258
rect 28014 15206 28066 15258
rect 28078 15206 28130 15258
rect 28142 15206 28194 15258
rect 28206 15206 28258 15258
rect 37950 15206 38002 15258
rect 38014 15206 38066 15258
rect 38078 15206 38130 15258
rect 38142 15206 38194 15258
rect 38206 15206 38258 15258
rect 47950 15206 48002 15258
rect 48014 15206 48066 15258
rect 48078 15206 48130 15258
rect 48142 15206 48194 15258
rect 48206 15206 48258 15258
rect 19340 15104 19392 15156
rect 25044 15104 25096 15156
rect 29184 15104 29236 15156
rect 29644 15104 29696 15156
rect 37648 15104 37700 15156
rect 24584 15036 24636 15088
rect 27804 15036 27856 15088
rect 29460 15036 29512 15088
rect 29920 15079 29972 15088
rect 29920 15045 29929 15079
rect 29929 15045 29963 15079
rect 29963 15045 29972 15079
rect 29920 15036 29972 15045
rect 31484 15036 31536 15088
rect 36820 15036 36872 15088
rect 17868 14968 17920 15020
rect 22468 15011 22520 15020
rect 22468 14977 22477 15011
rect 22477 14977 22511 15011
rect 22511 14977 22520 15011
rect 22468 14968 22520 14977
rect 25688 14968 25740 15020
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 27620 14968 27672 14977
rect 32220 14968 32272 15020
rect 41788 15011 41840 15020
rect 41788 14977 41797 15011
rect 41797 14977 41831 15011
rect 41831 14977 41840 15011
rect 41788 14968 41840 14977
rect 46756 14968 46808 15020
rect 21180 14900 21232 14952
rect 26148 14900 26200 14952
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 26608 14900 26660 14952
rect 27896 14943 27948 14952
rect 27896 14909 27905 14943
rect 27905 14909 27939 14943
rect 27939 14909 27948 14943
rect 27896 14900 27948 14909
rect 32128 14900 32180 14952
rect 32864 14943 32916 14952
rect 32864 14909 32873 14943
rect 32873 14909 32907 14943
rect 32907 14909 32916 14943
rect 32864 14900 32916 14909
rect 36912 14900 36964 14952
rect 49148 14943 49200 14952
rect 49148 14909 49157 14943
rect 49157 14909 49191 14943
rect 49191 14909 49200 14943
rect 49148 14900 49200 14909
rect 30012 14764 30064 14816
rect 30196 14764 30248 14816
rect 38292 14832 38344 14884
rect 33784 14764 33836 14816
rect 41236 14764 41288 14816
rect 44180 14764 44232 14816
rect 2950 14662 3002 14714
rect 3014 14662 3066 14714
rect 3078 14662 3130 14714
rect 3142 14662 3194 14714
rect 3206 14662 3258 14714
rect 12950 14662 13002 14714
rect 13014 14662 13066 14714
rect 13078 14662 13130 14714
rect 13142 14662 13194 14714
rect 13206 14662 13258 14714
rect 22950 14662 23002 14714
rect 23014 14662 23066 14714
rect 23078 14662 23130 14714
rect 23142 14662 23194 14714
rect 23206 14662 23258 14714
rect 32950 14662 33002 14714
rect 33014 14662 33066 14714
rect 33078 14662 33130 14714
rect 33142 14662 33194 14714
rect 33206 14662 33258 14714
rect 42950 14662 43002 14714
rect 43014 14662 43066 14714
rect 43078 14662 43130 14714
rect 43142 14662 43194 14714
rect 43206 14662 43258 14714
rect 20444 14560 20496 14612
rect 26332 14560 26384 14612
rect 27896 14560 27948 14612
rect 25688 14424 25740 14476
rect 32220 14603 32272 14612
rect 32220 14569 32229 14603
rect 32229 14569 32263 14603
rect 32263 14569 32272 14603
rect 32220 14560 32272 14569
rect 34336 14492 34388 14544
rect 41328 14492 41380 14544
rect 31760 14424 31812 14476
rect 33968 14424 34020 14476
rect 34520 14424 34572 14476
rect 37740 14467 37792 14476
rect 37740 14433 37749 14467
rect 37749 14433 37783 14467
rect 37783 14433 37792 14467
rect 37740 14424 37792 14433
rect 30196 14399 30248 14408
rect 30196 14365 30205 14399
rect 30205 14365 30239 14399
rect 30239 14365 30248 14399
rect 30196 14356 30248 14365
rect 30288 14356 30340 14408
rect 34244 14356 34296 14408
rect 40040 14356 40092 14408
rect 40224 14399 40276 14408
rect 40224 14365 40233 14399
rect 40233 14365 40267 14399
rect 40267 14365 40276 14399
rect 40224 14356 40276 14365
rect 26148 14331 26200 14340
rect 26148 14297 26157 14331
rect 26157 14297 26191 14331
rect 26191 14297 26200 14331
rect 26148 14288 26200 14297
rect 29460 14288 29512 14340
rect 29920 14220 29972 14272
rect 35164 14331 35216 14340
rect 35164 14297 35173 14331
rect 35173 14297 35207 14331
rect 35207 14297 35216 14331
rect 35164 14288 35216 14297
rect 37740 14288 37792 14340
rect 36912 14220 36964 14272
rect 42800 14220 42852 14272
rect 7950 14118 8002 14170
rect 8014 14118 8066 14170
rect 8078 14118 8130 14170
rect 8142 14118 8194 14170
rect 8206 14118 8258 14170
rect 17950 14118 18002 14170
rect 18014 14118 18066 14170
rect 18078 14118 18130 14170
rect 18142 14118 18194 14170
rect 18206 14118 18258 14170
rect 27950 14118 28002 14170
rect 28014 14118 28066 14170
rect 28078 14118 28130 14170
rect 28142 14118 28194 14170
rect 28206 14118 28258 14170
rect 37950 14118 38002 14170
rect 38014 14118 38066 14170
rect 38078 14118 38130 14170
rect 38142 14118 38194 14170
rect 38206 14118 38258 14170
rect 47950 14118 48002 14170
rect 48014 14118 48066 14170
rect 48078 14118 48130 14170
rect 48142 14118 48194 14170
rect 48206 14118 48258 14170
rect 26332 13948 26384 14000
rect 34888 14016 34940 14068
rect 35900 14016 35952 14068
rect 43720 14016 43772 14068
rect 5632 13880 5684 13932
rect 29276 13880 29328 13932
rect 34704 13948 34756 14000
rect 36544 13948 36596 14000
rect 37740 13991 37792 14000
rect 37740 13957 37749 13991
rect 37749 13957 37783 13991
rect 37783 13957 37792 13991
rect 37740 13948 37792 13957
rect 38384 13948 38436 14000
rect 38936 13948 38988 14000
rect 42708 13948 42760 14000
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 2780 13812 2832 13821
rect 29736 13812 29788 13864
rect 35532 13812 35584 13864
rect 36912 13923 36964 13932
rect 36912 13889 36921 13923
rect 36921 13889 36955 13923
rect 36955 13889 36964 13923
rect 36912 13880 36964 13889
rect 38476 13855 38528 13864
rect 38476 13821 38485 13855
rect 38485 13821 38519 13855
rect 38519 13821 38528 13855
rect 38476 13812 38528 13821
rect 39120 13923 39172 13932
rect 39120 13889 39129 13923
rect 39129 13889 39163 13923
rect 39163 13889 39172 13923
rect 39120 13880 39172 13889
rect 40132 13880 40184 13932
rect 46664 13880 46716 13932
rect 40592 13812 40644 13864
rect 38936 13787 38988 13796
rect 38936 13753 38945 13787
rect 38945 13753 38979 13787
rect 38979 13753 38988 13787
rect 38936 13744 38988 13753
rect 44364 13812 44416 13864
rect 49148 13855 49200 13864
rect 49148 13821 49157 13855
rect 49157 13821 49191 13855
rect 49191 13821 49200 13855
rect 49148 13812 49200 13821
rect 35440 13676 35492 13728
rect 2950 13574 3002 13626
rect 3014 13574 3066 13626
rect 3078 13574 3130 13626
rect 3142 13574 3194 13626
rect 3206 13574 3258 13626
rect 12950 13574 13002 13626
rect 13014 13574 13066 13626
rect 13078 13574 13130 13626
rect 13142 13574 13194 13626
rect 13206 13574 13258 13626
rect 22950 13574 23002 13626
rect 23014 13574 23066 13626
rect 23078 13574 23130 13626
rect 23142 13574 23194 13626
rect 23206 13574 23258 13626
rect 32950 13574 33002 13626
rect 33014 13574 33066 13626
rect 33078 13574 33130 13626
rect 33142 13574 33194 13626
rect 33206 13574 33258 13626
rect 42950 13574 43002 13626
rect 43014 13574 43066 13626
rect 43078 13574 43130 13626
rect 43142 13574 43194 13626
rect 43206 13574 43258 13626
rect 27804 13472 27856 13524
rect 33968 13472 34020 13524
rect 27344 13336 27396 13388
rect 27804 13336 27856 13388
rect 28448 13336 28500 13388
rect 34888 13379 34940 13388
rect 34888 13345 34897 13379
rect 34897 13345 34931 13379
rect 34931 13345 34940 13379
rect 34888 13336 34940 13345
rect 37648 13336 37700 13388
rect 25412 13268 25464 13320
rect 28908 13268 28960 13320
rect 33508 13268 33560 13320
rect 37096 13268 37148 13320
rect 37280 13268 37332 13320
rect 38292 13268 38344 13320
rect 40592 13311 40644 13320
rect 40592 13277 40601 13311
rect 40601 13277 40635 13311
rect 40635 13277 40644 13311
rect 40592 13268 40644 13277
rect 44824 13268 44876 13320
rect 25780 13175 25832 13184
rect 25780 13141 25789 13175
rect 25789 13141 25823 13175
rect 25823 13141 25832 13175
rect 25780 13132 25832 13141
rect 33692 13200 33744 13252
rect 31760 13132 31812 13184
rect 32588 13132 32640 13184
rect 34244 13175 34296 13184
rect 34244 13141 34253 13175
rect 34253 13141 34287 13175
rect 34287 13141 34296 13175
rect 34244 13132 34296 13141
rect 34704 13132 34756 13184
rect 36544 13200 36596 13252
rect 37372 13243 37424 13252
rect 37372 13209 37381 13243
rect 37381 13209 37415 13243
rect 37415 13209 37424 13243
rect 37372 13200 37424 13209
rect 49148 13243 49200 13252
rect 49148 13209 49157 13243
rect 49157 13209 49191 13243
rect 49191 13209 49200 13243
rect 49148 13200 49200 13209
rect 39856 13132 39908 13184
rect 46756 13132 46808 13184
rect 7950 13030 8002 13082
rect 8014 13030 8066 13082
rect 8078 13030 8130 13082
rect 8142 13030 8194 13082
rect 8206 13030 8258 13082
rect 17950 13030 18002 13082
rect 18014 13030 18066 13082
rect 18078 13030 18130 13082
rect 18142 13030 18194 13082
rect 18206 13030 18258 13082
rect 27950 13030 28002 13082
rect 28014 13030 28066 13082
rect 28078 13030 28130 13082
rect 28142 13030 28194 13082
rect 28206 13030 28258 13082
rect 37950 13030 38002 13082
rect 38014 13030 38066 13082
rect 38078 13030 38130 13082
rect 38142 13030 38194 13082
rect 38206 13030 38258 13082
rect 47950 13030 48002 13082
rect 48014 13030 48066 13082
rect 48078 13030 48130 13082
rect 48142 13030 48194 13082
rect 48206 13030 48258 13082
rect 27528 12928 27580 12980
rect 29276 12971 29328 12980
rect 29276 12937 29285 12971
rect 29285 12937 29319 12971
rect 29319 12937 29328 12971
rect 29276 12928 29328 12937
rect 30288 12928 30340 12980
rect 30564 12928 30616 12980
rect 26516 12860 26568 12912
rect 28356 12860 28408 12912
rect 32404 12860 32456 12912
rect 28448 12792 28500 12844
rect 34796 12928 34848 12980
rect 35440 12971 35492 12980
rect 35440 12937 35449 12971
rect 35449 12937 35483 12971
rect 35483 12937 35492 12971
rect 35440 12928 35492 12937
rect 33968 12903 34020 12912
rect 33968 12869 33977 12903
rect 33977 12869 34011 12903
rect 34011 12869 34020 12903
rect 33968 12860 34020 12869
rect 34704 12860 34756 12912
rect 37280 12928 37332 12980
rect 29552 12724 29604 12776
rect 27160 12656 27212 12708
rect 30012 12699 30064 12708
rect 30012 12665 30021 12699
rect 30021 12665 30055 12699
rect 30055 12665 30064 12699
rect 30012 12656 30064 12665
rect 25228 12588 25280 12640
rect 34336 12724 34388 12776
rect 43720 12903 43772 12912
rect 43720 12869 43729 12903
rect 43729 12869 43763 12903
rect 43763 12869 43772 12903
rect 43720 12860 43772 12869
rect 46756 12792 46808 12844
rect 49148 12767 49200 12776
rect 49148 12733 49157 12767
rect 49157 12733 49191 12767
rect 49191 12733 49200 12767
rect 49148 12724 49200 12733
rect 36084 12656 36136 12708
rect 36820 12656 36872 12708
rect 44732 12656 44784 12708
rect 39948 12588 40000 12640
rect 2950 12486 3002 12538
rect 3014 12486 3066 12538
rect 3078 12486 3130 12538
rect 3142 12486 3194 12538
rect 3206 12486 3258 12538
rect 12950 12486 13002 12538
rect 13014 12486 13066 12538
rect 13078 12486 13130 12538
rect 13142 12486 13194 12538
rect 13206 12486 13258 12538
rect 22950 12486 23002 12538
rect 23014 12486 23066 12538
rect 23078 12486 23130 12538
rect 23142 12486 23194 12538
rect 23206 12486 23258 12538
rect 32950 12486 33002 12538
rect 33014 12486 33066 12538
rect 33078 12486 33130 12538
rect 33142 12486 33194 12538
rect 33206 12486 33258 12538
rect 42950 12486 43002 12538
rect 43014 12486 43066 12538
rect 43078 12486 43130 12538
rect 43142 12486 43194 12538
rect 43206 12486 43258 12538
rect 3332 12316 3384 12368
rect 9496 12316 9548 12368
rect 39856 12248 39908 12300
rect 28908 12180 28960 12232
rect 38936 12223 38988 12232
rect 38936 12189 38945 12223
rect 38945 12189 38979 12223
rect 38979 12189 38988 12223
rect 38936 12180 38988 12189
rect 41236 12223 41288 12232
rect 41236 12189 41245 12223
rect 41245 12189 41279 12223
rect 41279 12189 41288 12223
rect 41236 12180 41288 12189
rect 44732 12180 44784 12232
rect 29184 12112 29236 12164
rect 41880 12112 41932 12164
rect 49148 12155 49200 12164
rect 49148 12121 49157 12155
rect 49157 12121 49191 12155
rect 49191 12121 49200 12155
rect 49148 12112 49200 12121
rect 43352 12044 43404 12096
rect 44272 12087 44324 12096
rect 44272 12053 44281 12087
rect 44281 12053 44315 12087
rect 44315 12053 44324 12087
rect 44272 12044 44324 12053
rect 7950 11942 8002 11994
rect 8014 11942 8066 11994
rect 8078 11942 8130 11994
rect 8142 11942 8194 11994
rect 8206 11942 8258 11994
rect 17950 11942 18002 11994
rect 18014 11942 18066 11994
rect 18078 11942 18130 11994
rect 18142 11942 18194 11994
rect 18206 11942 18258 11994
rect 27950 11942 28002 11994
rect 28014 11942 28066 11994
rect 28078 11942 28130 11994
rect 28142 11942 28194 11994
rect 28206 11942 28258 11994
rect 37950 11942 38002 11994
rect 38014 11942 38066 11994
rect 38078 11942 38130 11994
rect 38142 11942 38194 11994
rect 38206 11942 38258 11994
rect 47950 11942 48002 11994
rect 48014 11942 48066 11994
rect 48078 11942 48130 11994
rect 48142 11942 48194 11994
rect 48206 11942 48258 11994
rect 44180 11772 44232 11824
rect 41328 11704 41380 11756
rect 42708 11704 42760 11756
rect 42800 11636 42852 11688
rect 45652 11568 45704 11620
rect 46848 11568 46900 11620
rect 44180 11500 44232 11552
rect 46388 11543 46440 11552
rect 46388 11509 46397 11543
rect 46397 11509 46431 11543
rect 46431 11509 46440 11543
rect 46388 11500 46440 11509
rect 2950 11398 3002 11450
rect 3014 11398 3066 11450
rect 3078 11398 3130 11450
rect 3142 11398 3194 11450
rect 3206 11398 3258 11450
rect 12950 11398 13002 11450
rect 13014 11398 13066 11450
rect 13078 11398 13130 11450
rect 13142 11398 13194 11450
rect 13206 11398 13258 11450
rect 22950 11398 23002 11450
rect 23014 11398 23066 11450
rect 23078 11398 23130 11450
rect 23142 11398 23194 11450
rect 23206 11398 23258 11450
rect 32950 11398 33002 11450
rect 33014 11398 33066 11450
rect 33078 11398 33130 11450
rect 33142 11398 33194 11450
rect 33206 11398 33258 11450
rect 42950 11398 43002 11450
rect 43014 11398 43066 11450
rect 43078 11398 43130 11450
rect 43142 11398 43194 11450
rect 43206 11398 43258 11450
rect 17868 11296 17920 11348
rect 19708 11160 19760 11212
rect 44272 11092 44324 11144
rect 49148 11135 49200 11144
rect 49148 11101 49157 11135
rect 49157 11101 49191 11135
rect 49191 11101 49200 11135
rect 49148 11092 49200 11101
rect 7564 11024 7616 11076
rect 44364 11024 44416 11076
rect 46480 11067 46532 11076
rect 46480 11033 46489 11067
rect 46489 11033 46523 11067
rect 46523 11033 46532 11067
rect 46480 11024 46532 11033
rect 7950 10854 8002 10906
rect 8014 10854 8066 10906
rect 8078 10854 8130 10906
rect 8142 10854 8194 10906
rect 8206 10854 8258 10906
rect 17950 10854 18002 10906
rect 18014 10854 18066 10906
rect 18078 10854 18130 10906
rect 18142 10854 18194 10906
rect 18206 10854 18258 10906
rect 27950 10854 28002 10906
rect 28014 10854 28066 10906
rect 28078 10854 28130 10906
rect 28142 10854 28194 10906
rect 28206 10854 28258 10906
rect 37950 10854 38002 10906
rect 38014 10854 38066 10906
rect 38078 10854 38130 10906
rect 38142 10854 38194 10906
rect 38206 10854 38258 10906
rect 47950 10854 48002 10906
rect 48014 10854 48066 10906
rect 48078 10854 48130 10906
rect 48142 10854 48194 10906
rect 48206 10854 48258 10906
rect 24216 10684 24268 10736
rect 39948 10616 40000 10668
rect 47584 10616 47636 10668
rect 49148 10591 49200 10600
rect 49148 10557 49157 10591
rect 49157 10557 49191 10591
rect 49191 10557 49200 10591
rect 49148 10548 49200 10557
rect 25136 10480 25188 10532
rect 42708 10412 42760 10464
rect 2950 10310 3002 10362
rect 3014 10310 3066 10362
rect 3078 10310 3130 10362
rect 3142 10310 3194 10362
rect 3206 10310 3258 10362
rect 12950 10310 13002 10362
rect 13014 10310 13066 10362
rect 13078 10310 13130 10362
rect 13142 10310 13194 10362
rect 13206 10310 13258 10362
rect 22950 10310 23002 10362
rect 23014 10310 23066 10362
rect 23078 10310 23130 10362
rect 23142 10310 23194 10362
rect 23206 10310 23258 10362
rect 32950 10310 33002 10362
rect 33014 10310 33066 10362
rect 33078 10310 33130 10362
rect 33142 10310 33194 10362
rect 33206 10310 33258 10362
rect 42950 10310 43002 10362
rect 43014 10310 43066 10362
rect 43078 10310 43130 10362
rect 43142 10310 43194 10362
rect 43206 10310 43258 10362
rect 28540 10004 28592 10056
rect 31852 10047 31904 10056
rect 31852 10013 31861 10047
rect 31861 10013 31895 10047
rect 31895 10013 31904 10047
rect 31852 10004 31904 10013
rect 45652 10004 45704 10056
rect 30104 9936 30156 9988
rect 49148 9979 49200 9988
rect 49148 9945 49157 9979
rect 49157 9945 49191 9979
rect 49191 9945 49200 9979
rect 49148 9936 49200 9945
rect 29920 9868 29972 9920
rect 7950 9766 8002 9818
rect 8014 9766 8066 9818
rect 8078 9766 8130 9818
rect 8142 9766 8194 9818
rect 8206 9766 8258 9818
rect 17950 9766 18002 9818
rect 18014 9766 18066 9818
rect 18078 9766 18130 9818
rect 18142 9766 18194 9818
rect 18206 9766 18258 9818
rect 27950 9766 28002 9818
rect 28014 9766 28066 9818
rect 28078 9766 28130 9818
rect 28142 9766 28194 9818
rect 28206 9766 28258 9818
rect 37950 9766 38002 9818
rect 38014 9766 38066 9818
rect 38078 9766 38130 9818
rect 38142 9766 38194 9818
rect 38206 9766 38258 9818
rect 47950 9766 48002 9818
rect 48014 9766 48066 9818
rect 48078 9766 48130 9818
rect 48142 9766 48194 9818
rect 48206 9766 48258 9818
rect 31944 9596 31996 9648
rect 34980 9596 35032 9648
rect 44180 9528 44232 9580
rect 46848 9528 46900 9580
rect 47768 9460 47820 9512
rect 48688 9460 48740 9512
rect 49148 9503 49200 9512
rect 49148 9469 49157 9503
rect 49157 9469 49191 9503
rect 49191 9469 49200 9503
rect 49148 9460 49200 9469
rect 33968 9392 34020 9444
rect 37280 9392 37332 9444
rect 47768 9324 47820 9376
rect 2950 9222 3002 9274
rect 3014 9222 3066 9274
rect 3078 9222 3130 9274
rect 3142 9222 3194 9274
rect 3206 9222 3258 9274
rect 12950 9222 13002 9274
rect 13014 9222 13066 9274
rect 13078 9222 13130 9274
rect 13142 9222 13194 9274
rect 13206 9222 13258 9274
rect 22950 9222 23002 9274
rect 23014 9222 23066 9274
rect 23078 9222 23130 9274
rect 23142 9222 23194 9274
rect 23206 9222 23258 9274
rect 32950 9222 33002 9274
rect 33014 9222 33066 9274
rect 33078 9222 33130 9274
rect 33142 9222 33194 9274
rect 33206 9222 33258 9274
rect 42950 9222 43002 9274
rect 43014 9222 43066 9274
rect 43078 9222 43130 9274
rect 43142 9222 43194 9274
rect 43206 9222 43258 9274
rect 3332 9052 3384 9104
rect 9404 9052 9456 9104
rect 43352 8916 43404 8968
rect 47676 8916 47728 8968
rect 46204 8891 46256 8900
rect 46204 8857 46213 8891
rect 46213 8857 46247 8891
rect 46247 8857 46256 8891
rect 46204 8848 46256 8857
rect 47124 8848 47176 8900
rect 48412 8848 48464 8900
rect 48688 8891 48740 8900
rect 48688 8857 48697 8891
rect 48697 8857 48731 8891
rect 48731 8857 48740 8891
rect 48688 8848 48740 8857
rect 47860 8780 47912 8832
rect 7950 8678 8002 8730
rect 8014 8678 8066 8730
rect 8078 8678 8130 8730
rect 8142 8678 8194 8730
rect 8206 8678 8258 8730
rect 17950 8678 18002 8730
rect 18014 8678 18066 8730
rect 18078 8678 18130 8730
rect 18142 8678 18194 8730
rect 18206 8678 18258 8730
rect 27950 8678 28002 8730
rect 28014 8678 28066 8730
rect 28078 8678 28130 8730
rect 28142 8678 28194 8730
rect 28206 8678 28258 8730
rect 37950 8678 38002 8730
rect 38014 8678 38066 8730
rect 38078 8678 38130 8730
rect 38142 8678 38194 8730
rect 38206 8678 38258 8730
rect 47950 8678 48002 8730
rect 48014 8678 48066 8730
rect 48078 8678 48130 8730
rect 48142 8678 48194 8730
rect 48206 8678 48258 8730
rect 5540 8508 5592 8560
rect 16488 8508 16540 8560
rect 19248 8508 19300 8560
rect 32312 8508 32364 8560
rect 37832 8551 37884 8560
rect 37832 8517 37841 8551
rect 37841 8517 37875 8551
rect 37875 8517 37884 8551
rect 37832 8508 37884 8517
rect 42708 8508 42760 8560
rect 18604 8440 18656 8492
rect 46480 8440 46532 8492
rect 23388 8372 23440 8424
rect 42616 8372 42668 8424
rect 49148 8415 49200 8424
rect 49148 8381 49157 8415
rect 49157 8381 49191 8415
rect 49191 8381 49200 8415
rect 49148 8372 49200 8381
rect 16488 8304 16540 8356
rect 37648 8304 37700 8356
rect 45928 8347 45980 8356
rect 45928 8313 45937 8347
rect 45937 8313 45971 8347
rect 45971 8313 45980 8347
rect 45928 8304 45980 8313
rect 2950 8134 3002 8186
rect 3014 8134 3066 8186
rect 3078 8134 3130 8186
rect 3142 8134 3194 8186
rect 3206 8134 3258 8186
rect 12950 8134 13002 8186
rect 13014 8134 13066 8186
rect 13078 8134 13130 8186
rect 13142 8134 13194 8186
rect 13206 8134 13258 8186
rect 22950 8134 23002 8186
rect 23014 8134 23066 8186
rect 23078 8134 23130 8186
rect 23142 8134 23194 8186
rect 23206 8134 23258 8186
rect 32950 8134 33002 8186
rect 33014 8134 33066 8186
rect 33078 8134 33130 8186
rect 33142 8134 33194 8186
rect 33206 8134 33258 8186
rect 42950 8134 43002 8186
rect 43014 8134 43066 8186
rect 43078 8134 43130 8186
rect 43142 8134 43194 8186
rect 43206 8134 43258 8186
rect 46388 7828 46440 7880
rect 49148 7803 49200 7812
rect 49148 7769 49157 7803
rect 49157 7769 49191 7803
rect 49191 7769 49200 7803
rect 49148 7760 49200 7769
rect 7950 7590 8002 7642
rect 8014 7590 8066 7642
rect 8078 7590 8130 7642
rect 8142 7590 8194 7642
rect 8206 7590 8258 7642
rect 17950 7590 18002 7642
rect 18014 7590 18066 7642
rect 18078 7590 18130 7642
rect 18142 7590 18194 7642
rect 18206 7590 18258 7642
rect 27950 7590 28002 7642
rect 28014 7590 28066 7642
rect 28078 7590 28130 7642
rect 28142 7590 28194 7642
rect 28206 7590 28258 7642
rect 37950 7590 38002 7642
rect 38014 7590 38066 7642
rect 38078 7590 38130 7642
rect 38142 7590 38194 7642
rect 38206 7590 38258 7642
rect 47950 7590 48002 7642
rect 48014 7590 48066 7642
rect 48078 7590 48130 7642
rect 48142 7590 48194 7642
rect 48206 7590 48258 7642
rect 31760 7420 31812 7472
rect 29644 7352 29696 7404
rect 47768 7352 47820 7404
rect 41420 7284 41472 7336
rect 49148 7327 49200 7336
rect 49148 7293 49157 7327
rect 49157 7293 49191 7327
rect 49191 7293 49200 7327
rect 49148 7284 49200 7293
rect 45192 7216 45244 7268
rect 47584 7216 47636 7268
rect 47768 7216 47820 7268
rect 2950 7046 3002 7098
rect 3014 7046 3066 7098
rect 3078 7046 3130 7098
rect 3142 7046 3194 7098
rect 3206 7046 3258 7098
rect 12950 7046 13002 7098
rect 13014 7046 13066 7098
rect 13078 7046 13130 7098
rect 13142 7046 13194 7098
rect 13206 7046 13258 7098
rect 22950 7046 23002 7098
rect 23014 7046 23066 7098
rect 23078 7046 23130 7098
rect 23142 7046 23194 7098
rect 23206 7046 23258 7098
rect 32950 7046 33002 7098
rect 33014 7046 33066 7098
rect 33078 7046 33130 7098
rect 33142 7046 33194 7098
rect 33206 7046 33258 7098
rect 42950 7046 43002 7098
rect 43014 7046 43066 7098
rect 43078 7046 43130 7098
rect 43142 7046 43194 7098
rect 43206 7046 43258 7098
rect 36820 6740 36872 6792
rect 32404 6672 32456 6724
rect 40132 6740 40184 6792
rect 45928 6740 45980 6792
rect 44456 6672 44508 6724
rect 49148 6715 49200 6724
rect 49148 6681 49157 6715
rect 49157 6681 49191 6715
rect 49191 6681 49200 6715
rect 49148 6672 49200 6681
rect 3424 6604 3476 6656
rect 8944 6604 8996 6656
rect 7950 6502 8002 6554
rect 8014 6502 8066 6554
rect 8078 6502 8130 6554
rect 8142 6502 8194 6554
rect 8206 6502 8258 6554
rect 17950 6502 18002 6554
rect 18014 6502 18066 6554
rect 18078 6502 18130 6554
rect 18142 6502 18194 6554
rect 18206 6502 18258 6554
rect 27950 6502 28002 6554
rect 28014 6502 28066 6554
rect 28078 6502 28130 6554
rect 28142 6502 28194 6554
rect 28206 6502 28258 6554
rect 37950 6502 38002 6554
rect 38014 6502 38066 6554
rect 38078 6502 38130 6554
rect 38142 6502 38194 6554
rect 38206 6502 38258 6554
rect 47950 6502 48002 6554
rect 48014 6502 48066 6554
rect 48078 6502 48130 6554
rect 48142 6502 48194 6554
rect 48206 6502 48258 6554
rect 2950 5958 3002 6010
rect 3014 5958 3066 6010
rect 3078 5958 3130 6010
rect 3142 5958 3194 6010
rect 3206 5958 3258 6010
rect 12950 5958 13002 6010
rect 13014 5958 13066 6010
rect 13078 5958 13130 6010
rect 13142 5958 13194 6010
rect 13206 5958 13258 6010
rect 22950 5958 23002 6010
rect 23014 5958 23066 6010
rect 23078 5958 23130 6010
rect 23142 5958 23194 6010
rect 23206 5958 23258 6010
rect 32950 5958 33002 6010
rect 33014 5958 33066 6010
rect 33078 5958 33130 6010
rect 33142 5958 33194 6010
rect 33206 5958 33258 6010
rect 42950 5958 43002 6010
rect 43014 5958 43066 6010
rect 43078 5958 43130 6010
rect 43142 5958 43194 6010
rect 43206 5958 43258 6010
rect 46204 5652 46256 5704
rect 49148 5695 49200 5704
rect 49148 5661 49157 5695
rect 49157 5661 49191 5695
rect 49191 5661 49200 5695
rect 49148 5652 49200 5661
rect 7950 5414 8002 5466
rect 8014 5414 8066 5466
rect 8078 5414 8130 5466
rect 8142 5414 8194 5466
rect 8206 5414 8258 5466
rect 17950 5414 18002 5466
rect 18014 5414 18066 5466
rect 18078 5414 18130 5466
rect 18142 5414 18194 5466
rect 18206 5414 18258 5466
rect 27950 5414 28002 5466
rect 28014 5414 28066 5466
rect 28078 5414 28130 5466
rect 28142 5414 28194 5466
rect 28206 5414 28258 5466
rect 37950 5414 38002 5466
rect 38014 5414 38066 5466
rect 38078 5414 38130 5466
rect 38142 5414 38194 5466
rect 38206 5414 38258 5466
rect 47950 5414 48002 5466
rect 48014 5414 48066 5466
rect 48078 5414 48130 5466
rect 48142 5414 48194 5466
rect 48206 5414 48258 5466
rect 3424 5244 3476 5296
rect 9036 5244 9088 5296
rect 29460 5015 29512 5024
rect 29460 4981 29469 5015
rect 29469 4981 29503 5015
rect 29503 4981 29512 5015
rect 29460 4972 29512 4981
rect 47768 4972 47820 5024
rect 49332 5015 49384 5024
rect 49332 4981 49341 5015
rect 49341 4981 49375 5015
rect 49375 4981 49384 5015
rect 49332 4972 49384 4981
rect 2950 4870 3002 4922
rect 3014 4870 3066 4922
rect 3078 4870 3130 4922
rect 3142 4870 3194 4922
rect 3206 4870 3258 4922
rect 12950 4870 13002 4922
rect 13014 4870 13066 4922
rect 13078 4870 13130 4922
rect 13142 4870 13194 4922
rect 13206 4870 13258 4922
rect 22950 4870 23002 4922
rect 23014 4870 23066 4922
rect 23078 4870 23130 4922
rect 23142 4870 23194 4922
rect 23206 4870 23258 4922
rect 32950 4870 33002 4922
rect 33014 4870 33066 4922
rect 33078 4870 33130 4922
rect 33142 4870 33194 4922
rect 33206 4870 33258 4922
rect 42950 4870 43002 4922
rect 43014 4870 43066 4922
rect 43078 4870 43130 4922
rect 43142 4870 43194 4922
rect 43206 4870 43258 4922
rect 10048 4768 10100 4820
rect 29460 4768 29512 4820
rect 24768 4564 24820 4616
rect 49148 4539 49200 4548
rect 49148 4505 49157 4539
rect 49157 4505 49191 4539
rect 49191 4505 49200 4539
rect 49148 4496 49200 4505
rect 7950 4326 8002 4378
rect 8014 4326 8066 4378
rect 8078 4326 8130 4378
rect 8142 4326 8194 4378
rect 8206 4326 8258 4378
rect 17950 4326 18002 4378
rect 18014 4326 18066 4378
rect 18078 4326 18130 4378
rect 18142 4326 18194 4378
rect 18206 4326 18258 4378
rect 27950 4326 28002 4378
rect 28014 4326 28066 4378
rect 28078 4326 28130 4378
rect 28142 4326 28194 4378
rect 28206 4326 28258 4378
rect 37950 4326 38002 4378
rect 38014 4326 38066 4378
rect 38078 4326 38130 4378
rect 38142 4326 38194 4378
rect 38206 4326 38258 4378
rect 47950 4326 48002 4378
rect 48014 4326 48066 4378
rect 48078 4326 48130 4378
rect 48142 4326 48194 4378
rect 48206 4326 48258 4378
rect 33968 4131 34020 4140
rect 33968 4097 33977 4131
rect 33977 4097 34011 4131
rect 34011 4097 34020 4131
rect 33968 4088 34020 4097
rect 38476 4088 38528 4140
rect 40132 4088 40184 4140
rect 46020 4131 46072 4140
rect 46020 4097 46029 4131
rect 46029 4097 46063 4131
rect 46063 4097 46072 4131
rect 46020 4088 46072 4097
rect 48596 4088 48648 4140
rect 33876 4020 33928 4072
rect 39028 4020 39080 4072
rect 43444 4020 43496 4072
rect 36544 3952 36596 4004
rect 46020 3952 46072 4004
rect 48872 3995 48924 4004
rect 48872 3961 48881 3995
rect 48881 3961 48915 3995
rect 48915 3961 48924 3995
rect 48872 3952 48924 3961
rect 47768 3884 47820 3936
rect 2950 3782 3002 3834
rect 3014 3782 3066 3834
rect 3078 3782 3130 3834
rect 3142 3782 3194 3834
rect 3206 3782 3258 3834
rect 12950 3782 13002 3834
rect 13014 3782 13066 3834
rect 13078 3782 13130 3834
rect 13142 3782 13194 3834
rect 13206 3782 13258 3834
rect 22950 3782 23002 3834
rect 23014 3782 23066 3834
rect 23078 3782 23130 3834
rect 23142 3782 23194 3834
rect 23206 3782 23258 3834
rect 32950 3782 33002 3834
rect 33014 3782 33066 3834
rect 33078 3782 33130 3834
rect 33142 3782 33194 3834
rect 33206 3782 33258 3834
rect 42950 3782 43002 3834
rect 43014 3782 43066 3834
rect 43078 3782 43130 3834
rect 43142 3782 43194 3834
rect 43206 3782 43258 3834
rect 5540 3680 5592 3732
rect 18328 3612 18380 3664
rect 26884 3612 26936 3664
rect 24308 3544 24360 3596
rect 29460 3544 29512 3596
rect 30932 3544 30984 3596
rect 34612 3544 34664 3596
rect 36084 3544 36136 3596
rect 39764 3544 39816 3596
rect 41236 3544 41288 3596
rect 44180 3544 44232 3596
rect 2780 3476 2832 3528
rect 25780 3476 25832 3528
rect 29736 3519 29788 3528
rect 29736 3485 29745 3519
rect 29745 3485 29779 3519
rect 29779 3485 29788 3519
rect 29736 3476 29788 3485
rect 30104 3476 30156 3528
rect 34244 3476 34296 3528
rect 36728 3519 36780 3528
rect 36728 3485 36737 3519
rect 36737 3485 36771 3519
rect 36771 3485 36780 3519
rect 36728 3476 36780 3485
rect 37280 3476 37332 3528
rect 41880 3519 41932 3528
rect 41880 3485 41889 3519
rect 41889 3485 41923 3519
rect 41923 3485 41932 3519
rect 41880 3476 41932 3485
rect 45192 3519 45244 3528
rect 45192 3485 45201 3519
rect 45201 3485 45235 3519
rect 45235 3485 45244 3519
rect 45192 3476 45244 3485
rect 47676 3476 47728 3528
rect 49332 3408 49384 3460
rect 12900 3340 12952 3392
rect 26792 3340 26844 3392
rect 7950 3238 8002 3290
rect 8014 3238 8066 3290
rect 8078 3238 8130 3290
rect 8142 3238 8194 3290
rect 8206 3238 8258 3290
rect 17950 3238 18002 3290
rect 18014 3238 18066 3290
rect 18078 3238 18130 3290
rect 18142 3238 18194 3290
rect 18206 3238 18258 3290
rect 27950 3238 28002 3290
rect 28014 3238 28066 3290
rect 28078 3238 28130 3290
rect 28142 3238 28194 3290
rect 28206 3238 28258 3290
rect 37950 3238 38002 3290
rect 38014 3238 38066 3290
rect 38078 3238 38130 3290
rect 38142 3238 38194 3290
rect 38206 3238 38258 3290
rect 47950 3238 48002 3290
rect 48014 3238 48066 3290
rect 48078 3238 48130 3290
rect 48142 3238 48194 3290
rect 48206 3238 48258 3290
rect 14464 3136 14516 3188
rect 7564 3068 7616 3120
rect 1492 3000 1544 3052
rect 756 2932 808 2984
rect 3700 3000 3752 3052
rect 5172 3000 5224 3052
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 6644 3000 6696 3052
rect 10324 3000 10376 3052
rect 12532 3000 12584 3052
rect 12900 3111 12952 3120
rect 12900 3077 12909 3111
rect 12909 3077 12943 3111
rect 12943 3077 12952 3111
rect 12900 3068 12952 3077
rect 19984 3136 20036 3188
rect 14004 3000 14056 3052
rect 18420 3068 18472 3120
rect 17684 3000 17736 3052
rect 18328 3000 18380 3052
rect 30564 3136 30616 3188
rect 47124 3179 47176 3188
rect 47124 3145 47133 3179
rect 47133 3145 47167 3179
rect 47167 3145 47176 3179
rect 47124 3136 47176 3145
rect 25596 3068 25648 3120
rect 37372 3068 37424 3120
rect 24676 3000 24728 3052
rect 25136 3043 25188 3052
rect 25136 3009 25145 3043
rect 25145 3009 25179 3043
rect 25179 3009 25188 3043
rect 25136 3000 25188 3009
rect 29092 3000 29144 3052
rect 29184 3043 29236 3052
rect 29184 3009 29193 3043
rect 29193 3009 29227 3043
rect 29227 3009 29236 3043
rect 29184 3000 29236 3009
rect 32036 3000 32088 3052
rect 34152 3043 34204 3052
rect 34152 3009 34161 3043
rect 34161 3009 34195 3043
rect 34195 3009 34204 3043
rect 34152 3000 34204 3009
rect 37648 3043 37700 3052
rect 37648 3009 37657 3043
rect 37657 3009 37691 3043
rect 37691 3009 37700 3043
rect 37648 3000 37700 3009
rect 47860 3068 47912 3120
rect 42616 3043 42668 3052
rect 42616 3009 42625 3043
rect 42625 3009 42659 3043
rect 42659 3009 42668 3043
rect 42616 3000 42668 3009
rect 44456 3043 44508 3052
rect 44456 3009 44465 3043
rect 44465 3009 44499 3043
rect 44499 3009 44508 3043
rect 44456 3000 44508 3009
rect 47124 3000 47176 3052
rect 19156 2932 19208 2984
rect 17224 2864 17276 2916
rect 18788 2864 18840 2916
rect 20628 2975 20680 2984
rect 20628 2941 20637 2975
rect 20637 2941 20671 2975
rect 20671 2941 20680 2975
rect 20628 2932 20680 2941
rect 22100 2932 22152 2984
rect 23572 2932 23624 2984
rect 25044 2932 25096 2984
rect 27252 2932 27304 2984
rect 28724 2932 28776 2984
rect 31668 2932 31720 2984
rect 28356 2864 28408 2916
rect 32404 2864 32456 2916
rect 36820 2932 36872 2984
rect 37556 2864 37608 2916
rect 41972 2932 42024 2984
rect 42708 2864 42760 2916
rect 47860 2932 47912 2984
rect 46388 2796 46440 2848
rect 48320 2796 48372 2848
rect 2950 2694 3002 2746
rect 3014 2694 3066 2746
rect 3078 2694 3130 2746
rect 3142 2694 3194 2746
rect 3206 2694 3258 2746
rect 12950 2694 13002 2746
rect 13014 2694 13066 2746
rect 13078 2694 13130 2746
rect 13142 2694 13194 2746
rect 13206 2694 13258 2746
rect 22950 2694 23002 2746
rect 23014 2694 23066 2746
rect 23078 2694 23130 2746
rect 23142 2694 23194 2746
rect 23206 2694 23258 2746
rect 32950 2694 33002 2746
rect 33014 2694 33066 2746
rect 33078 2694 33130 2746
rect 33142 2694 33194 2746
rect 33206 2694 33258 2746
rect 42950 2694 43002 2746
rect 43014 2694 43066 2746
rect 43078 2694 43130 2746
rect 43142 2694 43194 2746
rect 43206 2694 43258 2746
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 11152 2592 11204 2644
rect 13636 2635 13688 2644
rect 13636 2601 13645 2635
rect 13645 2601 13679 2635
rect 13679 2601 13688 2635
rect 13636 2592 13688 2601
rect 18696 2592 18748 2644
rect 27804 2592 27856 2644
rect 46020 2592 46072 2644
rect 27712 2524 27764 2576
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 18420 2456 18472 2508
rect 21364 2456 21416 2508
rect 22836 2456 22888 2508
rect 25780 2499 25832 2508
rect 25780 2465 25789 2499
rect 25789 2465 25823 2499
rect 25823 2465 25832 2499
rect 25780 2456 25832 2465
rect 26516 2456 26568 2508
rect 28356 2456 28408 2508
rect 30288 2456 30340 2508
rect 35348 2456 35400 2508
rect 38292 2456 38344 2508
rect 40592 2456 40644 2508
rect 48320 2499 48372 2508
rect 48320 2465 48329 2499
rect 48329 2465 48363 2499
rect 48363 2465 48372 2499
rect 48320 2456 48372 2465
rect 2228 2388 2280 2440
rect 7380 2388 7432 2440
rect 9588 2388 9640 2440
rect 14740 2388 14792 2440
rect 2964 2320 3016 2372
rect 4436 2320 4488 2372
rect 4988 2363 5040 2372
rect 4988 2329 4997 2363
rect 4997 2329 5031 2363
rect 5031 2329 5040 2363
rect 4988 2320 5040 2329
rect 5908 2320 5960 2372
rect 6000 2363 6052 2372
rect 6000 2329 6009 2363
rect 6009 2329 6043 2363
rect 6043 2329 6052 2363
rect 6000 2320 6052 2329
rect 7840 2320 7892 2372
rect 8852 2320 8904 2372
rect 11060 2320 11112 2372
rect 11796 2320 11848 2372
rect 13268 2320 13320 2372
rect 15476 2320 15528 2372
rect 16212 2320 16264 2372
rect 16304 2363 16356 2372
rect 16304 2329 16313 2363
rect 16313 2329 16347 2363
rect 16347 2329 16356 2363
rect 16304 2320 16356 2329
rect 16948 2320 17000 2372
rect 19892 2388 19944 2440
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 25228 2431 25280 2440
rect 25228 2397 25237 2431
rect 25237 2397 25271 2431
rect 25271 2397 25280 2431
rect 25228 2388 25280 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29920 2431 29972 2440
rect 29920 2397 29929 2431
rect 29929 2397 29963 2431
rect 29963 2397 29972 2431
rect 29920 2388 29972 2397
rect 32220 2388 32272 2440
rect 33784 2388 33836 2440
rect 35256 2388 35308 2440
rect 40040 2431 40092 2440
rect 40040 2397 40049 2431
rect 40049 2397 40083 2431
rect 40083 2397 40092 2431
rect 40040 2388 40092 2397
rect 41420 2388 41472 2440
rect 47768 2431 47820 2440
rect 47768 2397 47777 2431
rect 47777 2397 47811 2431
rect 47811 2397 47820 2431
rect 47768 2388 47820 2397
rect 2412 2295 2464 2304
rect 2412 2261 2421 2295
rect 2421 2261 2455 2295
rect 2455 2261 2464 2295
rect 2412 2252 2464 2261
rect 3332 2295 3384 2304
rect 3332 2261 3341 2295
rect 3341 2261 3375 2295
rect 3375 2261 3384 2295
rect 3332 2252 3384 2261
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 17316 2252 17368 2304
rect 17408 2295 17460 2304
rect 17408 2261 17417 2295
rect 17417 2261 17451 2295
rect 17451 2261 17460 2295
rect 17408 2252 17460 2261
rect 29276 2320 29328 2372
rect 28816 2252 28868 2304
rect 33140 2252 33192 2304
rect 45652 2320 45704 2372
rect 7950 2150 8002 2202
rect 8014 2150 8066 2202
rect 8078 2150 8130 2202
rect 8142 2150 8194 2202
rect 8206 2150 8258 2202
rect 17950 2150 18002 2202
rect 18014 2150 18066 2202
rect 18078 2150 18130 2202
rect 18142 2150 18194 2202
rect 18206 2150 18258 2202
rect 27950 2150 28002 2202
rect 28014 2150 28066 2202
rect 28078 2150 28130 2202
rect 28142 2150 28194 2202
rect 28206 2150 28258 2202
rect 37950 2150 38002 2202
rect 38014 2150 38066 2202
rect 38078 2150 38130 2202
rect 38142 2150 38194 2202
rect 38206 2150 38258 2202
rect 47950 2150 48002 2202
rect 48014 2150 48066 2202
rect 48078 2150 48130 2202
rect 48142 2150 48194 2202
rect 48206 2150 48258 2202
rect 16304 2048 16356 2100
rect 28448 2048 28500 2100
rect 6000 1980 6052 2032
rect 17132 1980 17184 2032
rect 7564 1912 7616 1964
rect 23756 1980 23808 2032
rect 17316 1912 17368 1964
rect 26792 1912 26844 1964
rect 2412 1844 2464 1896
rect 17408 1844 17460 1896
rect 28632 1844 28684 1896
rect 19524 1776 19576 1828
rect 8484 1708 8536 1760
rect 22284 1708 22336 1760
rect 3332 1640 3384 1692
rect 20720 1640 20772 1692
rect 17132 1572 17184 1624
rect 25320 1572 25372 1624
<< metal2 >>
rect 386 56200 442 57000
rect 1122 56200 1178 57000
rect 1858 56200 1914 57000
rect 2594 56200 2650 57000
rect 3330 56200 3386 57000
rect 4066 56200 4122 57000
rect 4802 56200 4858 57000
rect 5538 56200 5594 57000
rect 6274 56200 6330 57000
rect 7010 56200 7066 57000
rect 7746 56200 7802 57000
rect 8482 56200 8538 57000
rect 9218 56200 9274 57000
rect 9954 56200 10010 57000
rect 10690 56200 10746 57000
rect 11426 56200 11482 57000
rect 12162 56200 12218 57000
rect 12898 56200 12954 57000
rect 13634 56200 13690 57000
rect 14370 56200 14426 57000
rect 15106 56200 15162 57000
rect 15842 56200 15898 57000
rect 16578 56200 16634 57000
rect 17314 56200 17370 57000
rect 18050 56200 18106 57000
rect 18156 56222 18368 56250
rect 400 55758 428 56200
rect 388 55752 440 55758
rect 388 55694 440 55700
rect 940 53100 992 53106
rect 940 53042 992 53048
rect 952 52737 980 53042
rect 938 52728 994 52737
rect 938 52663 994 52672
rect 1136 52562 1164 56200
rect 1872 53650 1900 56200
rect 1860 53644 1912 53650
rect 1860 53586 1912 53592
rect 2608 53038 2636 56200
rect 2872 55752 2924 55758
rect 2872 55694 2924 55700
rect 2778 55040 2834 55049
rect 2778 54975 2834 54984
rect 2792 54194 2820 54975
rect 2780 54188 2832 54194
rect 2780 54130 2832 54136
rect 2596 53032 2648 53038
rect 2596 52974 2648 52980
rect 1676 52896 1728 52902
rect 1676 52838 1728 52844
rect 1124 52556 1176 52562
rect 1124 52498 1176 52504
rect 1584 52012 1636 52018
rect 1584 51954 1636 51960
rect 940 50924 992 50930
rect 940 50866 992 50872
rect 952 50425 980 50866
rect 938 50416 994 50425
rect 938 50351 994 50360
rect 938 48104 994 48113
rect 938 48039 940 48048
rect 992 48039 994 48048
rect 940 48010 992 48016
rect 940 45892 992 45898
rect 940 45834 992 45840
rect 952 45801 980 45834
rect 938 45792 994 45801
rect 938 45727 994 45736
rect 940 43784 992 43790
rect 940 43726 992 43732
rect 952 43489 980 43726
rect 938 43480 994 43489
rect 938 43415 994 43424
rect 1596 42090 1624 51954
rect 1688 43330 1716 52838
rect 2884 52086 2912 55694
rect 3344 54262 3372 56200
rect 3332 54256 3384 54262
rect 3332 54198 3384 54204
rect 3976 53984 4028 53990
rect 3976 53926 4028 53932
rect 2950 53884 3258 53893
rect 2950 53882 2956 53884
rect 3012 53882 3036 53884
rect 3092 53882 3116 53884
rect 3172 53882 3196 53884
rect 3252 53882 3258 53884
rect 3012 53830 3014 53882
rect 3194 53830 3196 53882
rect 2950 53828 2956 53830
rect 3012 53828 3036 53830
rect 3092 53828 3116 53830
rect 3172 53828 3196 53830
rect 3252 53828 3258 53830
rect 2950 53819 3258 53828
rect 2950 52796 3258 52805
rect 2950 52794 2956 52796
rect 3012 52794 3036 52796
rect 3092 52794 3116 52796
rect 3172 52794 3196 52796
rect 3252 52794 3258 52796
rect 3012 52742 3014 52794
rect 3194 52742 3196 52794
rect 2950 52740 2956 52742
rect 3012 52740 3036 52742
rect 3092 52740 3116 52742
rect 3172 52740 3196 52742
rect 3252 52740 3258 52742
rect 2950 52731 3258 52740
rect 2872 52080 2924 52086
rect 2872 52022 2924 52028
rect 2950 51708 3258 51717
rect 2950 51706 2956 51708
rect 3012 51706 3036 51708
rect 3092 51706 3116 51708
rect 3172 51706 3196 51708
rect 3252 51706 3258 51708
rect 3012 51654 3014 51706
rect 3194 51654 3196 51706
rect 2950 51652 2956 51654
rect 3012 51652 3036 51654
rect 3092 51652 3116 51654
rect 3172 51652 3196 51654
rect 3252 51652 3258 51654
rect 2950 51643 3258 51652
rect 1952 50788 2004 50794
rect 1952 50730 2004 50736
rect 1860 48068 1912 48074
rect 1860 48010 1912 48016
rect 1768 45824 1820 45830
rect 1768 45766 1820 45772
rect 1780 45626 1808 45766
rect 1768 45620 1820 45626
rect 1768 45562 1820 45568
rect 1688 43302 1808 43330
rect 1584 42084 1636 42090
rect 1584 42026 1636 42032
rect 1676 41540 1728 41546
rect 1676 41482 1728 41488
rect 1688 41177 1716 41482
rect 1674 41168 1730 41177
rect 1674 41103 1730 41112
rect 1780 41070 1808 43302
rect 1768 41064 1820 41070
rect 1768 41006 1820 41012
rect 1872 39302 1900 48010
rect 1860 39296 1912 39302
rect 1860 39238 1912 39244
rect 1964 38962 1992 50730
rect 2950 50620 3258 50629
rect 2950 50618 2956 50620
rect 3012 50618 3036 50620
rect 3092 50618 3116 50620
rect 3172 50618 3196 50620
rect 3252 50618 3258 50620
rect 3012 50566 3014 50618
rect 3194 50566 3196 50618
rect 2950 50564 2956 50566
rect 3012 50564 3036 50566
rect 3092 50564 3116 50566
rect 3172 50564 3196 50566
rect 3252 50564 3258 50566
rect 2950 50555 3258 50564
rect 2950 49532 3258 49541
rect 2950 49530 2956 49532
rect 3012 49530 3036 49532
rect 3092 49530 3116 49532
rect 3172 49530 3196 49532
rect 3252 49530 3258 49532
rect 3012 49478 3014 49530
rect 3194 49478 3196 49530
rect 2950 49476 2956 49478
rect 3012 49476 3036 49478
rect 3092 49476 3116 49478
rect 3172 49476 3196 49478
rect 3252 49476 3258 49478
rect 2950 49467 3258 49476
rect 2950 48444 3258 48453
rect 2950 48442 2956 48444
rect 3012 48442 3036 48444
rect 3092 48442 3116 48444
rect 3172 48442 3196 48444
rect 3252 48442 3258 48444
rect 3012 48390 3014 48442
rect 3194 48390 3196 48442
rect 2950 48388 2956 48390
rect 3012 48388 3036 48390
rect 3092 48388 3116 48390
rect 3172 48388 3196 48390
rect 3252 48388 3258 48390
rect 2950 48379 3258 48388
rect 3988 48074 4016 53926
rect 4080 52562 4108 56200
rect 4816 55214 4844 56200
rect 4816 55186 4936 55214
rect 4908 53038 4936 55186
rect 5552 53650 5580 56200
rect 6288 54262 6316 56200
rect 6276 54256 6328 54262
rect 6276 54198 6328 54204
rect 7024 53650 7052 56200
rect 5540 53644 5592 53650
rect 5540 53586 5592 53592
rect 7012 53644 7064 53650
rect 7012 53586 7064 53592
rect 6368 53508 6420 53514
rect 6368 53450 6420 53456
rect 6276 53168 6328 53174
rect 6276 53110 6328 53116
rect 4896 53032 4948 53038
rect 4896 52974 4948 52980
rect 5816 52624 5868 52630
rect 5816 52566 5868 52572
rect 4068 52556 4120 52562
rect 4068 52498 4120 52504
rect 3976 48068 4028 48074
rect 3976 48010 4028 48016
rect 2950 47356 3258 47365
rect 2950 47354 2956 47356
rect 3012 47354 3036 47356
rect 3092 47354 3116 47356
rect 3172 47354 3196 47356
rect 3252 47354 3258 47356
rect 3012 47302 3014 47354
rect 3194 47302 3196 47354
rect 2950 47300 2956 47302
rect 3012 47300 3036 47302
rect 3092 47300 3116 47302
rect 3172 47300 3196 47302
rect 3252 47300 3258 47302
rect 2950 47291 3258 47300
rect 2950 46268 3258 46277
rect 2950 46266 2956 46268
rect 3012 46266 3036 46268
rect 3092 46266 3116 46268
rect 3172 46266 3196 46268
rect 3252 46266 3258 46268
rect 3012 46214 3014 46266
rect 3194 46214 3196 46266
rect 2950 46212 2956 46214
rect 3012 46212 3036 46214
rect 3092 46212 3116 46214
rect 3172 46212 3196 46214
rect 3252 46212 3258 46214
rect 2950 46203 3258 46212
rect 2950 45180 3258 45189
rect 2950 45178 2956 45180
rect 3012 45178 3036 45180
rect 3092 45178 3116 45180
rect 3172 45178 3196 45180
rect 3252 45178 3258 45180
rect 3012 45126 3014 45178
rect 3194 45126 3196 45178
rect 2950 45124 2956 45126
rect 3012 45124 3036 45126
rect 3092 45124 3116 45126
rect 3172 45124 3196 45126
rect 3252 45124 3258 45126
rect 2950 45115 3258 45124
rect 2950 44092 3258 44101
rect 2950 44090 2956 44092
rect 3012 44090 3036 44092
rect 3092 44090 3116 44092
rect 3172 44090 3196 44092
rect 3252 44090 3258 44092
rect 3012 44038 3014 44090
rect 3194 44038 3196 44090
rect 2950 44036 2956 44038
rect 3012 44036 3036 44038
rect 3092 44036 3116 44038
rect 3172 44036 3196 44038
rect 3252 44036 3258 44038
rect 2950 44027 3258 44036
rect 2044 43648 2096 43654
rect 2044 43590 2096 43596
rect 2056 43450 2084 43590
rect 2044 43444 2096 43450
rect 2044 43386 2096 43392
rect 2950 43004 3258 43013
rect 2950 43002 2956 43004
rect 3012 43002 3036 43004
rect 3092 43002 3116 43004
rect 3172 43002 3196 43004
rect 3252 43002 3258 43004
rect 3012 42950 3014 43002
rect 3194 42950 3196 43002
rect 2950 42948 2956 42950
rect 3012 42948 3036 42950
rect 3092 42948 3116 42950
rect 3172 42948 3196 42950
rect 3252 42948 3258 42950
rect 2950 42939 3258 42948
rect 2950 41916 3258 41925
rect 2950 41914 2956 41916
rect 3012 41914 3036 41916
rect 3092 41914 3116 41916
rect 3172 41914 3196 41916
rect 3252 41914 3258 41916
rect 3012 41862 3014 41914
rect 3194 41862 3196 41914
rect 2950 41860 2956 41862
rect 3012 41860 3036 41862
rect 3092 41860 3116 41862
rect 3172 41860 3196 41862
rect 3252 41860 3258 41862
rect 2950 41851 3258 41860
rect 5828 41274 5856 52566
rect 6288 42294 6316 53110
rect 6380 42362 6408 53450
rect 7760 53038 7788 56200
rect 7950 54428 8258 54437
rect 7950 54426 7956 54428
rect 8012 54426 8036 54428
rect 8092 54426 8116 54428
rect 8172 54426 8196 54428
rect 8252 54426 8258 54428
rect 8012 54374 8014 54426
rect 8194 54374 8196 54426
rect 7950 54372 7956 54374
rect 8012 54372 8036 54374
rect 8092 54372 8116 54374
rect 8172 54372 8196 54374
rect 8252 54372 8258 54374
rect 7950 54363 8258 54372
rect 8496 54262 8524 56200
rect 8484 54256 8536 54262
rect 8484 54198 8536 54204
rect 8944 53576 8996 53582
rect 8944 53518 8996 53524
rect 7950 53340 8258 53349
rect 7950 53338 7956 53340
rect 8012 53338 8036 53340
rect 8092 53338 8116 53340
rect 8172 53338 8196 53340
rect 8252 53338 8258 53340
rect 8012 53286 8014 53338
rect 8194 53286 8196 53338
rect 7950 53284 7956 53286
rect 8012 53284 8036 53286
rect 8092 53284 8116 53286
rect 8172 53284 8196 53286
rect 8252 53284 8258 53286
rect 7950 53275 8258 53284
rect 7748 53032 7800 53038
rect 7748 52974 7800 52980
rect 7950 52252 8258 52261
rect 7950 52250 7956 52252
rect 8012 52250 8036 52252
rect 8092 52250 8116 52252
rect 8172 52250 8196 52252
rect 8252 52250 8258 52252
rect 8012 52198 8014 52250
rect 8194 52198 8196 52250
rect 7950 52196 7956 52198
rect 8012 52196 8036 52198
rect 8092 52196 8116 52198
rect 8172 52196 8196 52198
rect 8252 52196 8258 52198
rect 7950 52187 8258 52196
rect 7950 51164 8258 51173
rect 7950 51162 7956 51164
rect 8012 51162 8036 51164
rect 8092 51162 8116 51164
rect 8172 51162 8196 51164
rect 8252 51162 8258 51164
rect 8012 51110 8014 51162
rect 8194 51110 8196 51162
rect 7950 51108 7956 51110
rect 8012 51108 8036 51110
rect 8092 51108 8116 51110
rect 8172 51108 8196 51110
rect 8252 51108 8258 51110
rect 7950 51099 8258 51108
rect 7950 50076 8258 50085
rect 7950 50074 7956 50076
rect 8012 50074 8036 50076
rect 8092 50074 8116 50076
rect 8172 50074 8196 50076
rect 8252 50074 8258 50076
rect 8012 50022 8014 50074
rect 8194 50022 8196 50074
rect 7950 50020 7956 50022
rect 8012 50020 8036 50022
rect 8092 50020 8116 50022
rect 8172 50020 8196 50022
rect 8252 50020 8258 50022
rect 7950 50011 8258 50020
rect 7950 48988 8258 48997
rect 7950 48986 7956 48988
rect 8012 48986 8036 48988
rect 8092 48986 8116 48988
rect 8172 48986 8196 48988
rect 8252 48986 8258 48988
rect 8012 48934 8014 48986
rect 8194 48934 8196 48986
rect 7950 48932 7956 48934
rect 8012 48932 8036 48934
rect 8092 48932 8116 48934
rect 8172 48932 8196 48934
rect 8252 48932 8258 48934
rect 7950 48923 8258 48932
rect 7950 47900 8258 47909
rect 7950 47898 7956 47900
rect 8012 47898 8036 47900
rect 8092 47898 8116 47900
rect 8172 47898 8196 47900
rect 8252 47898 8258 47900
rect 8012 47846 8014 47898
rect 8194 47846 8196 47898
rect 7950 47844 7956 47846
rect 8012 47844 8036 47846
rect 8092 47844 8116 47846
rect 8172 47844 8196 47846
rect 8252 47844 8258 47846
rect 7950 47835 8258 47844
rect 7950 46812 8258 46821
rect 7950 46810 7956 46812
rect 8012 46810 8036 46812
rect 8092 46810 8116 46812
rect 8172 46810 8196 46812
rect 8252 46810 8258 46812
rect 8012 46758 8014 46810
rect 8194 46758 8196 46810
rect 7950 46756 7956 46758
rect 8012 46756 8036 46758
rect 8092 46756 8116 46758
rect 8172 46756 8196 46758
rect 8252 46756 8258 46758
rect 7950 46747 8258 46756
rect 7950 45724 8258 45733
rect 7950 45722 7956 45724
rect 8012 45722 8036 45724
rect 8092 45722 8116 45724
rect 8172 45722 8196 45724
rect 8252 45722 8258 45724
rect 8012 45670 8014 45722
rect 8194 45670 8196 45722
rect 7950 45668 7956 45670
rect 8012 45668 8036 45670
rect 8092 45668 8116 45670
rect 8172 45668 8196 45670
rect 8252 45668 8258 45670
rect 7950 45659 8258 45668
rect 7950 44636 8258 44645
rect 7950 44634 7956 44636
rect 8012 44634 8036 44636
rect 8092 44634 8116 44636
rect 8172 44634 8196 44636
rect 8252 44634 8258 44636
rect 8012 44582 8014 44634
rect 8194 44582 8196 44634
rect 7950 44580 7956 44582
rect 8012 44580 8036 44582
rect 8092 44580 8116 44582
rect 8172 44580 8196 44582
rect 8252 44580 8258 44582
rect 7950 44571 8258 44580
rect 7950 43548 8258 43557
rect 7950 43546 7956 43548
rect 8012 43546 8036 43548
rect 8092 43546 8116 43548
rect 8172 43546 8196 43548
rect 8252 43546 8258 43548
rect 8012 43494 8014 43546
rect 8194 43494 8196 43546
rect 7950 43492 7956 43494
rect 8012 43492 8036 43494
rect 8092 43492 8116 43494
rect 8172 43492 8196 43494
rect 8252 43492 8258 43494
rect 7950 43483 8258 43492
rect 8956 43450 8984 53518
rect 9232 52630 9260 56200
rect 9864 53168 9916 53174
rect 9864 53110 9916 53116
rect 9772 53100 9824 53106
rect 9772 53042 9824 53048
rect 9220 52624 9272 52630
rect 9220 52566 9272 52572
rect 9220 52488 9272 52494
rect 9220 52430 9272 52436
rect 8944 43444 8996 43450
rect 8944 43386 8996 43392
rect 7950 42460 8258 42469
rect 7950 42458 7956 42460
rect 8012 42458 8036 42460
rect 8092 42458 8116 42460
rect 8172 42458 8196 42460
rect 8252 42458 8258 42460
rect 8012 42406 8014 42458
rect 8194 42406 8196 42458
rect 7950 42404 7956 42406
rect 8012 42404 8036 42406
rect 8092 42404 8116 42406
rect 8172 42404 8196 42406
rect 8252 42404 8258 42406
rect 7950 42395 8258 42404
rect 9232 42362 9260 52430
rect 9784 44538 9812 53042
rect 9772 44532 9824 44538
rect 9772 44474 9824 44480
rect 6368 42356 6420 42362
rect 6368 42298 6420 42304
rect 9220 42356 9272 42362
rect 9220 42298 9272 42304
rect 6276 42288 6328 42294
rect 6276 42230 6328 42236
rect 7196 42220 7248 42226
rect 7196 42162 7248 42168
rect 9128 42220 9180 42226
rect 9128 42162 9180 42168
rect 5816 41268 5868 41274
rect 5816 41210 5868 41216
rect 5724 41132 5776 41138
rect 5724 41074 5776 41080
rect 2950 40828 3258 40837
rect 2950 40826 2956 40828
rect 3012 40826 3036 40828
rect 3092 40826 3116 40828
rect 3172 40826 3196 40828
rect 3252 40826 3258 40828
rect 3012 40774 3014 40826
rect 3194 40774 3196 40826
rect 2950 40772 2956 40774
rect 3012 40772 3036 40774
rect 3092 40772 3116 40774
rect 3172 40772 3196 40774
rect 3252 40772 3258 40774
rect 2950 40763 3258 40772
rect 2950 39740 3258 39749
rect 2950 39738 2956 39740
rect 3012 39738 3036 39740
rect 3092 39738 3116 39740
rect 3172 39738 3196 39740
rect 3252 39738 3258 39740
rect 3012 39686 3014 39738
rect 3194 39686 3196 39738
rect 2950 39684 2956 39686
rect 3012 39684 3036 39686
rect 3092 39684 3116 39686
rect 3172 39684 3196 39686
rect 3252 39684 3258 39686
rect 2950 39675 3258 39684
rect 940 38956 992 38962
rect 940 38898 992 38904
rect 1952 38956 2004 38962
rect 1952 38898 2004 38904
rect 952 38865 980 38898
rect 938 38856 994 38865
rect 938 38791 994 38800
rect 2950 38652 3258 38661
rect 2950 38650 2956 38652
rect 3012 38650 3036 38652
rect 3092 38650 3116 38652
rect 3172 38650 3196 38652
rect 3252 38650 3258 38652
rect 3012 38598 3014 38650
rect 3194 38598 3196 38650
rect 2950 38596 2956 38598
rect 3012 38596 3036 38598
rect 3092 38596 3116 38598
rect 3172 38596 3196 38598
rect 3252 38596 3258 38598
rect 2950 38587 3258 38596
rect 2950 37564 3258 37573
rect 2950 37562 2956 37564
rect 3012 37562 3036 37564
rect 3092 37562 3116 37564
rect 3172 37562 3196 37564
rect 3252 37562 3258 37564
rect 3012 37510 3014 37562
rect 3194 37510 3196 37562
rect 2950 37508 2956 37510
rect 3012 37508 3036 37510
rect 3092 37508 3116 37510
rect 3172 37508 3196 37510
rect 3252 37508 3258 37510
rect 2950 37499 3258 37508
rect 940 36780 992 36786
rect 940 36722 992 36728
rect 952 36553 980 36722
rect 938 36544 994 36553
rect 938 36479 994 36488
rect 2950 36476 3258 36485
rect 2950 36474 2956 36476
rect 3012 36474 3036 36476
rect 3092 36474 3116 36476
rect 3172 36474 3196 36476
rect 3252 36474 3258 36476
rect 3012 36422 3014 36474
rect 3194 36422 3196 36474
rect 2950 36420 2956 36422
rect 3012 36420 3036 36422
rect 3092 36420 3116 36422
rect 3172 36420 3196 36422
rect 3252 36420 3258 36422
rect 2950 36411 3258 36420
rect 2950 35388 3258 35397
rect 2950 35386 2956 35388
rect 3012 35386 3036 35388
rect 3092 35386 3116 35388
rect 3172 35386 3196 35388
rect 3252 35386 3258 35388
rect 3012 35334 3014 35386
rect 3194 35334 3196 35386
rect 2950 35332 2956 35334
rect 3012 35332 3036 35334
rect 3092 35332 3116 35334
rect 3172 35332 3196 35334
rect 3252 35332 3258 35334
rect 2950 35323 3258 35332
rect 1768 34604 1820 34610
rect 1768 34546 1820 34552
rect 1780 34241 1808 34546
rect 2950 34300 3258 34309
rect 2950 34298 2956 34300
rect 3012 34298 3036 34300
rect 3092 34298 3116 34300
rect 3172 34298 3196 34300
rect 3252 34298 3258 34300
rect 3012 34246 3014 34298
rect 3194 34246 3196 34298
rect 2950 34244 2956 34246
rect 3012 34244 3036 34246
rect 3092 34244 3116 34246
rect 3172 34244 3196 34246
rect 3252 34244 3258 34246
rect 1766 34232 1822 34241
rect 2950 34235 3258 34244
rect 1766 34167 1822 34176
rect 2950 33212 3258 33221
rect 2950 33210 2956 33212
rect 3012 33210 3036 33212
rect 3092 33210 3116 33212
rect 3172 33210 3196 33212
rect 3252 33210 3258 33212
rect 3012 33158 3014 33210
rect 3194 33158 3196 33210
rect 2950 33156 2956 33158
rect 3012 33156 3036 33158
rect 3092 33156 3116 33158
rect 3172 33156 3196 33158
rect 3252 33156 3258 33158
rect 2950 33147 3258 33156
rect 940 32428 992 32434
rect 940 32370 992 32376
rect 952 31929 980 32370
rect 5736 32366 5764 41074
rect 5724 32360 5776 32366
rect 5724 32302 5776 32308
rect 2950 32124 3258 32133
rect 2950 32122 2956 32124
rect 3012 32122 3036 32124
rect 3092 32122 3116 32124
rect 3172 32122 3196 32124
rect 3252 32122 3258 32124
rect 3012 32070 3014 32122
rect 3194 32070 3196 32122
rect 2950 32068 2956 32070
rect 3012 32068 3036 32070
rect 3092 32068 3116 32070
rect 3172 32068 3196 32070
rect 3252 32068 3258 32070
rect 2950 32059 3258 32068
rect 938 31920 994 31929
rect 938 31855 994 31864
rect 2950 31036 3258 31045
rect 2950 31034 2956 31036
rect 3012 31034 3036 31036
rect 3092 31034 3116 31036
rect 3172 31034 3196 31036
rect 3252 31034 3258 31036
rect 3012 30982 3014 31034
rect 3194 30982 3196 31034
rect 2950 30980 2956 30982
rect 3012 30980 3036 30982
rect 3092 30980 3116 30982
rect 3172 30980 3196 30982
rect 3252 30980 3258 30982
rect 2950 30971 3258 30980
rect 2950 29948 3258 29957
rect 2950 29946 2956 29948
rect 3012 29946 3036 29948
rect 3092 29946 3116 29948
rect 3172 29946 3196 29948
rect 3252 29946 3258 29948
rect 3012 29894 3014 29946
rect 3194 29894 3196 29946
rect 2950 29892 2956 29894
rect 3012 29892 3036 29894
rect 3092 29892 3116 29894
rect 3172 29892 3196 29894
rect 3252 29892 3258 29894
rect 2950 29883 3258 29892
rect 1308 29708 1360 29714
rect 1308 29650 1360 29656
rect 1320 29617 1348 29650
rect 4896 29640 4948 29646
rect 1306 29608 1362 29617
rect 4896 29582 4948 29588
rect 1306 29543 1362 29552
rect 2950 28860 3258 28869
rect 2950 28858 2956 28860
rect 3012 28858 3036 28860
rect 3092 28858 3116 28860
rect 3172 28858 3196 28860
rect 3252 28858 3258 28860
rect 3012 28806 3014 28858
rect 3194 28806 3196 28858
rect 2950 28804 2956 28806
rect 3012 28804 3036 28806
rect 3092 28804 3116 28806
rect 3172 28804 3196 28806
rect 3252 28804 3258 28806
rect 2950 28795 3258 28804
rect 4908 28218 4936 29582
rect 7208 28558 7236 42162
rect 7950 41372 8258 41381
rect 7950 41370 7956 41372
rect 8012 41370 8036 41372
rect 8092 41370 8116 41372
rect 8172 41370 8196 41372
rect 8252 41370 8258 41372
rect 8012 41318 8014 41370
rect 8194 41318 8196 41370
rect 7950 41316 7956 41318
rect 8012 41316 8036 41318
rect 8092 41316 8116 41318
rect 8172 41316 8196 41318
rect 8252 41316 8258 41318
rect 7950 41307 8258 41316
rect 7950 40284 8258 40293
rect 7950 40282 7956 40284
rect 8012 40282 8036 40284
rect 8092 40282 8116 40284
rect 8172 40282 8196 40284
rect 8252 40282 8258 40284
rect 8012 40230 8014 40282
rect 8194 40230 8196 40282
rect 7950 40228 7956 40230
rect 8012 40228 8036 40230
rect 8092 40228 8116 40230
rect 8172 40228 8196 40230
rect 8252 40228 8258 40230
rect 7950 40219 8258 40228
rect 7950 39196 8258 39205
rect 7950 39194 7956 39196
rect 8012 39194 8036 39196
rect 8092 39194 8116 39196
rect 8172 39194 8196 39196
rect 8252 39194 8258 39196
rect 8012 39142 8014 39194
rect 8194 39142 8196 39194
rect 7950 39140 7956 39142
rect 8012 39140 8036 39142
rect 8092 39140 8116 39142
rect 8172 39140 8196 39142
rect 8252 39140 8258 39142
rect 7950 39131 8258 39140
rect 7380 38752 7432 38758
rect 7380 38694 7432 38700
rect 7392 30258 7420 38694
rect 7950 38108 8258 38117
rect 7950 38106 7956 38108
rect 8012 38106 8036 38108
rect 8092 38106 8116 38108
rect 8172 38106 8196 38108
rect 8252 38106 8258 38108
rect 8012 38054 8014 38106
rect 8194 38054 8196 38106
rect 7950 38052 7956 38054
rect 8012 38052 8036 38054
rect 8092 38052 8116 38054
rect 8172 38052 8196 38054
rect 8252 38052 8258 38054
rect 7950 38043 8258 38052
rect 7950 37020 8258 37029
rect 7950 37018 7956 37020
rect 8012 37018 8036 37020
rect 8092 37018 8116 37020
rect 8172 37018 8196 37020
rect 8252 37018 8258 37020
rect 8012 36966 8014 37018
rect 8194 36966 8196 37018
rect 7950 36964 7956 36966
rect 8012 36964 8036 36966
rect 8092 36964 8116 36966
rect 8172 36964 8196 36966
rect 8252 36964 8258 36966
rect 7950 36955 8258 36964
rect 7564 36576 7616 36582
rect 7564 36518 7616 36524
rect 7472 32224 7524 32230
rect 7472 32166 7524 32172
rect 7380 30252 7432 30258
rect 7380 30194 7432 30200
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 4896 28212 4948 28218
rect 4896 28154 4948 28160
rect 2950 27772 3258 27781
rect 2950 27770 2956 27772
rect 3012 27770 3036 27772
rect 3092 27770 3116 27772
rect 3172 27770 3196 27772
rect 3252 27770 3258 27772
rect 3012 27718 3014 27770
rect 3194 27718 3196 27770
rect 2950 27716 2956 27718
rect 3012 27716 3036 27718
rect 3092 27716 3116 27718
rect 3172 27716 3196 27718
rect 3252 27716 3258 27718
rect 2950 27707 3258 27716
rect 1308 27532 1360 27538
rect 1308 27474 1360 27480
rect 1320 27305 1348 27474
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 5448 27464 5500 27470
rect 5448 27406 5500 27412
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 2950 26684 3258 26693
rect 2950 26682 2956 26684
rect 3012 26682 3036 26684
rect 3092 26682 3116 26684
rect 3172 26682 3196 26684
rect 3252 26682 3258 26684
rect 3012 26630 3014 26682
rect 3194 26630 3196 26682
rect 2950 26628 2956 26630
rect 3012 26628 3036 26630
rect 3092 26628 3116 26630
rect 3172 26628 3196 26630
rect 3252 26628 3258 26630
rect 2950 26619 3258 26628
rect 2950 25596 3258 25605
rect 2950 25594 2956 25596
rect 3012 25594 3036 25596
rect 3092 25594 3116 25596
rect 3172 25594 3196 25596
rect 3252 25594 3258 25596
rect 3012 25542 3014 25594
rect 3194 25542 3196 25594
rect 2950 25540 2956 25542
rect 3012 25540 3036 25542
rect 3092 25540 3116 25542
rect 3172 25540 3196 25542
rect 3252 25540 3258 25542
rect 2950 25531 3258 25540
rect 4908 25498 4936 27406
rect 5460 26314 5488 27406
rect 4988 26308 5040 26314
rect 4988 26250 5040 26256
rect 5448 26308 5500 26314
rect 5448 26250 5500 26256
rect 4896 25492 4948 25498
rect 4896 25434 4948 25440
rect 1308 25356 1360 25362
rect 1308 25298 1360 25304
rect 1320 24993 1348 25298
rect 4160 25288 4212 25294
rect 4160 25230 4212 25236
rect 1306 24984 1362 24993
rect 1306 24919 1362 24928
rect 2950 24508 3258 24517
rect 2950 24506 2956 24508
rect 3012 24506 3036 24508
rect 3092 24506 3116 24508
rect 3172 24506 3196 24508
rect 3252 24506 3258 24508
rect 3012 24454 3014 24506
rect 3194 24454 3196 24506
rect 2950 24452 2956 24454
rect 3012 24452 3036 24454
rect 3092 24452 3116 24454
rect 3172 24452 3196 24454
rect 3252 24452 3258 24454
rect 2950 24443 3258 24452
rect 2950 23420 3258 23429
rect 2950 23418 2956 23420
rect 3012 23418 3036 23420
rect 3092 23418 3116 23420
rect 3172 23418 3196 23420
rect 3252 23418 3258 23420
rect 3012 23366 3014 23418
rect 3194 23366 3196 23418
rect 2950 23364 2956 23366
rect 3012 23364 3036 23366
rect 3092 23364 3116 23366
rect 3172 23364 3196 23366
rect 3252 23364 3258 23366
rect 2950 23355 3258 23364
rect 4172 23322 4200 25230
rect 4160 23316 4212 23322
rect 4160 23258 4212 23264
rect 1308 23180 1360 23186
rect 1308 23122 1360 23128
rect 1320 22681 1348 23122
rect 5000 23118 5028 26250
rect 7484 26234 7512 32166
rect 7576 28082 7604 36518
rect 7950 35932 8258 35941
rect 7950 35930 7956 35932
rect 8012 35930 8036 35932
rect 8092 35930 8116 35932
rect 8172 35930 8196 35932
rect 8252 35930 8258 35932
rect 8012 35878 8014 35930
rect 8194 35878 8196 35930
rect 7950 35876 7956 35878
rect 8012 35876 8036 35878
rect 8092 35876 8116 35878
rect 8172 35876 8196 35878
rect 8252 35876 8258 35878
rect 7950 35867 8258 35876
rect 7950 34844 8258 34853
rect 7950 34842 7956 34844
rect 8012 34842 8036 34844
rect 8092 34842 8116 34844
rect 8172 34842 8196 34844
rect 8252 34842 8258 34844
rect 8012 34790 8014 34842
rect 8194 34790 8196 34842
rect 7950 34788 7956 34790
rect 8012 34788 8036 34790
rect 8092 34788 8116 34790
rect 8172 34788 8196 34790
rect 8252 34788 8258 34790
rect 7950 34779 8258 34788
rect 7840 34740 7892 34746
rect 7840 34682 7892 34688
rect 7656 30184 7708 30190
rect 7656 30126 7708 30132
rect 7564 28076 7616 28082
rect 7564 28018 7616 28024
rect 7668 27606 7696 30126
rect 7748 28008 7800 28014
rect 7748 27950 7800 27956
rect 7656 27600 7708 27606
rect 7656 27542 7708 27548
rect 7760 26586 7788 27950
rect 7852 26994 7880 34682
rect 7950 33756 8258 33765
rect 7950 33754 7956 33756
rect 8012 33754 8036 33756
rect 8092 33754 8116 33756
rect 8172 33754 8196 33756
rect 8252 33754 8258 33756
rect 8012 33702 8014 33754
rect 8194 33702 8196 33754
rect 7950 33700 7956 33702
rect 8012 33700 8036 33702
rect 8092 33700 8116 33702
rect 8172 33700 8196 33702
rect 8252 33700 8258 33702
rect 7950 33691 8258 33700
rect 7950 32668 8258 32677
rect 7950 32666 7956 32668
rect 8012 32666 8036 32668
rect 8092 32666 8116 32668
rect 8172 32666 8196 32668
rect 8252 32666 8258 32668
rect 8012 32614 8014 32666
rect 8194 32614 8196 32666
rect 7950 32612 7956 32614
rect 8012 32612 8036 32614
rect 8092 32612 8116 32614
rect 8172 32612 8196 32614
rect 8252 32612 8258 32614
rect 7950 32603 8258 32612
rect 7950 31580 8258 31589
rect 7950 31578 7956 31580
rect 8012 31578 8036 31580
rect 8092 31578 8116 31580
rect 8172 31578 8196 31580
rect 8252 31578 8258 31580
rect 8012 31526 8014 31578
rect 8194 31526 8196 31578
rect 7950 31524 7956 31526
rect 8012 31524 8036 31526
rect 8092 31524 8116 31526
rect 8172 31524 8196 31526
rect 8252 31524 8258 31526
rect 7950 31515 8258 31524
rect 9140 30666 9168 42162
rect 9876 41274 9904 53110
rect 9968 53038 9996 56200
rect 10048 54324 10100 54330
rect 10048 54266 10100 54272
rect 9956 53032 10008 53038
rect 9956 52974 10008 52980
rect 10060 51610 10088 54266
rect 10704 53650 10732 56200
rect 11440 54262 11468 56200
rect 11428 54256 11480 54262
rect 11428 54198 11480 54204
rect 11704 54188 11756 54194
rect 11704 54130 11756 54136
rect 10692 53644 10744 53650
rect 10692 53586 10744 53592
rect 10416 53576 10468 53582
rect 10416 53518 10468 53524
rect 10048 51604 10100 51610
rect 10048 51546 10100 51552
rect 10428 45558 10456 53518
rect 10784 53508 10836 53514
rect 10784 53450 10836 53456
rect 10416 45552 10468 45558
rect 10416 45494 10468 45500
rect 10600 41472 10652 41478
rect 10600 41414 10652 41420
rect 9864 41268 9916 41274
rect 9864 41210 9916 41216
rect 9772 41132 9824 41138
rect 9772 41074 9824 41080
rect 9784 31249 9812 41074
rect 9770 31240 9826 31249
rect 9770 31175 9826 31184
rect 9128 30660 9180 30666
rect 9128 30602 9180 30608
rect 7950 30492 8258 30501
rect 7950 30490 7956 30492
rect 8012 30490 8036 30492
rect 8092 30490 8116 30492
rect 8172 30490 8196 30492
rect 8252 30490 8258 30492
rect 8012 30438 8014 30490
rect 8194 30438 8196 30490
rect 7950 30436 7956 30438
rect 8012 30436 8036 30438
rect 8092 30436 8116 30438
rect 8172 30436 8196 30438
rect 8252 30436 8258 30438
rect 7950 30427 8258 30436
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 7950 29404 8258 29413
rect 7950 29402 7956 29404
rect 8012 29402 8036 29404
rect 8092 29402 8116 29404
rect 8172 29402 8196 29404
rect 8252 29402 8258 29404
rect 8012 29350 8014 29402
rect 8194 29350 8196 29402
rect 7950 29348 7956 29350
rect 8012 29348 8036 29350
rect 8092 29348 8116 29350
rect 8172 29348 8196 29350
rect 8252 29348 8258 29350
rect 7950 29339 8258 29348
rect 7950 28316 8258 28325
rect 7950 28314 7956 28316
rect 8012 28314 8036 28316
rect 8092 28314 8116 28316
rect 8172 28314 8196 28316
rect 8252 28314 8258 28316
rect 8012 28262 8014 28314
rect 8194 28262 8196 28314
rect 7950 28260 7956 28262
rect 8012 28260 8036 28262
rect 8092 28260 8116 28262
rect 8172 28260 8196 28262
rect 8252 28260 8258 28262
rect 7950 28251 8258 28260
rect 7950 27228 8258 27237
rect 7950 27226 7956 27228
rect 8012 27226 8036 27228
rect 8092 27226 8116 27228
rect 8172 27226 8196 27228
rect 8252 27226 8258 27228
rect 8012 27174 8014 27226
rect 8194 27174 8196 27226
rect 7950 27172 7956 27174
rect 8012 27172 8036 27174
rect 8092 27172 8116 27174
rect 8172 27172 8196 27174
rect 8252 27172 8258 27174
rect 7950 27163 8258 27172
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 8300 26920 8352 26926
rect 8300 26862 8352 26868
rect 8944 26920 8996 26926
rect 8944 26862 8996 26868
rect 7748 26580 7800 26586
rect 7748 26522 7800 26528
rect 7748 26376 7800 26382
rect 7748 26318 7800 26324
rect 7760 26234 7788 26318
rect 7484 26206 7696 26234
rect 7760 26206 7880 26234
rect 7668 25906 7696 26206
rect 7656 25900 7708 25906
rect 7656 25842 7708 25848
rect 6276 25288 6328 25294
rect 6276 25230 6328 25236
rect 6288 23866 6316 25230
rect 7852 24070 7880 26206
rect 7950 26140 8258 26149
rect 7950 26138 7956 26140
rect 8012 26138 8036 26140
rect 8092 26138 8116 26140
rect 8172 26138 8196 26140
rect 8252 26138 8258 26140
rect 8012 26086 8014 26138
rect 8194 26086 8196 26138
rect 7950 26084 7956 26086
rect 8012 26084 8036 26086
rect 8092 26084 8116 26086
rect 8172 26084 8196 26086
rect 8252 26084 8258 26086
rect 7950 26075 8258 26084
rect 7950 25052 8258 25061
rect 7950 25050 7956 25052
rect 8012 25050 8036 25052
rect 8092 25050 8116 25052
rect 8172 25050 8196 25052
rect 8252 25050 8258 25052
rect 8012 24998 8014 25050
rect 8194 24998 8196 25050
rect 7950 24996 7956 24998
rect 8012 24996 8036 24998
rect 8092 24996 8116 24998
rect 8172 24996 8196 24998
rect 8252 24996 8258 24998
rect 7950 24987 8258 24996
rect 8312 24750 8340 26862
rect 8850 24984 8906 24993
rect 8850 24919 8906 24928
rect 8300 24744 8352 24750
rect 8300 24686 8352 24692
rect 7840 24064 7892 24070
rect 7840 24006 7892 24012
rect 6276 23860 6328 23866
rect 6276 23802 6328 23808
rect 7852 23662 7880 24006
rect 7950 23964 8258 23973
rect 7950 23962 7956 23964
rect 8012 23962 8036 23964
rect 8092 23962 8116 23964
rect 8172 23962 8196 23964
rect 8252 23962 8258 23964
rect 8012 23910 8014 23962
rect 8194 23910 8196 23962
rect 7950 23908 7956 23910
rect 8012 23908 8036 23910
rect 8092 23908 8116 23910
rect 8172 23908 8196 23910
rect 8252 23908 8258 23910
rect 7950 23899 8258 23908
rect 7840 23656 7892 23662
rect 7840 23598 7892 23604
rect 5540 23180 5592 23186
rect 5540 23122 5592 23128
rect 4988 23112 5040 23118
rect 4988 23054 5040 23060
rect 2780 22976 2832 22982
rect 2780 22918 2832 22924
rect 1306 22672 1362 22681
rect 1306 22607 1362 22616
rect 2792 20466 2820 22918
rect 2950 22332 3258 22341
rect 2950 22330 2956 22332
rect 3012 22330 3036 22332
rect 3092 22330 3116 22332
rect 3172 22330 3196 22332
rect 3252 22330 3258 22332
rect 3012 22278 3014 22330
rect 3194 22278 3196 22330
rect 2950 22276 2956 22278
rect 3012 22276 3036 22278
rect 3092 22276 3116 22278
rect 3172 22276 3196 22278
rect 3252 22276 3258 22278
rect 2950 22267 3258 22276
rect 5552 22166 5580 23122
rect 5540 22160 5592 22166
rect 5540 22102 5592 22108
rect 2950 21244 3258 21253
rect 2950 21242 2956 21244
rect 3012 21242 3036 21244
rect 3092 21242 3116 21244
rect 3172 21242 3196 21244
rect 3252 21242 3258 21244
rect 3012 21190 3014 21242
rect 3194 21190 3196 21242
rect 2950 21188 2956 21190
rect 3012 21188 3036 21190
rect 3092 21188 3116 21190
rect 3172 21188 3196 21190
rect 3252 21188 3258 21190
rect 2950 21179 3258 21188
rect 7852 20942 7880 23598
rect 7950 22876 8258 22885
rect 7950 22874 7956 22876
rect 8012 22874 8036 22876
rect 8092 22874 8116 22876
rect 8172 22874 8196 22876
rect 8252 22874 8258 22876
rect 8012 22822 8014 22874
rect 8194 22822 8196 22874
rect 7950 22820 7956 22822
rect 8012 22820 8036 22822
rect 8092 22820 8116 22822
rect 8172 22820 8196 22822
rect 8252 22820 8258 22822
rect 7950 22811 8258 22820
rect 7950 21788 8258 21797
rect 7950 21786 7956 21788
rect 8012 21786 8036 21788
rect 8092 21786 8116 21788
rect 8172 21786 8196 21788
rect 8252 21786 8258 21788
rect 8012 21734 8014 21786
rect 8194 21734 8196 21786
rect 7950 21732 7956 21734
rect 8012 21732 8036 21734
rect 8092 21732 8116 21734
rect 8172 21732 8196 21734
rect 8252 21732 8258 21734
rect 7950 21723 8258 21732
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2780 20460 2832 20466
rect 2780 20402 2832 20408
rect 1308 20392 1360 20398
rect 1306 20360 1308 20369
rect 1360 20360 1362 20369
rect 1306 20295 1362 20304
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 1308 18216 1360 18222
rect 1308 18158 1360 18164
rect 1320 18057 1348 18158
rect 1306 18048 1362 18057
rect 1306 17983 1362 17992
rect 2792 16114 2820 18566
rect 2884 18290 2912 20742
rect 7950 20700 8258 20709
rect 7950 20698 7956 20700
rect 8012 20698 8036 20700
rect 8092 20698 8116 20700
rect 8172 20698 8196 20700
rect 8252 20698 8258 20700
rect 8012 20646 8014 20698
rect 8194 20646 8196 20698
rect 7950 20644 7956 20646
rect 8012 20644 8036 20646
rect 8092 20644 8116 20646
rect 8172 20644 8196 20646
rect 8252 20644 8258 20646
rect 7950 20635 8258 20644
rect 2950 20156 3258 20165
rect 2950 20154 2956 20156
rect 3012 20154 3036 20156
rect 3092 20154 3116 20156
rect 3172 20154 3196 20156
rect 3252 20154 3258 20156
rect 3012 20102 3014 20154
rect 3194 20102 3196 20154
rect 2950 20100 2956 20102
rect 3012 20100 3036 20102
rect 3092 20100 3116 20102
rect 3172 20100 3196 20102
rect 3252 20100 3258 20102
rect 2950 20091 3258 20100
rect 7950 19612 8258 19621
rect 7950 19610 7956 19612
rect 8012 19610 8036 19612
rect 8092 19610 8116 19612
rect 8172 19610 8196 19612
rect 8252 19610 8258 19612
rect 8012 19558 8014 19610
rect 8194 19558 8196 19610
rect 7950 19556 7956 19558
rect 8012 19556 8036 19558
rect 8092 19556 8116 19558
rect 8172 19556 8196 19558
rect 8252 19556 8258 19558
rect 7950 19547 8258 19556
rect 2950 19068 3258 19077
rect 2950 19066 2956 19068
rect 3012 19066 3036 19068
rect 3092 19066 3116 19068
rect 3172 19066 3196 19068
rect 3252 19066 3258 19068
rect 3012 19014 3014 19066
rect 3194 19014 3196 19066
rect 2950 19012 2956 19014
rect 3012 19012 3036 19014
rect 3092 19012 3116 19014
rect 3172 19012 3196 19014
rect 3252 19012 3258 19014
rect 2950 19003 3258 19012
rect 7950 18524 8258 18533
rect 7950 18522 7956 18524
rect 8012 18522 8036 18524
rect 8092 18522 8116 18524
rect 8172 18522 8196 18524
rect 8252 18522 8258 18524
rect 8012 18470 8014 18522
rect 8194 18470 8196 18522
rect 7950 18468 7956 18470
rect 8012 18468 8036 18470
rect 8092 18468 8116 18470
rect 8172 18468 8196 18470
rect 8252 18468 8258 18470
rect 7950 18459 8258 18468
rect 2872 18284 2924 18290
rect 2872 18226 2924 18232
rect 2950 17980 3258 17989
rect 2950 17978 2956 17980
rect 3012 17978 3036 17980
rect 3092 17978 3116 17980
rect 3172 17978 3196 17980
rect 3252 17978 3258 17980
rect 3012 17926 3014 17978
rect 3194 17926 3196 17978
rect 2950 17924 2956 17926
rect 3012 17924 3036 17926
rect 3092 17924 3116 17926
rect 3172 17924 3196 17926
rect 3252 17924 3258 17926
rect 2950 17915 3258 17924
rect 7950 17436 8258 17445
rect 7950 17434 7956 17436
rect 8012 17434 8036 17436
rect 8092 17434 8116 17436
rect 8172 17434 8196 17436
rect 8252 17434 8258 17436
rect 8012 17382 8014 17434
rect 8194 17382 8196 17434
rect 7950 17380 7956 17382
rect 8012 17380 8036 17382
rect 8092 17380 8116 17382
rect 8172 17380 8196 17382
rect 8252 17380 8258 17382
rect 7950 17371 8258 17380
rect 2950 16892 3258 16901
rect 2950 16890 2956 16892
rect 3012 16890 3036 16892
rect 3092 16890 3116 16892
rect 3172 16890 3196 16892
rect 3252 16890 3258 16892
rect 3012 16838 3014 16890
rect 3194 16838 3196 16890
rect 2950 16836 2956 16838
rect 3012 16836 3036 16838
rect 3092 16836 3116 16838
rect 3172 16836 3196 16838
rect 3252 16836 3258 16838
rect 2950 16827 3258 16836
rect 8864 16574 8892 24919
rect 8956 22681 8984 26862
rect 9036 25832 9088 25838
rect 9036 25774 9088 25780
rect 9048 23186 9076 25774
rect 9036 23180 9088 23186
rect 9036 23122 9088 23128
rect 8942 22672 8998 22681
rect 8942 22607 8998 22616
rect 8956 22137 8984 22607
rect 8942 22128 8998 22137
rect 8942 22063 8998 22072
rect 9140 22030 9168 30126
rect 9588 28008 9640 28014
rect 9588 27950 9640 27956
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9312 24812 9364 24818
rect 9312 24754 9364 24760
rect 9128 22024 9180 22030
rect 9128 21966 9180 21972
rect 8864 16546 8984 16574
rect 5632 16448 5684 16454
rect 5632 16390 5684 16396
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 1308 16040 1360 16046
rect 1308 15982 1360 15988
rect 1320 15745 1348 15982
rect 2950 15804 3258 15813
rect 2950 15802 2956 15804
rect 3012 15802 3036 15804
rect 3092 15802 3116 15804
rect 3172 15802 3196 15804
rect 3252 15802 3258 15804
rect 3012 15750 3014 15802
rect 3194 15750 3196 15802
rect 2950 15748 2956 15750
rect 3012 15748 3036 15750
rect 3092 15748 3116 15750
rect 3172 15748 3196 15750
rect 3252 15748 3258 15750
rect 1306 15736 1362 15745
rect 2950 15739 3258 15748
rect 1306 15671 1362 15680
rect 2950 14716 3258 14725
rect 2950 14714 2956 14716
rect 3012 14714 3036 14716
rect 3092 14714 3116 14716
rect 3172 14714 3196 14716
rect 3252 14714 3258 14716
rect 3012 14662 3014 14714
rect 3194 14662 3196 14714
rect 2950 14660 2956 14662
rect 3012 14660 3036 14662
rect 3092 14660 3116 14662
rect 3172 14660 3196 14662
rect 3252 14660 3258 14662
rect 2950 14651 3258 14660
rect 5644 13938 5672 16390
rect 7950 16348 8258 16357
rect 7950 16346 7956 16348
rect 8012 16346 8036 16348
rect 8092 16346 8116 16348
rect 8172 16346 8196 16348
rect 8252 16346 8258 16348
rect 8012 16294 8014 16346
rect 8194 16294 8196 16346
rect 7950 16292 7956 16294
rect 8012 16292 8036 16294
rect 8092 16292 8116 16294
rect 8172 16292 8196 16294
rect 8252 16292 8258 16294
rect 7950 16283 8258 16292
rect 7950 15260 8258 15269
rect 7950 15258 7956 15260
rect 8012 15258 8036 15260
rect 8092 15258 8116 15260
rect 8172 15258 8196 15260
rect 8252 15258 8258 15260
rect 8012 15206 8014 15258
rect 8194 15206 8196 15258
rect 7950 15204 7956 15206
rect 8012 15204 8036 15206
rect 8092 15204 8116 15206
rect 8172 15204 8196 15206
rect 8252 15204 8258 15206
rect 7950 15195 8258 15204
rect 7950 14172 8258 14181
rect 7950 14170 7956 14172
rect 8012 14170 8036 14172
rect 8092 14170 8116 14172
rect 8172 14170 8196 14172
rect 8252 14170 8258 14172
rect 8012 14118 8014 14170
rect 8194 14118 8196 14170
rect 7950 14116 7956 14118
rect 8012 14116 8036 14118
rect 8092 14116 8116 14118
rect 8172 14116 8196 14118
rect 8252 14116 8258 14118
rect 7950 14107 8258 14116
rect 5632 13932 5684 13938
rect 5632 13874 5684 13880
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13433 2820 13806
rect 2950 13628 3258 13637
rect 2950 13626 2956 13628
rect 3012 13626 3036 13628
rect 3092 13626 3116 13628
rect 3172 13626 3196 13628
rect 3252 13626 3258 13628
rect 3012 13574 3014 13626
rect 3194 13574 3196 13626
rect 2950 13572 2956 13574
rect 3012 13572 3036 13574
rect 3092 13572 3116 13574
rect 3172 13572 3196 13574
rect 3252 13572 3258 13574
rect 2950 13563 3258 13572
rect 2778 13424 2834 13433
rect 2778 13359 2834 13368
rect 7950 13084 8258 13093
rect 7950 13082 7956 13084
rect 8012 13082 8036 13084
rect 8092 13082 8116 13084
rect 8172 13082 8196 13084
rect 8252 13082 8258 13084
rect 8012 13030 8014 13082
rect 8194 13030 8196 13082
rect 7950 13028 7956 13030
rect 8012 13028 8036 13030
rect 8092 13028 8116 13030
rect 8172 13028 8196 13030
rect 8252 13028 8258 13030
rect 7950 13019 8258 13028
rect 2950 12540 3258 12549
rect 2950 12538 2956 12540
rect 3012 12538 3036 12540
rect 3092 12538 3116 12540
rect 3172 12538 3196 12540
rect 3252 12538 3258 12540
rect 3012 12486 3014 12538
rect 3194 12486 3196 12538
rect 2950 12484 2956 12486
rect 3012 12484 3036 12486
rect 3092 12484 3116 12486
rect 3172 12484 3196 12486
rect 3252 12484 3258 12486
rect 2950 12475 3258 12484
rect 3332 12368 3384 12374
rect 3332 12310 3384 12316
rect 2950 11452 3258 11461
rect 2950 11450 2956 11452
rect 3012 11450 3036 11452
rect 3092 11450 3116 11452
rect 3172 11450 3196 11452
rect 3252 11450 3258 11452
rect 3012 11398 3014 11450
rect 3194 11398 3196 11450
rect 2950 11396 2956 11398
rect 3012 11396 3036 11398
rect 3092 11396 3116 11398
rect 3172 11396 3196 11398
rect 3252 11396 3258 11398
rect 2950 11387 3258 11396
rect 3344 11121 3372 12310
rect 7950 11996 8258 12005
rect 7950 11994 7956 11996
rect 8012 11994 8036 11996
rect 8092 11994 8116 11996
rect 8172 11994 8196 11996
rect 8252 11994 8258 11996
rect 8012 11942 8014 11994
rect 8194 11942 8196 11994
rect 7950 11940 7956 11942
rect 8012 11940 8036 11942
rect 8092 11940 8116 11942
rect 8172 11940 8196 11942
rect 8252 11940 8258 11942
rect 7950 11931 8258 11940
rect 3330 11112 3386 11121
rect 3330 11047 3386 11056
rect 7564 11076 7616 11082
rect 7564 11018 7616 11024
rect 2950 10364 3258 10373
rect 2950 10362 2956 10364
rect 3012 10362 3036 10364
rect 3092 10362 3116 10364
rect 3172 10362 3196 10364
rect 3252 10362 3258 10364
rect 3012 10310 3014 10362
rect 3194 10310 3196 10362
rect 2950 10308 2956 10310
rect 3012 10308 3036 10310
rect 3092 10308 3116 10310
rect 3172 10308 3196 10310
rect 3252 10308 3258 10310
rect 2950 10299 3258 10308
rect 2950 9276 3258 9285
rect 2950 9274 2956 9276
rect 3012 9274 3036 9276
rect 3092 9274 3116 9276
rect 3172 9274 3196 9276
rect 3252 9274 3258 9276
rect 3012 9222 3014 9274
rect 3194 9222 3196 9274
rect 2950 9220 2956 9222
rect 3012 9220 3036 9222
rect 3092 9220 3116 9222
rect 3172 9220 3196 9222
rect 3252 9220 3258 9222
rect 2950 9211 3258 9220
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3344 8809 3372 9046
rect 3330 8800 3386 8809
rect 3330 8735 3386 8744
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 2950 8188 3258 8197
rect 2950 8186 2956 8188
rect 3012 8186 3036 8188
rect 3092 8186 3116 8188
rect 3172 8186 3196 8188
rect 3252 8186 3258 8188
rect 3012 8134 3014 8186
rect 3194 8134 3196 8186
rect 2950 8132 2956 8134
rect 3012 8132 3036 8134
rect 3092 8132 3116 8134
rect 3172 8132 3196 8134
rect 3252 8132 3258 8134
rect 2950 8123 3258 8132
rect 2950 7100 3258 7109
rect 2950 7098 2956 7100
rect 3012 7098 3036 7100
rect 3092 7098 3116 7100
rect 3172 7098 3196 7100
rect 3252 7098 3258 7100
rect 3012 7046 3014 7098
rect 3194 7046 3196 7098
rect 2950 7044 2956 7046
rect 3012 7044 3036 7046
rect 3092 7044 3116 7046
rect 3172 7044 3196 7046
rect 3252 7044 3258 7046
rect 2950 7035 3258 7044
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 6497 3464 6598
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2950 6012 3258 6021
rect 2950 6010 2956 6012
rect 3012 6010 3036 6012
rect 3092 6010 3116 6012
rect 3172 6010 3196 6012
rect 3252 6010 3258 6012
rect 3012 5958 3014 6010
rect 3194 5958 3196 6010
rect 2950 5956 2956 5958
rect 3012 5956 3036 5958
rect 3092 5956 3116 5958
rect 3172 5956 3196 5958
rect 3252 5956 3258 5958
rect 2950 5947 3258 5956
rect 3424 5296 3476 5302
rect 3424 5238 3476 5244
rect 2950 4924 3258 4933
rect 2950 4922 2956 4924
rect 3012 4922 3036 4924
rect 3092 4922 3116 4924
rect 3172 4922 3196 4924
rect 3252 4922 3258 4924
rect 3012 4870 3014 4922
rect 3194 4870 3196 4922
rect 2950 4868 2956 4870
rect 3012 4868 3036 4870
rect 3092 4868 3116 4870
rect 3172 4868 3196 4870
rect 3252 4868 3258 4870
rect 2950 4859 3258 4868
rect 3436 4185 3464 5238
rect 3422 4176 3478 4185
rect 3422 4111 3478 4120
rect 2950 3836 3258 3845
rect 2950 3834 2956 3836
rect 3012 3834 3036 3836
rect 3092 3834 3116 3836
rect 3172 3834 3196 3836
rect 3252 3834 3258 3836
rect 3012 3782 3014 3834
rect 3194 3782 3196 3834
rect 2950 3780 2956 3782
rect 3012 3780 3036 3782
rect 3092 3780 3116 3782
rect 3172 3780 3196 3782
rect 3252 3780 3258 3782
rect 2950 3771 3258 3780
rect 5552 3738 5580 8502
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 2780 3528 2832 3534
rect 2780 3470 2832 3476
rect 1492 3052 1544 3058
rect 1492 2994 1544 3000
rect 756 2984 808 2990
rect 756 2926 808 2932
rect 768 800 796 2926
rect 1504 800 1532 2994
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 2240 800 2268 2382
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 1902 2452 2246
rect 2412 1896 2464 1902
rect 2792 1873 2820 3470
rect 7576 3126 7604 11018
rect 7950 10908 8258 10917
rect 7950 10906 7956 10908
rect 8012 10906 8036 10908
rect 8092 10906 8116 10908
rect 8172 10906 8196 10908
rect 8252 10906 8258 10908
rect 8012 10854 8014 10906
rect 8194 10854 8196 10906
rect 7950 10852 7956 10854
rect 8012 10852 8036 10854
rect 8092 10852 8116 10854
rect 8172 10852 8196 10854
rect 8252 10852 8258 10854
rect 7950 10843 8258 10852
rect 7950 9820 8258 9829
rect 7950 9818 7956 9820
rect 8012 9818 8036 9820
rect 8092 9818 8116 9820
rect 8172 9818 8196 9820
rect 8252 9818 8258 9820
rect 8012 9766 8014 9818
rect 8194 9766 8196 9818
rect 7950 9764 7956 9766
rect 8012 9764 8036 9766
rect 8092 9764 8116 9766
rect 8172 9764 8196 9766
rect 8252 9764 8258 9766
rect 7950 9755 8258 9764
rect 7950 8732 8258 8741
rect 7950 8730 7956 8732
rect 8012 8730 8036 8732
rect 8092 8730 8116 8732
rect 8172 8730 8196 8732
rect 8252 8730 8258 8732
rect 8012 8678 8014 8730
rect 8194 8678 8196 8730
rect 7950 8676 7956 8678
rect 8012 8676 8036 8678
rect 8092 8676 8116 8678
rect 8172 8676 8196 8678
rect 8252 8676 8258 8678
rect 7950 8667 8258 8676
rect 7950 7644 8258 7653
rect 7950 7642 7956 7644
rect 8012 7642 8036 7644
rect 8092 7642 8116 7644
rect 8172 7642 8196 7644
rect 8252 7642 8258 7644
rect 8012 7590 8014 7642
rect 8194 7590 8196 7642
rect 7950 7588 7956 7590
rect 8012 7588 8036 7590
rect 8092 7588 8116 7590
rect 8172 7588 8196 7590
rect 8252 7588 8258 7590
rect 7950 7579 8258 7588
rect 8956 6662 8984 16546
rect 9140 6914 9168 21966
rect 9324 21894 9352 24754
rect 9402 22128 9458 22137
rect 9402 22063 9458 22072
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9324 20942 9352 21830
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 9324 18766 9352 20878
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 9416 9110 9444 22063
rect 9508 12374 9536 25774
rect 9600 25265 9628 27950
rect 9680 27940 9732 27946
rect 9680 27882 9732 27888
rect 9692 26586 9720 27882
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 10612 25294 10640 41414
rect 10796 41274 10824 53450
rect 11716 43994 11744 54130
rect 12176 53650 12204 56200
rect 12912 55214 12940 56200
rect 12820 55186 12940 55214
rect 12348 53984 12400 53990
rect 12348 53926 12400 53932
rect 12164 53644 12216 53650
rect 12164 53586 12216 53592
rect 12360 49978 12388 53926
rect 12820 53038 12848 55186
rect 13648 54262 13676 56200
rect 13636 54256 13688 54262
rect 13636 54198 13688 54204
rect 12950 53884 13258 53893
rect 12950 53882 12956 53884
rect 13012 53882 13036 53884
rect 13092 53882 13116 53884
rect 13172 53882 13196 53884
rect 13252 53882 13258 53884
rect 13012 53830 13014 53882
rect 13194 53830 13196 53882
rect 12950 53828 12956 53830
rect 13012 53828 13036 53830
rect 13092 53828 13116 53830
rect 13172 53828 13196 53830
rect 13252 53828 13258 53830
rect 12950 53819 13258 53828
rect 12808 53032 12860 53038
rect 12808 52974 12860 52980
rect 12440 52964 12492 52970
rect 12440 52906 12492 52912
rect 12348 49972 12400 49978
rect 12348 49914 12400 49920
rect 11980 48068 12032 48074
rect 11980 48010 12032 48016
rect 11704 43988 11756 43994
rect 11704 43930 11756 43936
rect 11992 43314 12020 48010
rect 12452 43926 12480 52906
rect 12950 52796 13258 52805
rect 12950 52794 12956 52796
rect 13012 52794 13036 52796
rect 13092 52794 13116 52796
rect 13172 52794 13196 52796
rect 13252 52794 13258 52796
rect 13012 52742 13014 52794
rect 13194 52742 13196 52794
rect 12950 52740 12956 52742
rect 13012 52740 13036 52742
rect 13092 52740 13116 52742
rect 13172 52740 13196 52742
rect 13252 52740 13258 52742
rect 12950 52731 13258 52740
rect 14384 52562 14412 56200
rect 14556 54188 14608 54194
rect 14556 54130 14608 54136
rect 14372 52556 14424 52562
rect 14372 52498 14424 52504
rect 14464 52488 14516 52494
rect 14464 52430 14516 52436
rect 12950 51708 13258 51717
rect 12950 51706 12956 51708
rect 13012 51706 13036 51708
rect 13092 51706 13116 51708
rect 13172 51706 13196 51708
rect 13252 51706 13258 51708
rect 13012 51654 13014 51706
rect 13194 51654 13196 51706
rect 12950 51652 12956 51654
rect 13012 51652 13036 51654
rect 13092 51652 13116 51654
rect 13172 51652 13196 51654
rect 13252 51652 13258 51654
rect 12950 51643 13258 51652
rect 14476 51610 14504 52430
rect 14464 51604 14516 51610
rect 14464 51546 14516 51552
rect 14280 51332 14332 51338
rect 14280 51274 14332 51280
rect 12950 50620 13258 50629
rect 12950 50618 12956 50620
rect 13012 50618 13036 50620
rect 13092 50618 13116 50620
rect 13172 50618 13196 50620
rect 13252 50618 13258 50620
rect 13012 50566 13014 50618
rect 13194 50566 13196 50618
rect 12950 50564 12956 50566
rect 13012 50564 13036 50566
rect 13092 50564 13116 50566
rect 13172 50564 13196 50566
rect 13252 50564 13258 50566
rect 12950 50555 13258 50564
rect 12950 49532 13258 49541
rect 12950 49530 12956 49532
rect 13012 49530 13036 49532
rect 13092 49530 13116 49532
rect 13172 49530 13196 49532
rect 13252 49530 13258 49532
rect 13012 49478 13014 49530
rect 13194 49478 13196 49530
rect 12950 49476 12956 49478
rect 13012 49476 13036 49478
rect 13092 49476 13116 49478
rect 13172 49476 13196 49478
rect 13252 49476 13258 49478
rect 12950 49467 13258 49476
rect 12950 48444 13258 48453
rect 12950 48442 12956 48444
rect 13012 48442 13036 48444
rect 13092 48442 13116 48444
rect 13172 48442 13196 48444
rect 13252 48442 13258 48444
rect 13012 48390 13014 48442
rect 13194 48390 13196 48442
rect 12950 48388 12956 48390
rect 13012 48388 13036 48390
rect 13092 48388 13116 48390
rect 13172 48388 13196 48390
rect 13252 48388 13258 48390
rect 12950 48379 13258 48388
rect 12950 47356 13258 47365
rect 12950 47354 12956 47356
rect 13012 47354 13036 47356
rect 13092 47354 13116 47356
rect 13172 47354 13196 47356
rect 13252 47354 13258 47356
rect 13012 47302 13014 47354
rect 13194 47302 13196 47354
rect 12950 47300 12956 47302
rect 13012 47300 13036 47302
rect 13092 47300 13116 47302
rect 13172 47300 13196 47302
rect 13252 47300 13258 47302
rect 12950 47291 13258 47300
rect 12950 46268 13258 46277
rect 12950 46266 12956 46268
rect 13012 46266 13036 46268
rect 13092 46266 13116 46268
rect 13172 46266 13196 46268
rect 13252 46266 13258 46268
rect 13012 46214 13014 46266
rect 13194 46214 13196 46266
rect 12950 46212 12956 46214
rect 13012 46212 13036 46214
rect 13092 46212 13116 46214
rect 13172 46212 13196 46214
rect 13252 46212 13258 46214
rect 12950 46203 13258 46212
rect 14292 45898 14320 51274
rect 14280 45892 14332 45898
rect 14280 45834 14332 45840
rect 12950 45180 13258 45189
rect 12950 45178 12956 45180
rect 13012 45178 13036 45180
rect 13092 45178 13116 45180
rect 13172 45178 13196 45180
rect 13252 45178 13258 45180
rect 13012 45126 13014 45178
rect 13194 45126 13196 45178
rect 12950 45124 12956 45126
rect 13012 45124 13036 45126
rect 13092 45124 13116 45126
rect 13172 45124 13196 45126
rect 13252 45124 13258 45126
rect 12950 45115 13258 45124
rect 14464 44396 14516 44402
rect 14464 44338 14516 44344
rect 12950 44092 13258 44101
rect 12950 44090 12956 44092
rect 13012 44090 13036 44092
rect 13092 44090 13116 44092
rect 13172 44090 13196 44092
rect 13252 44090 13258 44092
rect 13012 44038 13014 44090
rect 13194 44038 13196 44090
rect 12950 44036 12956 44038
rect 13012 44036 13036 44038
rect 13092 44036 13116 44038
rect 13172 44036 13196 44038
rect 13252 44036 13258 44038
rect 12950 44027 13258 44036
rect 12440 43920 12492 43926
rect 12440 43862 12492 43868
rect 13452 43716 13504 43722
rect 13452 43658 13504 43664
rect 11980 43308 12032 43314
rect 11980 43250 12032 43256
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 11992 41546 12020 43250
rect 12084 42906 12112 43250
rect 13464 43178 13492 43658
rect 13452 43172 13504 43178
rect 13452 43114 13504 43120
rect 12950 43004 13258 43013
rect 12950 43002 12956 43004
rect 13012 43002 13036 43004
rect 13092 43002 13116 43004
rect 13172 43002 13196 43004
rect 13252 43002 13258 43004
rect 13012 42950 13014 43002
rect 13194 42950 13196 43002
rect 12950 42948 12956 42950
rect 13012 42948 13036 42950
rect 13092 42948 13116 42950
rect 13172 42948 13196 42950
rect 13252 42948 13258 42950
rect 12950 42939 13258 42948
rect 12072 42900 12124 42906
rect 12072 42842 12124 42848
rect 12950 41916 13258 41925
rect 12950 41914 12956 41916
rect 13012 41914 13036 41916
rect 13092 41914 13116 41916
rect 13172 41914 13196 41916
rect 13252 41914 13258 41916
rect 13012 41862 13014 41914
rect 13194 41862 13196 41914
rect 12950 41860 12956 41862
rect 13012 41860 13036 41862
rect 13092 41860 13116 41862
rect 13172 41860 13196 41862
rect 13252 41860 13258 41862
rect 12950 41851 13258 41860
rect 11980 41540 12032 41546
rect 11980 41482 12032 41488
rect 10784 41268 10836 41274
rect 10784 41210 10836 41216
rect 10692 41132 10744 41138
rect 10692 41074 10744 41080
rect 10704 30326 10732 41074
rect 12950 40828 13258 40837
rect 12950 40826 12956 40828
rect 13012 40826 13036 40828
rect 13092 40826 13116 40828
rect 13172 40826 13196 40828
rect 13252 40826 13258 40828
rect 13012 40774 13014 40826
rect 13194 40774 13196 40826
rect 12950 40772 12956 40774
rect 13012 40772 13036 40774
rect 13092 40772 13116 40774
rect 13172 40772 13196 40774
rect 13252 40772 13258 40774
rect 12950 40763 13258 40772
rect 12950 39740 13258 39749
rect 12950 39738 12956 39740
rect 13012 39738 13036 39740
rect 13092 39738 13116 39740
rect 13172 39738 13196 39740
rect 13252 39738 13258 39740
rect 13012 39686 13014 39738
rect 13194 39686 13196 39738
rect 12950 39684 12956 39686
rect 13012 39684 13036 39686
rect 13092 39684 13116 39686
rect 13172 39684 13196 39686
rect 13252 39684 13258 39686
rect 12950 39675 13258 39684
rect 12950 38652 13258 38661
rect 12950 38650 12956 38652
rect 13012 38650 13036 38652
rect 13092 38650 13116 38652
rect 13172 38650 13196 38652
rect 13252 38650 13258 38652
rect 13012 38598 13014 38650
rect 13194 38598 13196 38650
rect 12950 38596 12956 38598
rect 13012 38596 13036 38598
rect 13092 38596 13116 38598
rect 13172 38596 13196 38598
rect 13252 38596 13258 38598
rect 12950 38587 13258 38596
rect 12950 37564 13258 37573
rect 12950 37562 12956 37564
rect 13012 37562 13036 37564
rect 13092 37562 13116 37564
rect 13172 37562 13196 37564
rect 13252 37562 13258 37564
rect 13012 37510 13014 37562
rect 13194 37510 13196 37562
rect 12950 37508 12956 37510
rect 13012 37508 13036 37510
rect 13092 37508 13116 37510
rect 13172 37508 13196 37510
rect 13252 37508 13258 37510
rect 12950 37499 13258 37508
rect 14476 37194 14504 44338
rect 14568 42362 14596 54130
rect 14648 54052 14700 54058
rect 14648 53994 14700 54000
rect 14660 43994 14688 53994
rect 14740 53576 14792 53582
rect 14740 53518 14792 53524
rect 14752 49978 14780 53518
rect 15120 53038 15148 56200
rect 15856 53718 15884 56200
rect 16592 54262 16620 56200
rect 16580 54256 16632 54262
rect 16580 54198 16632 54204
rect 15844 53712 15896 53718
rect 15844 53654 15896 53660
rect 16948 53168 17000 53174
rect 16948 53110 17000 53116
rect 15200 53100 15252 53106
rect 15200 53042 15252 53048
rect 15108 53032 15160 53038
rect 15108 52974 15160 52980
rect 14740 49972 14792 49978
rect 14740 49914 14792 49920
rect 15212 49434 15240 53042
rect 15936 51332 15988 51338
rect 15936 51274 15988 51280
rect 15200 49428 15252 49434
rect 15200 49370 15252 49376
rect 15948 46170 15976 51274
rect 16856 49836 16908 49842
rect 16856 49778 16908 49784
rect 15936 46164 15988 46170
rect 15936 46106 15988 46112
rect 14924 45484 14976 45490
rect 14924 45426 14976 45432
rect 14648 43988 14700 43994
rect 14648 43930 14700 43936
rect 14556 42356 14608 42362
rect 14556 42298 14608 42304
rect 14464 37188 14516 37194
rect 14464 37130 14516 37136
rect 12950 36476 13258 36485
rect 12950 36474 12956 36476
rect 13012 36474 13036 36476
rect 13092 36474 13116 36476
rect 13172 36474 13196 36476
rect 13252 36474 13258 36476
rect 13012 36422 13014 36474
rect 13194 36422 13196 36474
rect 12950 36420 12956 36422
rect 13012 36420 13036 36422
rect 13092 36420 13116 36422
rect 13172 36420 13196 36422
rect 13252 36420 13258 36422
rect 12950 36411 13258 36420
rect 12950 35388 13258 35397
rect 12950 35386 12956 35388
rect 13012 35386 13036 35388
rect 13092 35386 13116 35388
rect 13172 35386 13196 35388
rect 13252 35386 13258 35388
rect 13012 35334 13014 35386
rect 13194 35334 13196 35386
rect 12950 35332 12956 35334
rect 13012 35332 13036 35334
rect 13092 35332 13116 35334
rect 13172 35332 13196 35334
rect 13252 35332 13258 35334
rect 12950 35323 13258 35332
rect 12950 34300 13258 34309
rect 12950 34298 12956 34300
rect 13012 34298 13036 34300
rect 13092 34298 13116 34300
rect 13172 34298 13196 34300
rect 13252 34298 13258 34300
rect 13012 34246 13014 34298
rect 13194 34246 13196 34298
rect 12950 34244 12956 34246
rect 13012 34244 13036 34246
rect 13092 34244 13116 34246
rect 13172 34244 13196 34246
rect 13252 34244 13258 34246
rect 12950 34235 13258 34244
rect 12950 33212 13258 33221
rect 12950 33210 12956 33212
rect 13012 33210 13036 33212
rect 13092 33210 13116 33212
rect 13172 33210 13196 33212
rect 13252 33210 13258 33212
rect 13012 33158 13014 33210
rect 13194 33158 13196 33210
rect 12950 33156 12956 33158
rect 13012 33156 13036 33158
rect 13092 33156 13116 33158
rect 13172 33156 13196 33158
rect 13252 33156 13258 33158
rect 12950 33147 13258 33156
rect 12950 32124 13258 32133
rect 12950 32122 12956 32124
rect 13012 32122 13036 32124
rect 13092 32122 13116 32124
rect 13172 32122 13196 32124
rect 13252 32122 13258 32124
rect 13012 32070 13014 32122
rect 13194 32070 13196 32122
rect 12950 32068 12956 32070
rect 13012 32068 13036 32070
rect 13092 32068 13116 32070
rect 13172 32068 13196 32070
rect 13252 32068 13258 32070
rect 12950 32059 13258 32068
rect 12950 31036 13258 31045
rect 12950 31034 12956 31036
rect 13012 31034 13036 31036
rect 13092 31034 13116 31036
rect 13172 31034 13196 31036
rect 13252 31034 13258 31036
rect 13012 30982 13014 31034
rect 13194 30982 13196 31034
rect 12950 30980 12956 30982
rect 13012 30980 13036 30982
rect 13092 30980 13116 30982
rect 13172 30980 13196 30982
rect 13252 30980 13258 30982
rect 12950 30971 13258 30980
rect 10692 30320 10744 30326
rect 10692 30262 10744 30268
rect 12950 29948 13258 29957
rect 12950 29946 12956 29948
rect 13012 29946 13036 29948
rect 13092 29946 13116 29948
rect 13172 29946 13196 29948
rect 13252 29946 13258 29948
rect 13012 29894 13014 29946
rect 13194 29894 13196 29946
rect 12950 29892 12956 29894
rect 13012 29892 13036 29894
rect 13092 29892 13116 29894
rect 13172 29892 13196 29894
rect 13252 29892 13258 29894
rect 12950 29883 13258 29892
rect 12950 28860 13258 28869
rect 12950 28858 12956 28860
rect 13012 28858 13036 28860
rect 13092 28858 13116 28860
rect 13172 28858 13196 28860
rect 13252 28858 13258 28860
rect 13012 28806 13014 28858
rect 13194 28806 13196 28858
rect 12950 28804 12956 28806
rect 13012 28804 13036 28806
rect 13092 28804 13116 28806
rect 13172 28804 13196 28806
rect 13252 28804 13258 28806
rect 12950 28795 13258 28804
rect 12950 27772 13258 27781
rect 12950 27770 12956 27772
rect 13012 27770 13036 27772
rect 13092 27770 13116 27772
rect 13172 27770 13196 27772
rect 13252 27770 13258 27772
rect 13012 27718 13014 27770
rect 13194 27718 13196 27770
rect 12950 27716 12956 27718
rect 13012 27716 13036 27718
rect 13092 27716 13116 27718
rect 13172 27716 13196 27718
rect 13252 27716 13258 27718
rect 12950 27707 13258 27716
rect 12950 26684 13258 26693
rect 12950 26682 12956 26684
rect 13012 26682 13036 26684
rect 13092 26682 13116 26684
rect 13172 26682 13196 26684
rect 13252 26682 13258 26684
rect 13012 26630 13014 26682
rect 13194 26630 13196 26682
rect 12950 26628 12956 26630
rect 13012 26628 13036 26630
rect 13092 26628 13116 26630
rect 13172 26628 13196 26630
rect 13252 26628 13258 26630
rect 12950 26619 13258 26628
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 10888 25430 10916 26386
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10980 25498 11008 26318
rect 12950 25596 13258 25605
rect 12950 25594 12956 25596
rect 13012 25594 13036 25596
rect 13092 25594 13116 25596
rect 13172 25594 13196 25596
rect 13252 25594 13258 25596
rect 13012 25542 13014 25594
rect 13194 25542 13196 25594
rect 12950 25540 12956 25542
rect 13012 25540 13036 25542
rect 13092 25540 13116 25542
rect 13172 25540 13196 25542
rect 13252 25540 13258 25542
rect 12950 25531 13258 25540
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10876 25424 10928 25430
rect 10876 25366 10928 25372
rect 12348 25356 12400 25362
rect 12348 25298 12400 25304
rect 10600 25288 10652 25294
rect 9586 25256 9642 25265
rect 10600 25230 10652 25236
rect 9586 25191 9642 25200
rect 9600 24993 9628 25191
rect 9586 24984 9642 24993
rect 9586 24919 9642 24928
rect 10612 24206 10640 25230
rect 12360 24410 12388 25298
rect 12950 24508 13258 24517
rect 12950 24506 12956 24508
rect 13012 24506 13036 24508
rect 13092 24506 13116 24508
rect 13172 24506 13196 24508
rect 13252 24506 13258 24508
rect 13012 24454 13014 24506
rect 13194 24454 13196 24506
rect 12950 24452 12956 24454
rect 13012 24452 13036 24454
rect 13092 24452 13116 24454
rect 13172 24452 13196 24454
rect 13252 24452 13258 24454
rect 12950 24443 13258 24452
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 10600 24200 10652 24206
rect 10600 24142 10652 24148
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 9772 23112 9824 23118
rect 9772 23054 9824 23060
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9692 21146 9720 22986
rect 9784 21486 9812 23054
rect 10232 21956 10284 21962
rect 10232 21898 10284 21904
rect 10244 21690 10272 21898
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9680 21140 9732 21146
rect 9680 21082 9732 21088
rect 9784 18902 9812 21422
rect 10968 21004 11020 21010
rect 10968 20946 11020 20952
rect 10980 20058 11008 20946
rect 10968 20052 11020 20058
rect 10968 19994 11020 20000
rect 9772 18896 9824 18902
rect 9772 18838 9824 18844
rect 9784 16522 9812 18838
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9496 12368 9548 12374
rect 9496 12310 9548 12316
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9048 6886 9168 6914
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 7950 6556 8258 6565
rect 7950 6554 7956 6556
rect 8012 6554 8036 6556
rect 8092 6554 8116 6556
rect 8172 6554 8196 6556
rect 8252 6554 8258 6556
rect 8012 6502 8014 6554
rect 8194 6502 8196 6554
rect 7950 6500 7956 6502
rect 8012 6500 8036 6502
rect 8092 6500 8116 6502
rect 8172 6500 8196 6502
rect 8252 6500 8258 6502
rect 7950 6491 8258 6500
rect 7950 5468 8258 5477
rect 7950 5466 7956 5468
rect 8012 5466 8036 5468
rect 8092 5466 8116 5468
rect 8172 5466 8196 5468
rect 8252 5466 8258 5468
rect 8012 5414 8014 5466
rect 8194 5414 8196 5466
rect 7950 5412 7956 5414
rect 8012 5412 8036 5414
rect 8092 5412 8116 5414
rect 8172 5412 8196 5414
rect 8252 5412 8258 5414
rect 7950 5403 8258 5412
rect 9048 5302 9076 6886
rect 9036 5296 9088 5302
rect 9036 5238 9088 5244
rect 10048 4820 10100 4826
rect 10048 4762 10100 4768
rect 7950 4380 8258 4389
rect 7950 4378 7956 4380
rect 8012 4378 8036 4380
rect 8092 4378 8116 4380
rect 8172 4378 8196 4380
rect 8252 4378 8258 4380
rect 8012 4326 8014 4378
rect 8194 4326 8196 4378
rect 7950 4324 7956 4326
rect 8012 4324 8036 4326
rect 8092 4324 8116 4326
rect 8172 4324 8196 4326
rect 8252 4324 8258 4326
rect 7950 4315 8258 4324
rect 7950 3292 8258 3301
rect 7950 3290 7956 3292
rect 8012 3290 8036 3292
rect 8092 3290 8116 3292
rect 8172 3290 8196 3292
rect 8252 3290 8258 3292
rect 8012 3238 8014 3290
rect 8194 3238 8196 3290
rect 7950 3236 7956 3238
rect 8012 3236 8036 3238
rect 8092 3236 8116 3238
rect 8172 3236 8196 3238
rect 8252 3236 8258 3238
rect 7950 3227 8258 3236
rect 7564 3120 7616 3126
rect 7564 3062 7616 3068
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 2950 2748 3258 2757
rect 2950 2746 2956 2748
rect 3012 2746 3036 2748
rect 3092 2746 3116 2748
rect 3172 2746 3196 2748
rect 3252 2746 3258 2748
rect 3012 2694 3014 2746
rect 3194 2694 3196 2746
rect 2950 2692 2956 2694
rect 3012 2692 3036 2694
rect 3092 2692 3116 2694
rect 3172 2692 3196 2694
rect 3252 2692 3258 2694
rect 2950 2683 3258 2692
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2412 1838 2464 1844
rect 2778 1864 2834 1873
rect 2778 1799 2834 1808
rect 2976 800 3004 2314
rect 3332 2304 3384 2310
rect 3332 2246 3384 2252
rect 3344 1698 3372 2246
rect 3332 1692 3384 1698
rect 3332 1634 3384 1640
rect 3712 800 3740 2994
rect 4986 2408 5042 2417
rect 4436 2372 4488 2378
rect 4986 2343 4988 2352
rect 4436 2314 4488 2320
rect 5040 2343 5042 2352
rect 4988 2314 5040 2320
rect 4448 800 4476 2314
rect 5184 800 5212 2994
rect 5736 2961 5764 2994
rect 5722 2952 5778 2961
rect 5722 2887 5778 2896
rect 5908 2372 5960 2378
rect 5908 2314 5960 2320
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5920 800 5948 2314
rect 6012 2038 6040 2314
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6656 800 6684 2994
rect 10060 2650 10088 4762
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9494 2544 9550 2553
rect 9494 2479 9496 2488
rect 9548 2479 9550 2488
rect 9496 2450 9548 2456
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 7392 800 7420 2382
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 8852 2372 8904 2378
rect 8852 2314 8904 2320
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 1970 7604 2246
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 754 0 810 800
rect 1490 0 1546 800
rect 2226 0 2282 800
rect 2962 0 3018 800
rect 3698 0 3754 800
rect 4434 0 4490 800
rect 5170 0 5226 800
rect 5906 0 5962 800
rect 6642 0 6698 800
rect 7378 0 7434 800
rect 7852 762 7880 2314
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 7950 2204 8258 2213
rect 7950 2202 7956 2204
rect 8012 2202 8036 2204
rect 8092 2202 8116 2204
rect 8172 2202 8196 2204
rect 8252 2202 8258 2204
rect 8012 2150 8014 2202
rect 8194 2150 8196 2202
rect 7950 2148 7956 2150
rect 8012 2148 8036 2150
rect 8092 2148 8116 2150
rect 8172 2148 8196 2150
rect 8252 2148 8258 2150
rect 7950 2139 8258 2148
rect 8496 1766 8524 2246
rect 8484 1760 8536 1766
rect 8484 1702 8536 1708
rect 8036 870 8156 898
rect 8036 762 8064 870
rect 8128 800 8156 870
rect 8864 800 8892 2314
rect 9600 800 9628 2382
rect 10336 800 10364 2994
rect 11164 2650 11192 24006
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12268 21418 12296 23666
rect 12360 23662 12388 24346
rect 12532 24200 12584 24206
rect 12532 24142 12584 24148
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12544 22030 12572 24142
rect 12950 23420 13258 23429
rect 12950 23418 12956 23420
rect 13012 23418 13036 23420
rect 13092 23418 13116 23420
rect 13172 23418 13196 23420
rect 13252 23418 13258 23420
rect 13012 23366 13014 23418
rect 13194 23366 13196 23418
rect 12950 23364 12956 23366
rect 13012 23364 13036 23366
rect 13092 23364 13116 23366
rect 13172 23364 13196 23366
rect 13252 23364 13258 23366
rect 12950 23355 13258 23364
rect 12950 22332 13258 22341
rect 12950 22330 12956 22332
rect 13012 22330 13036 22332
rect 13092 22330 13116 22332
rect 13172 22330 13196 22332
rect 13252 22330 13258 22332
rect 13012 22278 13014 22330
rect 13194 22278 13196 22330
rect 12950 22276 12956 22278
rect 13012 22276 13036 22278
rect 13092 22276 13116 22278
rect 13172 22276 13196 22278
rect 13252 22276 13258 22278
rect 12950 22267 13258 22276
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 13636 22024 13688 22030
rect 13636 21966 13688 21972
rect 12256 21412 12308 21418
rect 12256 21354 12308 21360
rect 12544 18766 12572 21966
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21554 13492 21830
rect 13648 21690 13676 21966
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 12950 21244 13258 21253
rect 12950 21242 12956 21244
rect 13012 21242 13036 21244
rect 13092 21242 13116 21244
rect 13172 21242 13196 21244
rect 13252 21242 13258 21244
rect 13012 21190 13014 21242
rect 13194 21190 13196 21242
rect 12950 21188 12956 21190
rect 13012 21188 13036 21190
rect 13092 21188 13116 21190
rect 13172 21188 13196 21190
rect 13252 21188 13258 21190
rect 12950 21179 13258 21188
rect 12950 20156 13258 20165
rect 12950 20154 12956 20156
rect 13012 20154 13036 20156
rect 13092 20154 13116 20156
rect 13172 20154 13196 20156
rect 13252 20154 13258 20156
rect 13012 20102 13014 20154
rect 13194 20102 13196 20154
rect 12950 20100 12956 20102
rect 13012 20100 13036 20102
rect 13092 20100 13116 20102
rect 13172 20100 13196 20102
rect 13252 20100 13258 20102
rect 12950 20091 13258 20100
rect 12950 19068 13258 19077
rect 12950 19066 12956 19068
rect 13012 19066 13036 19068
rect 13092 19066 13116 19068
rect 13172 19066 13196 19068
rect 13252 19066 13258 19068
rect 13012 19014 13014 19066
rect 13194 19014 13196 19066
rect 12950 19012 12956 19014
rect 13012 19012 13036 19014
rect 13092 19012 13116 19014
rect 13172 19012 13196 19014
rect 13252 19012 13258 19014
rect 12950 19003 13258 19012
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12950 17980 13258 17989
rect 12950 17978 12956 17980
rect 13012 17978 13036 17980
rect 13092 17978 13116 17980
rect 13172 17978 13196 17980
rect 13252 17978 13258 17980
rect 13012 17926 13014 17978
rect 13194 17926 13196 17978
rect 12950 17924 12956 17926
rect 13012 17924 13036 17926
rect 13092 17924 13116 17926
rect 13172 17924 13196 17926
rect 13252 17924 13258 17926
rect 12950 17915 13258 17924
rect 12950 16892 13258 16901
rect 12950 16890 12956 16892
rect 13012 16890 13036 16892
rect 13092 16890 13116 16892
rect 13172 16890 13196 16892
rect 13252 16890 13258 16892
rect 13012 16838 13014 16890
rect 13194 16838 13196 16890
rect 12950 16836 12956 16838
rect 13012 16836 13036 16838
rect 13092 16836 13116 16838
rect 13172 16836 13196 16838
rect 13252 16836 13258 16838
rect 12950 16827 13258 16836
rect 12950 15804 13258 15813
rect 12950 15802 12956 15804
rect 13012 15802 13036 15804
rect 13092 15802 13116 15804
rect 13172 15802 13196 15804
rect 13252 15802 13258 15804
rect 13012 15750 13014 15802
rect 13194 15750 13196 15802
rect 12950 15748 12956 15750
rect 13012 15748 13036 15750
rect 13092 15748 13116 15750
rect 13172 15748 13196 15750
rect 13252 15748 13258 15750
rect 12950 15739 13258 15748
rect 12950 14716 13258 14725
rect 12950 14714 12956 14716
rect 13012 14714 13036 14716
rect 13092 14714 13116 14716
rect 13172 14714 13196 14716
rect 13252 14714 13258 14716
rect 13012 14662 13014 14714
rect 13194 14662 13196 14714
rect 12950 14660 12956 14662
rect 13012 14660 13036 14662
rect 13092 14660 13116 14662
rect 13172 14660 13196 14662
rect 13252 14660 13258 14662
rect 12950 14651 13258 14660
rect 12950 13628 13258 13637
rect 12950 13626 12956 13628
rect 13012 13626 13036 13628
rect 13092 13626 13116 13628
rect 13172 13626 13196 13628
rect 13252 13626 13258 13628
rect 13012 13574 13014 13626
rect 13194 13574 13196 13626
rect 12950 13572 12956 13574
rect 13012 13572 13036 13574
rect 13092 13572 13116 13574
rect 13172 13572 13196 13574
rect 13252 13572 13258 13574
rect 12950 13563 13258 13572
rect 12950 12540 13258 12549
rect 12950 12538 12956 12540
rect 13012 12538 13036 12540
rect 13092 12538 13116 12540
rect 13172 12538 13196 12540
rect 13252 12538 13258 12540
rect 13012 12486 13014 12538
rect 13194 12486 13196 12538
rect 12950 12484 12956 12486
rect 13012 12484 13036 12486
rect 13092 12484 13116 12486
rect 13172 12484 13196 12486
rect 13252 12484 13258 12486
rect 12950 12475 13258 12484
rect 12950 11452 13258 11461
rect 12950 11450 12956 11452
rect 13012 11450 13036 11452
rect 13092 11450 13116 11452
rect 13172 11450 13196 11452
rect 13252 11450 13258 11452
rect 13012 11398 13014 11450
rect 13194 11398 13196 11450
rect 12950 11396 12956 11398
rect 13012 11396 13036 11398
rect 13092 11396 13116 11398
rect 13172 11396 13196 11398
rect 13252 11396 13258 11398
rect 12950 11387 13258 11396
rect 12950 10364 13258 10373
rect 12950 10362 12956 10364
rect 13012 10362 13036 10364
rect 13092 10362 13116 10364
rect 13172 10362 13196 10364
rect 13252 10362 13258 10364
rect 13012 10310 13014 10362
rect 13194 10310 13196 10362
rect 12950 10308 12956 10310
rect 13012 10308 13036 10310
rect 13092 10308 13116 10310
rect 13172 10308 13196 10310
rect 13252 10308 13258 10310
rect 12950 10299 13258 10308
rect 12950 9276 13258 9285
rect 12950 9274 12956 9276
rect 13012 9274 13036 9276
rect 13092 9274 13116 9276
rect 13172 9274 13196 9276
rect 13252 9274 13258 9276
rect 13012 9222 13014 9274
rect 13194 9222 13196 9274
rect 12950 9220 12956 9222
rect 13012 9220 13036 9222
rect 13092 9220 13116 9222
rect 13172 9220 13196 9222
rect 13252 9220 13258 9222
rect 12950 9211 13258 9220
rect 12950 8188 13258 8197
rect 12950 8186 12956 8188
rect 13012 8186 13036 8188
rect 13092 8186 13116 8188
rect 13172 8186 13196 8188
rect 13252 8186 13258 8188
rect 13012 8134 13014 8186
rect 13194 8134 13196 8186
rect 12950 8132 12956 8134
rect 13012 8132 13036 8134
rect 13092 8132 13116 8134
rect 13172 8132 13196 8134
rect 13252 8132 13258 8134
rect 12950 8123 13258 8132
rect 12950 7100 13258 7109
rect 12950 7098 12956 7100
rect 13012 7098 13036 7100
rect 13092 7098 13116 7100
rect 13172 7098 13196 7100
rect 13252 7098 13258 7100
rect 13012 7046 13014 7098
rect 13194 7046 13196 7098
rect 12950 7044 12956 7046
rect 13012 7044 13036 7046
rect 13092 7044 13116 7046
rect 13172 7044 13196 7046
rect 13252 7044 13258 7046
rect 12950 7035 13258 7044
rect 12950 6012 13258 6021
rect 12950 6010 12956 6012
rect 13012 6010 13036 6012
rect 13092 6010 13116 6012
rect 13172 6010 13196 6012
rect 13252 6010 13258 6012
rect 13012 5958 13014 6010
rect 13194 5958 13196 6010
rect 12950 5956 12956 5958
rect 13012 5956 13036 5958
rect 13092 5956 13116 5958
rect 13172 5956 13196 5958
rect 13252 5956 13258 5958
rect 12950 5947 13258 5956
rect 12950 4924 13258 4933
rect 12950 4922 12956 4924
rect 13012 4922 13036 4924
rect 13092 4922 13116 4924
rect 13172 4922 13196 4924
rect 13252 4922 13258 4924
rect 13012 4870 13014 4922
rect 13194 4870 13196 4922
rect 12950 4868 12956 4870
rect 13012 4868 13036 4870
rect 13092 4868 13116 4870
rect 13172 4868 13196 4870
rect 13252 4868 13258 4870
rect 12950 4859 13258 4868
rect 12950 3836 13258 3845
rect 12950 3834 12956 3836
rect 13012 3834 13036 3836
rect 13092 3834 13116 3836
rect 13172 3834 13196 3836
rect 13252 3834 13258 3836
rect 13012 3782 13014 3834
rect 13194 3782 13196 3834
rect 12950 3780 12956 3782
rect 13012 3780 13036 3782
rect 13092 3780 13116 3782
rect 13172 3780 13196 3782
rect 13252 3780 13258 3782
rect 12950 3771 13258 3780
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3126 12940 3334
rect 14476 3194 14504 37130
rect 14936 37126 14964 45426
rect 16868 43450 16896 49778
rect 16960 43994 16988 53110
rect 17328 53038 17356 56200
rect 18064 56114 18092 56200
rect 18156 56114 18184 56222
rect 18064 56086 18184 56114
rect 17950 54428 18258 54437
rect 17950 54426 17956 54428
rect 18012 54426 18036 54428
rect 18092 54426 18116 54428
rect 18172 54426 18196 54428
rect 18252 54426 18258 54428
rect 18012 54374 18014 54426
rect 18194 54374 18196 54426
rect 17950 54372 17956 54374
rect 18012 54372 18036 54374
rect 18092 54372 18116 54374
rect 18172 54372 18196 54374
rect 18252 54372 18258 54374
rect 17950 54363 18258 54372
rect 17684 54188 17736 54194
rect 17684 54130 17736 54136
rect 17316 53032 17368 53038
rect 17316 52974 17368 52980
rect 17696 50522 17724 54130
rect 18340 53650 18368 56222
rect 18786 56200 18842 57000
rect 19522 56200 19578 57000
rect 20258 56200 20314 57000
rect 20994 56200 21050 57000
rect 21730 56200 21786 57000
rect 22466 56200 22522 57000
rect 23202 56200 23258 57000
rect 23938 56200 23994 57000
rect 24674 56200 24730 57000
rect 25410 56200 25466 57000
rect 26146 56200 26202 57000
rect 26882 56200 26938 57000
rect 27618 56200 27674 57000
rect 28354 56200 28410 57000
rect 29090 56200 29146 57000
rect 29826 56200 29882 57000
rect 30562 56200 30618 57000
rect 31298 56200 31354 57000
rect 32034 56200 32090 57000
rect 32770 56200 32826 57000
rect 33506 56200 33562 57000
rect 34242 56200 34298 57000
rect 34978 56200 35034 57000
rect 35714 56200 35770 57000
rect 36450 56200 36506 57000
rect 37186 56200 37242 57000
rect 37922 56200 37978 57000
rect 38658 56200 38714 57000
rect 39394 56200 39450 57000
rect 40130 56200 40186 57000
rect 40866 56200 40922 57000
rect 41602 56200 41658 57000
rect 42338 56200 42394 57000
rect 43074 56200 43130 57000
rect 43810 56200 43866 57000
rect 43916 56222 44128 56250
rect 18800 54262 18828 56200
rect 18788 54256 18840 54262
rect 18788 54198 18840 54204
rect 18328 53644 18380 53650
rect 18328 53586 18380 53592
rect 18420 53576 18472 53582
rect 18420 53518 18472 53524
rect 17950 53340 18258 53349
rect 17950 53338 17956 53340
rect 18012 53338 18036 53340
rect 18092 53338 18116 53340
rect 18172 53338 18196 53340
rect 18252 53338 18258 53340
rect 18012 53286 18014 53338
rect 18194 53286 18196 53338
rect 17950 53284 17956 53286
rect 18012 53284 18036 53286
rect 18092 53284 18116 53286
rect 18172 53284 18196 53286
rect 18252 53284 18258 53286
rect 17950 53275 18258 53284
rect 17950 52252 18258 52261
rect 17950 52250 17956 52252
rect 18012 52250 18036 52252
rect 18092 52250 18116 52252
rect 18172 52250 18196 52252
rect 18252 52250 18258 52252
rect 18012 52198 18014 52250
rect 18194 52198 18196 52250
rect 17950 52196 17956 52198
rect 18012 52196 18036 52198
rect 18092 52196 18116 52198
rect 18172 52196 18196 52198
rect 18252 52196 18258 52198
rect 17950 52187 18258 52196
rect 17950 51164 18258 51173
rect 17950 51162 17956 51164
rect 18012 51162 18036 51164
rect 18092 51162 18116 51164
rect 18172 51162 18196 51164
rect 18252 51162 18258 51164
rect 18012 51110 18014 51162
rect 18194 51110 18196 51162
rect 17950 51108 17956 51110
rect 18012 51108 18036 51110
rect 18092 51108 18116 51110
rect 18172 51108 18196 51110
rect 18252 51108 18258 51110
rect 17950 51099 18258 51108
rect 17684 50516 17736 50522
rect 17684 50458 17736 50464
rect 17950 50076 18258 50085
rect 17950 50074 17956 50076
rect 18012 50074 18036 50076
rect 18092 50074 18116 50076
rect 18172 50074 18196 50076
rect 18252 50074 18258 50076
rect 18012 50022 18014 50074
rect 18194 50022 18196 50074
rect 17950 50020 17956 50022
rect 18012 50020 18036 50022
rect 18092 50020 18116 50022
rect 18172 50020 18196 50022
rect 18252 50020 18258 50022
rect 17950 50011 18258 50020
rect 18432 49434 18460 53518
rect 19536 53038 19564 56200
rect 20168 54120 20220 54126
rect 20168 54062 20220 54068
rect 19616 53100 19668 53106
rect 19616 53042 19668 53048
rect 19524 53032 19576 53038
rect 19524 52974 19576 52980
rect 19156 52488 19208 52494
rect 19156 52430 19208 52436
rect 18420 49428 18472 49434
rect 18420 49370 18472 49376
rect 17950 48988 18258 48997
rect 17950 48986 17956 48988
rect 18012 48986 18036 48988
rect 18092 48986 18116 48988
rect 18172 48986 18196 48988
rect 18252 48986 18258 48988
rect 18012 48934 18014 48986
rect 18194 48934 18196 48986
rect 17950 48932 17956 48934
rect 18012 48932 18036 48934
rect 18092 48932 18116 48934
rect 18172 48932 18196 48934
rect 18252 48932 18258 48934
rect 17950 48923 18258 48932
rect 17950 47900 18258 47909
rect 17950 47898 17956 47900
rect 18012 47898 18036 47900
rect 18092 47898 18116 47900
rect 18172 47898 18196 47900
rect 18252 47898 18258 47900
rect 18012 47846 18014 47898
rect 18194 47846 18196 47898
rect 17950 47844 17956 47846
rect 18012 47844 18036 47846
rect 18092 47844 18116 47846
rect 18172 47844 18196 47846
rect 18252 47844 18258 47846
rect 17950 47835 18258 47844
rect 17950 46812 18258 46821
rect 17950 46810 17956 46812
rect 18012 46810 18036 46812
rect 18092 46810 18116 46812
rect 18172 46810 18196 46812
rect 18252 46810 18258 46812
rect 18012 46758 18014 46810
rect 18194 46758 18196 46810
rect 17950 46756 17956 46758
rect 18012 46756 18036 46758
rect 18092 46756 18116 46758
rect 18172 46756 18196 46758
rect 18252 46756 18258 46758
rect 17950 46747 18258 46756
rect 17950 45724 18258 45733
rect 17950 45722 17956 45724
rect 18012 45722 18036 45724
rect 18092 45722 18116 45724
rect 18172 45722 18196 45724
rect 18252 45722 18258 45724
rect 18012 45670 18014 45722
rect 18194 45670 18196 45722
rect 17950 45668 17956 45670
rect 18012 45668 18036 45670
rect 18092 45668 18116 45670
rect 18172 45668 18196 45670
rect 18252 45668 18258 45670
rect 17950 45659 18258 45668
rect 17950 44636 18258 44645
rect 17950 44634 17956 44636
rect 18012 44634 18036 44636
rect 18092 44634 18116 44636
rect 18172 44634 18196 44636
rect 18252 44634 18258 44636
rect 18012 44582 18014 44634
rect 18194 44582 18196 44634
rect 17950 44580 17956 44582
rect 18012 44580 18036 44582
rect 18092 44580 18116 44582
rect 18172 44580 18196 44582
rect 18252 44580 18258 44582
rect 17950 44571 18258 44580
rect 16948 43988 17000 43994
rect 16948 43930 17000 43936
rect 17950 43548 18258 43557
rect 17950 43546 17956 43548
rect 18012 43546 18036 43548
rect 18092 43546 18116 43548
rect 18172 43546 18196 43548
rect 18252 43546 18258 43548
rect 18012 43494 18014 43546
rect 18194 43494 18196 43546
rect 17950 43492 17956 43494
rect 18012 43492 18036 43494
rect 18092 43492 18116 43494
rect 18172 43492 18196 43494
rect 18252 43492 18258 43494
rect 17950 43483 18258 43492
rect 19168 43450 19196 52430
rect 19628 43926 19656 53042
rect 20180 45554 20208 54062
rect 20272 53650 20300 56200
rect 21008 54262 21036 56200
rect 20996 54256 21048 54262
rect 20996 54198 21048 54204
rect 20352 54188 20404 54194
rect 20352 54130 20404 54136
rect 20260 53644 20312 53650
rect 20260 53586 20312 53592
rect 20364 50998 20392 54130
rect 21744 53650 21772 56200
rect 22480 54126 22508 56200
rect 23216 55214 23244 56200
rect 23216 55186 23336 55214
rect 22744 54188 22796 54194
rect 22744 54130 22796 54136
rect 22468 54120 22520 54126
rect 22468 54062 22520 54068
rect 21732 53644 21784 53650
rect 21732 53586 21784 53592
rect 22192 53508 22244 53514
rect 22192 53450 22244 53456
rect 20444 53440 20496 53446
rect 20444 53382 20496 53388
rect 20352 50992 20404 50998
rect 20352 50934 20404 50940
rect 20180 45526 20392 45554
rect 19616 43920 19668 43926
rect 19616 43862 19668 43868
rect 19984 43716 20036 43722
rect 19984 43658 20036 43664
rect 16856 43444 16908 43450
rect 16856 43386 16908 43392
rect 19156 43444 19208 43450
rect 19156 43386 19208 43392
rect 19064 43308 19116 43314
rect 19064 43250 19116 43256
rect 17950 42460 18258 42469
rect 17950 42458 17956 42460
rect 18012 42458 18036 42460
rect 18092 42458 18116 42460
rect 18172 42458 18196 42460
rect 18252 42458 18258 42460
rect 18012 42406 18014 42458
rect 18194 42406 18196 42458
rect 17950 42404 17956 42406
rect 18012 42404 18036 42406
rect 18092 42404 18116 42406
rect 18172 42404 18196 42406
rect 18252 42404 18258 42406
rect 17950 42395 18258 42404
rect 17408 42220 17460 42226
rect 17408 42162 17460 42168
rect 17316 42152 17368 42158
rect 17316 42094 17368 42100
rect 14924 37120 14976 37126
rect 14924 37062 14976 37068
rect 17224 36780 17276 36786
rect 17224 36722 17276 36728
rect 17236 32570 17264 36722
rect 17224 32564 17276 32570
rect 17224 32506 17276 32512
rect 17328 29306 17356 42094
rect 17316 29300 17368 29306
rect 17316 29242 17368 29248
rect 17420 29186 17448 42162
rect 17950 41372 18258 41381
rect 17950 41370 17956 41372
rect 18012 41370 18036 41372
rect 18092 41370 18116 41372
rect 18172 41370 18196 41372
rect 18252 41370 18258 41372
rect 18012 41318 18014 41370
rect 18194 41318 18196 41370
rect 17950 41316 17956 41318
rect 18012 41316 18036 41318
rect 18092 41316 18116 41318
rect 18172 41316 18196 41318
rect 18252 41316 18258 41318
rect 17950 41307 18258 41316
rect 17950 40284 18258 40293
rect 17950 40282 17956 40284
rect 18012 40282 18036 40284
rect 18092 40282 18116 40284
rect 18172 40282 18196 40284
rect 18252 40282 18258 40284
rect 18012 40230 18014 40282
rect 18194 40230 18196 40282
rect 17950 40228 17956 40230
rect 18012 40228 18036 40230
rect 18092 40228 18116 40230
rect 18172 40228 18196 40230
rect 18252 40228 18258 40230
rect 17950 40219 18258 40228
rect 17950 39196 18258 39205
rect 17950 39194 17956 39196
rect 18012 39194 18036 39196
rect 18092 39194 18116 39196
rect 18172 39194 18196 39196
rect 18252 39194 18258 39196
rect 18012 39142 18014 39194
rect 18194 39142 18196 39194
rect 17950 39140 17956 39142
rect 18012 39140 18036 39142
rect 18092 39140 18116 39142
rect 18172 39140 18196 39142
rect 18252 39140 18258 39142
rect 17950 39131 18258 39140
rect 17950 38108 18258 38117
rect 17950 38106 17956 38108
rect 18012 38106 18036 38108
rect 18092 38106 18116 38108
rect 18172 38106 18196 38108
rect 18252 38106 18258 38108
rect 18012 38054 18014 38106
rect 18194 38054 18196 38106
rect 17950 38052 17956 38054
rect 18012 38052 18036 38054
rect 18092 38052 18116 38054
rect 18172 38052 18196 38054
rect 18252 38052 18258 38054
rect 17950 38043 18258 38052
rect 17950 37020 18258 37029
rect 17950 37018 17956 37020
rect 18012 37018 18036 37020
rect 18092 37018 18116 37020
rect 18172 37018 18196 37020
rect 18252 37018 18258 37020
rect 18012 36966 18014 37018
rect 18194 36966 18196 37018
rect 17950 36964 17956 36966
rect 18012 36964 18036 36966
rect 18092 36964 18116 36966
rect 18172 36964 18196 36966
rect 18252 36964 18258 36966
rect 17950 36955 18258 36964
rect 17950 35932 18258 35941
rect 17950 35930 17956 35932
rect 18012 35930 18036 35932
rect 18092 35930 18116 35932
rect 18172 35930 18196 35932
rect 18252 35930 18258 35932
rect 18012 35878 18014 35930
rect 18194 35878 18196 35930
rect 17950 35876 17956 35878
rect 18012 35876 18036 35878
rect 18092 35876 18116 35878
rect 18172 35876 18196 35878
rect 18252 35876 18258 35878
rect 17950 35867 18258 35876
rect 17868 35624 17920 35630
rect 17868 35566 17920 35572
rect 17880 32366 17908 35566
rect 17950 34844 18258 34853
rect 17950 34842 17956 34844
rect 18012 34842 18036 34844
rect 18092 34842 18116 34844
rect 18172 34842 18196 34844
rect 18252 34842 18258 34844
rect 18012 34790 18014 34842
rect 18194 34790 18196 34842
rect 17950 34788 17956 34790
rect 18012 34788 18036 34790
rect 18092 34788 18116 34790
rect 18172 34788 18196 34790
rect 18252 34788 18258 34790
rect 17950 34779 18258 34788
rect 17950 33756 18258 33765
rect 17950 33754 17956 33756
rect 18012 33754 18036 33756
rect 18092 33754 18116 33756
rect 18172 33754 18196 33756
rect 18252 33754 18258 33756
rect 18012 33702 18014 33754
rect 18194 33702 18196 33754
rect 17950 33700 17956 33702
rect 18012 33700 18036 33702
rect 18092 33700 18116 33702
rect 18172 33700 18196 33702
rect 18252 33700 18258 33702
rect 17950 33691 18258 33700
rect 17950 32668 18258 32677
rect 17950 32666 17956 32668
rect 18012 32666 18036 32668
rect 18092 32666 18116 32668
rect 18172 32666 18196 32668
rect 18252 32666 18258 32668
rect 18012 32614 18014 32666
rect 18194 32614 18196 32666
rect 17950 32612 17956 32614
rect 18012 32612 18036 32614
rect 18092 32612 18116 32614
rect 18172 32612 18196 32614
rect 18252 32612 18258 32614
rect 17950 32603 18258 32612
rect 17868 32360 17920 32366
rect 17868 32302 17920 32308
rect 18512 32224 18564 32230
rect 18512 32166 18564 32172
rect 17950 31580 18258 31589
rect 17950 31578 17956 31580
rect 18012 31578 18036 31580
rect 18092 31578 18116 31580
rect 18172 31578 18196 31580
rect 18252 31578 18258 31580
rect 18012 31526 18014 31578
rect 18194 31526 18196 31578
rect 17950 31524 17956 31526
rect 18012 31524 18036 31526
rect 18092 31524 18116 31526
rect 18172 31524 18196 31526
rect 18252 31524 18258 31526
rect 17950 31515 18258 31524
rect 17950 30492 18258 30501
rect 17950 30490 17956 30492
rect 18012 30490 18036 30492
rect 18092 30490 18116 30492
rect 18172 30490 18196 30492
rect 18252 30490 18258 30492
rect 18012 30438 18014 30490
rect 18194 30438 18196 30490
rect 17950 30436 17956 30438
rect 18012 30436 18036 30438
rect 18092 30436 18116 30438
rect 18172 30436 18196 30438
rect 18252 30436 18258 30438
rect 17950 30427 18258 30436
rect 17950 29404 18258 29413
rect 17950 29402 17956 29404
rect 18012 29402 18036 29404
rect 18092 29402 18116 29404
rect 18172 29402 18196 29404
rect 18252 29402 18258 29404
rect 18012 29350 18014 29402
rect 18194 29350 18196 29402
rect 17950 29348 17956 29350
rect 18012 29348 18036 29350
rect 18092 29348 18116 29350
rect 18172 29348 18196 29350
rect 18252 29348 18258 29350
rect 17950 29339 18258 29348
rect 17236 29170 17448 29186
rect 17236 29164 17460 29170
rect 17236 29158 17408 29164
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14568 23662 14596 24278
rect 15292 24268 15344 24274
rect 15292 24210 15344 24216
rect 15200 24132 15252 24138
rect 15200 24074 15252 24080
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14568 22166 14596 23598
rect 15212 22642 15240 24074
rect 15304 23866 15332 24210
rect 15384 24132 15436 24138
rect 15384 24074 15436 24080
rect 15292 23860 15344 23866
rect 15292 23802 15344 23808
rect 15304 23186 15332 23802
rect 15396 23798 15424 24074
rect 16500 23866 16528 25230
rect 16488 23860 16540 23866
rect 16488 23802 16540 23808
rect 15384 23792 15436 23798
rect 15384 23734 15436 23740
rect 15292 23180 15344 23186
rect 15292 23122 15344 23128
rect 15396 22982 15424 23734
rect 15384 22976 15436 22982
rect 15384 22918 15436 22924
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 14752 22234 15148 22250
rect 14740 22228 15160 22234
rect 14792 22222 15108 22228
rect 14740 22170 14792 22176
rect 15108 22170 15160 22176
rect 14556 22160 14608 22166
rect 14556 22102 14608 22108
rect 15396 22094 15424 22918
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 15396 22066 15516 22094
rect 15488 21962 15516 22066
rect 15476 21956 15528 21962
rect 15476 21898 15528 21904
rect 16500 21672 16528 22170
rect 16408 21644 16528 21672
rect 16408 16182 16436 21644
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16500 19514 16528 21490
rect 16488 19508 16540 19514
rect 16488 19450 16540 19456
rect 16396 16176 16448 16182
rect 16396 16118 16448 16124
rect 16488 8560 16540 8566
rect 16488 8502 16540 8508
rect 16500 8362 16528 8502
rect 16488 8356 16540 8362
rect 16488 8298 16540 8304
rect 14464 3188 14516 3194
rect 14464 3130 14516 3136
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 11060 2372 11112 2378
rect 11060 2314 11112 2320
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11072 800 11100 2314
rect 11808 800 11836 2314
rect 12544 800 12572 2994
rect 12950 2748 13258 2757
rect 12950 2746 12956 2748
rect 13012 2746 13036 2748
rect 13092 2746 13116 2748
rect 13172 2746 13196 2748
rect 13252 2746 13258 2748
rect 13012 2694 13014 2746
rect 13194 2694 13196 2746
rect 12950 2692 12956 2694
rect 13012 2692 13036 2694
rect 13092 2692 13116 2694
rect 13172 2692 13196 2694
rect 13252 2692 13258 2694
rect 12950 2683 13258 2692
rect 13634 2680 13690 2689
rect 13634 2615 13636 2624
rect 13688 2615 13690 2624
rect 13636 2586 13688 2592
rect 13268 2372 13320 2378
rect 13268 2314 13320 2320
rect 13280 800 13308 2314
rect 14016 800 14044 2994
rect 17236 2922 17264 29158
rect 17408 29106 17460 29112
rect 17950 28316 18258 28325
rect 17950 28314 17956 28316
rect 18012 28314 18036 28316
rect 18092 28314 18116 28316
rect 18172 28314 18196 28316
rect 18252 28314 18258 28316
rect 18012 28262 18014 28314
rect 18194 28262 18196 28314
rect 17950 28260 17956 28262
rect 18012 28260 18036 28262
rect 18092 28260 18116 28262
rect 18172 28260 18196 28262
rect 18252 28260 18258 28262
rect 17950 28251 18258 28260
rect 17950 27228 18258 27237
rect 17950 27226 17956 27228
rect 18012 27226 18036 27228
rect 18092 27226 18116 27228
rect 18172 27226 18196 27228
rect 18252 27226 18258 27228
rect 18012 27174 18014 27226
rect 18194 27174 18196 27226
rect 17950 27172 17956 27174
rect 18012 27172 18036 27174
rect 18092 27172 18116 27174
rect 18172 27172 18196 27174
rect 18252 27172 18258 27174
rect 17950 27163 18258 27172
rect 17950 26140 18258 26149
rect 17950 26138 17956 26140
rect 18012 26138 18036 26140
rect 18092 26138 18116 26140
rect 18172 26138 18196 26140
rect 18252 26138 18258 26140
rect 18012 26086 18014 26138
rect 18194 26086 18196 26138
rect 17950 26084 17956 26086
rect 18012 26084 18036 26086
rect 18092 26084 18116 26086
rect 18172 26084 18196 26086
rect 18252 26084 18258 26086
rect 17950 26075 18258 26084
rect 17950 25052 18258 25061
rect 17950 25050 17956 25052
rect 18012 25050 18036 25052
rect 18092 25050 18116 25052
rect 18172 25050 18196 25052
rect 18252 25050 18258 25052
rect 18012 24998 18014 25050
rect 18194 24998 18196 25050
rect 17950 24996 17956 24998
rect 18012 24996 18036 24998
rect 18092 24996 18116 24998
rect 18172 24996 18196 24998
rect 18252 24996 18258 24998
rect 17950 24987 18258 24996
rect 17950 23964 18258 23973
rect 17950 23962 17956 23964
rect 18012 23962 18036 23964
rect 18092 23962 18116 23964
rect 18172 23962 18196 23964
rect 18252 23962 18258 23964
rect 18012 23910 18014 23962
rect 18194 23910 18196 23962
rect 17950 23908 17956 23910
rect 18012 23908 18036 23910
rect 18092 23908 18116 23910
rect 18172 23908 18196 23910
rect 18252 23908 18258 23910
rect 17950 23899 18258 23908
rect 17408 23044 17460 23050
rect 17408 22986 17460 22992
rect 17420 22710 17448 22986
rect 17950 22876 18258 22885
rect 17950 22874 17956 22876
rect 18012 22874 18036 22876
rect 18092 22874 18116 22876
rect 18172 22874 18196 22876
rect 18252 22874 18258 22876
rect 18012 22822 18014 22874
rect 18194 22822 18196 22874
rect 17950 22820 17956 22822
rect 18012 22820 18036 22822
rect 18092 22820 18116 22822
rect 18172 22820 18196 22822
rect 18252 22820 18258 22822
rect 17950 22811 18258 22820
rect 17408 22704 17460 22710
rect 17408 22646 17460 22652
rect 17408 22432 17460 22438
rect 17408 22374 17460 22380
rect 17420 21690 17448 22374
rect 18524 22094 18552 32166
rect 19076 31754 19104 43250
rect 19432 43240 19484 43246
rect 19432 43182 19484 43188
rect 19444 36922 19472 43182
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19996 34746 20024 43658
rect 20364 43450 20392 45526
rect 20456 43994 20484 53382
rect 21272 53168 21324 53174
rect 21272 53110 21324 53116
rect 20904 49904 20956 49910
rect 20904 49846 20956 49852
rect 20628 49224 20680 49230
rect 20628 49166 20680 49172
rect 20536 45892 20588 45898
rect 20536 45834 20588 45840
rect 20444 43988 20496 43994
rect 20444 43930 20496 43936
rect 20444 43716 20496 43722
rect 20444 43658 20496 43664
rect 20352 43444 20404 43450
rect 20352 43386 20404 43392
rect 20260 43308 20312 43314
rect 20260 43250 20312 43256
rect 19984 34740 20036 34746
rect 19984 34682 20036 34688
rect 18708 31726 19104 31754
rect 18708 30054 18736 31726
rect 20272 30394 20300 43250
rect 20456 34406 20484 43658
rect 20548 40730 20576 45834
rect 20640 42362 20668 49166
rect 20916 43450 20944 49846
rect 21088 48204 21140 48210
rect 21088 48146 21140 48152
rect 20996 43648 21048 43654
rect 20996 43590 21048 43596
rect 21008 43450 21036 43590
rect 20904 43444 20956 43450
rect 20904 43386 20956 43392
rect 20996 43444 21048 43450
rect 20996 43386 21048 43392
rect 20628 42356 20680 42362
rect 20628 42298 20680 42304
rect 20812 42220 20864 42226
rect 20812 42162 20864 42168
rect 20536 40724 20588 40730
rect 20536 40666 20588 40672
rect 20444 34400 20496 34406
rect 20444 34342 20496 34348
rect 20824 34202 20852 42162
rect 21100 39982 21128 48146
rect 21284 43994 21312 53110
rect 22204 51066 22232 53450
rect 22756 52154 22784 54130
rect 22950 53884 23258 53893
rect 22950 53882 22956 53884
rect 23012 53882 23036 53884
rect 23092 53882 23116 53884
rect 23172 53882 23196 53884
rect 23252 53882 23258 53884
rect 23012 53830 23014 53882
rect 23194 53830 23196 53882
rect 22950 53828 22956 53830
rect 23012 53828 23036 53830
rect 23092 53828 23116 53830
rect 23172 53828 23196 53830
rect 23252 53828 23258 53830
rect 22950 53819 23258 53828
rect 23308 53582 23336 55186
rect 23952 53582 23980 56200
rect 24688 54194 24716 56200
rect 25424 54194 25452 56200
rect 26160 54210 26188 56200
rect 26160 54194 26280 54210
rect 26896 54194 26924 56200
rect 27632 54194 27660 56200
rect 27950 54428 28258 54437
rect 27950 54426 27956 54428
rect 28012 54426 28036 54428
rect 28092 54426 28116 54428
rect 28172 54426 28196 54428
rect 28252 54426 28258 54428
rect 28012 54374 28014 54426
rect 28194 54374 28196 54426
rect 27950 54372 27956 54374
rect 28012 54372 28036 54374
rect 28092 54372 28116 54374
rect 28172 54372 28196 54374
rect 28252 54372 28258 54374
rect 27950 54363 28258 54372
rect 28368 54262 28396 56200
rect 28356 54256 28408 54262
rect 28356 54198 28408 54204
rect 24676 54188 24728 54194
rect 24676 54130 24728 54136
rect 25412 54188 25464 54194
rect 26160 54188 26292 54194
rect 26160 54182 26240 54188
rect 25412 54130 25464 54136
rect 26240 54130 26292 54136
rect 26884 54188 26936 54194
rect 26884 54130 26936 54136
rect 27620 54188 27672 54194
rect 27620 54130 27672 54136
rect 24952 53984 25004 53990
rect 24950 53952 24952 53961
rect 25688 53984 25740 53990
rect 25004 53952 25006 53961
rect 25688 53926 25740 53932
rect 26240 53984 26292 53990
rect 26240 53926 26292 53932
rect 27436 53984 27488 53990
rect 27436 53926 27488 53932
rect 28540 53984 28592 53990
rect 28540 53926 28592 53932
rect 24950 53887 25006 53896
rect 22836 53576 22888 53582
rect 22836 53518 22888 53524
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 23940 53576 23992 53582
rect 23940 53518 23992 53524
rect 22744 52148 22796 52154
rect 22744 52090 22796 52096
rect 22848 51610 22876 53518
rect 24952 53508 25004 53514
rect 24952 53450 25004 53456
rect 22950 52796 23258 52805
rect 22950 52794 22956 52796
rect 23012 52794 23036 52796
rect 23092 52794 23116 52796
rect 23172 52794 23196 52796
rect 23252 52794 23258 52796
rect 23012 52742 23014 52794
rect 23194 52742 23196 52794
rect 22950 52740 22956 52742
rect 23012 52740 23036 52742
rect 23092 52740 23116 52742
rect 23172 52740 23196 52742
rect 23252 52740 23258 52742
rect 22950 52731 23258 52740
rect 23756 52012 23808 52018
rect 23756 51954 23808 51960
rect 22950 51708 23258 51717
rect 22950 51706 22956 51708
rect 23012 51706 23036 51708
rect 23092 51706 23116 51708
rect 23172 51706 23196 51708
rect 23252 51706 23258 51708
rect 23012 51654 23014 51706
rect 23194 51654 23196 51706
rect 22950 51652 22956 51654
rect 23012 51652 23036 51654
rect 23092 51652 23116 51654
rect 23172 51652 23196 51654
rect 23252 51652 23258 51654
rect 22950 51643 23258 51652
rect 22836 51604 22888 51610
rect 22836 51546 22888 51552
rect 22192 51060 22244 51066
rect 22192 51002 22244 51008
rect 22744 50924 22796 50930
rect 22744 50866 22796 50872
rect 22284 50244 22336 50250
rect 22284 50186 22336 50192
rect 22192 49156 22244 49162
rect 22192 49098 22244 49104
rect 22100 48068 22152 48074
rect 22100 48010 22152 48016
rect 22008 45960 22060 45966
rect 22008 45902 22060 45908
rect 21272 43988 21324 43994
rect 21272 43930 21324 43936
rect 21916 43784 21968 43790
rect 21916 43726 21968 43732
rect 21732 43308 21784 43314
rect 21732 43250 21784 43256
rect 21548 42900 21600 42906
rect 21548 42842 21600 42848
rect 21088 39976 21140 39982
rect 21088 39918 21140 39924
rect 21100 38418 21128 39918
rect 21088 38412 21140 38418
rect 21088 38354 21140 38360
rect 21100 35834 21128 38354
rect 21364 38276 21416 38282
rect 21364 38218 21416 38224
rect 21376 36718 21404 38218
rect 21364 36712 21416 36718
rect 21364 36654 21416 36660
rect 21376 35834 21404 36654
rect 21088 35828 21140 35834
rect 21088 35770 21140 35776
rect 21364 35828 21416 35834
rect 21364 35770 21416 35776
rect 21100 35630 21128 35770
rect 21088 35624 21140 35630
rect 21088 35566 21140 35572
rect 20812 34196 20864 34202
rect 20812 34138 20864 34144
rect 21456 33516 21508 33522
rect 21456 33458 21508 33464
rect 21468 30938 21496 33458
rect 21560 32774 21588 42842
rect 21744 36106 21772 43250
rect 21824 36780 21876 36786
rect 21824 36722 21876 36728
rect 21732 36100 21784 36106
rect 21732 36042 21784 36048
rect 21836 35290 21864 36722
rect 21928 36378 21956 43726
rect 22020 40662 22048 45902
rect 22112 41562 22140 48010
rect 22204 42362 22232 49098
rect 22296 43994 22324 50186
rect 22468 45620 22520 45626
rect 22468 45562 22520 45568
rect 22284 43988 22336 43994
rect 22284 43930 22336 43936
rect 22192 42356 22244 42362
rect 22192 42298 22244 42304
rect 22376 42220 22428 42226
rect 22376 42162 22428 42168
rect 22112 41534 22232 41562
rect 22100 41472 22152 41478
rect 22100 41414 22152 41420
rect 22112 41274 22140 41414
rect 22100 41268 22152 41274
rect 22100 41210 22152 41216
rect 22204 41206 22232 41534
rect 22388 41414 22416 42162
rect 22480 41698 22508 45562
rect 22756 45082 22784 50866
rect 22950 50620 23258 50629
rect 22950 50618 22956 50620
rect 23012 50618 23036 50620
rect 23092 50618 23116 50620
rect 23172 50618 23196 50620
rect 23252 50618 23258 50620
rect 23012 50566 23014 50618
rect 23194 50566 23196 50618
rect 22950 50564 22956 50566
rect 23012 50564 23036 50566
rect 23092 50564 23116 50566
rect 23172 50564 23196 50566
rect 23252 50564 23258 50566
rect 22950 50555 23258 50564
rect 22950 49532 23258 49541
rect 22950 49530 22956 49532
rect 23012 49530 23036 49532
rect 23092 49530 23116 49532
rect 23172 49530 23196 49532
rect 23252 49530 23258 49532
rect 23012 49478 23014 49530
rect 23194 49478 23196 49530
rect 22950 49476 22956 49478
rect 23012 49476 23036 49478
rect 23092 49476 23116 49478
rect 23172 49476 23196 49478
rect 23252 49476 23258 49478
rect 22950 49467 23258 49476
rect 22950 48444 23258 48453
rect 22950 48442 22956 48444
rect 23012 48442 23036 48444
rect 23092 48442 23116 48444
rect 23172 48442 23196 48444
rect 23252 48442 23258 48444
rect 23012 48390 23014 48442
rect 23194 48390 23196 48442
rect 22950 48388 22956 48390
rect 23012 48388 23036 48390
rect 23092 48388 23116 48390
rect 23172 48388 23196 48390
rect 23252 48388 23258 48390
rect 22950 48379 23258 48388
rect 23768 47802 23796 51954
rect 24124 50924 24176 50930
rect 24124 50866 24176 50872
rect 23756 47796 23808 47802
rect 23756 47738 23808 47744
rect 22950 47356 23258 47365
rect 22950 47354 22956 47356
rect 23012 47354 23036 47356
rect 23092 47354 23116 47356
rect 23172 47354 23196 47356
rect 23252 47354 23258 47356
rect 23012 47302 23014 47354
rect 23194 47302 23196 47354
rect 22950 47300 22956 47302
rect 23012 47300 23036 47302
rect 23092 47300 23116 47302
rect 23172 47300 23196 47302
rect 23252 47300 23258 47302
rect 22950 47291 23258 47300
rect 22950 46268 23258 46277
rect 22950 46266 22956 46268
rect 23012 46266 23036 46268
rect 23092 46266 23116 46268
rect 23172 46266 23196 46268
rect 23252 46266 23258 46268
rect 23012 46214 23014 46266
rect 23194 46214 23196 46266
rect 22950 46212 22956 46214
rect 23012 46212 23036 46214
rect 23092 46212 23116 46214
rect 23172 46212 23196 46214
rect 23252 46212 23258 46214
rect 22950 46203 23258 46212
rect 22950 45180 23258 45189
rect 22950 45178 22956 45180
rect 23012 45178 23036 45180
rect 23092 45178 23116 45180
rect 23172 45178 23196 45180
rect 23252 45178 23258 45180
rect 23012 45126 23014 45178
rect 23194 45126 23196 45178
rect 22950 45124 22956 45126
rect 23012 45124 23036 45126
rect 23092 45124 23116 45126
rect 23172 45124 23196 45126
rect 23252 45124 23258 45126
rect 22950 45115 23258 45124
rect 24136 45082 24164 50866
rect 24860 47660 24912 47666
rect 24860 47602 24912 47608
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 24124 45076 24176 45082
rect 24124 45018 24176 45024
rect 24492 44872 24544 44878
rect 24492 44814 24544 44820
rect 22950 44092 23258 44101
rect 22950 44090 22956 44092
rect 23012 44090 23036 44092
rect 23092 44090 23116 44092
rect 23172 44090 23196 44092
rect 23252 44090 23258 44092
rect 23012 44038 23014 44090
rect 23194 44038 23196 44090
rect 22950 44036 22956 44038
rect 23012 44036 23036 44038
rect 23092 44036 23116 44038
rect 23172 44036 23196 44038
rect 23252 44036 23258 44038
rect 22950 44027 23258 44036
rect 23296 43784 23348 43790
rect 23296 43726 23348 43732
rect 22950 43004 23258 43013
rect 22950 43002 22956 43004
rect 23012 43002 23036 43004
rect 23092 43002 23116 43004
rect 23172 43002 23196 43004
rect 23252 43002 23258 43004
rect 23012 42950 23014 43002
rect 23194 42950 23196 43002
rect 22950 42948 22956 42950
rect 23012 42948 23036 42950
rect 23092 42948 23116 42950
rect 23172 42948 23196 42950
rect 23252 42948 23258 42950
rect 22950 42939 23258 42948
rect 22950 41916 23258 41925
rect 22950 41914 22956 41916
rect 23012 41914 23036 41916
rect 23092 41914 23116 41916
rect 23172 41914 23196 41916
rect 23252 41914 23258 41916
rect 23012 41862 23014 41914
rect 23194 41862 23196 41914
rect 22950 41860 22956 41862
rect 23012 41860 23036 41862
rect 23092 41860 23116 41862
rect 23172 41860 23196 41862
rect 23252 41860 23258 41862
rect 22950 41851 23258 41860
rect 22480 41670 22600 41698
rect 22468 41540 22520 41546
rect 22468 41482 22520 41488
rect 22296 41386 22416 41414
rect 22192 41200 22244 41206
rect 22192 41142 22244 41148
rect 22008 40656 22060 40662
rect 22008 40598 22060 40604
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 22112 37466 22140 40326
rect 22192 39432 22244 39438
rect 22192 39374 22244 39380
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 21916 36372 21968 36378
rect 21916 36314 21968 36320
rect 22008 35624 22060 35630
rect 22008 35566 22060 35572
rect 21824 35284 21876 35290
rect 21824 35226 21876 35232
rect 22020 35154 22048 35566
rect 22008 35148 22060 35154
rect 22008 35090 22060 35096
rect 22020 34066 22048 35090
rect 22100 35012 22152 35018
rect 22204 35000 22232 39374
rect 22152 34972 22232 35000
rect 22100 34954 22152 34960
rect 22008 34060 22060 34066
rect 22008 34002 22060 34008
rect 21548 32768 21600 32774
rect 21548 32710 21600 32716
rect 21824 31816 21876 31822
rect 21824 31758 21876 31764
rect 21456 30932 21508 30938
rect 21456 30874 21508 30880
rect 21836 30734 21864 31758
rect 22112 30802 22140 34954
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22100 30796 22152 30802
rect 22100 30738 22152 30744
rect 21824 30728 21876 30734
rect 21824 30670 21876 30676
rect 21916 30660 21968 30666
rect 21916 30602 21968 30608
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18432 22066 18552 22094
rect 17950 21788 18258 21797
rect 17950 21786 17956 21788
rect 18012 21786 18036 21788
rect 18092 21786 18116 21788
rect 18172 21786 18196 21788
rect 18252 21786 18258 21788
rect 18012 21734 18014 21786
rect 18194 21734 18196 21786
rect 17950 21732 17956 21734
rect 18012 21732 18036 21734
rect 18092 21732 18116 21734
rect 18172 21732 18196 21734
rect 18252 21732 18258 21734
rect 17950 21723 18258 21732
rect 17408 21684 17460 21690
rect 17408 21626 17460 21632
rect 17950 20700 18258 20709
rect 17950 20698 17956 20700
rect 18012 20698 18036 20700
rect 18092 20698 18116 20700
rect 18172 20698 18196 20700
rect 18252 20698 18258 20700
rect 18012 20646 18014 20698
rect 18194 20646 18196 20698
rect 17950 20644 17956 20646
rect 18012 20644 18036 20646
rect 18092 20644 18116 20646
rect 18172 20644 18196 20646
rect 18252 20644 18258 20646
rect 17950 20635 18258 20644
rect 17868 19848 17920 19854
rect 17868 19790 17920 19796
rect 17880 17882 17908 19790
rect 18432 19718 18460 22066
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 17950 19612 18258 19621
rect 17950 19610 17956 19612
rect 18012 19610 18036 19612
rect 18092 19610 18116 19612
rect 18172 19610 18196 19612
rect 18252 19610 18258 19612
rect 18012 19558 18014 19610
rect 18194 19558 18196 19610
rect 17950 19556 17956 19558
rect 18012 19556 18036 19558
rect 18092 19556 18116 19558
rect 18172 19556 18196 19558
rect 18252 19556 18258 19558
rect 17950 19547 18258 19556
rect 17950 18524 18258 18533
rect 17950 18522 17956 18524
rect 18012 18522 18036 18524
rect 18092 18522 18116 18524
rect 18172 18522 18196 18524
rect 18252 18522 18258 18524
rect 18012 18470 18014 18522
rect 18194 18470 18196 18522
rect 17950 18468 17956 18470
rect 18012 18468 18036 18470
rect 18092 18468 18116 18470
rect 18172 18468 18196 18470
rect 18252 18468 18258 18470
rect 17950 18459 18258 18468
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17950 17436 18258 17445
rect 17950 17434 17956 17436
rect 18012 17434 18036 17436
rect 18092 17434 18116 17436
rect 18172 17434 18196 17436
rect 18252 17434 18258 17436
rect 18012 17382 18014 17434
rect 18194 17382 18196 17434
rect 17950 17380 17956 17382
rect 18012 17380 18036 17382
rect 18092 17380 18116 17382
rect 18172 17380 18196 17382
rect 18252 17380 18258 17382
rect 17950 17371 18258 17380
rect 17950 16348 18258 16357
rect 17950 16346 17956 16348
rect 18012 16346 18036 16348
rect 18092 16346 18116 16348
rect 18172 16346 18196 16348
rect 18252 16346 18258 16348
rect 18012 16294 18014 16346
rect 18194 16294 18196 16346
rect 17950 16292 17956 16294
rect 18012 16292 18036 16294
rect 18092 16292 18116 16294
rect 18172 16292 18196 16294
rect 18252 16292 18258 16294
rect 17950 16283 18258 16292
rect 17950 15260 18258 15269
rect 17950 15258 17956 15260
rect 18012 15258 18036 15260
rect 18092 15258 18116 15260
rect 18172 15258 18196 15260
rect 18252 15258 18258 15260
rect 18012 15206 18014 15258
rect 18194 15206 18196 15258
rect 17950 15204 17956 15206
rect 18012 15204 18036 15206
rect 18092 15204 18116 15206
rect 18172 15204 18196 15206
rect 18252 15204 18258 15206
rect 17950 15195 18258 15204
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17880 11354 17908 14962
rect 17950 14172 18258 14181
rect 17950 14170 17956 14172
rect 18012 14170 18036 14172
rect 18092 14170 18116 14172
rect 18172 14170 18196 14172
rect 18252 14170 18258 14172
rect 18012 14118 18014 14170
rect 18194 14118 18196 14170
rect 17950 14116 17956 14118
rect 18012 14116 18036 14118
rect 18092 14116 18116 14118
rect 18172 14116 18196 14118
rect 18252 14116 18258 14118
rect 17950 14107 18258 14116
rect 17950 13084 18258 13093
rect 17950 13082 17956 13084
rect 18012 13082 18036 13084
rect 18092 13082 18116 13084
rect 18172 13082 18196 13084
rect 18252 13082 18258 13084
rect 18012 13030 18014 13082
rect 18194 13030 18196 13082
rect 17950 13028 17956 13030
rect 18012 13028 18036 13030
rect 18092 13028 18116 13030
rect 18172 13028 18196 13030
rect 18252 13028 18258 13030
rect 17950 13019 18258 13028
rect 17950 11996 18258 12005
rect 17950 11994 17956 11996
rect 18012 11994 18036 11996
rect 18092 11994 18116 11996
rect 18172 11994 18196 11996
rect 18252 11994 18258 11996
rect 18012 11942 18014 11994
rect 18194 11942 18196 11994
rect 17950 11940 17956 11942
rect 18012 11940 18036 11942
rect 18092 11940 18116 11942
rect 18172 11940 18196 11942
rect 18252 11940 18258 11942
rect 17950 11931 18258 11940
rect 17868 11348 17920 11354
rect 17868 11290 17920 11296
rect 17950 10908 18258 10917
rect 17950 10906 17956 10908
rect 18012 10906 18036 10908
rect 18092 10906 18116 10908
rect 18172 10906 18196 10908
rect 18252 10906 18258 10908
rect 18012 10854 18014 10906
rect 18194 10854 18196 10906
rect 17950 10852 17956 10854
rect 18012 10852 18036 10854
rect 18092 10852 18116 10854
rect 18172 10852 18196 10854
rect 18252 10852 18258 10854
rect 17950 10843 18258 10852
rect 17950 9820 18258 9829
rect 17950 9818 17956 9820
rect 18012 9818 18036 9820
rect 18092 9818 18116 9820
rect 18172 9818 18196 9820
rect 18252 9818 18258 9820
rect 18012 9766 18014 9818
rect 18194 9766 18196 9818
rect 17950 9764 17956 9766
rect 18012 9764 18036 9766
rect 18092 9764 18116 9766
rect 18172 9764 18196 9766
rect 18252 9764 18258 9766
rect 17950 9755 18258 9764
rect 17950 8732 18258 8741
rect 17950 8730 17956 8732
rect 18012 8730 18036 8732
rect 18092 8730 18116 8732
rect 18172 8730 18196 8732
rect 18252 8730 18258 8732
rect 18012 8678 18014 8730
rect 18194 8678 18196 8730
rect 17950 8676 17956 8678
rect 18012 8676 18036 8678
rect 18092 8676 18116 8678
rect 18172 8676 18196 8678
rect 18252 8676 18258 8678
rect 17950 8667 18258 8676
rect 17950 7644 18258 7653
rect 17950 7642 17956 7644
rect 18012 7642 18036 7644
rect 18092 7642 18116 7644
rect 18172 7642 18196 7644
rect 18252 7642 18258 7644
rect 18012 7590 18014 7642
rect 18194 7590 18196 7642
rect 17950 7588 17956 7590
rect 18012 7588 18036 7590
rect 18092 7588 18116 7590
rect 18172 7588 18196 7590
rect 18252 7588 18258 7590
rect 17950 7579 18258 7588
rect 17950 6556 18258 6565
rect 17950 6554 17956 6556
rect 18012 6554 18036 6556
rect 18092 6554 18116 6556
rect 18172 6554 18196 6556
rect 18252 6554 18258 6556
rect 18012 6502 18014 6554
rect 18194 6502 18196 6554
rect 17950 6500 17956 6502
rect 18012 6500 18036 6502
rect 18092 6500 18116 6502
rect 18172 6500 18196 6502
rect 18252 6500 18258 6502
rect 17950 6491 18258 6500
rect 17950 5468 18258 5477
rect 17950 5466 17956 5468
rect 18012 5466 18036 5468
rect 18092 5466 18116 5468
rect 18172 5466 18196 5468
rect 18252 5466 18258 5468
rect 18012 5414 18014 5466
rect 18194 5414 18196 5466
rect 17950 5412 17956 5414
rect 18012 5412 18036 5414
rect 18092 5412 18116 5414
rect 18172 5412 18196 5414
rect 18252 5412 18258 5414
rect 17950 5403 18258 5412
rect 17950 4380 18258 4389
rect 17950 4378 17956 4380
rect 18012 4378 18036 4380
rect 18092 4378 18116 4380
rect 18172 4378 18196 4380
rect 18252 4378 18258 4380
rect 18012 4326 18014 4378
rect 18194 4326 18196 4378
rect 17950 4324 17956 4326
rect 18012 4324 18036 4326
rect 18092 4324 18116 4326
rect 18172 4324 18196 4326
rect 18252 4324 18258 4326
rect 17950 4315 18258 4324
rect 18328 3664 18380 3670
rect 18328 3606 18380 3612
rect 17950 3292 18258 3301
rect 17950 3290 17956 3292
rect 18012 3290 18036 3292
rect 18092 3290 18116 3292
rect 18172 3290 18196 3292
rect 18252 3290 18258 3292
rect 18012 3238 18014 3290
rect 18194 3238 18196 3290
rect 17950 3236 17956 3238
rect 18012 3236 18036 3238
rect 18092 3236 18116 3238
rect 18172 3236 18196 3238
rect 18252 3236 18258 3238
rect 17950 3227 18258 3236
rect 18340 3058 18368 3606
rect 18432 3126 18460 19654
rect 18604 16652 18656 16658
rect 18604 16594 18656 16600
rect 18616 8498 18644 16594
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 17684 3052 17736 3058
rect 17684 2994 17736 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14752 800 14780 2382
rect 15476 2372 15528 2378
rect 15476 2314 15528 2320
rect 16212 2372 16264 2378
rect 16212 2314 16264 2320
rect 16304 2372 16356 2378
rect 16304 2314 16356 2320
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 15488 800 15516 2314
rect 16224 800 16252 2314
rect 16316 2106 16344 2314
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16960 800 16988 2314
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 17132 2032 17184 2038
rect 17132 1974 17184 1980
rect 17144 1630 17172 1974
rect 17328 1970 17356 2246
rect 17316 1964 17368 1970
rect 17316 1906 17368 1912
rect 17420 1902 17448 2246
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17132 1624 17184 1630
rect 17132 1566 17184 1572
rect 17696 800 17724 2994
rect 18708 2650 18736 29990
rect 19524 28620 19576 28626
rect 19524 28562 19576 28568
rect 18880 22976 18932 22982
rect 18880 22918 18932 22924
rect 18892 22642 18920 22918
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 19432 22092 19484 22098
rect 19432 22034 19484 22040
rect 19340 19984 19392 19990
rect 19340 19926 19392 19932
rect 18788 18964 18840 18970
rect 18788 18906 18840 18912
rect 18800 18154 18828 18906
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 19248 17672 19300 17678
rect 19248 17614 19300 17620
rect 18788 17536 18840 17542
rect 18788 17478 18840 17484
rect 18800 16250 18828 17478
rect 19260 17134 19288 17614
rect 19248 17128 19300 17134
rect 19248 17070 19300 17076
rect 19260 16658 19288 17070
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19248 16448 19300 16454
rect 19248 16390 19300 16396
rect 18788 16244 18840 16250
rect 18788 16186 18840 16192
rect 18800 2922 18828 16186
rect 19260 8566 19288 16390
rect 19352 15162 19380 19926
rect 19444 19922 19472 22034
rect 19536 21554 19564 28562
rect 21640 28552 21692 28558
rect 21692 28500 21864 28506
rect 21640 28494 21864 28500
rect 21652 28490 21864 28494
rect 21652 28484 21876 28490
rect 21652 28478 21824 28484
rect 21824 28426 21876 28432
rect 20996 24880 21048 24886
rect 20996 24822 21048 24828
rect 19708 24744 19760 24750
rect 19708 24686 19760 24692
rect 19720 24274 19748 24686
rect 19708 24268 19760 24274
rect 19708 24210 19760 24216
rect 19720 23186 19748 24210
rect 19708 23180 19760 23186
rect 19708 23122 19760 23128
rect 21008 23050 21036 24822
rect 21272 24744 21324 24750
rect 21272 24686 21324 24692
rect 21284 24070 21312 24686
rect 21928 24682 21956 30602
rect 22112 30161 22140 30738
rect 22098 30152 22154 30161
rect 22098 30087 22154 30096
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22008 28620 22060 28626
rect 22008 28562 22060 28568
rect 22020 28422 22048 28562
rect 22008 28416 22060 28422
rect 22008 28358 22060 28364
rect 22008 28076 22060 28082
rect 22008 28018 22060 28024
rect 21732 24676 21784 24682
rect 21732 24618 21784 24624
rect 21916 24676 21968 24682
rect 21916 24618 21968 24624
rect 21456 24608 21508 24614
rect 21456 24550 21508 24556
rect 21364 24132 21416 24138
rect 21364 24074 21416 24080
rect 21272 24064 21324 24070
rect 21272 24006 21324 24012
rect 21284 23662 21312 24006
rect 21180 23656 21232 23662
rect 21180 23598 21232 23604
rect 21272 23656 21324 23662
rect 21272 23598 21324 23604
rect 19984 23044 20036 23050
rect 19984 22986 20036 22992
rect 20996 23044 21048 23050
rect 20996 22986 21048 22992
rect 19800 22568 19852 22574
rect 19800 22510 19852 22516
rect 19812 21690 19840 22510
rect 19800 21684 19852 21690
rect 19800 21626 19852 21632
rect 19524 21548 19576 21554
rect 19524 21490 19576 21496
rect 19432 19916 19484 19922
rect 19432 19858 19484 19864
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19444 16794 19472 19722
rect 19432 16788 19484 16794
rect 19432 16730 19484 16736
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 18788 2916 18840 2922
rect 18788 2858 18840 2864
rect 18696 2644 18748 2650
rect 18696 2586 18748 2592
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 17950 2204 18258 2213
rect 17950 2202 17956 2204
rect 18012 2202 18036 2204
rect 18092 2202 18116 2204
rect 18172 2202 18196 2204
rect 18252 2202 18258 2204
rect 18012 2150 18014 2202
rect 18194 2150 18196 2202
rect 17950 2148 17956 2150
rect 18012 2148 18036 2150
rect 18092 2148 18116 2150
rect 18172 2148 18196 2150
rect 18252 2148 18258 2150
rect 17950 2139 18258 2148
rect 18432 800 18460 2450
rect 19168 800 19196 2926
rect 19536 1834 19564 21490
rect 19996 21486 20024 22986
rect 20168 22092 20220 22098
rect 20168 22034 20220 22040
rect 19892 21480 19944 21486
rect 19892 21422 19944 21428
rect 19984 21480 20036 21486
rect 19984 21422 20036 21428
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 19812 18426 19840 20198
rect 19904 18970 19932 21422
rect 20180 19786 20208 22034
rect 21008 22030 21036 22986
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 19800 18420 19852 18426
rect 19800 18362 19852 18368
rect 20076 18216 20128 18222
rect 20076 18158 20128 18164
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 19812 17542 19840 18022
rect 19892 17808 19944 17814
rect 19944 17756 20024 17762
rect 19892 17750 20024 17756
rect 19904 17734 20024 17750
rect 19996 17542 20024 17734
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19892 17536 19944 17542
rect 19892 17478 19944 17484
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19904 17082 19932 17478
rect 20088 17134 20116 18158
rect 20076 17128 20128 17134
rect 19904 17054 20024 17082
rect 20076 17070 20128 17076
rect 19996 16998 20024 17054
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 20088 16794 20116 17070
rect 19708 16788 19760 16794
rect 19708 16730 19760 16736
rect 20076 16788 20128 16794
rect 20076 16730 20128 16736
rect 19720 11218 19748 16730
rect 20548 15502 20576 18634
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20640 18426 20668 18566
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20720 17264 20772 17270
rect 20720 17206 20772 17212
rect 20732 17134 20760 17206
rect 20720 17128 20772 17134
rect 20720 17070 20772 17076
rect 20732 16454 20760 17070
rect 20720 16448 20772 16454
rect 20720 16390 20772 16396
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 19708 11212 19760 11218
rect 19708 11154 19760 11160
rect 19904 6914 19932 15438
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14618 20484 14758
rect 20444 14612 20496 14618
rect 20444 14554 20496 14560
rect 20824 12434 20852 20402
rect 21008 19854 21036 21966
rect 21192 21690 21220 23598
rect 21272 22976 21324 22982
rect 21272 22918 21324 22924
rect 21284 22574 21312 22918
rect 21272 22568 21324 22574
rect 21272 22510 21324 22516
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20996 18216 21048 18222
rect 20996 18158 21048 18164
rect 21008 17678 21036 18158
rect 20996 17672 21048 17678
rect 20996 17614 21048 17620
rect 21100 17490 21128 21490
rect 21376 21486 21404 24074
rect 21468 23798 21496 24550
rect 21456 23792 21508 23798
rect 21456 23734 21508 23740
rect 21640 22432 21692 22438
rect 21640 22374 21692 22380
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21376 20534 21404 21422
rect 21652 20602 21680 22374
rect 21744 21622 21772 24618
rect 22020 24290 22048 28018
rect 22112 25838 22140 29174
rect 22204 28694 22232 34682
rect 22296 34048 22324 41386
rect 22480 41274 22508 41482
rect 22468 41268 22520 41274
rect 22468 41210 22520 41216
rect 22376 41132 22428 41138
rect 22376 41074 22428 41080
rect 22388 39302 22416 41074
rect 22572 40934 22600 41670
rect 22744 41064 22796 41070
rect 22744 41006 22796 41012
rect 22560 40928 22612 40934
rect 22560 40870 22612 40876
rect 22756 40526 22784 41006
rect 22836 40928 22888 40934
rect 22836 40870 22888 40876
rect 22744 40520 22796 40526
rect 22744 40462 22796 40468
rect 22468 39840 22520 39846
rect 22468 39782 22520 39788
rect 22480 39506 22508 39782
rect 22468 39500 22520 39506
rect 22468 39442 22520 39448
rect 22376 39296 22428 39302
rect 22376 39238 22428 39244
rect 22388 39001 22416 39238
rect 22374 38992 22430 39001
rect 22374 38927 22430 38936
rect 22468 37664 22520 37670
rect 22468 37606 22520 37612
rect 22480 37262 22508 37606
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22560 36712 22612 36718
rect 22560 36654 22612 36660
rect 22572 35154 22600 36654
rect 22756 36242 22784 40462
rect 22848 39030 22876 40870
rect 22950 40828 23258 40837
rect 22950 40826 22956 40828
rect 23012 40826 23036 40828
rect 23092 40826 23116 40828
rect 23172 40826 23196 40828
rect 23252 40826 23258 40828
rect 23012 40774 23014 40826
rect 23194 40774 23196 40826
rect 22950 40772 22956 40774
rect 23012 40772 23036 40774
rect 23092 40772 23116 40774
rect 23172 40772 23196 40774
rect 23252 40772 23258 40774
rect 22950 40763 23258 40772
rect 22950 39740 23258 39749
rect 22950 39738 22956 39740
rect 23012 39738 23036 39740
rect 23092 39738 23116 39740
rect 23172 39738 23196 39740
rect 23252 39738 23258 39740
rect 23012 39686 23014 39738
rect 23194 39686 23196 39738
rect 22950 39684 22956 39686
rect 23012 39684 23036 39686
rect 23092 39684 23116 39686
rect 23172 39684 23196 39686
rect 23252 39684 23258 39686
rect 22950 39675 23258 39684
rect 22836 39024 22888 39030
rect 22836 38966 22888 38972
rect 22950 38652 23258 38661
rect 22950 38650 22956 38652
rect 23012 38650 23036 38652
rect 23092 38650 23116 38652
rect 23172 38650 23196 38652
rect 23252 38650 23258 38652
rect 23012 38598 23014 38650
rect 23194 38598 23196 38650
rect 22950 38596 22956 38598
rect 23012 38596 23036 38598
rect 23092 38596 23116 38598
rect 23172 38596 23196 38598
rect 23252 38596 23258 38598
rect 22950 38587 23258 38596
rect 23308 38554 23336 43726
rect 24216 43648 24268 43654
rect 24216 43590 24268 43596
rect 24032 43172 24084 43178
rect 24032 43114 24084 43120
rect 23756 42084 23808 42090
rect 23756 42026 23808 42032
rect 23768 41614 23796 42026
rect 23756 41608 23808 41614
rect 23756 41550 23808 41556
rect 23388 40452 23440 40458
rect 23388 40394 23440 40400
rect 23296 38548 23348 38554
rect 23296 38490 23348 38496
rect 22950 37564 23258 37573
rect 22950 37562 22956 37564
rect 23012 37562 23036 37564
rect 23092 37562 23116 37564
rect 23172 37562 23196 37564
rect 23252 37562 23258 37564
rect 23012 37510 23014 37562
rect 23194 37510 23196 37562
rect 22950 37508 22956 37510
rect 23012 37508 23036 37510
rect 23092 37508 23116 37510
rect 23172 37508 23196 37510
rect 23252 37508 23258 37510
rect 22950 37499 23258 37508
rect 23400 37126 23428 40394
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 23584 39302 23612 39918
rect 23572 39296 23624 39302
rect 23572 39238 23624 39244
rect 23584 37330 23612 39238
rect 23848 38412 23900 38418
rect 23848 38354 23900 38360
rect 23664 38208 23716 38214
rect 23664 38150 23716 38156
rect 23572 37324 23624 37330
rect 23572 37266 23624 37272
rect 23388 37120 23440 37126
rect 23388 37062 23440 37068
rect 22836 36576 22888 36582
rect 22836 36518 22888 36524
rect 22652 36236 22704 36242
rect 22652 36178 22704 36184
rect 22744 36236 22796 36242
rect 22744 36178 22796 36184
rect 22664 36038 22692 36178
rect 22848 36174 22876 36518
rect 22950 36476 23258 36485
rect 22950 36474 22956 36476
rect 23012 36474 23036 36476
rect 23092 36474 23116 36476
rect 23172 36474 23196 36476
rect 23252 36474 23258 36476
rect 23012 36422 23014 36474
rect 23194 36422 23196 36474
rect 22950 36420 22956 36422
rect 23012 36420 23036 36422
rect 23092 36420 23116 36422
rect 23172 36420 23196 36422
rect 23252 36420 23258 36422
rect 22950 36411 23258 36420
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22572 34542 22600 35090
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 22376 34060 22428 34066
rect 22296 34020 22376 34048
rect 22376 34002 22428 34008
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22192 28688 22244 28694
rect 22192 28630 22244 28636
rect 22296 28626 22324 32846
rect 22572 32230 22600 34478
rect 22560 32224 22612 32230
rect 22560 32166 22612 32172
rect 22572 32026 22600 32166
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22468 31272 22520 31278
rect 22466 31240 22468 31249
rect 22520 31240 22522 31249
rect 22466 31175 22522 31184
rect 22572 29714 22600 31962
rect 22664 29782 22692 35974
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 22950 35388 23258 35397
rect 22950 35386 22956 35388
rect 23012 35386 23036 35388
rect 23092 35386 23116 35388
rect 23172 35386 23196 35388
rect 23252 35386 23258 35388
rect 23012 35334 23014 35386
rect 23194 35334 23196 35386
rect 22950 35332 22956 35334
rect 23012 35332 23036 35334
rect 23092 35332 23116 35334
rect 23172 35332 23196 35334
rect 23252 35332 23258 35334
rect 22950 35323 23258 35332
rect 23308 35018 23336 35634
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 23400 35154 23428 35430
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 22950 34300 23258 34309
rect 22950 34298 22956 34300
rect 23012 34298 23036 34300
rect 23092 34298 23116 34300
rect 23172 34298 23196 34300
rect 23252 34298 23258 34300
rect 23012 34246 23014 34298
rect 23194 34246 23196 34298
rect 22950 34244 22956 34246
rect 23012 34244 23036 34246
rect 23092 34244 23116 34246
rect 23172 34244 23196 34246
rect 23252 34244 23258 34246
rect 22950 34235 23258 34244
rect 23308 33998 23336 34954
rect 23400 34134 23428 35090
rect 23388 34128 23440 34134
rect 23388 34070 23440 34076
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 23296 33992 23348 33998
rect 23296 33934 23348 33940
rect 22848 32842 22876 33934
rect 23480 33924 23532 33930
rect 23480 33866 23532 33872
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 22950 33212 23258 33221
rect 22950 33210 22956 33212
rect 23012 33210 23036 33212
rect 23092 33210 23116 33212
rect 23172 33210 23196 33212
rect 23252 33210 23258 33212
rect 23012 33158 23014 33210
rect 23194 33158 23196 33210
rect 22950 33156 22956 33158
rect 23012 33156 23036 33158
rect 23092 33156 23116 33158
rect 23172 33156 23196 33158
rect 23252 33156 23258 33158
rect 22950 33147 23258 33156
rect 22836 32836 22888 32842
rect 22836 32778 22888 32784
rect 22848 32502 22876 32778
rect 22836 32496 22888 32502
rect 22836 32438 22888 32444
rect 22848 31754 22876 32438
rect 22950 32124 23258 32133
rect 22950 32122 22956 32124
rect 23012 32122 23036 32124
rect 23092 32122 23116 32124
rect 23172 32122 23196 32124
rect 23252 32122 23258 32124
rect 23012 32070 23014 32122
rect 23194 32070 23196 32122
rect 22950 32068 22956 32070
rect 23012 32068 23036 32070
rect 23092 32068 23116 32070
rect 23172 32068 23196 32070
rect 23252 32068 23258 32070
rect 22950 32059 23258 32068
rect 22836 31748 22888 31754
rect 22836 31690 22888 31696
rect 22836 31272 22888 31278
rect 22836 31214 22888 31220
rect 22652 29776 22704 29782
rect 22652 29718 22704 29724
rect 22560 29708 22612 29714
rect 22560 29650 22612 29656
rect 22468 29572 22520 29578
rect 22468 29514 22520 29520
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22296 28082 22324 28562
rect 22376 28552 22428 28558
rect 22376 28494 22428 28500
rect 22388 28422 22416 28494
rect 22480 28490 22508 29514
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22468 28484 22520 28490
rect 22468 28426 22520 28432
rect 22376 28416 22428 28422
rect 22572 28370 22600 28494
rect 22376 28358 22428 28364
rect 22480 28342 22600 28370
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22100 25832 22152 25838
rect 22100 25774 22152 25780
rect 22376 25832 22428 25838
rect 22376 25774 22428 25780
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 21836 24274 22048 24290
rect 21824 24268 22048 24274
rect 21876 24262 22048 24268
rect 21824 24210 21876 24216
rect 22020 23730 22048 24262
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22100 23520 22152 23526
rect 22100 23462 22152 23468
rect 21916 22704 21968 22710
rect 21916 22646 21968 22652
rect 21732 21616 21784 21622
rect 21732 21558 21784 21564
rect 21640 20596 21692 20602
rect 21640 20538 21692 20544
rect 21824 20596 21876 20602
rect 21824 20538 21876 20544
rect 21364 20528 21416 20534
rect 21364 20470 21416 20476
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21548 19984 21600 19990
rect 21548 19926 21600 19932
rect 21180 19440 21232 19446
rect 21180 19382 21232 19388
rect 21192 18902 21220 19382
rect 21560 19310 21588 19926
rect 21548 19304 21600 19310
rect 21548 19246 21600 19252
rect 21180 18896 21232 18902
rect 21180 18838 21232 18844
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 21468 18358 21496 18634
rect 21560 18358 21588 19246
rect 21456 18352 21508 18358
rect 21456 18294 21508 18300
rect 21548 18352 21600 18358
rect 21548 18294 21600 18300
rect 21272 17740 21324 17746
rect 21272 17682 21324 17688
rect 21364 17740 21416 17746
rect 21364 17682 21416 17688
rect 20732 12406 20852 12434
rect 21008 17462 21128 17490
rect 21008 12434 21036 17462
rect 21284 17338 21312 17682
rect 21376 17610 21404 17682
rect 21364 17604 21416 17610
rect 21364 17546 21416 17552
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21744 17134 21772 20334
rect 21836 19922 21864 20538
rect 21824 19916 21876 19922
rect 21824 19858 21876 19864
rect 21836 18834 21864 19858
rect 21928 19174 21956 22646
rect 22112 21894 22140 23462
rect 22192 23316 22244 23322
rect 22192 23258 22244 23264
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 22112 18970 22140 21558
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 21824 18828 21876 18834
rect 21824 18770 21876 18776
rect 22112 18630 22140 18906
rect 22100 18624 22152 18630
rect 22100 18566 22152 18572
rect 22100 18284 22152 18290
rect 22100 18226 22152 18232
rect 21916 18148 21968 18154
rect 21916 18090 21968 18096
rect 21928 17882 21956 18090
rect 21916 17876 21968 17882
rect 21916 17818 21968 17824
rect 22008 17876 22060 17882
rect 22008 17818 22060 17824
rect 22020 17542 22048 17818
rect 22008 17536 22060 17542
rect 22008 17478 22060 17484
rect 22112 17338 22140 18226
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 21732 17128 21784 17134
rect 21732 17070 21784 17076
rect 21916 17128 21968 17134
rect 21916 17070 21968 17076
rect 21928 16522 21956 17070
rect 22008 16992 22060 16998
rect 22008 16934 22060 16940
rect 21916 16516 21968 16522
rect 21916 16458 21968 16464
rect 21180 16448 21232 16454
rect 22020 16436 22048 16934
rect 22100 16448 22152 16454
rect 22020 16408 22100 16436
rect 21180 16390 21232 16396
rect 22100 16390 22152 16396
rect 21192 14958 21220 16390
rect 21180 14952 21232 14958
rect 21180 14894 21232 14900
rect 22204 12434 22232 23258
rect 22296 22778 22324 25094
rect 22284 22772 22336 22778
rect 22284 22714 22336 22720
rect 22388 22094 22416 25774
rect 22480 23633 22508 28342
rect 22664 25786 22692 29718
rect 22848 29306 22876 31214
rect 22950 31036 23258 31045
rect 22950 31034 22956 31036
rect 23012 31034 23036 31036
rect 23092 31034 23116 31036
rect 23172 31034 23196 31036
rect 23252 31034 23258 31036
rect 23012 30982 23014 31034
rect 23194 30982 23196 31034
rect 22950 30980 22956 30982
rect 23012 30980 23036 30982
rect 23092 30980 23116 30982
rect 23172 30980 23196 30982
rect 23252 30980 23258 30982
rect 22950 30971 23258 30980
rect 23400 30938 23428 33798
rect 23492 31482 23520 33866
rect 23676 33658 23704 38150
rect 23756 37324 23808 37330
rect 23756 37266 23808 37272
rect 23768 36922 23796 37266
rect 23756 36916 23808 36922
rect 23756 36858 23808 36864
rect 23860 35834 23888 38354
rect 23940 37324 23992 37330
rect 23940 37266 23992 37272
rect 23848 35828 23900 35834
rect 23848 35770 23900 35776
rect 23860 34542 23888 35770
rect 23952 35630 23980 37266
rect 23940 35624 23992 35630
rect 23940 35566 23992 35572
rect 23952 35222 23980 35566
rect 23940 35216 23992 35222
rect 23940 35158 23992 35164
rect 23848 34536 23900 34542
rect 23848 34478 23900 34484
rect 23940 34060 23992 34066
rect 23940 34002 23992 34008
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23664 33652 23716 33658
rect 23664 33594 23716 33600
rect 23768 33046 23796 33798
rect 23756 33040 23808 33046
rect 23756 32982 23808 32988
rect 23860 32910 23888 33934
rect 23952 32978 23980 34002
rect 23940 32972 23992 32978
rect 23940 32914 23992 32920
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23952 32026 23980 32914
rect 24044 32774 24072 43114
rect 24124 42696 24176 42702
rect 24124 42638 24176 42644
rect 24136 42158 24164 42638
rect 24124 42152 24176 42158
rect 24124 42094 24176 42100
rect 24136 41682 24164 42094
rect 24124 41676 24176 41682
rect 24124 41618 24176 41624
rect 24136 41138 24164 41618
rect 24124 41132 24176 41138
rect 24124 41074 24176 41080
rect 24228 38654 24256 43590
rect 24400 43444 24452 43450
rect 24400 43386 24452 43392
rect 24308 42288 24360 42294
rect 24308 42230 24360 42236
rect 24320 40526 24348 42230
rect 24308 40520 24360 40526
rect 24308 40462 24360 40468
rect 24228 38626 24348 38654
rect 24216 35216 24268 35222
rect 24216 35158 24268 35164
rect 24228 33454 24256 35158
rect 24216 33448 24268 33454
rect 24216 33390 24268 33396
rect 24320 32978 24348 38626
rect 24412 35329 24440 43386
rect 24504 39098 24532 44814
rect 24872 43450 24900 47602
rect 24860 43444 24912 43450
rect 24860 43386 24912 43392
rect 24860 42288 24912 42294
rect 24860 42230 24912 42236
rect 24872 41274 24900 42230
rect 24964 41414 24992 53450
rect 24964 41386 25452 41414
rect 24860 41268 24912 41274
rect 24860 41210 24912 41216
rect 24584 41132 24636 41138
rect 24584 41074 24636 41080
rect 24596 39506 24624 41074
rect 24872 40118 24900 41210
rect 25044 41064 25096 41070
rect 25044 41006 25096 41012
rect 25056 40594 25084 41006
rect 25044 40588 25096 40594
rect 25044 40530 25096 40536
rect 25056 40186 25084 40530
rect 25044 40180 25096 40186
rect 25044 40122 25096 40128
rect 24860 40112 24912 40118
rect 24860 40054 24912 40060
rect 24676 39908 24728 39914
rect 24676 39850 24728 39856
rect 24584 39500 24636 39506
rect 24584 39442 24636 39448
rect 24492 39092 24544 39098
rect 24492 39034 24544 39040
rect 24584 39092 24636 39098
rect 24584 39034 24636 39040
rect 24596 38894 24624 39034
rect 24688 39030 24716 39850
rect 24872 39370 24900 40054
rect 25228 39500 25280 39506
rect 25228 39442 25280 39448
rect 24860 39364 24912 39370
rect 24860 39306 24912 39312
rect 25044 39092 25096 39098
rect 25044 39034 25096 39040
rect 24676 39024 24728 39030
rect 24676 38966 24728 38972
rect 24860 39024 24912 39030
rect 24860 38966 24912 38972
rect 24584 38888 24636 38894
rect 24584 38830 24636 38836
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24688 37942 24716 38218
rect 24676 37936 24728 37942
rect 24676 37878 24728 37884
rect 24688 36854 24716 37878
rect 24676 36848 24728 36854
rect 24676 36790 24728 36796
rect 24688 35562 24716 36790
rect 24676 35556 24728 35562
rect 24676 35498 24728 35504
rect 24398 35320 24454 35329
rect 24398 35255 24454 35264
rect 24584 34944 24636 34950
rect 24584 34886 24636 34892
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24214 32872 24270 32881
rect 24214 32807 24270 32816
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 24228 32366 24256 32807
rect 24492 32768 24544 32774
rect 24492 32710 24544 32716
rect 24216 32360 24268 32366
rect 24216 32302 24268 32308
rect 23940 32020 23992 32026
rect 23940 31962 23992 31968
rect 23848 31884 23900 31890
rect 23848 31826 23900 31832
rect 23480 31476 23532 31482
rect 23480 31418 23532 31424
rect 23388 30932 23440 30938
rect 23388 30874 23440 30880
rect 23860 30802 23888 31826
rect 24228 31278 24256 32302
rect 24216 31272 24268 31278
rect 24216 31214 24268 31220
rect 23848 30796 23900 30802
rect 23848 30738 23900 30744
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23296 30660 23348 30666
rect 23296 30602 23348 30608
rect 22950 29948 23258 29957
rect 22950 29946 22956 29948
rect 23012 29946 23036 29948
rect 23092 29946 23116 29948
rect 23172 29946 23196 29948
rect 23252 29946 23258 29948
rect 23012 29894 23014 29946
rect 23194 29894 23196 29946
rect 22950 29892 22956 29894
rect 23012 29892 23036 29894
rect 23092 29892 23116 29894
rect 23172 29892 23196 29894
rect 23252 29892 23258 29894
rect 22950 29883 23258 29892
rect 22836 29300 22888 29306
rect 22836 29242 22888 29248
rect 22950 28860 23258 28869
rect 22950 28858 22956 28860
rect 23012 28858 23036 28860
rect 23092 28858 23116 28860
rect 23172 28858 23196 28860
rect 23252 28858 23258 28860
rect 23012 28806 23014 28858
rect 23194 28806 23196 28858
rect 22950 28804 22956 28806
rect 23012 28804 23036 28806
rect 23092 28804 23116 28806
rect 23172 28804 23196 28806
rect 23252 28804 23258 28806
rect 22950 28795 23258 28804
rect 23308 28762 23336 30602
rect 23296 28756 23348 28762
rect 23296 28698 23348 28704
rect 23204 28688 23256 28694
rect 23204 28630 23256 28636
rect 23216 28490 23244 28630
rect 23400 28626 23428 30670
rect 23572 30592 23624 30598
rect 23572 30534 23624 30540
rect 23584 30258 23612 30534
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23388 28620 23440 28626
rect 23388 28562 23440 28568
rect 23204 28484 23256 28490
rect 23204 28426 23256 28432
rect 23296 28416 23348 28422
rect 23296 28358 23348 28364
rect 22950 27772 23258 27781
rect 22950 27770 22956 27772
rect 23012 27770 23036 27772
rect 23092 27770 23116 27772
rect 23172 27770 23196 27772
rect 23252 27770 23258 27772
rect 23012 27718 23014 27770
rect 23194 27718 23196 27770
rect 22950 27716 22956 27718
rect 23012 27716 23036 27718
rect 23092 27716 23116 27718
rect 23172 27716 23196 27718
rect 23252 27716 23258 27718
rect 22950 27707 23258 27716
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23124 27130 23152 27406
rect 23308 27130 23336 28358
rect 23388 28212 23440 28218
rect 23388 28154 23440 28160
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23296 27124 23348 27130
rect 23296 27066 23348 27072
rect 23400 26926 23428 28154
rect 23756 28076 23808 28082
rect 23756 28018 23808 28024
rect 23768 27334 23796 28018
rect 24400 27872 24452 27878
rect 24400 27814 24452 27820
rect 23480 27328 23532 27334
rect 23480 27270 23532 27276
rect 23756 27328 23808 27334
rect 23756 27270 23808 27276
rect 23388 26920 23440 26926
rect 23388 26862 23440 26868
rect 22950 26684 23258 26693
rect 22950 26682 22956 26684
rect 23012 26682 23036 26684
rect 23092 26682 23116 26684
rect 23172 26682 23196 26684
rect 23252 26682 23258 26684
rect 23012 26630 23014 26682
rect 23194 26630 23196 26682
rect 22950 26628 22956 26630
rect 23012 26628 23036 26630
rect 23092 26628 23116 26630
rect 23172 26628 23196 26630
rect 23252 26628 23258 26630
rect 22950 26619 23258 26628
rect 23492 26382 23520 27270
rect 24124 26784 24176 26790
rect 24124 26726 24176 26732
rect 24216 26784 24268 26790
rect 24216 26726 24268 26732
rect 23572 26512 23624 26518
rect 23572 26454 23624 26460
rect 23940 26512 23992 26518
rect 23940 26454 23992 26460
rect 23480 26376 23532 26382
rect 23480 26318 23532 26324
rect 23584 26330 23612 26454
rect 22664 25758 22784 25786
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22664 25294 22692 25638
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22560 24064 22612 24070
rect 22560 24006 22612 24012
rect 22466 23624 22522 23633
rect 22466 23559 22522 23568
rect 22572 22166 22600 24006
rect 22756 23322 22784 25758
rect 22950 25596 23258 25605
rect 22950 25594 22956 25596
rect 23012 25594 23036 25596
rect 23092 25594 23116 25596
rect 23172 25594 23196 25596
rect 23252 25594 23258 25596
rect 23012 25542 23014 25594
rect 23194 25542 23196 25594
rect 22950 25540 22956 25542
rect 23012 25540 23036 25542
rect 23092 25540 23116 25542
rect 23172 25540 23196 25542
rect 23252 25540 23258 25542
rect 22950 25531 23258 25540
rect 23296 25152 23348 25158
rect 23296 25094 23348 25100
rect 22950 24508 23258 24517
rect 22950 24506 22956 24508
rect 23012 24506 23036 24508
rect 23092 24506 23116 24508
rect 23172 24506 23196 24508
rect 23252 24506 23258 24508
rect 23012 24454 23014 24506
rect 23194 24454 23196 24506
rect 22950 24452 22956 24454
rect 23012 24452 23036 24454
rect 23092 24452 23116 24454
rect 23172 24452 23196 24454
rect 23252 24452 23258 24454
rect 22950 24443 23258 24452
rect 22836 24268 22888 24274
rect 22836 24210 22888 24216
rect 22744 23316 22796 23322
rect 22744 23258 22796 23264
rect 22652 22976 22704 22982
rect 22652 22918 22704 22924
rect 22560 22160 22612 22166
rect 22560 22102 22612 22108
rect 22296 22066 22416 22094
rect 22296 20466 22324 22066
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22480 21690 22508 21830
rect 22468 21684 22520 21690
rect 22468 21626 22520 21632
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22284 20460 22336 20466
rect 22284 20402 22336 20408
rect 22388 19514 22416 21490
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22480 20602 22508 21422
rect 22468 20596 22520 20602
rect 22468 20538 22520 20544
rect 22558 20496 22614 20505
rect 22558 20431 22614 20440
rect 22468 19916 22520 19922
rect 22468 19858 22520 19864
rect 22480 19530 22508 19858
rect 22572 19786 22600 20431
rect 22560 19780 22612 19786
rect 22560 19722 22612 19728
rect 22376 19508 22428 19514
rect 22480 19502 22600 19530
rect 22376 19450 22428 19456
rect 22468 19372 22520 19378
rect 22468 19314 22520 19320
rect 22480 18970 22508 19314
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22284 18692 22336 18698
rect 22284 18634 22336 18640
rect 22296 18290 22324 18634
rect 22284 18284 22336 18290
rect 22284 18226 22336 18232
rect 22388 17814 22416 18906
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 17882 22508 18702
rect 22572 18154 22600 19502
rect 22560 18148 22612 18154
rect 22560 18090 22612 18096
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22376 17808 22428 17814
rect 22376 17750 22428 17756
rect 22664 17746 22692 22918
rect 22848 21622 22876 24210
rect 23308 23866 23336 25094
rect 23492 24138 23520 26318
rect 23584 26314 23704 26330
rect 23584 26308 23716 26314
rect 23584 26302 23664 26308
rect 23480 24132 23532 24138
rect 23480 24074 23532 24080
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23492 23662 23520 24074
rect 23480 23656 23532 23662
rect 23386 23624 23442 23633
rect 23480 23598 23532 23604
rect 23386 23559 23388 23568
rect 23440 23559 23442 23568
rect 23388 23530 23440 23536
rect 23386 23488 23442 23497
rect 22950 23420 23258 23429
rect 23386 23423 23442 23432
rect 22950 23418 22956 23420
rect 23012 23418 23036 23420
rect 23092 23418 23116 23420
rect 23172 23418 23196 23420
rect 23252 23418 23258 23420
rect 23012 23366 23014 23418
rect 23194 23366 23196 23418
rect 22950 23364 22956 23366
rect 23012 23364 23036 23366
rect 23092 23364 23116 23366
rect 23172 23364 23196 23366
rect 23252 23364 23258 23366
rect 22950 23355 23258 23364
rect 23400 23118 23428 23423
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22950 22332 23258 22341
rect 22950 22330 22956 22332
rect 23012 22330 23036 22332
rect 23092 22330 23116 22332
rect 23172 22330 23196 22332
rect 23252 22330 23258 22332
rect 23012 22278 23014 22330
rect 23194 22278 23196 22330
rect 22950 22276 22956 22278
rect 23012 22276 23036 22278
rect 23092 22276 23116 22278
rect 23172 22276 23196 22278
rect 23252 22276 23258 22278
rect 22950 22267 23258 22276
rect 23308 22234 23336 22578
rect 23388 22432 23440 22438
rect 23388 22374 23440 22380
rect 23296 22228 23348 22234
rect 23296 22170 23348 22176
rect 23296 22092 23348 22098
rect 23296 22034 23348 22040
rect 23308 21622 23336 22034
rect 22836 21616 22888 21622
rect 22836 21558 22888 21564
rect 23296 21616 23348 21622
rect 23296 21558 23348 21564
rect 22950 21244 23258 21253
rect 22950 21242 22956 21244
rect 23012 21242 23036 21244
rect 23092 21242 23116 21244
rect 23172 21242 23196 21244
rect 23252 21242 23258 21244
rect 23012 21190 23014 21242
rect 23194 21190 23196 21242
rect 22950 21188 22956 21190
rect 23012 21188 23036 21190
rect 23092 21188 23116 21190
rect 23172 21188 23196 21190
rect 23252 21188 23258 21190
rect 22950 21179 23258 21188
rect 23308 20534 23336 21558
rect 23296 20528 23348 20534
rect 23294 20496 23296 20505
rect 23348 20496 23350 20505
rect 23294 20431 23350 20440
rect 23296 20392 23348 20398
rect 23296 20334 23348 20340
rect 22950 20156 23258 20165
rect 22950 20154 22956 20156
rect 23012 20154 23036 20156
rect 23092 20154 23116 20156
rect 23172 20154 23196 20156
rect 23252 20154 23258 20156
rect 23012 20102 23014 20154
rect 23194 20102 23196 20154
rect 22950 20100 22956 20102
rect 23012 20100 23036 20102
rect 23092 20100 23116 20102
rect 23172 20100 23196 20102
rect 23252 20100 23258 20102
rect 22950 20091 23258 20100
rect 23204 19984 23256 19990
rect 22848 19944 23204 19972
rect 22848 19938 22876 19944
rect 22756 19922 22876 19938
rect 23204 19926 23256 19932
rect 22744 19916 22876 19922
rect 22796 19910 22876 19916
rect 22744 19858 22796 19864
rect 23308 19310 23336 20334
rect 23296 19304 23348 19310
rect 23296 19246 23348 19252
rect 22744 19168 22796 19174
rect 22744 19110 22796 19116
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22756 18970 22784 19110
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22848 18873 22876 19110
rect 22950 19068 23258 19077
rect 22950 19066 22956 19068
rect 23012 19066 23036 19068
rect 23092 19066 23116 19068
rect 23172 19066 23196 19068
rect 23252 19066 23258 19068
rect 23012 19014 23014 19066
rect 23194 19014 23196 19066
rect 22950 19012 22956 19014
rect 23012 19012 23036 19014
rect 23092 19012 23116 19014
rect 23172 19012 23196 19014
rect 23252 19012 23258 19014
rect 22950 19003 23258 19012
rect 22834 18864 22890 18873
rect 22834 18799 22890 18808
rect 22950 17980 23258 17989
rect 22950 17978 22956 17980
rect 23012 17978 23036 17980
rect 23092 17978 23116 17980
rect 23172 17978 23196 17980
rect 23252 17978 23258 17980
rect 23012 17926 23014 17978
rect 23194 17926 23196 17978
rect 22950 17924 22956 17926
rect 23012 17924 23036 17926
rect 23092 17924 23116 17926
rect 23172 17924 23196 17926
rect 23252 17924 23258 17926
rect 22950 17915 23258 17924
rect 23308 17762 23336 19246
rect 23400 18630 23428 22374
rect 23492 22098 23520 23598
rect 23584 22166 23612 26302
rect 23664 26250 23716 26256
rect 23848 24064 23900 24070
rect 23848 24006 23900 24012
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23676 23186 23704 23598
rect 23664 23180 23716 23186
rect 23664 23122 23716 23128
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23676 22778 23704 22986
rect 23664 22772 23716 22778
rect 23664 22714 23716 22720
rect 23756 22704 23808 22710
rect 23756 22646 23808 22652
rect 23572 22160 23624 22166
rect 23572 22102 23624 22108
rect 23480 22092 23532 22098
rect 23480 22034 23532 22040
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23584 20058 23612 21830
rect 23572 20052 23624 20058
rect 23572 19994 23624 20000
rect 23480 19916 23532 19922
rect 23480 19858 23532 19864
rect 23492 18834 23520 19858
rect 23480 18828 23532 18834
rect 23480 18770 23532 18776
rect 23388 18624 23440 18630
rect 23388 18566 23440 18572
rect 22652 17740 22704 17746
rect 23308 17734 23428 17762
rect 22652 17682 22704 17688
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 22284 17604 22336 17610
rect 22284 17546 22336 17552
rect 22296 17270 22324 17546
rect 23308 17338 23336 17614
rect 23296 17332 23348 17338
rect 23296 17274 23348 17280
rect 22284 17264 22336 17270
rect 22284 17206 22336 17212
rect 22950 16892 23258 16901
rect 22950 16890 22956 16892
rect 23012 16890 23036 16892
rect 23092 16890 23116 16892
rect 23172 16890 23196 16892
rect 23252 16890 23258 16892
rect 23012 16838 23014 16890
rect 23194 16838 23196 16890
rect 22950 16836 22956 16838
rect 23012 16836 23036 16838
rect 23092 16836 23116 16838
rect 23172 16836 23196 16838
rect 23252 16836 23258 16838
rect 22950 16827 23258 16836
rect 22468 16652 22520 16658
rect 22468 16594 22520 16600
rect 22480 16114 22508 16594
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22480 15026 22508 16050
rect 22950 15804 23258 15813
rect 22950 15802 22956 15804
rect 23012 15802 23036 15804
rect 23092 15802 23116 15804
rect 23172 15802 23196 15804
rect 23252 15802 23258 15804
rect 23012 15750 23014 15802
rect 23194 15750 23196 15802
rect 22950 15748 22956 15750
rect 23012 15748 23036 15750
rect 23092 15748 23116 15750
rect 23172 15748 23196 15750
rect 23252 15748 23258 15750
rect 22950 15739 23258 15748
rect 23400 15570 23428 17734
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 22652 15360 22704 15366
rect 22652 15302 22704 15308
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 21008 12406 21220 12434
rect 22204 12406 22324 12434
rect 19904 6886 20024 6914
rect 19996 3194 20024 6886
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19524 1828 19576 1834
rect 19524 1770 19576 1776
rect 19904 800 19932 2382
rect 20640 800 20668 2926
rect 20732 1698 20760 12406
rect 21192 6914 21220 12406
rect 21100 6886 21220 6914
rect 21100 2417 21128 6886
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21364 2508 21416 2514
rect 21364 2450 21416 2456
rect 21086 2408 21142 2417
rect 21086 2343 21142 2352
rect 20720 1692 20772 1698
rect 20720 1634 20772 1640
rect 21376 800 21404 2450
rect 22112 800 22140 2926
rect 22296 1766 22324 12406
rect 22664 2446 22692 15302
rect 22950 14716 23258 14725
rect 22950 14714 22956 14716
rect 23012 14714 23036 14716
rect 23092 14714 23116 14716
rect 23172 14714 23196 14716
rect 23252 14714 23258 14716
rect 23012 14662 23014 14714
rect 23194 14662 23196 14714
rect 22950 14660 22956 14662
rect 23012 14660 23036 14662
rect 23092 14660 23116 14662
rect 23172 14660 23196 14662
rect 23252 14660 23258 14662
rect 22950 14651 23258 14660
rect 22950 13628 23258 13637
rect 22950 13626 22956 13628
rect 23012 13626 23036 13628
rect 23092 13626 23116 13628
rect 23172 13626 23196 13628
rect 23252 13626 23258 13628
rect 23012 13574 23014 13626
rect 23194 13574 23196 13626
rect 22950 13572 22956 13574
rect 23012 13572 23036 13574
rect 23092 13572 23116 13574
rect 23172 13572 23196 13574
rect 23252 13572 23258 13574
rect 22950 13563 23258 13572
rect 22950 12540 23258 12549
rect 22950 12538 22956 12540
rect 23012 12538 23036 12540
rect 23092 12538 23116 12540
rect 23172 12538 23196 12540
rect 23252 12538 23258 12540
rect 23012 12486 23014 12538
rect 23194 12486 23196 12538
rect 22950 12484 22956 12486
rect 23012 12484 23036 12486
rect 23092 12484 23116 12486
rect 23172 12484 23196 12486
rect 23252 12484 23258 12486
rect 22950 12475 23258 12484
rect 22950 11452 23258 11461
rect 22950 11450 22956 11452
rect 23012 11450 23036 11452
rect 23092 11450 23116 11452
rect 23172 11450 23196 11452
rect 23252 11450 23258 11452
rect 23012 11398 23014 11450
rect 23194 11398 23196 11450
rect 22950 11396 22956 11398
rect 23012 11396 23036 11398
rect 23092 11396 23116 11398
rect 23172 11396 23196 11398
rect 23252 11396 23258 11398
rect 22950 11387 23258 11396
rect 22950 10364 23258 10373
rect 22950 10362 22956 10364
rect 23012 10362 23036 10364
rect 23092 10362 23116 10364
rect 23172 10362 23196 10364
rect 23252 10362 23258 10364
rect 23012 10310 23014 10362
rect 23194 10310 23196 10362
rect 22950 10308 22956 10310
rect 23012 10308 23036 10310
rect 23092 10308 23116 10310
rect 23172 10308 23196 10310
rect 23252 10308 23258 10310
rect 22950 10299 23258 10308
rect 22950 9276 23258 9285
rect 22950 9274 22956 9276
rect 23012 9274 23036 9276
rect 23092 9274 23116 9276
rect 23172 9274 23196 9276
rect 23252 9274 23258 9276
rect 23012 9222 23014 9274
rect 23194 9222 23196 9274
rect 22950 9220 22956 9222
rect 23012 9220 23036 9222
rect 23092 9220 23116 9222
rect 23172 9220 23196 9222
rect 23252 9220 23258 9222
rect 22950 9211 23258 9220
rect 23400 8430 23428 15506
rect 23388 8424 23440 8430
rect 23388 8366 23440 8372
rect 22950 8188 23258 8197
rect 22950 8186 22956 8188
rect 23012 8186 23036 8188
rect 23092 8186 23116 8188
rect 23172 8186 23196 8188
rect 23252 8186 23258 8188
rect 23012 8134 23014 8186
rect 23194 8134 23196 8186
rect 22950 8132 22956 8134
rect 23012 8132 23036 8134
rect 23092 8132 23116 8134
rect 23172 8132 23196 8134
rect 23252 8132 23258 8134
rect 22950 8123 23258 8132
rect 22950 7100 23258 7109
rect 22950 7098 22956 7100
rect 23012 7098 23036 7100
rect 23092 7098 23116 7100
rect 23172 7098 23196 7100
rect 23252 7098 23258 7100
rect 23012 7046 23014 7098
rect 23194 7046 23196 7098
rect 22950 7044 22956 7046
rect 23012 7044 23036 7046
rect 23092 7044 23116 7046
rect 23172 7044 23196 7046
rect 23252 7044 23258 7046
rect 22950 7035 23258 7044
rect 22950 6012 23258 6021
rect 22950 6010 22956 6012
rect 23012 6010 23036 6012
rect 23092 6010 23116 6012
rect 23172 6010 23196 6012
rect 23252 6010 23258 6012
rect 23012 5958 23014 6010
rect 23194 5958 23196 6010
rect 22950 5956 22956 5958
rect 23012 5956 23036 5958
rect 23092 5956 23116 5958
rect 23172 5956 23196 5958
rect 23252 5956 23258 5958
rect 22950 5947 23258 5956
rect 22950 4924 23258 4933
rect 22950 4922 22956 4924
rect 23012 4922 23036 4924
rect 23092 4922 23116 4924
rect 23172 4922 23196 4924
rect 23252 4922 23258 4924
rect 23012 4870 23014 4922
rect 23194 4870 23196 4922
rect 22950 4868 22956 4870
rect 23012 4868 23036 4870
rect 23092 4868 23116 4870
rect 23172 4868 23196 4870
rect 23252 4868 23258 4870
rect 22950 4859 23258 4868
rect 22950 3836 23258 3845
rect 22950 3834 22956 3836
rect 23012 3834 23036 3836
rect 23092 3834 23116 3836
rect 23172 3834 23196 3836
rect 23252 3834 23258 3836
rect 23012 3782 23014 3834
rect 23194 3782 23196 3834
rect 22950 3780 22956 3782
rect 23012 3780 23036 3782
rect 23092 3780 23116 3782
rect 23172 3780 23196 3782
rect 23252 3780 23258 3782
rect 22950 3771 23258 3780
rect 23572 2984 23624 2990
rect 23572 2926 23624 2932
rect 22950 2748 23258 2757
rect 22950 2746 22956 2748
rect 23012 2746 23036 2748
rect 23092 2746 23116 2748
rect 23172 2746 23196 2748
rect 23252 2746 23258 2748
rect 23012 2694 23014 2746
rect 23194 2694 23196 2746
rect 22950 2692 22956 2694
rect 23012 2692 23036 2694
rect 23092 2692 23116 2694
rect 23172 2692 23196 2694
rect 23252 2692 23258 2694
rect 22950 2683 23258 2692
rect 22836 2508 22888 2514
rect 22836 2450 22888 2456
rect 22652 2440 22704 2446
rect 22652 2382 22704 2388
rect 22284 1760 22336 1766
rect 22284 1702 22336 1708
rect 22848 800 22876 2450
rect 23584 800 23612 2926
rect 23768 2038 23796 22646
rect 23860 21962 23888 24006
rect 23848 21956 23900 21962
rect 23848 21898 23900 21904
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 23860 19514 23888 19790
rect 23952 19718 23980 26454
rect 24136 26042 24164 26726
rect 24124 26036 24176 26042
rect 24124 25978 24176 25984
rect 23940 19712 23992 19718
rect 23940 19654 23992 19660
rect 23848 19508 23900 19514
rect 23848 19450 23900 19456
rect 24228 17338 24256 26726
rect 24412 26586 24440 27814
rect 24400 26580 24452 26586
rect 24400 26522 24452 26528
rect 24412 25838 24440 26522
rect 24308 25832 24360 25838
rect 24308 25774 24360 25780
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 24320 25498 24348 25774
rect 24308 25492 24360 25498
rect 24308 25434 24360 25440
rect 24308 25356 24360 25362
rect 24308 25298 24360 25304
rect 24320 22098 24348 25298
rect 24308 22092 24360 22098
rect 24308 22034 24360 22040
rect 24320 21350 24348 22034
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24320 18834 24348 21286
rect 24504 19378 24532 32710
rect 24596 30122 24624 34886
rect 24688 34678 24716 35498
rect 24872 34746 24900 38966
rect 24952 38888 25004 38894
rect 24952 38830 25004 38836
rect 24964 37670 24992 38830
rect 25056 37670 25084 39034
rect 25240 38486 25268 39442
rect 25228 38480 25280 38486
rect 25228 38422 25280 38428
rect 24952 37664 25004 37670
rect 24952 37606 25004 37612
rect 25044 37664 25096 37670
rect 25044 37606 25096 37612
rect 24964 36718 24992 37606
rect 24952 36712 25004 36718
rect 24952 36654 25004 36660
rect 25056 35766 25084 37606
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 24860 34740 24912 34746
rect 24860 34682 24912 34688
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24952 34604 25004 34610
rect 24952 34546 25004 34552
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 24688 32366 24716 32438
rect 24676 32360 24728 32366
rect 24676 32302 24728 32308
rect 24860 32224 24912 32230
rect 24860 32166 24912 32172
rect 24768 31816 24820 31822
rect 24768 31758 24820 31764
rect 24780 31482 24808 31758
rect 24768 31476 24820 31482
rect 24768 31418 24820 31424
rect 24872 31346 24900 32166
rect 24860 31340 24912 31346
rect 24860 31282 24912 31288
rect 24964 31142 24992 34546
rect 25056 31414 25084 35702
rect 25136 34536 25188 34542
rect 25136 34478 25188 34484
rect 25148 34406 25176 34478
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 25044 31408 25096 31414
rect 25044 31350 25096 31356
rect 25148 31278 25176 34342
rect 25228 34060 25280 34066
rect 25228 34002 25280 34008
rect 25240 32570 25268 34002
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 25424 31482 25452 41386
rect 25504 38208 25556 38214
rect 25504 38150 25556 38156
rect 25516 37466 25544 38150
rect 25504 37460 25556 37466
rect 25504 37402 25556 37408
rect 25596 37120 25648 37126
rect 25596 37062 25648 37068
rect 25504 36576 25556 36582
rect 25504 36518 25556 36524
rect 25412 31476 25464 31482
rect 25412 31418 25464 31424
rect 25136 31272 25188 31278
rect 25136 31214 25188 31220
rect 24952 31136 25004 31142
rect 24952 31078 25004 31084
rect 24860 30728 24912 30734
rect 24860 30670 24912 30676
rect 24584 30116 24636 30122
rect 24584 30058 24636 30064
rect 24872 27878 24900 30670
rect 25044 30184 25096 30190
rect 25044 30126 25096 30132
rect 25056 29850 25084 30126
rect 25044 29844 25096 29850
rect 25044 29786 25096 29792
rect 25148 29102 25176 31214
rect 25136 29096 25188 29102
rect 25136 29038 25188 29044
rect 24952 28144 25004 28150
rect 24952 28086 25004 28092
rect 24860 27872 24912 27878
rect 24860 27814 24912 27820
rect 24872 27470 24900 27814
rect 24860 27464 24912 27470
rect 24860 27406 24912 27412
rect 24872 27062 24900 27406
rect 24964 27334 24992 28086
rect 25424 27962 25452 31418
rect 25056 27934 25452 27962
rect 24952 27328 25004 27334
rect 24952 27270 25004 27276
rect 24860 27056 24912 27062
rect 24860 26998 24912 27004
rect 24872 26450 24900 26998
rect 25056 26586 25084 27934
rect 25136 27396 25188 27402
rect 25136 27338 25188 27344
rect 25044 26580 25096 26586
rect 25044 26522 25096 26528
rect 25056 26450 25084 26522
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 25044 26444 25096 26450
rect 25044 26386 25096 26392
rect 25148 25498 25176 27338
rect 25516 26994 25544 36518
rect 25608 36009 25636 37062
rect 25594 36000 25650 36009
rect 25594 35935 25650 35944
rect 25596 30320 25648 30326
rect 25596 30262 25648 30268
rect 25504 26988 25556 26994
rect 25504 26930 25556 26936
rect 25228 26580 25280 26586
rect 25228 26522 25280 26528
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 24676 23656 24728 23662
rect 24676 23598 24728 23604
rect 24584 22976 24636 22982
rect 24584 22918 24636 22924
rect 24596 22778 24624 22918
rect 24584 22772 24636 22778
rect 24584 22714 24636 22720
rect 24688 22094 24716 23598
rect 24952 23520 25004 23526
rect 24952 23462 25004 23468
rect 24964 23118 24992 23462
rect 24952 23112 25004 23118
rect 24952 23054 25004 23060
rect 25044 22976 25096 22982
rect 25042 22944 25044 22953
rect 25096 22944 25098 22953
rect 25042 22879 25098 22888
rect 25136 22568 25188 22574
rect 25136 22510 25188 22516
rect 25044 22432 25096 22438
rect 25044 22374 25096 22380
rect 24596 22066 24716 22094
rect 24492 19372 24544 19378
rect 24492 19314 24544 19320
rect 24596 19242 24624 22066
rect 24676 20596 24728 20602
rect 24676 20538 24728 20544
rect 24688 19428 24716 20538
rect 24768 19440 24820 19446
rect 24688 19400 24768 19428
rect 24584 19236 24636 19242
rect 24584 19178 24636 19184
rect 24688 19122 24716 19400
rect 24768 19382 24820 19388
rect 24860 19304 24912 19310
rect 24596 19094 24716 19122
rect 24780 19252 24860 19258
rect 24780 19246 24912 19252
rect 24780 19230 24900 19246
rect 24308 18828 24360 18834
rect 24308 18770 24360 18776
rect 24596 18358 24624 19094
rect 24780 18970 24808 19230
rect 24768 18964 24820 18970
rect 24768 18906 24820 18912
rect 24860 18624 24912 18630
rect 24860 18566 24912 18572
rect 24952 18624 25004 18630
rect 24952 18566 25004 18572
rect 24872 18358 24900 18566
rect 24964 18426 24992 18566
rect 24952 18420 25004 18426
rect 24952 18362 25004 18368
rect 24584 18352 24636 18358
rect 24584 18294 24636 18300
rect 24860 18352 24912 18358
rect 24860 18294 24912 18300
rect 24596 17542 24624 18294
rect 25056 18290 25084 22374
rect 25148 20398 25176 22510
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19990 25176 20334
rect 25136 19984 25188 19990
rect 25136 19926 25188 19932
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24768 18080 24820 18086
rect 24768 18022 24820 18028
rect 24584 17536 24636 17542
rect 24584 17478 24636 17484
rect 24216 17332 24268 17338
rect 24216 17274 24268 17280
rect 24228 10742 24256 17274
rect 24596 16590 24624 17478
rect 24676 16788 24728 16794
rect 24676 16730 24728 16736
rect 24584 16584 24636 16590
rect 24584 16526 24636 16532
rect 24596 16182 24624 16526
rect 24584 16176 24636 16182
rect 24584 16118 24636 16124
rect 24596 15094 24624 16118
rect 24584 15088 24636 15094
rect 24584 15030 24636 15036
rect 24216 10736 24268 10742
rect 24216 10678 24268 10684
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23756 2032 23808 2038
rect 23756 1974 23808 1980
rect 24320 800 24348 3538
rect 24688 3058 24716 16730
rect 24780 16182 24808 18022
rect 25056 17270 25084 18226
rect 25044 17264 25096 17270
rect 25044 17206 25096 17212
rect 25056 17134 25084 17206
rect 25044 17128 25096 17134
rect 25044 17070 25096 17076
rect 25044 16652 25096 16658
rect 25044 16594 25096 16600
rect 24768 16176 24820 16182
rect 24768 16118 24820 16124
rect 24780 4622 24808 16118
rect 25056 15162 25084 16594
rect 25240 15434 25268 26522
rect 25412 26240 25464 26246
rect 25412 26182 25464 26188
rect 25424 25226 25452 26182
rect 25412 25220 25464 25226
rect 25412 25162 25464 25168
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25044 15156 25096 15162
rect 25044 15098 25096 15104
rect 25228 12640 25280 12646
rect 25228 12582 25280 12588
rect 25136 10532 25188 10538
rect 25136 10474 25188 10480
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 25148 3058 25176 10474
rect 24676 3052 24728 3058
rect 24676 2994 24728 3000
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 25044 2984 25096 2990
rect 25044 2926 25096 2932
rect 25056 800 25084 2926
rect 25240 2446 25268 12582
rect 25228 2440 25280 2446
rect 25228 2382 25280 2388
rect 25332 1630 25360 24686
rect 25424 13326 25452 25162
rect 25608 24750 25636 30262
rect 25700 29730 25728 53926
rect 26252 43790 26280 53926
rect 27068 53712 27120 53718
rect 27068 53654 27120 53660
rect 26700 51400 26752 51406
rect 26700 51342 26752 51348
rect 26712 46170 26740 51342
rect 26700 46164 26752 46170
rect 26700 46106 26752 46112
rect 26240 43784 26292 43790
rect 26240 43726 26292 43732
rect 25964 43308 26016 43314
rect 25964 43250 26016 43256
rect 25872 42628 25924 42634
rect 25872 42570 25924 42576
rect 25884 42362 25912 42570
rect 25872 42356 25924 42362
rect 25872 42298 25924 42304
rect 25884 42022 25912 42298
rect 25872 42016 25924 42022
rect 25872 41958 25924 41964
rect 25976 41426 26004 43250
rect 26332 43240 26384 43246
rect 26332 43182 26384 43188
rect 26148 42628 26200 42634
rect 26148 42570 26200 42576
rect 25884 41398 26004 41426
rect 26160 41414 26188 42570
rect 26344 41818 26372 43182
rect 26516 42016 26568 42022
rect 26516 41958 26568 41964
rect 26332 41812 26384 41818
rect 26332 41754 26384 41760
rect 26528 41682 26556 41958
rect 26516 41676 26568 41682
rect 26516 41618 26568 41624
rect 26424 41608 26476 41614
rect 26424 41550 26476 41556
rect 25884 39098 25912 41398
rect 26068 41386 26188 41414
rect 26068 41274 26096 41386
rect 26056 41268 26108 41274
rect 26056 41210 26108 41216
rect 26056 39840 26108 39846
rect 26056 39782 26108 39788
rect 25964 39636 26016 39642
rect 25964 39578 26016 39584
rect 25872 39092 25924 39098
rect 25872 39034 25924 39040
rect 25976 37126 26004 39578
rect 26068 39574 26096 39782
rect 26056 39568 26108 39574
rect 26056 39510 26108 39516
rect 26148 39432 26200 39438
rect 26148 39374 26200 39380
rect 26160 38962 26188 39374
rect 26148 38956 26200 38962
rect 26148 38898 26200 38904
rect 26240 38956 26292 38962
rect 26240 38898 26292 38904
rect 26056 38820 26108 38826
rect 26056 38762 26108 38768
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 25964 37120 26016 37126
rect 25964 37062 26016 37068
rect 25780 36712 25832 36718
rect 25780 36654 25832 36660
rect 25792 35737 25820 36654
rect 25884 36310 25912 37062
rect 25872 36304 25924 36310
rect 25872 36246 25924 36252
rect 25778 35728 25834 35737
rect 25778 35663 25834 35672
rect 26068 35290 26096 38762
rect 26252 36378 26280 38898
rect 26332 37800 26384 37806
rect 26332 37742 26384 37748
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26240 36032 26292 36038
rect 26240 35974 26292 35980
rect 26056 35284 26108 35290
rect 26056 35226 26108 35232
rect 26252 35086 26280 35974
rect 26344 35630 26372 37742
rect 26436 36718 26464 41550
rect 26528 38894 26556 41618
rect 27080 40526 27108 53654
rect 27160 44872 27212 44878
rect 27160 44814 27212 44820
rect 27068 40520 27120 40526
rect 27068 40462 27120 40468
rect 26608 40384 26660 40390
rect 26608 40326 26660 40332
rect 26700 40384 26752 40390
rect 26700 40326 26752 40332
rect 27068 40384 27120 40390
rect 27068 40326 27120 40332
rect 26516 38888 26568 38894
rect 26516 38830 26568 38836
rect 26620 38486 26648 40326
rect 26608 38480 26660 38486
rect 26608 38422 26660 38428
rect 26424 36712 26476 36718
rect 26424 36654 26476 36660
rect 26332 35624 26384 35630
rect 26332 35566 26384 35572
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26344 34542 26372 35566
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26528 35086 26556 35430
rect 26608 35284 26660 35290
rect 26608 35226 26660 35232
rect 26516 35080 26568 35086
rect 26516 35022 26568 35028
rect 25872 34536 25924 34542
rect 25872 34478 25924 34484
rect 26332 34536 26384 34542
rect 26332 34478 26384 34484
rect 25780 33516 25832 33522
rect 25780 33458 25832 33464
rect 25792 30054 25820 33458
rect 25884 30190 25912 34478
rect 26620 33930 26648 35226
rect 26608 33924 26660 33930
rect 26608 33866 26660 33872
rect 26712 33522 26740 40326
rect 27080 40089 27108 40326
rect 27066 40080 27122 40089
rect 27066 40015 27122 40024
rect 26976 39364 27028 39370
rect 26976 39306 27028 39312
rect 26988 39098 27016 39306
rect 27172 39098 27200 44814
rect 27344 43240 27396 43246
rect 27344 43182 27396 43188
rect 27356 42906 27384 43182
rect 27344 42900 27396 42906
rect 27344 42842 27396 42848
rect 27252 42560 27304 42566
rect 27252 42502 27304 42508
rect 27264 42022 27292 42502
rect 27356 42294 27384 42842
rect 27344 42288 27396 42294
rect 27344 42230 27396 42236
rect 27344 42152 27396 42158
rect 27344 42094 27396 42100
rect 27252 42016 27304 42022
rect 27252 41958 27304 41964
rect 27264 41138 27292 41958
rect 27252 41132 27304 41138
rect 27252 41074 27304 41080
rect 27252 40588 27304 40594
rect 27252 40530 27304 40536
rect 26976 39092 27028 39098
rect 26976 39034 27028 39040
rect 27160 39092 27212 39098
rect 27160 39034 27212 39040
rect 27068 39024 27120 39030
rect 27068 38966 27120 38972
rect 26792 38956 26844 38962
rect 26792 38898 26844 38904
rect 26804 38826 26832 38898
rect 26792 38820 26844 38826
rect 26792 38762 26844 38768
rect 26976 38752 27028 38758
rect 26976 38694 27028 38700
rect 26988 38214 27016 38694
rect 27080 38554 27108 38966
rect 27068 38548 27120 38554
rect 27068 38490 27120 38496
rect 27068 38412 27120 38418
rect 27068 38354 27120 38360
rect 26976 38208 27028 38214
rect 26976 38150 27028 38156
rect 27080 37806 27108 38354
rect 27160 38344 27212 38350
rect 27160 38286 27212 38292
rect 27172 38010 27200 38286
rect 27160 38004 27212 38010
rect 27160 37946 27212 37952
rect 27172 37874 27200 37946
rect 27160 37868 27212 37874
rect 27160 37810 27212 37816
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 27172 37330 27200 37810
rect 27160 37324 27212 37330
rect 27160 37266 27212 37272
rect 27068 37188 27120 37194
rect 27068 37130 27120 37136
rect 27080 35766 27108 37130
rect 27172 35834 27200 37266
rect 27160 35828 27212 35834
rect 27160 35770 27212 35776
rect 27068 35760 27120 35766
rect 27068 35702 27120 35708
rect 27080 35154 27108 35702
rect 27172 35698 27200 35770
rect 27160 35692 27212 35698
rect 27160 35634 27212 35640
rect 27172 35154 27200 35634
rect 27264 35290 27292 40530
rect 27356 36961 27384 42094
rect 27342 36952 27398 36961
rect 27342 36887 27398 36896
rect 27448 36802 27476 53926
rect 27950 53340 28258 53349
rect 27950 53338 27956 53340
rect 28012 53338 28036 53340
rect 28092 53338 28116 53340
rect 28172 53338 28196 53340
rect 28252 53338 28258 53340
rect 28012 53286 28014 53338
rect 28194 53286 28196 53338
rect 27950 53284 27956 53286
rect 28012 53284 28036 53286
rect 28092 53284 28116 53286
rect 28172 53284 28196 53286
rect 28252 53284 28258 53286
rect 27950 53275 28258 53284
rect 27950 52252 28258 52261
rect 27950 52250 27956 52252
rect 28012 52250 28036 52252
rect 28092 52250 28116 52252
rect 28172 52250 28196 52252
rect 28252 52250 28258 52252
rect 28012 52198 28014 52250
rect 28194 52198 28196 52250
rect 27950 52196 27956 52198
rect 28012 52196 28036 52198
rect 28092 52196 28116 52198
rect 28172 52196 28196 52198
rect 28252 52196 28258 52198
rect 27950 52187 28258 52196
rect 27950 51164 28258 51173
rect 27950 51162 27956 51164
rect 28012 51162 28036 51164
rect 28092 51162 28116 51164
rect 28172 51162 28196 51164
rect 28252 51162 28258 51164
rect 28012 51110 28014 51162
rect 28194 51110 28196 51162
rect 27950 51108 27956 51110
rect 28012 51108 28036 51110
rect 28092 51108 28116 51110
rect 28172 51108 28196 51110
rect 28252 51108 28258 51110
rect 27950 51099 28258 51108
rect 27950 50076 28258 50085
rect 27950 50074 27956 50076
rect 28012 50074 28036 50076
rect 28092 50074 28116 50076
rect 28172 50074 28196 50076
rect 28252 50074 28258 50076
rect 28012 50022 28014 50074
rect 28194 50022 28196 50074
rect 27950 50020 27956 50022
rect 28012 50020 28036 50022
rect 28092 50020 28116 50022
rect 28172 50020 28196 50022
rect 28252 50020 28258 50022
rect 27950 50011 28258 50020
rect 27950 48988 28258 48997
rect 27950 48986 27956 48988
rect 28012 48986 28036 48988
rect 28092 48986 28116 48988
rect 28172 48986 28196 48988
rect 28252 48986 28258 48988
rect 28012 48934 28014 48986
rect 28194 48934 28196 48986
rect 27950 48932 27956 48934
rect 28012 48932 28036 48934
rect 28092 48932 28116 48934
rect 28172 48932 28196 48934
rect 28252 48932 28258 48934
rect 27950 48923 28258 48932
rect 27950 47900 28258 47909
rect 27950 47898 27956 47900
rect 28012 47898 28036 47900
rect 28092 47898 28116 47900
rect 28172 47898 28196 47900
rect 28252 47898 28258 47900
rect 28012 47846 28014 47898
rect 28194 47846 28196 47898
rect 27950 47844 27956 47846
rect 28012 47844 28036 47846
rect 28092 47844 28116 47846
rect 28172 47844 28196 47846
rect 28252 47844 28258 47846
rect 27950 47835 28258 47844
rect 27950 46812 28258 46821
rect 27950 46810 27956 46812
rect 28012 46810 28036 46812
rect 28092 46810 28116 46812
rect 28172 46810 28196 46812
rect 28252 46810 28258 46812
rect 28012 46758 28014 46810
rect 28194 46758 28196 46810
rect 27950 46756 27956 46758
rect 28012 46756 28036 46758
rect 28092 46756 28116 46758
rect 28172 46756 28196 46758
rect 28252 46756 28258 46758
rect 27950 46747 28258 46756
rect 27712 45960 27764 45966
rect 27712 45902 27764 45908
rect 27724 41274 27752 45902
rect 27950 45724 28258 45733
rect 27950 45722 27956 45724
rect 28012 45722 28036 45724
rect 28092 45722 28116 45724
rect 28172 45722 28196 45724
rect 28252 45722 28258 45724
rect 28012 45670 28014 45722
rect 28194 45670 28196 45722
rect 27950 45668 27956 45670
rect 28012 45668 28036 45670
rect 28092 45668 28116 45670
rect 28172 45668 28196 45670
rect 28252 45668 28258 45670
rect 27950 45659 28258 45668
rect 27950 44636 28258 44645
rect 27950 44634 27956 44636
rect 28012 44634 28036 44636
rect 28092 44634 28116 44636
rect 28172 44634 28196 44636
rect 28252 44634 28258 44636
rect 28012 44582 28014 44634
rect 28194 44582 28196 44634
rect 27950 44580 27956 44582
rect 28012 44580 28036 44582
rect 28092 44580 28116 44582
rect 28172 44580 28196 44582
rect 28252 44580 28258 44582
rect 27950 44571 28258 44580
rect 27950 43548 28258 43557
rect 27950 43546 27956 43548
rect 28012 43546 28036 43548
rect 28092 43546 28116 43548
rect 28172 43546 28196 43548
rect 28252 43546 28258 43548
rect 28012 43494 28014 43546
rect 28194 43494 28196 43546
rect 27950 43492 27956 43494
rect 28012 43492 28036 43494
rect 28092 43492 28116 43494
rect 28172 43492 28196 43494
rect 28252 43492 28258 43494
rect 27950 43483 28258 43492
rect 27950 42460 28258 42469
rect 27950 42458 27956 42460
rect 28012 42458 28036 42460
rect 28092 42458 28116 42460
rect 28172 42458 28196 42460
rect 28252 42458 28258 42460
rect 28012 42406 28014 42458
rect 28194 42406 28196 42458
rect 27950 42404 27956 42406
rect 28012 42404 28036 42406
rect 28092 42404 28116 42406
rect 28172 42404 28196 42406
rect 28252 42404 28258 42406
rect 27950 42395 28258 42404
rect 28552 41414 28580 53926
rect 29104 53582 29132 56200
rect 29840 54194 29868 56200
rect 30576 54194 30604 56200
rect 31312 54194 31340 56200
rect 29828 54188 29880 54194
rect 29828 54130 29880 54136
rect 30564 54188 30616 54194
rect 30564 54130 30616 54136
rect 31300 54188 31352 54194
rect 31300 54130 31352 54136
rect 29644 54052 29696 54058
rect 29644 53994 29696 54000
rect 29092 53576 29144 53582
rect 29092 53518 29144 53524
rect 28816 43920 28868 43926
rect 28816 43862 28868 43868
rect 28632 43784 28684 43790
rect 28632 43726 28684 43732
rect 28644 43246 28672 43726
rect 28828 43450 28856 43862
rect 28920 43858 29040 43874
rect 28920 43852 29052 43858
rect 28920 43846 29000 43852
rect 28816 43444 28868 43450
rect 28816 43386 28868 43392
rect 28632 43240 28684 43246
rect 28632 43182 28684 43188
rect 28644 42022 28672 43182
rect 28632 42016 28684 42022
rect 28828 41970 28856 43386
rect 28920 43110 28948 43846
rect 29000 43794 29052 43800
rect 28908 43104 28960 43110
rect 28908 43046 28960 43052
rect 28632 41958 28684 41964
rect 28368 41386 28580 41414
rect 28736 41942 28856 41970
rect 27950 41372 28258 41381
rect 27950 41370 27956 41372
rect 28012 41370 28036 41372
rect 28092 41370 28116 41372
rect 28172 41370 28196 41372
rect 28252 41370 28258 41372
rect 28012 41318 28014 41370
rect 28194 41318 28196 41370
rect 27950 41316 27956 41318
rect 28012 41316 28036 41318
rect 28092 41316 28116 41318
rect 28172 41316 28196 41318
rect 28252 41316 28258 41318
rect 27950 41307 28258 41316
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 27988 41200 28040 41206
rect 27988 41142 28040 41148
rect 28000 41070 28028 41142
rect 27528 41064 27580 41070
rect 27528 41006 27580 41012
rect 27988 41064 28040 41070
rect 27988 41006 28040 41012
rect 27540 38842 27568 41006
rect 27950 40284 28258 40293
rect 27950 40282 27956 40284
rect 28012 40282 28036 40284
rect 28092 40282 28116 40284
rect 28172 40282 28196 40284
rect 28252 40282 28258 40284
rect 28012 40230 28014 40282
rect 28194 40230 28196 40282
rect 27950 40228 27956 40230
rect 28012 40228 28036 40230
rect 28092 40228 28116 40230
rect 28172 40228 28196 40230
rect 28252 40228 28258 40230
rect 27950 40219 28258 40228
rect 27712 39908 27764 39914
rect 27712 39850 27764 39856
rect 27540 38814 27660 38842
rect 27632 38298 27660 38814
rect 27540 38270 27660 38298
rect 27540 38010 27568 38270
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 27540 37466 27568 37946
rect 27528 37460 27580 37466
rect 27528 37402 27580 37408
rect 27620 37324 27672 37330
rect 27620 37266 27672 37272
rect 27344 36780 27396 36786
rect 27448 36774 27568 36802
rect 27344 36722 27396 36728
rect 27356 36378 27384 36722
rect 27436 36712 27488 36718
rect 27436 36654 27488 36660
rect 27448 36378 27476 36654
rect 27344 36372 27396 36378
rect 27344 36314 27396 36320
rect 27436 36372 27488 36378
rect 27436 36314 27488 36320
rect 27252 35284 27304 35290
rect 27252 35226 27304 35232
rect 27068 35148 27120 35154
rect 27068 35090 27120 35096
rect 27160 35148 27212 35154
rect 27160 35090 27212 35096
rect 27172 34610 27200 35090
rect 27160 34604 27212 34610
rect 27160 34546 27212 34552
rect 27172 34066 27200 34546
rect 27160 34060 27212 34066
rect 27160 34002 27212 34008
rect 27540 33946 27568 36774
rect 27632 35630 27660 37266
rect 27620 35624 27672 35630
rect 27620 35566 27672 35572
rect 27724 35494 27752 39850
rect 27950 39196 28258 39205
rect 27950 39194 27956 39196
rect 28012 39194 28036 39196
rect 28092 39194 28116 39196
rect 28172 39194 28196 39196
rect 28252 39194 28258 39196
rect 28012 39142 28014 39194
rect 28194 39142 28196 39194
rect 27950 39140 27956 39142
rect 28012 39140 28036 39142
rect 28092 39140 28116 39142
rect 28172 39140 28196 39142
rect 28252 39140 28258 39142
rect 27950 39131 28258 39140
rect 27986 38992 28042 39001
rect 27986 38927 28042 38936
rect 28000 38894 28028 38927
rect 27896 38888 27948 38894
rect 27896 38830 27948 38836
rect 27988 38888 28040 38894
rect 27988 38830 28040 38836
rect 27908 38298 27936 38830
rect 27816 38270 27936 38298
rect 27816 37806 27844 38270
rect 27950 38108 28258 38117
rect 27950 38106 27956 38108
rect 28012 38106 28036 38108
rect 28092 38106 28116 38108
rect 28172 38106 28196 38108
rect 28252 38106 28258 38108
rect 28012 38054 28014 38106
rect 28194 38054 28196 38106
rect 27950 38052 27956 38054
rect 28012 38052 28036 38054
rect 28092 38052 28116 38054
rect 28172 38052 28196 38054
rect 28252 38052 28258 38054
rect 27950 38043 28258 38052
rect 28172 37936 28224 37942
rect 28172 37878 28224 37884
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27816 37466 27844 37742
rect 27804 37460 27856 37466
rect 27804 37402 27856 37408
rect 28184 37262 28212 37878
rect 28172 37256 28224 37262
rect 28172 37198 28224 37204
rect 27950 37020 28258 37029
rect 27950 37018 27956 37020
rect 28012 37018 28036 37020
rect 28092 37018 28116 37020
rect 28172 37018 28196 37020
rect 28252 37018 28258 37020
rect 28012 36966 28014 37018
rect 28194 36966 28196 37018
rect 27950 36964 27956 36966
rect 28012 36964 28036 36966
rect 28092 36964 28116 36966
rect 28172 36964 28196 36966
rect 28252 36964 28258 36966
rect 27802 36952 27858 36961
rect 27950 36955 28258 36964
rect 27802 36887 27858 36896
rect 27816 36786 27844 36887
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 28172 36168 28224 36174
rect 28170 36136 28172 36145
rect 28224 36136 28226 36145
rect 28170 36071 28226 36080
rect 27950 35932 28258 35941
rect 27950 35930 27956 35932
rect 28012 35930 28036 35932
rect 28092 35930 28116 35932
rect 28172 35930 28196 35932
rect 28252 35930 28258 35932
rect 28012 35878 28014 35930
rect 28194 35878 28196 35930
rect 27950 35876 27956 35878
rect 28012 35876 28036 35878
rect 28092 35876 28116 35878
rect 28172 35876 28196 35878
rect 28252 35876 28258 35878
rect 27950 35867 28258 35876
rect 27712 35488 27764 35494
rect 27712 35430 27764 35436
rect 27710 35320 27766 35329
rect 27710 35255 27766 35264
rect 27172 33918 27568 33946
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 26700 33516 26752 33522
rect 26700 33458 26752 33464
rect 26974 33280 27030 33289
rect 26974 33215 27030 33224
rect 26988 32978 27016 33215
rect 26976 32972 27028 32978
rect 26976 32914 27028 32920
rect 26698 32872 26754 32881
rect 26424 32836 26476 32842
rect 26698 32807 26754 32816
rect 26424 32778 26476 32784
rect 26056 32564 26108 32570
rect 26056 32506 26108 32512
rect 26068 31890 26096 32506
rect 26240 32360 26292 32366
rect 26240 32302 26292 32308
rect 26056 31884 26108 31890
rect 26056 31826 26108 31832
rect 26252 31346 26280 32302
rect 26240 31340 26292 31346
rect 26240 31282 26292 31288
rect 26054 30424 26110 30433
rect 26054 30359 26110 30368
rect 25872 30184 25924 30190
rect 25872 30126 25924 30132
rect 25780 30048 25832 30054
rect 25780 29990 25832 29996
rect 25872 29776 25924 29782
rect 25700 29724 25872 29730
rect 25700 29718 25924 29724
rect 25700 29702 25912 29718
rect 25700 26246 25728 29702
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25688 25968 25740 25974
rect 25688 25910 25740 25916
rect 25700 25702 25728 25910
rect 25688 25696 25740 25702
rect 25688 25638 25740 25644
rect 25780 25696 25832 25702
rect 25780 25638 25832 25644
rect 25688 25356 25740 25362
rect 25688 25298 25740 25304
rect 25596 24744 25648 24750
rect 25596 24686 25648 24692
rect 25504 24404 25556 24410
rect 25504 24346 25556 24352
rect 25516 24313 25544 24346
rect 25502 24304 25558 24313
rect 25502 24239 25558 24248
rect 25516 24206 25544 24239
rect 25504 24200 25556 24206
rect 25504 24142 25556 24148
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25608 21622 25636 21830
rect 25596 21616 25648 21622
rect 25596 21558 25648 21564
rect 25700 21486 25728 25298
rect 25792 24954 25820 25638
rect 25780 24948 25832 24954
rect 25780 24890 25832 24896
rect 25872 23520 25924 23526
rect 25872 23462 25924 23468
rect 25884 21690 25912 23462
rect 25962 22536 26018 22545
rect 25962 22471 26018 22480
rect 25976 22030 26004 22471
rect 25964 22024 26016 22030
rect 25964 21966 26016 21972
rect 25872 21684 25924 21690
rect 25872 21626 25924 21632
rect 25688 21480 25740 21486
rect 25688 21422 25740 21428
rect 25700 20262 25728 21422
rect 25688 20256 25740 20262
rect 25688 20198 25740 20204
rect 25780 20256 25832 20262
rect 25780 20198 25832 20204
rect 25700 19922 25728 20198
rect 25688 19916 25740 19922
rect 25688 19858 25740 19864
rect 25596 19712 25648 19718
rect 25596 19654 25648 19660
rect 25608 17882 25636 19654
rect 25792 18766 25820 20198
rect 25780 18760 25832 18766
rect 25780 18702 25832 18708
rect 25872 18624 25924 18630
rect 25872 18566 25924 18572
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25596 17876 25648 17882
rect 25596 17818 25648 17824
rect 25688 16992 25740 16998
rect 25688 16934 25740 16940
rect 25596 15360 25648 15366
rect 25596 15302 25648 15308
rect 25412 13320 25464 13326
rect 25412 13262 25464 13268
rect 25608 3126 25636 15302
rect 25700 15026 25728 16934
rect 25780 16516 25832 16522
rect 25780 16458 25832 16464
rect 25792 16250 25820 16458
rect 25884 16250 25912 18566
rect 25976 16590 26004 18566
rect 26068 16590 26096 30359
rect 26436 26450 26464 32778
rect 26516 32768 26568 32774
rect 26516 32710 26568 32716
rect 26608 32768 26660 32774
rect 26608 32710 26660 32716
rect 26528 32502 26556 32710
rect 26516 32496 26568 32502
rect 26516 32438 26568 32444
rect 26620 32298 26648 32710
rect 26608 32292 26660 32298
rect 26608 32234 26660 32240
rect 26712 31482 26740 32807
rect 26700 31476 26752 31482
rect 26700 31418 26752 31424
rect 26884 31136 26936 31142
rect 26884 31078 26936 31084
rect 26896 30666 26924 31078
rect 26884 30660 26936 30666
rect 26884 30602 26936 30608
rect 26608 28008 26660 28014
rect 26608 27950 26660 27956
rect 26620 27334 26648 27950
rect 26700 27396 26752 27402
rect 26700 27338 26752 27344
rect 26608 27328 26660 27334
rect 26608 27270 26660 27276
rect 26516 26784 26568 26790
rect 26516 26726 26568 26732
rect 26424 26444 26476 26450
rect 26424 26386 26476 26392
rect 26436 26330 26464 26386
rect 26344 26302 26464 26330
rect 26148 25152 26200 25158
rect 26148 25094 26200 25100
rect 26160 24857 26188 25094
rect 26146 24848 26202 24857
rect 26146 24783 26202 24792
rect 26240 24064 26292 24070
rect 26240 24006 26292 24012
rect 26252 23633 26280 24006
rect 26238 23624 26294 23633
rect 26238 23559 26294 23568
rect 26148 23520 26200 23526
rect 26148 23462 26200 23468
rect 26160 20602 26188 23462
rect 26344 22710 26372 26302
rect 26424 26240 26476 26246
rect 26424 26182 26476 26188
rect 26436 25906 26464 26182
rect 26424 25900 26476 25906
rect 26424 25842 26476 25848
rect 26332 22704 26384 22710
rect 26332 22646 26384 22652
rect 26528 22506 26556 26726
rect 26712 25226 26740 27338
rect 26988 26874 27016 32914
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 27080 30802 27108 31962
rect 27172 31414 27200 33918
rect 27342 33824 27398 33833
rect 27342 33759 27398 33768
rect 27356 33454 27384 33759
rect 27344 33448 27396 33454
rect 27344 33390 27396 33396
rect 27252 33380 27304 33386
rect 27252 33322 27304 33328
rect 27264 32978 27292 33322
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27252 31884 27304 31890
rect 27252 31826 27304 31832
rect 27160 31408 27212 31414
rect 27160 31350 27212 31356
rect 27068 30796 27120 30802
rect 27068 30738 27120 30744
rect 27080 30326 27108 30738
rect 27068 30320 27120 30326
rect 27068 30262 27120 30268
rect 27080 29170 27108 30262
rect 27068 29164 27120 29170
rect 27068 29106 27120 29112
rect 27068 28484 27120 28490
rect 27068 28426 27120 28432
rect 27080 27713 27108 28426
rect 27066 27704 27122 27713
rect 27066 27639 27122 27648
rect 27172 27418 27200 31350
rect 27264 30598 27292 31826
rect 27356 30666 27384 33390
rect 27632 33130 27660 33934
rect 27540 33102 27660 33130
rect 27540 31754 27568 33102
rect 27528 31748 27580 31754
rect 27528 31690 27580 31696
rect 27540 31142 27568 31690
rect 27724 31686 27752 35255
rect 27950 34844 28258 34853
rect 27950 34842 27956 34844
rect 28012 34842 28036 34844
rect 28092 34842 28116 34844
rect 28172 34842 28196 34844
rect 28252 34842 28258 34844
rect 28012 34790 28014 34842
rect 28194 34790 28196 34842
rect 27950 34788 27956 34790
rect 28012 34788 28036 34790
rect 28092 34788 28116 34790
rect 28172 34788 28196 34790
rect 28252 34788 28258 34790
rect 27950 34779 28258 34788
rect 28172 34468 28224 34474
rect 28172 34410 28224 34416
rect 28184 34202 28212 34410
rect 28172 34196 28224 34202
rect 28172 34138 28224 34144
rect 27986 33960 28042 33969
rect 27986 33895 28042 33904
rect 28000 33862 28028 33895
rect 27804 33856 27856 33862
rect 27804 33798 27856 33804
rect 27988 33856 28040 33862
rect 27988 33798 28040 33804
rect 27816 33114 27844 33798
rect 27950 33756 28258 33765
rect 27950 33754 27956 33756
rect 28012 33754 28036 33756
rect 28092 33754 28116 33756
rect 28172 33754 28196 33756
rect 28252 33754 28258 33756
rect 28012 33702 28014 33754
rect 28194 33702 28196 33754
rect 27950 33700 27956 33702
rect 28012 33700 28036 33702
rect 28092 33700 28116 33702
rect 28172 33700 28196 33702
rect 28252 33700 28258 33702
rect 27950 33691 28258 33700
rect 27804 33108 27856 33114
rect 27804 33050 27856 33056
rect 27950 32668 28258 32677
rect 27950 32666 27956 32668
rect 28012 32666 28036 32668
rect 28092 32666 28116 32668
rect 28172 32666 28196 32668
rect 28252 32666 28258 32668
rect 28012 32614 28014 32666
rect 28194 32614 28196 32666
rect 27950 32612 27956 32614
rect 28012 32612 28036 32614
rect 28092 32612 28116 32614
rect 28172 32612 28196 32614
rect 28252 32612 28258 32614
rect 27950 32603 28258 32612
rect 27804 31748 27856 31754
rect 27804 31690 27856 31696
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27528 31136 27580 31142
rect 27528 31078 27580 31084
rect 27528 30932 27580 30938
rect 27528 30874 27580 30880
rect 27344 30660 27396 30666
rect 27344 30602 27396 30608
rect 27252 30592 27304 30598
rect 27252 30534 27304 30540
rect 27356 29714 27384 30602
rect 27436 30592 27488 30598
rect 27436 30534 27488 30540
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27448 28218 27476 30534
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 27172 27390 27384 27418
rect 27252 27328 27304 27334
rect 27252 27270 27304 27276
rect 26988 26846 27200 26874
rect 26700 25220 26752 25226
rect 26700 25162 26752 25168
rect 26712 24993 26740 25162
rect 26698 24984 26754 24993
rect 26698 24919 26754 24928
rect 26712 23594 26740 24919
rect 26884 24676 26936 24682
rect 26884 24618 26936 24624
rect 26896 24274 26924 24618
rect 26884 24268 26936 24274
rect 26884 24210 26936 24216
rect 26792 24064 26844 24070
rect 26792 24006 26844 24012
rect 26804 23798 26832 24006
rect 26792 23792 26844 23798
rect 26792 23734 26844 23740
rect 27068 23656 27120 23662
rect 27068 23598 27120 23604
rect 26700 23588 26752 23594
rect 26700 23530 26752 23536
rect 26516 22500 26568 22506
rect 26516 22442 26568 22448
rect 26148 20596 26200 20602
rect 26148 20538 26200 20544
rect 26424 19712 26476 19718
rect 26424 19654 26476 19660
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 25964 16584 26016 16590
rect 25964 16526 26016 16532
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 25780 16244 25832 16250
rect 25780 16186 25832 16192
rect 25872 16244 25924 16250
rect 25872 16186 25924 16192
rect 26056 16108 26108 16114
rect 26056 16050 26108 16056
rect 26068 15366 26096 16050
rect 26148 16040 26200 16046
rect 26148 15982 26200 15988
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 25700 14482 25728 14962
rect 26160 14958 26188 15982
rect 26436 15706 26464 19654
rect 26424 15700 26476 15706
rect 26424 15642 26476 15648
rect 26148 14952 26200 14958
rect 26148 14894 26200 14900
rect 25688 14476 25740 14482
rect 25688 14418 25740 14424
rect 26160 14346 26188 14894
rect 26332 14612 26384 14618
rect 26332 14554 26384 14560
rect 26148 14340 26200 14346
rect 26148 14282 26200 14288
rect 26344 14006 26372 14554
rect 26332 14000 26384 14006
rect 26332 13942 26384 13948
rect 25780 13184 25832 13190
rect 25780 13126 25832 13132
rect 25792 3534 25820 13126
rect 26528 12918 26556 22442
rect 26608 22432 26660 22438
rect 26608 22374 26660 22380
rect 26620 22166 26648 22374
rect 26608 22160 26660 22166
rect 26608 22102 26660 22108
rect 26700 21956 26752 21962
rect 26700 21898 26752 21904
rect 26608 20392 26660 20398
rect 26608 20334 26660 20340
rect 26620 19938 26648 20334
rect 26712 20058 26740 21898
rect 26700 20052 26752 20058
rect 26700 19994 26752 20000
rect 26620 19910 26740 19938
rect 26712 19446 26740 19910
rect 26976 19712 27028 19718
rect 26976 19654 27028 19660
rect 26700 19440 26752 19446
rect 26700 19382 26752 19388
rect 26792 19440 26844 19446
rect 26792 19382 26844 19388
rect 26608 18828 26660 18834
rect 26608 18770 26660 18776
rect 26620 17270 26648 18770
rect 26608 17264 26660 17270
rect 26608 17206 26660 17212
rect 26620 16998 26648 17206
rect 26608 16992 26660 16998
rect 26608 16934 26660 16940
rect 26620 14958 26648 16934
rect 26712 16658 26740 19382
rect 26804 18154 26832 19382
rect 26884 19168 26936 19174
rect 26884 19110 26936 19116
rect 26792 18148 26844 18154
rect 26792 18090 26844 18096
rect 26700 16652 26752 16658
rect 26700 16594 26752 16600
rect 26608 14952 26660 14958
rect 26608 14894 26660 14900
rect 26516 12912 26568 12918
rect 26516 12854 26568 12860
rect 25780 3528 25832 3534
rect 25780 3470 25832 3476
rect 26804 3398 26832 18090
rect 26896 3670 26924 19110
rect 26988 18834 27016 19654
rect 27080 19281 27108 23598
rect 27172 22094 27200 26846
rect 27264 25430 27292 27270
rect 27356 26790 27384 27390
rect 27344 26784 27396 26790
rect 27344 26726 27396 26732
rect 27540 25906 27568 30874
rect 27620 30388 27672 30394
rect 27620 30330 27672 30336
rect 27632 29714 27660 30330
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 27620 28688 27672 28694
rect 27620 28630 27672 28636
rect 27632 26994 27660 28630
rect 27724 28257 27752 31622
rect 27816 31346 27844 31690
rect 27950 31580 28258 31589
rect 27950 31578 27956 31580
rect 28012 31578 28036 31580
rect 28092 31578 28116 31580
rect 28172 31578 28196 31580
rect 28252 31578 28258 31580
rect 28012 31526 28014 31578
rect 28194 31526 28196 31578
rect 27950 31524 27956 31526
rect 28012 31524 28036 31526
rect 28092 31524 28116 31526
rect 28172 31524 28196 31526
rect 28252 31524 28258 31526
rect 27950 31515 28258 31524
rect 27804 31340 27856 31346
rect 27804 31282 27856 31288
rect 27950 30492 28258 30501
rect 27950 30490 27956 30492
rect 28012 30490 28036 30492
rect 28092 30490 28116 30492
rect 28172 30490 28196 30492
rect 28252 30490 28258 30492
rect 28012 30438 28014 30490
rect 28194 30438 28196 30490
rect 27950 30436 27956 30438
rect 28012 30436 28036 30438
rect 28092 30436 28116 30438
rect 28172 30436 28196 30438
rect 28252 30436 28258 30438
rect 27950 30427 28258 30436
rect 28264 30388 28316 30394
rect 28264 30330 28316 30336
rect 28276 30297 28304 30330
rect 28262 30288 28318 30297
rect 28262 30223 28318 30232
rect 28276 30122 28304 30223
rect 28264 30116 28316 30122
rect 28264 30058 28316 30064
rect 27950 29404 28258 29413
rect 27950 29402 27956 29404
rect 28012 29402 28036 29404
rect 28092 29402 28116 29404
rect 28172 29402 28196 29404
rect 28252 29402 28258 29404
rect 28012 29350 28014 29402
rect 28194 29350 28196 29402
rect 27950 29348 27956 29350
rect 28012 29348 28036 29350
rect 28092 29348 28116 29350
rect 28172 29348 28196 29350
rect 28252 29348 28258 29350
rect 27950 29339 28258 29348
rect 27950 28316 28258 28325
rect 27950 28314 27956 28316
rect 28012 28314 28036 28316
rect 28092 28314 28116 28316
rect 28172 28314 28196 28316
rect 28252 28314 28258 28316
rect 28012 28262 28014 28314
rect 28194 28262 28196 28314
rect 27950 28260 27956 28262
rect 28012 28260 28036 28262
rect 28092 28260 28116 28262
rect 28172 28260 28196 28262
rect 28252 28260 28258 28262
rect 27710 28248 27766 28257
rect 27950 28251 28258 28260
rect 27710 28183 27766 28192
rect 27712 28144 27764 28150
rect 27712 28086 27764 28092
rect 27620 26988 27672 26994
rect 27620 26930 27672 26936
rect 27632 26382 27660 26930
rect 27724 26450 27752 28086
rect 27804 28008 27856 28014
rect 27804 27950 27856 27956
rect 27816 27062 27844 27950
rect 27950 27228 28258 27237
rect 27950 27226 27956 27228
rect 28012 27226 28036 27228
rect 28092 27226 28116 27228
rect 28172 27226 28196 27228
rect 28252 27226 28258 27228
rect 28012 27174 28014 27226
rect 28194 27174 28196 27226
rect 27950 27172 27956 27174
rect 28012 27172 28036 27174
rect 28092 27172 28116 27174
rect 28172 27172 28196 27174
rect 28252 27172 28258 27174
rect 27950 27163 28258 27172
rect 27804 27056 27856 27062
rect 27804 26998 27856 27004
rect 28368 26450 28396 41386
rect 28736 39522 28764 41942
rect 28920 39982 28948 43046
rect 29184 42152 29236 42158
rect 29184 42094 29236 42100
rect 29092 42084 29144 42090
rect 29092 42026 29144 42032
rect 29104 41070 29132 42026
rect 29196 42022 29224 42094
rect 29184 42016 29236 42022
rect 29184 41958 29236 41964
rect 29656 41414 29684 53994
rect 30012 53984 30064 53990
rect 30012 53926 30064 53932
rect 30748 53984 30800 53990
rect 30748 53926 30800 53932
rect 31392 53984 31444 53990
rect 31392 53926 31444 53932
rect 29736 53440 29788 53446
rect 29736 53382 29788 53388
rect 29748 45490 29776 53382
rect 29736 45484 29788 45490
rect 29736 45426 29788 45432
rect 29828 42016 29880 42022
rect 29828 41958 29880 41964
rect 29380 41386 29684 41414
rect 29092 41064 29144 41070
rect 29092 41006 29144 41012
rect 29000 40928 29052 40934
rect 29000 40870 29052 40876
rect 29012 40662 29040 40870
rect 29000 40656 29052 40662
rect 29000 40598 29052 40604
rect 28908 39976 28960 39982
rect 28908 39918 28960 39924
rect 29184 39636 29236 39642
rect 29184 39578 29236 39584
rect 28448 39500 28500 39506
rect 28736 39494 28948 39522
rect 28448 39442 28500 39448
rect 28460 38962 28488 39442
rect 28724 39432 28776 39438
rect 28724 39374 28776 39380
rect 28448 38956 28500 38962
rect 28448 38898 28500 38904
rect 28736 38826 28764 39374
rect 28816 39296 28868 39302
rect 28816 39238 28868 39244
rect 28724 38820 28776 38826
rect 28724 38762 28776 38768
rect 28540 38752 28592 38758
rect 28540 38694 28592 38700
rect 28552 38418 28580 38694
rect 28540 38412 28592 38418
rect 28540 38354 28592 38360
rect 28632 36236 28684 36242
rect 28632 36178 28684 36184
rect 28448 34944 28500 34950
rect 28448 34886 28500 34892
rect 28540 34944 28592 34950
rect 28540 34886 28592 34892
rect 28460 32026 28488 34886
rect 28552 34678 28580 34886
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28540 34536 28592 34542
rect 28540 34478 28592 34484
rect 28552 32366 28580 34478
rect 28644 32978 28672 36178
rect 28736 36174 28764 38762
rect 28828 38486 28856 39238
rect 28816 38480 28868 38486
rect 28816 38422 28868 38428
rect 28816 38208 28868 38214
rect 28816 38150 28868 38156
rect 28828 37466 28856 38150
rect 28920 37738 28948 39494
rect 28908 37732 28960 37738
rect 28908 37674 28960 37680
rect 28816 37460 28868 37466
rect 28816 37402 28868 37408
rect 28724 36168 28776 36174
rect 28724 36110 28776 36116
rect 28920 35057 28948 37674
rect 29092 37324 29144 37330
rect 29092 37266 29144 37272
rect 29000 36780 29052 36786
rect 29000 36722 29052 36728
rect 28906 35048 28962 35057
rect 28906 34983 28962 34992
rect 28724 34740 28776 34746
rect 28724 34682 28776 34688
rect 28736 33017 28764 34682
rect 29012 33658 29040 36722
rect 29104 34542 29132 37266
rect 29092 34536 29144 34542
rect 29092 34478 29144 34484
rect 29092 33992 29144 33998
rect 29092 33934 29144 33940
rect 29104 33658 29132 33934
rect 29000 33652 29052 33658
rect 29000 33594 29052 33600
rect 29092 33652 29144 33658
rect 29092 33594 29144 33600
rect 29092 33448 29144 33454
rect 29092 33390 29144 33396
rect 28816 33312 28868 33318
rect 28954 33312 29006 33318
rect 28868 33272 28954 33300
rect 28816 33254 28868 33260
rect 28954 33254 29006 33260
rect 28722 33008 28778 33017
rect 28632 32972 28684 32978
rect 28722 32943 28778 32952
rect 28632 32914 28684 32920
rect 28540 32360 28592 32366
rect 28540 32302 28592 32308
rect 28538 32192 28594 32201
rect 28538 32127 28594 32136
rect 28448 32020 28500 32026
rect 28448 31962 28500 31968
rect 28448 27328 28500 27334
rect 28448 27270 28500 27276
rect 27712 26444 27764 26450
rect 27712 26386 27764 26392
rect 28356 26444 28408 26450
rect 28356 26386 28408 26392
rect 27620 26376 27672 26382
rect 27620 26318 27672 26324
rect 28356 26308 28408 26314
rect 28356 26250 28408 26256
rect 27950 26140 28258 26149
rect 27950 26138 27956 26140
rect 28012 26138 28036 26140
rect 28092 26138 28116 26140
rect 28172 26138 28196 26140
rect 28252 26138 28258 26140
rect 28012 26086 28014 26138
rect 28194 26086 28196 26138
rect 27950 26084 27956 26086
rect 28012 26084 28036 26086
rect 28092 26084 28116 26086
rect 28172 26084 28196 26086
rect 28252 26084 28258 26086
rect 27950 26075 28258 26084
rect 27804 26036 27856 26042
rect 27804 25978 27856 25984
rect 27528 25900 27580 25906
rect 27528 25842 27580 25848
rect 27344 25696 27396 25702
rect 27344 25638 27396 25644
rect 27436 25696 27488 25702
rect 27436 25638 27488 25644
rect 27252 25424 27304 25430
rect 27252 25366 27304 25372
rect 27172 22066 27292 22094
rect 27160 20460 27212 20466
rect 27160 20402 27212 20408
rect 27066 19272 27122 19281
rect 27172 19242 27200 20402
rect 27066 19207 27068 19216
rect 27120 19207 27122 19216
rect 27160 19236 27212 19242
rect 27068 19178 27120 19184
rect 27160 19178 27212 19184
rect 26976 18828 27028 18834
rect 26976 18770 27028 18776
rect 26884 3664 26936 3670
rect 26884 3606 26936 3612
rect 26792 3392 26844 3398
rect 26792 3334 26844 3340
rect 25596 3120 25648 3126
rect 25596 3062 25648 3068
rect 26988 2774 27016 18770
rect 27080 17814 27108 19178
rect 27264 19174 27292 22066
rect 27356 21078 27384 25638
rect 27448 24954 27476 25638
rect 27528 25356 27580 25362
rect 27528 25298 27580 25304
rect 27436 24948 27488 24954
rect 27436 24890 27488 24896
rect 27540 24886 27568 25298
rect 27620 25152 27672 25158
rect 27620 25094 27672 25100
rect 27632 24954 27660 25094
rect 27710 24984 27766 24993
rect 27620 24948 27672 24954
rect 27710 24919 27766 24928
rect 27620 24890 27672 24896
rect 27724 24886 27752 24919
rect 27528 24880 27580 24886
rect 27712 24880 27764 24886
rect 27528 24822 27580 24828
rect 27618 24848 27674 24857
rect 27540 24750 27568 24822
rect 27712 24822 27764 24828
rect 27618 24783 27674 24792
rect 27436 24744 27488 24750
rect 27436 24686 27488 24692
rect 27528 24744 27580 24750
rect 27528 24686 27580 24692
rect 27448 24274 27476 24686
rect 27436 24268 27488 24274
rect 27436 24210 27488 24216
rect 27436 23316 27488 23322
rect 27436 23258 27488 23264
rect 27448 22710 27476 23258
rect 27540 23186 27568 24686
rect 27528 23180 27580 23186
rect 27528 23122 27580 23128
rect 27528 23044 27580 23050
rect 27528 22986 27580 22992
rect 27436 22704 27488 22710
rect 27436 22646 27488 22652
rect 27540 22574 27568 22986
rect 27528 22568 27580 22574
rect 27528 22510 27580 22516
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27436 21412 27488 21418
rect 27436 21354 27488 21360
rect 27344 21072 27396 21078
rect 27344 21014 27396 21020
rect 27344 19916 27396 19922
rect 27344 19858 27396 19864
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27356 19122 27384 19858
rect 27448 19378 27476 21354
rect 27436 19372 27488 19378
rect 27436 19314 27488 19320
rect 27356 19094 27476 19122
rect 27252 18624 27304 18630
rect 27252 18566 27304 18572
rect 27344 18624 27396 18630
rect 27344 18566 27396 18572
rect 27160 18352 27212 18358
rect 27160 18294 27212 18300
rect 27068 17808 27120 17814
rect 27068 17750 27120 17756
rect 27172 16454 27200 18294
rect 27264 17338 27292 18566
rect 27356 18290 27384 18566
rect 27344 18284 27396 18290
rect 27344 18226 27396 18232
rect 27356 17542 27384 18226
rect 27448 18222 27476 19094
rect 27540 18766 27568 21830
rect 27632 18766 27660 24783
rect 27710 24168 27766 24177
rect 27710 24103 27766 24112
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27620 18760 27672 18766
rect 27620 18702 27672 18708
rect 27620 18420 27672 18426
rect 27620 18362 27672 18368
rect 27436 18216 27488 18222
rect 27436 18158 27488 18164
rect 27448 17746 27476 18158
rect 27436 17740 27488 17746
rect 27436 17682 27488 17688
rect 27344 17536 27396 17542
rect 27344 17478 27396 17484
rect 27252 17332 27304 17338
rect 27252 17274 27304 17280
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27252 16244 27304 16250
rect 27252 16186 27304 16192
rect 27264 15434 27292 16186
rect 27252 15428 27304 15434
rect 27252 15370 27304 15376
rect 27356 13394 27384 17478
rect 27448 16046 27476 17682
rect 27632 17678 27660 18362
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27724 17338 27752 24103
rect 27816 24070 27844 25978
rect 28368 25838 28396 26250
rect 28460 26042 28488 27270
rect 28448 26036 28500 26042
rect 28448 25978 28500 25984
rect 28356 25832 28408 25838
rect 28356 25774 28408 25780
rect 28264 25764 28316 25770
rect 28264 25706 28316 25712
rect 28276 25294 28304 25706
rect 28264 25288 28316 25294
rect 28264 25230 28316 25236
rect 27950 25052 28258 25061
rect 27950 25050 27956 25052
rect 28012 25050 28036 25052
rect 28092 25050 28116 25052
rect 28172 25050 28196 25052
rect 28252 25050 28258 25052
rect 28012 24998 28014 25050
rect 28194 24998 28196 25050
rect 27950 24996 27956 24998
rect 28012 24996 28036 24998
rect 28092 24996 28116 24998
rect 28172 24996 28196 24998
rect 28252 24996 28258 24998
rect 27950 24987 28258 24996
rect 28368 24834 28396 25774
rect 28552 25514 28580 32127
rect 28644 31890 28672 32914
rect 28724 32904 28776 32910
rect 28722 32872 28724 32881
rect 28776 32872 28778 32881
rect 28722 32807 28778 32816
rect 28906 32872 28962 32881
rect 28906 32807 28908 32816
rect 28960 32807 28962 32816
rect 29000 32836 29052 32842
rect 28908 32778 28960 32784
rect 29000 32778 29052 32784
rect 28724 32768 28776 32774
rect 29012 32722 29040 32778
rect 28724 32710 28776 32716
rect 28736 32298 28764 32710
rect 28966 32694 29040 32722
rect 28966 32586 28994 32694
rect 28920 32558 28994 32586
rect 28724 32292 28776 32298
rect 28724 32234 28776 32240
rect 28632 31884 28684 31890
rect 28632 31826 28684 31832
rect 28920 30870 28948 32558
rect 29104 32502 29132 33390
rect 29196 33318 29224 39578
rect 29276 37188 29328 37194
rect 29276 37130 29328 37136
rect 29184 33312 29236 33318
rect 29184 33254 29236 33260
rect 29288 32774 29316 37130
rect 29276 32768 29328 32774
rect 29276 32710 29328 32716
rect 29092 32496 29144 32502
rect 29092 32438 29144 32444
rect 29276 31136 29328 31142
rect 29276 31078 29328 31084
rect 28908 30864 28960 30870
rect 28908 30806 28960 30812
rect 29288 30802 29316 31078
rect 29276 30796 29328 30802
rect 29276 30738 29328 30744
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28828 30274 28856 30534
rect 28828 30258 29040 30274
rect 28828 30252 29052 30258
rect 28828 30246 29000 30252
rect 28828 29306 28856 30246
rect 29000 30194 29052 30200
rect 28908 30184 28960 30190
rect 28906 30152 28908 30161
rect 28960 30152 28962 30161
rect 28906 30087 28962 30096
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 28816 29300 28868 29306
rect 28816 29242 28868 29248
rect 28724 27396 28776 27402
rect 28724 27338 28776 27344
rect 28632 26376 28684 26382
rect 28632 26318 28684 26324
rect 28184 24806 28396 24834
rect 28460 25486 28580 25514
rect 28184 24750 28212 24806
rect 28172 24744 28224 24750
rect 28172 24686 28224 24692
rect 28460 24698 28488 25486
rect 28460 24670 28580 24698
rect 28448 24404 28500 24410
rect 28448 24346 28500 24352
rect 28080 24268 28132 24274
rect 28356 24268 28408 24274
rect 28132 24228 28356 24256
rect 28080 24210 28132 24216
rect 28356 24210 28408 24216
rect 28460 24206 28488 24346
rect 28448 24200 28500 24206
rect 28448 24142 28500 24148
rect 27804 24064 27856 24070
rect 27804 24006 27856 24012
rect 27816 22545 27844 24006
rect 27950 23964 28258 23973
rect 27950 23962 27956 23964
rect 28012 23962 28036 23964
rect 28092 23962 28116 23964
rect 28172 23962 28196 23964
rect 28252 23962 28258 23964
rect 28012 23910 28014 23962
rect 28194 23910 28196 23962
rect 27950 23908 27956 23910
rect 28012 23908 28036 23910
rect 28092 23908 28116 23910
rect 28172 23908 28196 23910
rect 28252 23908 28258 23910
rect 27950 23899 28258 23908
rect 27896 23588 27948 23594
rect 27896 23530 27948 23536
rect 27908 23186 27936 23530
rect 28552 23497 28580 24670
rect 28538 23488 28594 23497
rect 28538 23423 28594 23432
rect 28644 23338 28672 26318
rect 28736 24274 28764 27338
rect 28816 26444 28868 26450
rect 28816 26386 28868 26392
rect 28828 24993 28856 26386
rect 28920 25129 28948 29650
rect 29288 29238 29316 30738
rect 29380 29510 29408 41386
rect 29552 41268 29604 41274
rect 29552 41210 29604 41216
rect 29564 40730 29592 41210
rect 29840 41018 29868 41958
rect 29656 40990 29868 41018
rect 29920 40996 29972 41002
rect 29552 40724 29604 40730
rect 29552 40666 29604 40672
rect 29656 39642 29684 40990
rect 29920 40938 29972 40944
rect 29828 40928 29880 40934
rect 29828 40870 29880 40876
rect 29736 40520 29788 40526
rect 29736 40462 29788 40468
rect 29748 40118 29776 40462
rect 29736 40112 29788 40118
rect 29736 40054 29788 40060
rect 29840 39914 29868 40870
rect 29932 40390 29960 40938
rect 29920 40384 29972 40390
rect 29920 40326 29972 40332
rect 29828 39908 29880 39914
rect 29828 39850 29880 39856
rect 29644 39636 29696 39642
rect 29644 39578 29696 39584
rect 29828 39024 29880 39030
rect 29828 38966 29880 38972
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29642 37768 29698 37777
rect 29472 36689 29500 37742
rect 29642 37703 29698 37712
rect 29736 37732 29788 37738
rect 29458 36680 29514 36689
rect 29458 36615 29514 36624
rect 29656 36582 29684 37703
rect 29736 37674 29788 37680
rect 29748 37398 29776 37674
rect 29736 37392 29788 37398
rect 29736 37334 29788 37340
rect 29840 36922 29868 38966
rect 29932 38282 29960 40326
rect 29920 38276 29972 38282
rect 29920 38218 29972 38224
rect 29828 36916 29880 36922
rect 29828 36858 29880 36864
rect 29644 36576 29696 36582
rect 29644 36518 29696 36524
rect 29920 36576 29972 36582
rect 29920 36518 29972 36524
rect 29932 36106 29960 36518
rect 29920 36100 29972 36106
rect 29920 36042 29972 36048
rect 29460 35624 29512 35630
rect 29512 35584 29592 35612
rect 29460 35566 29512 35572
rect 29460 35216 29512 35222
rect 29460 35158 29512 35164
rect 29472 33454 29500 35158
rect 29460 33448 29512 33454
rect 29460 33390 29512 33396
rect 29564 29850 29592 35584
rect 29920 35148 29972 35154
rect 29920 35090 29972 35096
rect 29828 34944 29880 34950
rect 29828 34886 29880 34892
rect 29840 34610 29868 34886
rect 29828 34604 29880 34610
rect 29828 34546 29880 34552
rect 29932 34542 29960 35090
rect 29920 34536 29972 34542
rect 29920 34478 29972 34484
rect 30024 33810 30052 53926
rect 30656 43648 30708 43654
rect 30656 43590 30708 43596
rect 30196 39840 30248 39846
rect 30196 39782 30248 39788
rect 30288 39840 30340 39846
rect 30288 39782 30340 39788
rect 30104 39432 30156 39438
rect 30104 39374 30156 39380
rect 30116 38418 30144 39374
rect 30104 38412 30156 38418
rect 30104 38354 30156 38360
rect 30208 37398 30236 39782
rect 30300 39642 30328 39782
rect 30288 39636 30340 39642
rect 30288 39578 30340 39584
rect 30472 38276 30524 38282
rect 30472 38218 30524 38224
rect 30380 37868 30432 37874
rect 30380 37810 30432 37816
rect 30196 37392 30248 37398
rect 30196 37334 30248 37340
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 30116 34474 30144 35430
rect 30196 34944 30248 34950
rect 30196 34886 30248 34892
rect 30104 34468 30156 34474
rect 30104 34410 30156 34416
rect 29748 33782 30052 33810
rect 29644 33516 29696 33522
rect 29644 33458 29696 33464
rect 29552 29844 29604 29850
rect 29552 29786 29604 29792
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 29276 29232 29328 29238
rect 29276 29174 29328 29180
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 29012 25294 29040 28970
rect 29288 28082 29316 29174
rect 29276 28076 29328 28082
rect 29276 28018 29328 28024
rect 29184 27872 29236 27878
rect 29184 27814 29236 27820
rect 29196 26926 29224 27814
rect 29184 26920 29236 26926
rect 29184 26862 29236 26868
rect 29196 26586 29224 26862
rect 29184 26580 29236 26586
rect 29184 26522 29236 26528
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 29092 25288 29144 25294
rect 29092 25230 29144 25236
rect 29000 25152 29052 25158
rect 28906 25120 28962 25129
rect 29000 25094 29052 25100
rect 28906 25055 28962 25064
rect 28814 24984 28870 24993
rect 28814 24919 28870 24928
rect 28908 24948 28960 24954
rect 28908 24890 28960 24896
rect 28814 24712 28870 24721
rect 28814 24647 28870 24656
rect 28724 24268 28776 24274
rect 28724 24210 28776 24216
rect 28460 23310 28672 23338
rect 28736 23322 28764 24210
rect 28828 23712 28856 24647
rect 28920 24410 28948 24890
rect 29012 24614 29040 25094
rect 29000 24608 29052 24614
rect 29000 24550 29052 24556
rect 28908 24404 28960 24410
rect 28908 24346 28960 24352
rect 29104 24342 29132 25230
rect 29092 24336 29144 24342
rect 29092 24278 29144 24284
rect 29380 24154 29408 29446
rect 29460 29096 29512 29102
rect 29460 29038 29512 29044
rect 29472 28626 29500 29038
rect 29460 28620 29512 28626
rect 29460 28562 29512 28568
rect 29472 28218 29500 28562
rect 29460 28212 29512 28218
rect 29460 28154 29512 28160
rect 29460 28076 29512 28082
rect 29460 28018 29512 28024
rect 29472 27606 29500 28018
rect 29460 27600 29512 27606
rect 29460 27542 29512 27548
rect 29458 27296 29514 27305
rect 29458 27231 29514 27240
rect 29104 24126 29408 24154
rect 28908 23724 28960 23730
rect 28828 23684 28908 23712
rect 28724 23316 28776 23322
rect 27896 23180 27948 23186
rect 27896 23122 27948 23128
rect 27908 23050 27936 23122
rect 27896 23044 27948 23050
rect 27896 22986 27948 22992
rect 27950 22876 28258 22885
rect 27950 22874 27956 22876
rect 28012 22874 28036 22876
rect 28092 22874 28116 22876
rect 28172 22874 28196 22876
rect 28252 22874 28258 22876
rect 28012 22822 28014 22874
rect 28194 22822 28196 22874
rect 27950 22820 27956 22822
rect 28012 22820 28036 22822
rect 28092 22820 28116 22822
rect 28172 22820 28196 22822
rect 28252 22820 28258 22822
rect 27950 22811 28258 22820
rect 27802 22536 27858 22545
rect 27802 22471 27858 22480
rect 27804 22432 27856 22438
rect 27804 22374 27856 22380
rect 27816 21486 27844 22374
rect 27950 21788 28258 21797
rect 27950 21786 27956 21788
rect 28012 21786 28036 21788
rect 28092 21786 28116 21788
rect 28172 21786 28196 21788
rect 28252 21786 28258 21788
rect 28012 21734 28014 21786
rect 28194 21734 28196 21786
rect 27950 21732 27956 21734
rect 28012 21732 28036 21734
rect 28092 21732 28116 21734
rect 28172 21732 28196 21734
rect 28252 21732 28258 21734
rect 27950 21723 28258 21732
rect 28172 21548 28224 21554
rect 28172 21490 28224 21496
rect 27804 21480 27856 21486
rect 27804 21422 27856 21428
rect 27816 19514 27844 21422
rect 28184 21146 28212 21490
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 27950 20700 28258 20709
rect 27950 20698 27956 20700
rect 28012 20698 28036 20700
rect 28092 20698 28116 20700
rect 28172 20698 28196 20700
rect 28252 20698 28258 20700
rect 28012 20646 28014 20698
rect 28194 20646 28196 20698
rect 27950 20644 27956 20646
rect 28012 20644 28036 20646
rect 28092 20644 28116 20646
rect 28172 20644 28196 20646
rect 28252 20644 28258 20646
rect 27950 20635 28258 20644
rect 27950 19612 28258 19621
rect 27950 19610 27956 19612
rect 28012 19610 28036 19612
rect 28092 19610 28116 19612
rect 28172 19610 28196 19612
rect 28252 19610 28258 19612
rect 28012 19558 28014 19610
rect 28194 19558 28196 19610
rect 27950 19556 27956 19558
rect 28012 19556 28036 19558
rect 28092 19556 28116 19558
rect 28172 19556 28196 19558
rect 28252 19556 28258 19558
rect 27950 19547 28258 19556
rect 27804 19508 27856 19514
rect 27804 19450 27856 19456
rect 27804 19304 27856 19310
rect 27804 19246 27856 19252
rect 27816 18970 27844 19246
rect 27804 18964 27856 18970
rect 27804 18906 27856 18912
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 27950 18524 28258 18533
rect 27950 18522 27956 18524
rect 28012 18522 28036 18524
rect 28092 18522 28116 18524
rect 28172 18522 28196 18524
rect 28252 18522 28258 18524
rect 28012 18470 28014 18522
rect 28194 18470 28196 18522
rect 27950 18468 27956 18470
rect 28012 18468 28036 18470
rect 28092 18468 28116 18470
rect 28172 18468 28196 18470
rect 28252 18468 28258 18470
rect 27950 18459 28258 18468
rect 27950 17436 28258 17445
rect 27950 17434 27956 17436
rect 28012 17434 28036 17436
rect 28092 17434 28116 17436
rect 28172 17434 28196 17436
rect 28252 17434 28258 17436
rect 28012 17382 28014 17434
rect 28194 17382 28196 17434
rect 27950 17380 27956 17382
rect 28012 17380 28036 17382
rect 28092 17380 28116 17382
rect 28172 17380 28196 17382
rect 28252 17380 28258 17382
rect 27950 17371 28258 17380
rect 27712 17332 27764 17338
rect 27712 17274 27764 17280
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27436 16040 27488 16046
rect 27436 15982 27488 15988
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27540 12986 27568 16390
rect 27620 15972 27672 15978
rect 27620 15914 27672 15920
rect 27632 15026 27660 15914
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27528 12980 27580 12986
rect 27528 12922 27580 12928
rect 27160 12708 27212 12714
rect 27160 12650 27212 12656
rect 26804 2746 27016 2774
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 26516 2508 26568 2514
rect 26516 2450 26568 2456
rect 25320 1624 25372 1630
rect 25320 1566 25372 1572
rect 25792 800 25820 2450
rect 26528 800 26556 2450
rect 26804 1970 26832 2746
rect 27172 2446 27200 12650
rect 27252 2984 27304 2990
rect 27252 2926 27304 2932
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 26792 1964 26844 1970
rect 26792 1906 26844 1912
rect 27264 800 27292 2926
rect 27724 2582 27752 17274
rect 28264 17128 28316 17134
rect 28264 17070 28316 17076
rect 28276 16454 28304 17070
rect 28264 16448 28316 16454
rect 28264 16390 28316 16396
rect 27950 16348 28258 16357
rect 27950 16346 27956 16348
rect 28012 16346 28036 16348
rect 28092 16346 28116 16348
rect 28172 16346 28196 16348
rect 28252 16346 28258 16348
rect 28012 16294 28014 16346
rect 28194 16294 28196 16346
rect 27950 16292 27956 16294
rect 28012 16292 28036 16294
rect 28092 16292 28116 16294
rect 28172 16292 28196 16294
rect 28252 16292 28258 16294
rect 27950 16283 28258 16292
rect 27950 15260 28258 15269
rect 27950 15258 27956 15260
rect 28012 15258 28036 15260
rect 28092 15258 28116 15260
rect 28172 15258 28196 15260
rect 28252 15258 28258 15260
rect 28012 15206 28014 15258
rect 28194 15206 28196 15258
rect 27950 15204 27956 15206
rect 28012 15204 28036 15206
rect 28092 15204 28116 15206
rect 28172 15204 28196 15206
rect 28252 15204 28258 15206
rect 27950 15195 28258 15204
rect 27804 15088 27856 15094
rect 27804 15030 27856 15036
rect 27816 13530 27844 15030
rect 27896 14952 27948 14958
rect 27896 14894 27948 14900
rect 27908 14618 27936 14894
rect 27896 14612 27948 14618
rect 27896 14554 27948 14560
rect 27950 14172 28258 14181
rect 27950 14170 27956 14172
rect 28012 14170 28036 14172
rect 28092 14170 28116 14172
rect 28172 14170 28196 14172
rect 28252 14170 28258 14172
rect 28012 14118 28014 14170
rect 28194 14118 28196 14170
rect 27950 14116 27956 14118
rect 28012 14116 28036 14118
rect 28092 14116 28116 14118
rect 28172 14116 28196 14118
rect 28252 14116 28258 14118
rect 27950 14107 28258 14116
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27804 13388 27856 13394
rect 27804 13330 27856 13336
rect 27816 2650 27844 13330
rect 27950 13084 28258 13093
rect 27950 13082 27956 13084
rect 28012 13082 28036 13084
rect 28092 13082 28116 13084
rect 28172 13082 28196 13084
rect 28252 13082 28258 13084
rect 28012 13030 28014 13082
rect 28194 13030 28196 13082
rect 27950 13028 27956 13030
rect 28012 13028 28036 13030
rect 28092 13028 28116 13030
rect 28172 13028 28196 13030
rect 28252 13028 28258 13030
rect 27950 13019 28258 13028
rect 28368 12918 28396 18702
rect 28460 18698 28488 23310
rect 28724 23258 28776 23264
rect 28828 23202 28856 23684
rect 28908 23666 28960 23672
rect 28906 23624 28962 23633
rect 28906 23559 28908 23568
rect 28960 23559 28962 23568
rect 28908 23530 28960 23536
rect 28736 23174 28856 23202
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28552 22642 28580 23054
rect 28540 22636 28592 22642
rect 28540 22578 28592 22584
rect 28540 22092 28592 22098
rect 28540 22034 28592 22040
rect 28552 22001 28580 22034
rect 28538 21992 28594 22001
rect 28538 21927 28594 21936
rect 28552 21434 28580 21927
rect 28552 21406 28672 21434
rect 28538 19272 28594 19281
rect 28538 19207 28540 19216
rect 28592 19207 28594 19216
rect 28540 19178 28592 19184
rect 28540 18964 28592 18970
rect 28540 18906 28592 18912
rect 28448 18692 28500 18698
rect 28448 18634 28500 18640
rect 28460 18358 28488 18634
rect 28448 18352 28500 18358
rect 28448 18294 28500 18300
rect 28552 18170 28580 18906
rect 28460 18142 28580 18170
rect 28460 17202 28488 18142
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28540 17128 28592 17134
rect 28540 17070 28592 17076
rect 28448 16992 28500 16998
rect 28448 16934 28500 16940
rect 28460 16590 28488 16934
rect 28448 16584 28500 16590
rect 28448 16526 28500 16532
rect 28552 16454 28580 17070
rect 28448 16448 28500 16454
rect 28448 16390 28500 16396
rect 28540 16448 28592 16454
rect 28540 16390 28592 16396
rect 28460 13394 28488 16390
rect 28448 13388 28500 13394
rect 28448 13330 28500 13336
rect 28356 12912 28408 12918
rect 28356 12854 28408 12860
rect 28460 12850 28488 13330
rect 28448 12844 28500 12850
rect 28448 12786 28500 12792
rect 28552 12730 28580 16390
rect 28368 12702 28580 12730
rect 27950 11996 28258 12005
rect 27950 11994 27956 11996
rect 28012 11994 28036 11996
rect 28092 11994 28116 11996
rect 28172 11994 28196 11996
rect 28252 11994 28258 11996
rect 28012 11942 28014 11994
rect 28194 11942 28196 11994
rect 27950 11940 27956 11942
rect 28012 11940 28036 11942
rect 28092 11940 28116 11942
rect 28172 11940 28196 11942
rect 28252 11940 28258 11942
rect 27950 11931 28258 11940
rect 27950 10908 28258 10917
rect 27950 10906 27956 10908
rect 28012 10906 28036 10908
rect 28092 10906 28116 10908
rect 28172 10906 28196 10908
rect 28252 10906 28258 10908
rect 28012 10854 28014 10906
rect 28194 10854 28196 10906
rect 27950 10852 27956 10854
rect 28012 10852 28036 10854
rect 28092 10852 28116 10854
rect 28172 10852 28196 10854
rect 28252 10852 28258 10854
rect 27950 10843 28258 10852
rect 27950 9820 28258 9829
rect 27950 9818 27956 9820
rect 28012 9818 28036 9820
rect 28092 9818 28116 9820
rect 28172 9818 28196 9820
rect 28252 9818 28258 9820
rect 28012 9766 28014 9818
rect 28194 9766 28196 9818
rect 27950 9764 27956 9766
rect 28012 9764 28036 9766
rect 28092 9764 28116 9766
rect 28172 9764 28196 9766
rect 28252 9764 28258 9766
rect 27950 9755 28258 9764
rect 27950 8732 28258 8741
rect 27950 8730 27956 8732
rect 28012 8730 28036 8732
rect 28092 8730 28116 8732
rect 28172 8730 28196 8732
rect 28252 8730 28258 8732
rect 28012 8678 28014 8730
rect 28194 8678 28196 8730
rect 27950 8676 27956 8678
rect 28012 8676 28036 8678
rect 28092 8676 28116 8678
rect 28172 8676 28196 8678
rect 28252 8676 28258 8678
rect 27950 8667 28258 8676
rect 27950 7644 28258 7653
rect 27950 7642 27956 7644
rect 28012 7642 28036 7644
rect 28092 7642 28116 7644
rect 28172 7642 28196 7644
rect 28252 7642 28258 7644
rect 28012 7590 28014 7642
rect 28194 7590 28196 7642
rect 27950 7588 27956 7590
rect 28012 7588 28036 7590
rect 28092 7588 28116 7590
rect 28172 7588 28196 7590
rect 28252 7588 28258 7590
rect 27950 7579 28258 7588
rect 27950 6556 28258 6565
rect 27950 6554 27956 6556
rect 28012 6554 28036 6556
rect 28092 6554 28116 6556
rect 28172 6554 28196 6556
rect 28252 6554 28258 6556
rect 28012 6502 28014 6554
rect 28194 6502 28196 6554
rect 27950 6500 27956 6502
rect 28012 6500 28036 6502
rect 28092 6500 28116 6502
rect 28172 6500 28196 6502
rect 28252 6500 28258 6502
rect 27950 6491 28258 6500
rect 27950 5468 28258 5477
rect 27950 5466 27956 5468
rect 28012 5466 28036 5468
rect 28092 5466 28116 5468
rect 28172 5466 28196 5468
rect 28252 5466 28258 5468
rect 28012 5414 28014 5466
rect 28194 5414 28196 5466
rect 27950 5412 27956 5414
rect 28012 5412 28036 5414
rect 28092 5412 28116 5414
rect 28172 5412 28196 5414
rect 28252 5412 28258 5414
rect 27950 5403 28258 5412
rect 27950 4380 28258 4389
rect 27950 4378 27956 4380
rect 28012 4378 28036 4380
rect 28092 4378 28116 4380
rect 28172 4378 28196 4380
rect 28252 4378 28258 4380
rect 28012 4326 28014 4378
rect 28194 4326 28196 4378
rect 27950 4324 27956 4326
rect 28012 4324 28036 4326
rect 28092 4324 28116 4326
rect 28172 4324 28196 4326
rect 28252 4324 28258 4326
rect 27950 4315 28258 4324
rect 27950 3292 28258 3301
rect 27950 3290 27956 3292
rect 28012 3290 28036 3292
rect 28092 3290 28116 3292
rect 28172 3290 28196 3292
rect 28252 3290 28258 3292
rect 28012 3238 28014 3290
rect 28194 3238 28196 3290
rect 27950 3236 27956 3238
rect 28012 3236 28036 3238
rect 28092 3236 28116 3238
rect 28172 3236 28196 3238
rect 28252 3236 28258 3238
rect 27950 3227 28258 3236
rect 28368 2922 28396 12702
rect 28644 12594 28672 21406
rect 28460 12566 28672 12594
rect 28356 2916 28408 2922
rect 28356 2858 28408 2864
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 27712 2576 27764 2582
rect 27712 2518 27764 2524
rect 28356 2508 28408 2514
rect 28356 2450 28408 2456
rect 27950 2204 28258 2213
rect 27950 2202 27956 2204
rect 28012 2202 28036 2204
rect 28092 2202 28116 2204
rect 28172 2202 28196 2204
rect 28252 2202 28258 2204
rect 28012 2150 28014 2202
rect 28194 2150 28196 2202
rect 27950 2148 27956 2150
rect 28012 2148 28036 2150
rect 28092 2148 28116 2150
rect 28172 2148 28196 2150
rect 28252 2148 28258 2150
rect 27950 2139 28258 2148
rect 28000 870 28120 898
rect 28000 800 28028 870
rect 7852 734 8064 762
rect 8114 0 8170 800
rect 8850 0 8906 800
rect 9586 0 9642 800
rect 10322 0 10378 800
rect 11058 0 11114 800
rect 11794 0 11850 800
rect 12530 0 12586 800
rect 13266 0 13322 800
rect 14002 0 14058 800
rect 14738 0 14794 800
rect 15474 0 15530 800
rect 16210 0 16266 800
rect 16946 0 17002 800
rect 17682 0 17738 800
rect 18418 0 18474 800
rect 19154 0 19210 800
rect 19890 0 19946 800
rect 20626 0 20682 800
rect 21362 0 21418 800
rect 22098 0 22154 800
rect 22834 0 22890 800
rect 23570 0 23626 800
rect 24306 0 24362 800
rect 25042 0 25098 800
rect 25778 0 25834 800
rect 26514 0 26570 800
rect 27250 0 27306 800
rect 27986 0 28042 800
rect 28092 762 28120 870
rect 28368 762 28396 2450
rect 28460 2106 28488 12566
rect 28538 12472 28594 12481
rect 28736 12434 28764 23174
rect 29104 22094 29132 24126
rect 29276 23792 29328 23798
rect 29276 23734 29328 23740
rect 29184 22976 29236 22982
rect 29184 22918 29236 22924
rect 29012 22066 29132 22094
rect 28816 21888 28868 21894
rect 28816 21830 28868 21836
rect 28828 20874 28856 21830
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 28816 20868 28868 20874
rect 28816 20810 28868 20816
rect 28920 19854 28948 21354
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 28816 19508 28868 19514
rect 28816 19450 28868 19456
rect 28828 18834 28856 19450
rect 28816 18828 28868 18834
rect 28816 18770 28868 18776
rect 28814 17368 28870 17377
rect 28814 17303 28816 17312
rect 28868 17303 28870 17312
rect 28816 17274 28868 17280
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28828 15570 28856 16050
rect 28816 15564 28868 15570
rect 28816 15506 28868 15512
rect 28920 15450 28948 19790
rect 29012 15502 29040 22066
rect 29090 19408 29146 19417
rect 29090 19343 29092 19352
rect 29144 19343 29146 19352
rect 29092 19314 29144 19320
rect 29092 18080 29144 18086
rect 29090 18048 29092 18057
rect 29144 18048 29146 18057
rect 29196 18034 29224 22918
rect 29288 18630 29316 23734
rect 29472 22982 29500 27231
rect 29552 26036 29604 26042
rect 29552 25978 29604 25984
rect 29564 24274 29592 25978
rect 29552 24268 29604 24274
rect 29552 24210 29604 24216
rect 29460 22976 29512 22982
rect 29460 22918 29512 22924
rect 29656 22094 29684 33458
rect 29748 28490 29776 33782
rect 30104 33312 30156 33318
rect 30104 33254 30156 33260
rect 30012 30252 30064 30258
rect 30012 30194 30064 30200
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 29840 29646 29868 30126
rect 30024 29782 30052 30194
rect 30012 29776 30064 29782
rect 30012 29718 30064 29724
rect 30116 29714 30144 33254
rect 30208 32978 30236 34886
rect 30288 34536 30340 34542
rect 30288 34478 30340 34484
rect 30300 33114 30328 34478
rect 30288 33108 30340 33114
rect 30288 33050 30340 33056
rect 30196 32972 30248 32978
rect 30196 32914 30248 32920
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 30208 30705 30236 30874
rect 30194 30696 30250 30705
rect 30194 30631 30250 30640
rect 30208 30598 30236 30631
rect 30196 30592 30248 30598
rect 30196 30534 30248 30540
rect 30288 30388 30340 30394
rect 30288 30330 30340 30336
rect 30104 29708 30156 29714
rect 30104 29650 30156 29656
rect 29828 29640 29880 29646
rect 29828 29582 29880 29588
rect 30012 29640 30064 29646
rect 30012 29582 30064 29588
rect 29840 29102 29868 29582
rect 30024 29238 30052 29582
rect 30196 29572 30248 29578
rect 30196 29514 30248 29520
rect 30012 29232 30064 29238
rect 30012 29174 30064 29180
rect 29828 29096 29880 29102
rect 29828 29038 29880 29044
rect 30012 29028 30064 29034
rect 30012 28970 30064 28976
rect 29920 28552 29972 28558
rect 29920 28494 29972 28500
rect 29736 28484 29788 28490
rect 29736 28426 29788 28432
rect 29932 27470 29960 28494
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29828 25764 29880 25770
rect 29828 25706 29880 25712
rect 29840 24138 29868 25706
rect 29920 25696 29972 25702
rect 29920 25638 29972 25644
rect 29932 25344 29960 25638
rect 30024 25498 30052 28970
rect 30104 28008 30156 28014
rect 30104 27950 30156 27956
rect 30116 27062 30144 27950
rect 30208 27418 30236 29514
rect 30300 27538 30328 30330
rect 30392 28694 30420 37810
rect 30484 35698 30512 38218
rect 30472 35692 30524 35698
rect 30472 35634 30524 35640
rect 30484 35494 30512 35634
rect 30472 35488 30524 35494
rect 30524 35436 30604 35442
rect 30472 35430 30604 35436
rect 30484 35414 30604 35430
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 30484 34746 30512 35226
rect 30576 35154 30604 35414
rect 30564 35148 30616 35154
rect 30564 35090 30616 35096
rect 30472 34740 30524 34746
rect 30472 34682 30524 34688
rect 30576 34678 30604 35090
rect 30668 34746 30696 43590
rect 30760 40089 30788 53926
rect 31404 43450 31432 53926
rect 32048 53582 32076 56200
rect 32784 54262 32812 56200
rect 33520 54262 33548 56200
rect 32772 54256 32824 54262
rect 32772 54198 32824 54204
rect 33508 54256 33560 54262
rect 33508 54198 33560 54204
rect 34256 54194 34284 56200
rect 34244 54188 34296 54194
rect 34244 54130 34296 54136
rect 33324 54052 33376 54058
rect 33324 53994 33376 54000
rect 33968 54052 34020 54058
rect 33968 53994 34020 54000
rect 32950 53884 33258 53893
rect 32950 53882 32956 53884
rect 33012 53882 33036 53884
rect 33092 53882 33116 53884
rect 33172 53882 33196 53884
rect 33252 53882 33258 53884
rect 33012 53830 33014 53882
rect 33194 53830 33196 53882
rect 32950 53828 32956 53830
rect 33012 53828 33036 53830
rect 33092 53828 33116 53830
rect 33172 53828 33196 53830
rect 33252 53828 33258 53830
rect 32950 53819 33258 53828
rect 32036 53576 32088 53582
rect 32036 53518 32088 53524
rect 32128 53440 32180 53446
rect 32128 53382 32180 53388
rect 32140 45558 32168 53382
rect 32950 52796 33258 52805
rect 32950 52794 32956 52796
rect 33012 52794 33036 52796
rect 33092 52794 33116 52796
rect 33172 52794 33196 52796
rect 33252 52794 33258 52796
rect 33012 52742 33014 52794
rect 33194 52742 33196 52794
rect 32950 52740 32956 52742
rect 33012 52740 33036 52742
rect 33092 52740 33116 52742
rect 33172 52740 33196 52742
rect 33252 52740 33258 52742
rect 32950 52731 33258 52740
rect 32950 51708 33258 51717
rect 32950 51706 32956 51708
rect 33012 51706 33036 51708
rect 33092 51706 33116 51708
rect 33172 51706 33196 51708
rect 33252 51706 33258 51708
rect 33012 51654 33014 51706
rect 33194 51654 33196 51706
rect 32950 51652 32956 51654
rect 33012 51652 33036 51654
rect 33092 51652 33116 51654
rect 33172 51652 33196 51654
rect 33252 51652 33258 51654
rect 32950 51643 33258 51652
rect 32950 50620 33258 50629
rect 32950 50618 32956 50620
rect 33012 50618 33036 50620
rect 33092 50618 33116 50620
rect 33172 50618 33196 50620
rect 33252 50618 33258 50620
rect 33012 50566 33014 50618
rect 33194 50566 33196 50618
rect 32950 50564 32956 50566
rect 33012 50564 33036 50566
rect 33092 50564 33116 50566
rect 33172 50564 33196 50566
rect 33252 50564 33258 50566
rect 32950 50555 33258 50564
rect 32950 49532 33258 49541
rect 32950 49530 32956 49532
rect 33012 49530 33036 49532
rect 33092 49530 33116 49532
rect 33172 49530 33196 49532
rect 33252 49530 33258 49532
rect 33012 49478 33014 49530
rect 33194 49478 33196 49530
rect 32950 49476 32956 49478
rect 33012 49476 33036 49478
rect 33092 49476 33116 49478
rect 33172 49476 33196 49478
rect 33252 49476 33258 49478
rect 32950 49467 33258 49476
rect 32950 48444 33258 48453
rect 32950 48442 32956 48444
rect 33012 48442 33036 48444
rect 33092 48442 33116 48444
rect 33172 48442 33196 48444
rect 33252 48442 33258 48444
rect 33012 48390 33014 48442
rect 33194 48390 33196 48442
rect 32950 48388 32956 48390
rect 33012 48388 33036 48390
rect 33092 48388 33116 48390
rect 33172 48388 33196 48390
rect 33252 48388 33258 48390
rect 32950 48379 33258 48388
rect 32950 47356 33258 47365
rect 32950 47354 32956 47356
rect 33012 47354 33036 47356
rect 33092 47354 33116 47356
rect 33172 47354 33196 47356
rect 33252 47354 33258 47356
rect 33012 47302 33014 47354
rect 33194 47302 33196 47354
rect 32950 47300 32956 47302
rect 33012 47300 33036 47302
rect 33092 47300 33116 47302
rect 33172 47300 33196 47302
rect 33252 47300 33258 47302
rect 32950 47291 33258 47300
rect 32950 46268 33258 46277
rect 32950 46266 32956 46268
rect 33012 46266 33036 46268
rect 33092 46266 33116 46268
rect 33172 46266 33196 46268
rect 33252 46266 33258 46268
rect 33012 46214 33014 46266
rect 33194 46214 33196 46266
rect 32950 46212 32956 46214
rect 33012 46212 33036 46214
rect 33092 46212 33116 46214
rect 33172 46212 33196 46214
rect 33252 46212 33258 46214
rect 32950 46203 33258 46212
rect 32128 45552 32180 45558
rect 32128 45494 32180 45500
rect 33336 45554 33364 53994
rect 33980 45558 34008 53994
rect 34992 53582 35020 56200
rect 35728 54194 35756 56200
rect 36464 54194 36492 56200
rect 37200 54262 37228 56200
rect 37936 55214 37964 56200
rect 37844 55186 37964 55214
rect 37188 54256 37240 54262
rect 37188 54198 37240 54204
rect 35716 54188 35768 54194
rect 35716 54130 35768 54136
rect 36452 54188 36504 54194
rect 36452 54130 36504 54136
rect 35072 53984 35124 53990
rect 35072 53926 35124 53932
rect 36544 53984 36596 53990
rect 36544 53926 36596 53932
rect 36728 53984 36780 53990
rect 36728 53926 36780 53932
rect 37648 53984 37700 53990
rect 37648 53926 37700 53932
rect 34980 53576 35032 53582
rect 34980 53518 35032 53524
rect 33968 45554 34020 45558
rect 33336 45526 33732 45554
rect 33336 45490 33364 45526
rect 33324 45484 33376 45490
rect 33324 45426 33376 45432
rect 32864 45416 32916 45422
rect 32864 45358 32916 45364
rect 32680 45280 32732 45286
rect 32680 45222 32732 45228
rect 32404 44804 32456 44810
rect 32404 44746 32456 44752
rect 32036 43988 32088 43994
rect 32036 43930 32088 43936
rect 31668 43716 31720 43722
rect 31668 43658 31720 43664
rect 31392 43444 31444 43450
rect 31392 43386 31444 43392
rect 31680 43382 31708 43658
rect 31760 43648 31812 43654
rect 31760 43590 31812 43596
rect 31668 43376 31720 43382
rect 31668 43318 31720 43324
rect 31680 42294 31708 43318
rect 31772 42362 31800 43590
rect 31852 43240 31904 43246
rect 31852 43182 31904 43188
rect 31760 42356 31812 42362
rect 31760 42298 31812 42304
rect 31668 42288 31720 42294
rect 31668 42230 31720 42236
rect 31300 42152 31352 42158
rect 31300 42094 31352 42100
rect 31312 41614 31340 42094
rect 31392 42084 31444 42090
rect 31392 42026 31444 42032
rect 31404 41750 31432 42026
rect 31680 42022 31708 42230
rect 31864 42022 31892 43182
rect 31668 42016 31720 42022
rect 31668 41958 31720 41964
rect 31852 42016 31904 42022
rect 31852 41958 31904 41964
rect 31680 41818 31708 41958
rect 31668 41812 31720 41818
rect 31668 41754 31720 41760
rect 31392 41744 31444 41750
rect 31392 41686 31444 41692
rect 31300 41608 31352 41614
rect 31300 41550 31352 41556
rect 31208 41540 31260 41546
rect 31208 41482 31260 41488
rect 30840 41200 30892 41206
rect 30840 41142 30892 41148
rect 30746 40080 30802 40089
rect 30746 40015 30802 40024
rect 30748 39296 30800 39302
rect 30748 39238 30800 39244
rect 30656 34740 30708 34746
rect 30656 34682 30708 34688
rect 30564 34672 30616 34678
rect 30564 34614 30616 34620
rect 30760 34542 30788 39238
rect 30852 37126 30880 41142
rect 30944 40730 31064 40746
rect 30944 40724 31076 40730
rect 30944 40718 31024 40724
rect 30840 37120 30892 37126
rect 30840 37062 30892 37068
rect 30840 36712 30892 36718
rect 30840 36654 30892 36660
rect 30852 35834 30880 36654
rect 30840 35828 30892 35834
rect 30840 35770 30892 35776
rect 30748 34536 30800 34542
rect 30748 34478 30800 34484
rect 30944 34406 30972 40718
rect 31024 40666 31076 40672
rect 31024 40588 31076 40594
rect 31024 40530 31076 40536
rect 31036 39642 31064 40530
rect 31024 39636 31076 39642
rect 31024 39578 31076 39584
rect 31116 39500 31168 39506
rect 31116 39442 31168 39448
rect 31128 38758 31156 39442
rect 31116 38752 31168 38758
rect 31116 38694 31168 38700
rect 31022 36680 31078 36689
rect 31022 36615 31078 36624
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30932 34400 30984 34406
rect 30932 34342 30984 34348
rect 30576 33998 30604 34342
rect 30656 34196 30708 34202
rect 30656 34138 30708 34144
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30668 33318 30696 34138
rect 30656 33312 30708 33318
rect 30656 33254 30708 33260
rect 30564 30728 30616 30734
rect 30564 30670 30616 30676
rect 30576 30326 30604 30670
rect 30668 30326 30696 33254
rect 30564 30320 30616 30326
rect 30564 30262 30616 30268
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30668 30161 30696 30262
rect 31036 30190 31064 36615
rect 31128 35154 31156 38694
rect 31220 37330 31248 41482
rect 31312 40050 31340 41550
rect 31680 40458 31708 41754
rect 31668 40452 31720 40458
rect 31668 40394 31720 40400
rect 31680 40186 31708 40394
rect 31668 40180 31720 40186
rect 31668 40122 31720 40128
rect 31300 40044 31352 40050
rect 31300 39986 31352 39992
rect 31312 37942 31340 39986
rect 31576 39840 31628 39846
rect 31576 39782 31628 39788
rect 31484 39636 31536 39642
rect 31484 39578 31536 39584
rect 31300 37936 31352 37942
rect 31300 37878 31352 37884
rect 31300 37664 31352 37670
rect 31300 37606 31352 37612
rect 31392 37664 31444 37670
rect 31392 37606 31444 37612
rect 31208 37324 31260 37330
rect 31208 37266 31260 37272
rect 31312 37262 31340 37606
rect 31300 37256 31352 37262
rect 31300 37198 31352 37204
rect 31404 36786 31432 37606
rect 31496 37330 31524 39578
rect 31588 39574 31616 39782
rect 31576 39568 31628 39574
rect 31576 39510 31628 39516
rect 31576 39432 31628 39438
rect 31680 39386 31708 40122
rect 31628 39380 31708 39386
rect 31576 39374 31708 39380
rect 31588 39358 31708 39374
rect 31576 38820 31628 38826
rect 31576 38762 31628 38768
rect 31588 38282 31616 38762
rect 31864 38486 31892 41958
rect 31944 41268 31996 41274
rect 31944 41210 31996 41216
rect 31852 38480 31904 38486
rect 31852 38422 31904 38428
rect 31668 38344 31720 38350
rect 31668 38286 31720 38292
rect 31576 38276 31628 38282
rect 31576 38218 31628 38224
rect 31484 37324 31536 37330
rect 31484 37266 31536 37272
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 31392 36780 31444 36786
rect 31392 36722 31444 36728
rect 31116 35148 31168 35154
rect 31116 35090 31168 35096
rect 31496 34898 31524 37062
rect 31588 35630 31616 38218
rect 31680 37942 31708 38286
rect 31668 37936 31720 37942
rect 31668 37878 31720 37884
rect 31956 37194 31984 41210
rect 32048 37262 32076 43930
rect 32312 43784 32364 43790
rect 32312 43726 32364 43732
rect 32324 43450 32352 43726
rect 32312 43444 32364 43450
rect 32312 43386 32364 43392
rect 32324 43314 32352 43386
rect 32312 43308 32364 43314
rect 32312 43250 32364 43256
rect 32312 41064 32364 41070
rect 32312 41006 32364 41012
rect 32324 40050 32352 41006
rect 32312 40044 32364 40050
rect 32312 39986 32364 39992
rect 32220 39568 32272 39574
rect 32220 39510 32272 39516
rect 32232 39098 32260 39510
rect 32416 39250 32444 44746
rect 32496 42084 32548 42090
rect 32496 42026 32548 42032
rect 32324 39222 32444 39250
rect 32220 39092 32272 39098
rect 32220 39034 32272 39040
rect 32220 38276 32272 38282
rect 32220 38218 32272 38224
rect 32036 37256 32088 37262
rect 32036 37198 32088 37204
rect 31944 37188 31996 37194
rect 31944 37130 31996 37136
rect 31760 36780 31812 36786
rect 31760 36722 31812 36728
rect 31772 36174 31800 36722
rect 32128 36644 32180 36650
rect 32128 36586 32180 36592
rect 32140 36378 32168 36586
rect 32128 36372 32180 36378
rect 32128 36314 32180 36320
rect 31760 36168 31812 36174
rect 31760 36110 31812 36116
rect 31576 35624 31628 35630
rect 31576 35566 31628 35572
rect 31312 34870 31524 34898
rect 31116 33856 31168 33862
rect 31116 33798 31168 33804
rect 31208 33856 31260 33862
rect 31208 33798 31260 33804
rect 31128 33522 31156 33798
rect 31116 33516 31168 33522
rect 31116 33458 31168 33464
rect 31024 30184 31076 30190
rect 30654 30152 30710 30161
rect 30760 30122 30972 30138
rect 31024 30126 31076 30132
rect 30654 30087 30710 30096
rect 30748 30116 30984 30122
rect 30800 30110 30932 30116
rect 30748 30058 30800 30064
rect 30932 30058 30984 30064
rect 31220 29306 31248 33798
rect 31312 32978 31340 34870
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 31300 32972 31352 32978
rect 31300 32914 31352 32920
rect 31300 32768 31352 32774
rect 31300 32710 31352 32716
rect 31312 32570 31340 32710
rect 31300 32564 31352 32570
rect 31300 32506 31352 32512
rect 31404 31754 31432 34682
rect 31588 34105 31616 35566
rect 32232 35154 32260 38218
rect 31668 35148 31720 35154
rect 31668 35090 31720 35096
rect 32220 35148 32272 35154
rect 32220 35090 32272 35096
rect 31574 34096 31630 34105
rect 31574 34031 31630 34040
rect 31484 33108 31536 33114
rect 31484 33050 31536 33056
rect 31496 32978 31524 33050
rect 31484 32972 31536 32978
rect 31484 32914 31536 32920
rect 31680 31958 31708 35090
rect 32324 32910 32352 39222
rect 32404 39092 32456 39098
rect 32404 39034 32456 39040
rect 32416 36922 32444 39034
rect 32508 37670 32536 42026
rect 32588 41132 32640 41138
rect 32588 41074 32640 41080
rect 32600 39642 32628 41074
rect 32692 40594 32720 45222
rect 32876 43874 32904 45358
rect 33508 45280 33560 45286
rect 33508 45222 33560 45228
rect 32950 45180 33258 45189
rect 32950 45178 32956 45180
rect 33012 45178 33036 45180
rect 33092 45178 33116 45180
rect 33172 45178 33196 45180
rect 33252 45178 33258 45180
rect 33012 45126 33014 45178
rect 33194 45126 33196 45178
rect 32950 45124 32956 45126
rect 33012 45124 33036 45126
rect 33092 45124 33116 45126
rect 33172 45124 33196 45126
rect 33252 45124 33258 45126
rect 32950 45115 33258 45124
rect 32950 44092 33258 44101
rect 32950 44090 32956 44092
rect 33012 44090 33036 44092
rect 33092 44090 33116 44092
rect 33172 44090 33196 44092
rect 33252 44090 33258 44092
rect 33012 44038 33014 44090
rect 33194 44038 33196 44090
rect 32950 44036 32956 44038
rect 33012 44036 33036 44038
rect 33092 44036 33116 44038
rect 33172 44036 33196 44038
rect 33252 44036 33258 44038
rect 32950 44027 33258 44036
rect 32876 43858 32996 43874
rect 32876 43852 33008 43858
rect 32876 43846 32956 43852
rect 32956 43794 33008 43800
rect 33324 43648 33376 43654
rect 33324 43590 33376 43596
rect 33416 43648 33468 43654
rect 33416 43590 33468 43596
rect 32950 43004 33258 43013
rect 32950 43002 32956 43004
rect 33012 43002 33036 43004
rect 33092 43002 33116 43004
rect 33172 43002 33196 43004
rect 33252 43002 33258 43004
rect 33012 42950 33014 43002
rect 33194 42950 33196 43002
rect 32950 42948 32956 42950
rect 33012 42948 33036 42950
rect 33092 42948 33116 42950
rect 33172 42948 33196 42950
rect 33252 42948 33258 42950
rect 32950 42939 33258 42948
rect 32772 42356 32824 42362
rect 32772 42298 32824 42304
rect 32784 40594 32812 42298
rect 32950 41916 33258 41925
rect 32950 41914 32956 41916
rect 33012 41914 33036 41916
rect 33092 41914 33116 41916
rect 33172 41914 33196 41916
rect 33252 41914 33258 41916
rect 33012 41862 33014 41914
rect 33194 41862 33196 41914
rect 32950 41860 32956 41862
rect 33012 41860 33036 41862
rect 33092 41860 33116 41862
rect 33172 41860 33196 41862
rect 33252 41860 33258 41862
rect 32950 41851 33258 41860
rect 33048 41812 33100 41818
rect 33048 41754 33100 41760
rect 33060 41614 33088 41754
rect 33048 41608 33100 41614
rect 33048 41550 33100 41556
rect 32864 41200 32916 41206
rect 32864 41142 32916 41148
rect 32680 40588 32732 40594
rect 32680 40530 32732 40536
rect 32772 40588 32824 40594
rect 32772 40530 32824 40536
rect 32876 40474 32904 41142
rect 33060 40934 33088 41550
rect 33336 41478 33364 43590
rect 33324 41472 33376 41478
rect 33324 41414 33376 41420
rect 33048 40928 33100 40934
rect 33048 40870 33100 40876
rect 32950 40828 33258 40837
rect 32950 40826 32956 40828
rect 33012 40826 33036 40828
rect 33092 40826 33116 40828
rect 33172 40826 33196 40828
rect 33252 40826 33258 40828
rect 33012 40774 33014 40826
rect 33194 40774 33196 40826
rect 32950 40772 32956 40774
rect 33012 40772 33036 40774
rect 33092 40772 33116 40774
rect 33172 40772 33196 40774
rect 33252 40772 33258 40774
rect 32950 40763 33258 40772
rect 32784 40446 32904 40474
rect 33324 40452 33376 40458
rect 32784 40186 32812 40446
rect 33324 40394 33376 40400
rect 32772 40180 32824 40186
rect 32772 40122 32824 40128
rect 32588 39636 32640 39642
rect 32588 39578 32640 39584
rect 32588 38956 32640 38962
rect 32588 38898 32640 38904
rect 32496 37664 32548 37670
rect 32496 37606 32548 37612
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 32508 36281 32536 37062
rect 32494 36272 32550 36281
rect 32494 36207 32550 36216
rect 32508 34116 32536 36207
rect 32416 34088 32536 34116
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 32312 32904 32364 32910
rect 32312 32846 32364 32852
rect 31668 31952 31720 31958
rect 31668 31894 31720 31900
rect 31772 31890 31800 32846
rect 32220 32768 32272 32774
rect 32220 32710 32272 32716
rect 31944 32360 31996 32366
rect 31944 32302 31996 32308
rect 31760 31884 31812 31890
rect 31760 31826 31812 31832
rect 31404 31726 31524 31754
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31312 29306 31340 29446
rect 31208 29300 31260 29306
rect 31208 29242 31260 29248
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 30380 28688 30432 28694
rect 30380 28630 30432 28636
rect 30656 28416 30708 28422
rect 30656 28358 30708 28364
rect 31300 28416 31352 28422
rect 31300 28358 31352 28364
rect 30288 27532 30340 27538
rect 30288 27474 30340 27480
rect 30380 27464 30432 27470
rect 30208 27390 30328 27418
rect 30380 27406 30432 27412
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 30104 27056 30156 27062
rect 30104 26998 30156 27004
rect 30012 25492 30064 25498
rect 30012 25434 30064 25440
rect 30012 25356 30064 25362
rect 29932 25316 30012 25344
rect 29932 24886 29960 25316
rect 30012 25298 30064 25304
rect 29920 24880 29972 24886
rect 29920 24822 29972 24828
rect 30104 24744 30156 24750
rect 30104 24686 30156 24692
rect 29828 24132 29880 24138
rect 29828 24074 29880 24080
rect 30116 23662 30144 24686
rect 30208 24274 30236 27270
rect 30300 27130 30328 27390
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 30300 25838 30328 27066
rect 30392 26790 30420 27406
rect 30564 27328 30616 27334
rect 30564 27270 30616 27276
rect 30576 27130 30604 27270
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30564 26920 30616 26926
rect 30564 26862 30616 26868
rect 30380 26784 30432 26790
rect 30380 26726 30432 26732
rect 30472 26784 30524 26790
rect 30472 26726 30524 26732
rect 30288 25832 30340 25838
rect 30288 25774 30340 25780
rect 30196 24268 30248 24274
rect 30196 24210 30248 24216
rect 30104 23656 30156 23662
rect 30104 23598 30156 23604
rect 29918 23488 29974 23497
rect 29918 23423 29974 23432
rect 29472 22066 29684 22094
rect 29368 22024 29420 22030
rect 29368 21966 29420 21972
rect 29380 21690 29408 21966
rect 29368 21684 29420 21690
rect 29368 21626 29420 21632
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29196 18006 29316 18034
rect 29090 17983 29146 17992
rect 28828 15422 28948 15450
rect 29000 15496 29052 15502
rect 29000 15438 29052 15444
rect 28828 12617 28856 15422
rect 29104 15348 29132 17983
rect 29184 16040 29236 16046
rect 29184 15982 29236 15988
rect 29196 15434 29224 15982
rect 29184 15428 29236 15434
rect 29184 15370 29236 15376
rect 28920 15320 29132 15348
rect 28920 13410 28948 15320
rect 29196 15162 29224 15370
rect 29184 15156 29236 15162
rect 29184 15098 29236 15104
rect 29288 13938 29316 18006
rect 29472 16522 29500 22066
rect 29736 17536 29788 17542
rect 29736 17478 29788 17484
rect 29552 17128 29604 17134
rect 29552 17070 29604 17076
rect 29460 16516 29512 16522
rect 29460 16458 29512 16464
rect 29368 16176 29420 16182
rect 29420 16124 29500 16130
rect 29368 16118 29500 16124
rect 29380 16102 29500 16118
rect 29472 16046 29500 16102
rect 29460 16040 29512 16046
rect 29460 15982 29512 15988
rect 29460 15632 29512 15638
rect 29460 15574 29512 15580
rect 29472 15450 29500 15574
rect 29380 15422 29500 15450
rect 29276 13932 29328 13938
rect 29276 13874 29328 13880
rect 29380 13818 29408 15422
rect 29460 15360 29512 15366
rect 29460 15302 29512 15308
rect 29472 15094 29500 15302
rect 29460 15088 29512 15094
rect 29460 15030 29512 15036
rect 29472 14346 29500 15030
rect 29460 14340 29512 14346
rect 29460 14282 29512 14288
rect 29104 13790 29408 13818
rect 28920 13382 29040 13410
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 28814 12608 28870 12617
rect 28814 12543 28870 12552
rect 28920 12434 28948 13262
rect 28538 12407 28594 12416
rect 28552 10062 28580 12407
rect 28644 12406 28764 12434
rect 28828 12406 28948 12434
rect 28540 10056 28592 10062
rect 28540 9998 28592 10004
rect 28448 2100 28500 2106
rect 28448 2042 28500 2048
rect 28644 1902 28672 12406
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 28632 1896 28684 1902
rect 28632 1838 28684 1844
rect 28736 800 28764 2926
rect 28828 2310 28856 12406
rect 29012 12322 29040 13382
rect 28920 12294 29040 12322
rect 28920 12238 28948 12294
rect 28908 12232 28960 12238
rect 28908 12174 28960 12180
rect 29104 3058 29132 13790
rect 29276 12980 29328 12986
rect 29276 12922 29328 12928
rect 29184 12164 29236 12170
rect 29184 12106 29236 12112
rect 29196 3058 29224 12106
rect 29092 3052 29144 3058
rect 29092 2994 29144 3000
rect 29184 3052 29236 3058
rect 29184 2994 29236 3000
rect 29288 2378 29316 12922
rect 29564 12782 29592 17070
rect 29748 16250 29776 17478
rect 29736 16244 29788 16250
rect 29736 16186 29788 16192
rect 29644 15428 29696 15434
rect 29644 15370 29696 15376
rect 29656 15162 29684 15370
rect 29644 15156 29696 15162
rect 29644 15098 29696 15104
rect 29748 15042 29776 16186
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 29656 15014 29776 15042
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29656 7410 29684 15014
rect 29840 14362 29868 15846
rect 29932 15094 29960 23423
rect 30116 23186 30144 23598
rect 30104 23180 30156 23186
rect 30104 23122 30156 23128
rect 30484 22778 30512 26726
rect 30576 26450 30604 26862
rect 30668 26450 30696 28358
rect 31206 28112 31262 28121
rect 31206 28047 31262 28056
rect 30840 27872 30892 27878
rect 30840 27814 30892 27820
rect 30748 27056 30800 27062
rect 30748 26998 30800 27004
rect 30564 26444 30616 26450
rect 30564 26386 30616 26392
rect 30656 26444 30708 26450
rect 30656 26386 30708 26392
rect 30656 26240 30708 26246
rect 30656 26182 30708 26188
rect 30668 22982 30696 26182
rect 30760 25974 30788 26998
rect 30748 25968 30800 25974
rect 30748 25910 30800 25916
rect 30760 24818 30788 25910
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30852 24698 30880 27814
rect 30932 27396 30984 27402
rect 30932 27338 30984 27344
rect 30944 27305 30972 27338
rect 30930 27296 30986 27305
rect 30930 27231 30986 27240
rect 31220 27062 31248 28047
rect 31312 27062 31340 28358
rect 31496 27826 31524 31726
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31588 30394 31616 30602
rect 31576 30388 31628 30394
rect 31576 30330 31628 30336
rect 31772 29594 31800 31826
rect 31956 30802 31984 32302
rect 32128 32224 32180 32230
rect 32128 32166 32180 32172
rect 32036 31952 32088 31958
rect 32036 31894 32088 31900
rect 32048 31482 32076 31894
rect 32036 31476 32088 31482
rect 32036 31418 32088 31424
rect 32036 31272 32088 31278
rect 32036 31214 32088 31220
rect 31944 30796 31996 30802
rect 31944 30738 31996 30744
rect 31944 29776 31996 29782
rect 31944 29718 31996 29724
rect 31772 29566 31892 29594
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31576 27940 31628 27946
rect 31576 27882 31628 27888
rect 31588 27826 31616 27882
rect 31496 27798 31616 27826
rect 31392 27124 31444 27130
rect 31392 27066 31444 27072
rect 31208 27056 31260 27062
rect 31300 27056 31352 27062
rect 31208 26998 31260 27004
rect 31298 27024 31300 27033
rect 31352 27024 31354 27033
rect 31116 26852 31168 26858
rect 31116 26794 31168 26800
rect 31024 26512 31076 26518
rect 31024 26454 31076 26460
rect 31036 26353 31064 26454
rect 31022 26344 31078 26353
rect 31022 26279 31078 26288
rect 30932 25696 30984 25702
rect 30932 25638 30984 25644
rect 30944 24954 30972 25638
rect 30932 24948 30984 24954
rect 30932 24890 30984 24896
rect 31128 24750 31156 26794
rect 30760 24670 30880 24698
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 30656 22976 30708 22982
rect 30656 22918 30708 22924
rect 30472 22772 30524 22778
rect 30472 22714 30524 22720
rect 30380 22704 30432 22710
rect 30378 22672 30380 22681
rect 30432 22672 30434 22681
rect 30378 22607 30434 22616
rect 30656 21344 30708 21350
rect 30656 21286 30708 21292
rect 30668 20942 30696 21286
rect 30760 21146 30788 24670
rect 30840 24132 30892 24138
rect 30840 24074 30892 24080
rect 30852 23866 30880 24074
rect 30840 23860 30892 23866
rect 30840 23802 30892 23808
rect 31128 23322 31156 24686
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 30656 20936 30708 20942
rect 30656 20878 30708 20884
rect 30748 20936 30800 20942
rect 30748 20878 30800 20884
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 30012 18216 30064 18222
rect 30012 18158 30064 18164
rect 30024 17746 30052 18158
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30024 17134 30052 17682
rect 30300 17610 30328 20742
rect 30470 20632 30526 20641
rect 30470 20567 30472 20576
rect 30524 20567 30526 20576
rect 30472 20538 30524 20544
rect 30760 20534 30788 20878
rect 30748 20528 30800 20534
rect 30748 20470 30800 20476
rect 31220 18290 31248 26998
rect 31298 26959 31354 26968
rect 31300 25152 31352 25158
rect 31300 25094 31352 25100
rect 31312 20806 31340 25094
rect 31300 20800 31352 20806
rect 31300 20742 31352 20748
rect 31404 18834 31432 27066
rect 31496 23798 31524 27798
rect 31668 27464 31720 27470
rect 31574 27432 31630 27441
rect 31668 27406 31720 27412
rect 31574 27367 31630 27376
rect 31588 26994 31616 27367
rect 31576 26988 31628 26994
rect 31576 26930 31628 26936
rect 31680 26450 31708 27406
rect 31668 26444 31720 26450
rect 31668 26386 31720 26392
rect 31668 25424 31720 25430
rect 31668 25366 31720 25372
rect 31576 24676 31628 24682
rect 31576 24618 31628 24624
rect 31484 23792 31536 23798
rect 31484 23734 31536 23740
rect 31484 23588 31536 23594
rect 31484 23530 31536 23536
rect 31392 18828 31444 18834
rect 31392 18770 31444 18776
rect 31208 18284 31260 18290
rect 31208 18226 31260 18232
rect 30380 18216 30432 18222
rect 30380 18158 30432 18164
rect 30288 17604 30340 17610
rect 30288 17546 30340 17552
rect 30392 17490 30420 18158
rect 30932 17604 30984 17610
rect 30932 17546 30984 17552
rect 30300 17462 30420 17490
rect 30564 17536 30616 17542
rect 30564 17478 30616 17484
rect 30300 17134 30328 17462
rect 30576 17270 30604 17478
rect 30564 17264 30616 17270
rect 30484 17212 30564 17218
rect 30484 17206 30616 17212
rect 30484 17190 30604 17206
rect 30012 17128 30064 17134
rect 30012 17070 30064 17076
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30024 15570 30052 17070
rect 30196 15972 30248 15978
rect 30196 15914 30248 15920
rect 30104 15904 30156 15910
rect 30104 15846 30156 15852
rect 30012 15564 30064 15570
rect 30012 15506 30064 15512
rect 30116 15434 30144 15846
rect 30208 15706 30236 15914
rect 30196 15700 30248 15706
rect 30196 15642 30248 15648
rect 30104 15428 30156 15434
rect 30104 15370 30156 15376
rect 30300 15366 30328 17070
rect 30484 16998 30512 17190
rect 30944 17134 30972 17546
rect 30932 17128 30984 17134
rect 30932 17070 30984 17076
rect 30472 16992 30524 16998
rect 30472 16934 30524 16940
rect 30484 16182 30512 16934
rect 30564 16584 30616 16590
rect 30564 16526 30616 16532
rect 30472 16176 30524 16182
rect 30472 16118 30524 16124
rect 30484 15434 30512 16118
rect 30472 15428 30524 15434
rect 30472 15370 30524 15376
rect 30288 15360 30340 15366
rect 30288 15302 30340 15308
rect 29920 15088 29972 15094
rect 29920 15030 29972 15036
rect 30012 14816 30064 14822
rect 30012 14758 30064 14764
rect 30196 14816 30248 14822
rect 30196 14758 30248 14764
rect 29840 14334 29960 14362
rect 29932 14278 29960 14334
rect 29920 14272 29972 14278
rect 29920 14214 29972 14220
rect 29736 13864 29788 13870
rect 29736 13806 29788 13812
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29460 5024 29512 5030
rect 29460 4966 29512 4972
rect 29472 4826 29500 4966
rect 29460 4820 29512 4826
rect 29460 4762 29512 4768
rect 29460 3596 29512 3602
rect 29460 3538 29512 3544
rect 29276 2372 29328 2378
rect 29276 2314 29328 2320
rect 28816 2304 28868 2310
rect 28816 2246 28868 2252
rect 29472 800 29500 3538
rect 29748 3534 29776 13806
rect 30024 12714 30052 14758
rect 30208 14414 30236 14758
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30288 14408 30340 14414
rect 30288 14350 30340 14356
rect 30300 12986 30328 14350
rect 30576 12986 30604 16526
rect 31496 15094 31524 23530
rect 31588 23186 31616 24618
rect 31576 23180 31628 23186
rect 31576 23122 31628 23128
rect 31588 21622 31616 23122
rect 31680 21894 31708 25366
rect 31772 25294 31800 29446
rect 31864 27452 31892 29566
rect 31956 28694 31984 29718
rect 31944 28688 31996 28694
rect 31944 28630 31996 28636
rect 32048 28098 32076 31214
rect 32140 28218 32168 32166
rect 32232 29578 32260 32710
rect 32416 31278 32444 34088
rect 32600 31754 32628 38898
rect 32680 37664 32732 37670
rect 32680 37606 32732 37612
rect 32692 36242 32720 37606
rect 32784 37210 32812 40122
rect 32950 39740 33258 39749
rect 32950 39738 32956 39740
rect 33012 39738 33036 39740
rect 33092 39738 33116 39740
rect 33172 39738 33196 39740
rect 33252 39738 33258 39740
rect 33012 39686 33014 39738
rect 33194 39686 33196 39738
rect 32950 39684 32956 39686
rect 33012 39684 33036 39686
rect 33092 39684 33116 39686
rect 33172 39684 33196 39686
rect 33252 39684 33258 39686
rect 32950 39675 33258 39684
rect 32950 38652 33258 38661
rect 32950 38650 32956 38652
rect 33012 38650 33036 38652
rect 33092 38650 33116 38652
rect 33172 38650 33196 38652
rect 33252 38650 33258 38652
rect 33012 38598 33014 38650
rect 33194 38598 33196 38650
rect 32950 38596 32956 38598
rect 33012 38596 33036 38598
rect 33092 38596 33116 38598
rect 33172 38596 33196 38598
rect 33252 38596 33258 38598
rect 32950 38587 33258 38596
rect 33336 38418 33364 40394
rect 33324 38412 33376 38418
rect 33324 38354 33376 38360
rect 33232 38208 33284 38214
rect 33232 38150 33284 38156
rect 32864 38004 32916 38010
rect 32864 37946 32916 37952
rect 32876 37330 32904 37946
rect 32956 37800 33008 37806
rect 33244 37777 33272 38150
rect 32956 37742 33008 37748
rect 33230 37768 33286 37777
rect 32968 37670 32996 37742
rect 33230 37703 33286 37712
rect 32956 37664 33008 37670
rect 32956 37606 33008 37612
rect 32950 37564 33258 37573
rect 32950 37562 32956 37564
rect 33012 37562 33036 37564
rect 33092 37562 33116 37564
rect 33172 37562 33196 37564
rect 33252 37562 33258 37564
rect 33012 37510 33014 37562
rect 33194 37510 33196 37562
rect 32950 37508 32956 37510
rect 33012 37508 33036 37510
rect 33092 37508 33116 37510
rect 33172 37508 33196 37510
rect 33252 37508 33258 37510
rect 32950 37499 33258 37508
rect 32864 37324 32916 37330
rect 32864 37266 32916 37272
rect 32784 37182 32904 37210
rect 32680 36236 32732 36242
rect 32680 36178 32732 36184
rect 32876 35630 32904 37182
rect 32950 36476 33258 36485
rect 32950 36474 32956 36476
rect 33012 36474 33036 36476
rect 33092 36474 33116 36476
rect 33172 36474 33196 36476
rect 33252 36474 33258 36476
rect 33012 36422 33014 36474
rect 33194 36422 33196 36474
rect 32950 36420 32956 36422
rect 33012 36420 33036 36422
rect 33092 36420 33116 36422
rect 33172 36420 33196 36422
rect 33252 36420 33258 36422
rect 32950 36411 33258 36420
rect 33140 36100 33192 36106
rect 33140 36042 33192 36048
rect 33152 35834 33180 36042
rect 33140 35828 33192 35834
rect 33140 35770 33192 35776
rect 32772 35624 32824 35630
rect 32770 35592 32772 35601
rect 32864 35624 32916 35630
rect 32824 35592 32826 35601
rect 32864 35566 32916 35572
rect 32770 35527 32826 35536
rect 32950 35388 33258 35397
rect 32950 35386 32956 35388
rect 33012 35386 33036 35388
rect 33092 35386 33116 35388
rect 33172 35386 33196 35388
rect 33252 35386 33258 35388
rect 33012 35334 33014 35386
rect 33194 35334 33196 35386
rect 32950 35332 32956 35334
rect 33012 35332 33036 35334
rect 33092 35332 33116 35334
rect 33172 35332 33196 35334
rect 33252 35332 33258 35334
rect 32950 35323 33258 35332
rect 32680 34604 32732 34610
rect 32680 34546 32732 34552
rect 32692 34202 32720 34546
rect 32950 34300 33258 34309
rect 32950 34298 32956 34300
rect 33012 34298 33036 34300
rect 33092 34298 33116 34300
rect 33172 34298 33196 34300
rect 33252 34298 33258 34300
rect 33012 34246 33014 34298
rect 33194 34246 33196 34298
rect 32950 34244 32956 34246
rect 33012 34244 33036 34246
rect 33092 34244 33116 34246
rect 33172 34244 33196 34246
rect 33252 34244 33258 34246
rect 32950 34235 33258 34244
rect 32680 34196 32732 34202
rect 32680 34138 32732 34144
rect 32950 33212 33258 33221
rect 32950 33210 32956 33212
rect 33012 33210 33036 33212
rect 33092 33210 33116 33212
rect 33172 33210 33196 33212
rect 33252 33210 33258 33212
rect 33012 33158 33014 33210
rect 33194 33158 33196 33210
rect 32950 33156 32956 33158
rect 33012 33156 33036 33158
rect 33092 33156 33116 33158
rect 33172 33156 33196 33158
rect 33252 33156 33258 33158
rect 32950 33147 33258 33156
rect 32950 32124 33258 32133
rect 32950 32122 32956 32124
rect 33012 32122 33036 32124
rect 33092 32122 33116 32124
rect 33172 32122 33196 32124
rect 33252 32122 33258 32124
rect 33012 32070 33014 32122
rect 33194 32070 33196 32122
rect 32950 32068 32956 32070
rect 33012 32068 33036 32070
rect 33092 32068 33116 32070
rect 33172 32068 33196 32070
rect 33252 32068 33258 32070
rect 32950 32059 33258 32068
rect 32508 31726 32628 31754
rect 32404 31272 32456 31278
rect 32404 31214 32456 31220
rect 32312 30796 32364 30802
rect 32312 30738 32364 30744
rect 32220 29572 32272 29578
rect 32220 29514 32272 29520
rect 32324 28966 32352 30738
rect 32404 29504 32456 29510
rect 32404 29446 32456 29452
rect 32416 29306 32444 29446
rect 32404 29300 32456 29306
rect 32404 29242 32456 29248
rect 32312 28960 32364 28966
rect 32312 28902 32364 28908
rect 32220 28484 32272 28490
rect 32220 28426 32272 28432
rect 32128 28212 32180 28218
rect 32128 28154 32180 28160
rect 32048 28070 32168 28098
rect 31864 27424 32076 27452
rect 31944 27328 31996 27334
rect 31944 27270 31996 27276
rect 31852 25356 31904 25362
rect 31852 25298 31904 25304
rect 31760 25288 31812 25294
rect 31760 25230 31812 25236
rect 31864 23322 31892 25298
rect 31956 25294 31984 27270
rect 31944 25288 31996 25294
rect 31944 25230 31996 25236
rect 32048 23594 32076 27424
rect 32140 26353 32168 28070
rect 32232 27946 32260 28426
rect 32324 28082 32352 28902
rect 32404 28212 32456 28218
rect 32404 28154 32456 28160
rect 32312 28076 32364 28082
rect 32312 28018 32364 28024
rect 32220 27940 32272 27946
rect 32220 27882 32272 27888
rect 32220 27532 32272 27538
rect 32220 27474 32272 27480
rect 32126 26344 32182 26353
rect 32126 26279 32182 26288
rect 32232 25378 32260 27474
rect 32324 26314 32352 28018
rect 32416 26314 32444 28154
rect 32508 27130 32536 31726
rect 32680 31272 32732 31278
rect 32680 31214 32732 31220
rect 32588 30864 32640 30870
rect 32588 30806 32640 30812
rect 32600 27878 32628 30806
rect 32692 29782 32720 31214
rect 32864 31136 32916 31142
rect 32864 31078 32916 31084
rect 32772 30116 32824 30122
rect 32772 30058 32824 30064
rect 32680 29776 32732 29782
rect 32680 29718 32732 29724
rect 32680 29572 32732 29578
rect 32680 29514 32732 29520
rect 32588 27872 32640 27878
rect 32588 27814 32640 27820
rect 32692 27130 32720 29514
rect 32784 28506 32812 30058
rect 32876 28626 32904 31078
rect 32950 31036 33258 31045
rect 32950 31034 32956 31036
rect 33012 31034 33036 31036
rect 33092 31034 33116 31036
rect 33172 31034 33196 31036
rect 33252 31034 33258 31036
rect 33012 30982 33014 31034
rect 33194 30982 33196 31034
rect 32950 30980 32956 30982
rect 33012 30980 33036 30982
rect 33092 30980 33116 30982
rect 33172 30980 33196 30982
rect 33252 30980 33258 30982
rect 32950 30971 33258 30980
rect 33324 30728 33376 30734
rect 33324 30670 33376 30676
rect 32950 29948 33258 29957
rect 32950 29946 32956 29948
rect 33012 29946 33036 29948
rect 33092 29946 33116 29948
rect 33172 29946 33196 29948
rect 33252 29946 33258 29948
rect 33012 29894 33014 29946
rect 33194 29894 33196 29946
rect 32950 29892 32956 29894
rect 33012 29892 33036 29894
rect 33092 29892 33116 29894
rect 33172 29892 33196 29894
rect 33252 29892 33258 29894
rect 32950 29883 33258 29892
rect 32950 28860 33258 28869
rect 32950 28858 32956 28860
rect 33012 28858 33036 28860
rect 33092 28858 33116 28860
rect 33172 28858 33196 28860
rect 33252 28858 33258 28860
rect 33012 28806 33014 28858
rect 33194 28806 33196 28858
rect 32950 28804 32956 28806
rect 33012 28804 33036 28806
rect 33092 28804 33116 28806
rect 33172 28804 33196 28806
rect 33252 28804 33258 28806
rect 32950 28795 33258 28804
rect 33336 28762 33364 30670
rect 33428 30326 33456 43590
rect 33520 40594 33548 45222
rect 33600 43716 33652 43722
rect 33600 43658 33652 43664
rect 33612 43314 33640 43658
rect 33600 43308 33652 43314
rect 33600 43250 33652 43256
rect 33600 40928 33652 40934
rect 33600 40870 33652 40876
rect 33508 40588 33560 40594
rect 33508 40530 33560 40536
rect 33612 40118 33640 40870
rect 33600 40112 33652 40118
rect 33600 40054 33652 40060
rect 33600 39296 33652 39302
rect 33600 39238 33652 39244
rect 33612 39098 33640 39238
rect 33600 39092 33652 39098
rect 33600 39034 33652 39040
rect 33508 37868 33560 37874
rect 33508 37810 33560 37816
rect 33520 37194 33548 37810
rect 33508 37188 33560 37194
rect 33508 37130 33560 37136
rect 33704 36530 33732 45526
rect 33968 45552 34284 45554
rect 34020 45526 34284 45552
rect 33968 45494 34020 45500
rect 34152 45416 34204 45422
rect 34152 45358 34204 45364
rect 34164 43178 34192 45358
rect 34152 43172 34204 43178
rect 34152 43114 34204 43120
rect 34060 43104 34112 43110
rect 34060 43046 34112 43052
rect 34072 41698 34100 43046
rect 34072 41682 34192 41698
rect 34072 41676 34204 41682
rect 34072 41670 34152 41676
rect 34152 41618 34204 41624
rect 34060 41472 34112 41478
rect 34060 41414 34112 41420
rect 33966 40488 34022 40497
rect 33966 40423 33968 40432
rect 34020 40423 34022 40432
rect 33968 40394 34020 40400
rect 33876 40384 33928 40390
rect 33876 40326 33928 40332
rect 33784 39908 33836 39914
rect 33784 39850 33836 39856
rect 33520 36502 33732 36530
rect 33416 30320 33468 30326
rect 33416 30262 33468 30268
rect 33416 29028 33468 29034
rect 33416 28970 33468 28976
rect 33324 28756 33376 28762
rect 33324 28698 33376 28704
rect 32956 28688 33008 28694
rect 32956 28630 33008 28636
rect 32864 28620 32916 28626
rect 32864 28562 32916 28568
rect 32784 28478 32904 28506
rect 32772 28416 32824 28422
rect 32772 28358 32824 28364
rect 32496 27124 32548 27130
rect 32496 27066 32548 27072
rect 32680 27124 32732 27130
rect 32680 27066 32732 27072
rect 32588 26580 32640 26586
rect 32588 26522 32640 26528
rect 32312 26308 32364 26314
rect 32312 26250 32364 26256
rect 32404 26308 32456 26314
rect 32404 26250 32456 26256
rect 32416 25838 32444 26250
rect 32404 25832 32456 25838
rect 32404 25774 32456 25780
rect 32140 25350 32260 25378
rect 32036 23588 32088 23594
rect 32036 23530 32088 23536
rect 31852 23316 31904 23322
rect 31852 23258 31904 23264
rect 31760 23044 31812 23050
rect 31760 22986 31812 22992
rect 31668 21888 31720 21894
rect 31668 21830 31720 21836
rect 31576 21616 31628 21622
rect 31576 21558 31628 21564
rect 31772 21486 31800 22986
rect 31864 21554 31892 23258
rect 32140 23254 32168 25350
rect 32220 25220 32272 25226
rect 32220 25162 32272 25168
rect 32232 24886 32260 25162
rect 32220 24880 32272 24886
rect 32220 24822 32272 24828
rect 32600 24750 32628 26522
rect 32784 26194 32812 28358
rect 32876 27384 32904 28478
rect 32968 28014 32996 28630
rect 32956 28008 33008 28014
rect 32956 27950 33008 27956
rect 33324 28008 33376 28014
rect 33324 27950 33376 27956
rect 32950 27772 33258 27781
rect 32950 27770 32956 27772
rect 33012 27770 33036 27772
rect 33092 27770 33116 27772
rect 33172 27770 33196 27772
rect 33252 27770 33258 27772
rect 33012 27718 33014 27770
rect 33194 27718 33196 27770
rect 32950 27716 32956 27718
rect 33012 27716 33036 27718
rect 33092 27716 33116 27718
rect 33172 27716 33196 27718
rect 33252 27716 33258 27718
rect 32950 27707 33258 27716
rect 32956 27396 33008 27402
rect 32876 27356 32956 27384
rect 32876 26296 32904 27356
rect 32956 27338 33008 27344
rect 32950 26684 33258 26693
rect 32950 26682 32956 26684
rect 33012 26682 33036 26684
rect 33092 26682 33116 26684
rect 33172 26682 33196 26684
rect 33252 26682 33258 26684
rect 33012 26630 33014 26682
rect 33194 26630 33196 26682
rect 32950 26628 32956 26630
rect 33012 26628 33036 26630
rect 33092 26628 33116 26630
rect 33172 26628 33196 26630
rect 33252 26628 33258 26630
rect 32950 26619 33258 26628
rect 32876 26268 32996 26296
rect 32784 26166 32904 26194
rect 32680 26036 32732 26042
rect 32680 25978 32732 25984
rect 32692 25401 32720 25978
rect 32678 25392 32734 25401
rect 32678 25327 32734 25336
rect 32772 25152 32824 25158
rect 32772 25094 32824 25100
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32404 24608 32456 24614
rect 32404 24550 32456 24556
rect 32220 24336 32272 24342
rect 32220 24278 32272 24284
rect 32232 23526 32260 24278
rect 32312 23656 32364 23662
rect 32312 23598 32364 23604
rect 32220 23520 32272 23526
rect 32220 23462 32272 23468
rect 32128 23248 32180 23254
rect 32128 23190 32180 23196
rect 32140 22234 32168 23190
rect 32324 23186 32352 23598
rect 32312 23180 32364 23186
rect 32312 23122 32364 23128
rect 32312 22432 32364 22438
rect 32312 22374 32364 22380
rect 32128 22228 32180 22234
rect 32128 22170 32180 22176
rect 32140 22094 32168 22170
rect 32048 22066 32168 22094
rect 31852 21548 31904 21554
rect 31852 21490 31904 21496
rect 31760 21480 31812 21486
rect 31760 21422 31812 21428
rect 31772 21010 31800 21422
rect 31760 21004 31812 21010
rect 31760 20946 31812 20952
rect 31944 20800 31996 20806
rect 31944 20742 31996 20748
rect 31852 19984 31904 19990
rect 31852 19926 31904 19932
rect 31576 16516 31628 16522
rect 31576 16458 31628 16464
rect 31588 15366 31616 16458
rect 31576 15360 31628 15366
rect 31576 15302 31628 15308
rect 31760 15360 31812 15366
rect 31760 15302 31812 15308
rect 31484 15088 31536 15094
rect 31484 15030 31536 15036
rect 31772 14482 31800 15302
rect 31760 14476 31812 14482
rect 31760 14418 31812 14424
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 30288 12980 30340 12986
rect 30288 12922 30340 12928
rect 30564 12980 30616 12986
rect 30564 12922 30616 12928
rect 30012 12708 30064 12714
rect 30012 12650 30064 12656
rect 30104 9988 30156 9994
rect 30104 9930 30156 9936
rect 29920 9920 29972 9926
rect 29920 9862 29972 9868
rect 29736 3528 29788 3534
rect 29736 3470 29788 3476
rect 29932 2446 29960 9862
rect 30116 3534 30144 9930
rect 30104 3528 30156 3534
rect 30104 3470 30156 3476
rect 30576 3194 30604 12922
rect 31772 7478 31800 13126
rect 31864 10062 31892 19926
rect 31956 17338 31984 20742
rect 32048 19922 32076 22066
rect 32220 21480 32272 21486
rect 32220 21422 32272 21428
rect 32232 20398 32260 21422
rect 32220 20392 32272 20398
rect 32220 20334 32272 20340
rect 32036 19916 32088 19922
rect 32036 19858 32088 19864
rect 32324 19854 32352 22374
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32036 19780 32088 19786
rect 32036 19722 32088 19728
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31852 10056 31904 10062
rect 31852 9998 31904 10004
rect 31956 9654 31984 17274
rect 31944 9648 31996 9654
rect 31944 9590 31996 9596
rect 31760 7472 31812 7478
rect 31760 7414 31812 7420
rect 30932 3596 30984 3602
rect 30932 3538 30984 3544
rect 30564 3188 30616 3194
rect 30564 3130 30616 3136
rect 30288 2508 30340 2514
rect 30208 2468 30288 2496
rect 29920 2440 29972 2446
rect 29920 2382 29972 2388
rect 30208 800 30236 2468
rect 30288 2450 30340 2456
rect 30944 800 30972 3538
rect 32048 3058 32076 19722
rect 32312 19712 32364 19718
rect 32312 19654 32364 19660
rect 32324 18358 32352 19654
rect 32312 18352 32364 18358
rect 32312 18294 32364 18300
rect 32324 17082 32352 18294
rect 32416 17202 32444 24550
rect 32588 23860 32640 23866
rect 32588 23802 32640 23808
rect 32600 22574 32628 23802
rect 32680 23656 32732 23662
rect 32680 23598 32732 23604
rect 32692 22778 32720 23598
rect 32680 22772 32732 22778
rect 32680 22714 32732 22720
rect 32588 22568 32640 22574
rect 32588 22510 32640 22516
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32508 21690 32536 21966
rect 32496 21684 32548 21690
rect 32496 21626 32548 21632
rect 32508 21554 32536 21626
rect 32496 21548 32548 21554
rect 32496 21490 32548 21496
rect 32784 20584 32812 25094
rect 32876 24818 32904 26166
rect 32968 25974 32996 26268
rect 32956 25968 33008 25974
rect 32956 25910 33008 25916
rect 33336 25838 33364 27950
rect 33324 25832 33376 25838
rect 33324 25774 33376 25780
rect 32950 25596 33258 25605
rect 32950 25594 32956 25596
rect 33012 25594 33036 25596
rect 33092 25594 33116 25596
rect 33172 25594 33196 25596
rect 33252 25594 33258 25596
rect 33012 25542 33014 25594
rect 33194 25542 33196 25594
rect 32950 25540 32956 25542
rect 33012 25540 33036 25542
rect 33092 25540 33116 25542
rect 33172 25540 33196 25542
rect 33252 25540 33258 25542
rect 32950 25531 33258 25540
rect 32864 24812 32916 24818
rect 32864 24754 32916 24760
rect 33336 24750 33364 25774
rect 33324 24744 33376 24750
rect 33324 24686 33376 24692
rect 32950 24508 33258 24517
rect 32950 24506 32956 24508
rect 33012 24506 33036 24508
rect 33092 24506 33116 24508
rect 33172 24506 33196 24508
rect 33252 24506 33258 24508
rect 33012 24454 33014 24506
rect 33194 24454 33196 24506
rect 32950 24452 32956 24454
rect 33012 24452 33036 24454
rect 33092 24452 33116 24454
rect 33172 24452 33196 24454
rect 33252 24452 33258 24454
rect 32950 24443 33258 24452
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32876 21010 32904 24142
rect 32950 23420 33258 23429
rect 32950 23418 32956 23420
rect 33012 23418 33036 23420
rect 33092 23418 33116 23420
rect 33172 23418 33196 23420
rect 33252 23418 33258 23420
rect 33012 23366 33014 23418
rect 33194 23366 33196 23418
rect 32950 23364 32956 23366
rect 33012 23364 33036 23366
rect 33092 23364 33116 23366
rect 33172 23364 33196 23366
rect 33252 23364 33258 23366
rect 32950 23355 33258 23364
rect 32950 22332 33258 22341
rect 32950 22330 32956 22332
rect 33012 22330 33036 22332
rect 33092 22330 33116 22332
rect 33172 22330 33196 22332
rect 33252 22330 33258 22332
rect 33012 22278 33014 22330
rect 33194 22278 33196 22330
rect 32950 22276 32956 22278
rect 33012 22276 33036 22278
rect 33092 22276 33116 22278
rect 33172 22276 33196 22278
rect 33252 22276 33258 22278
rect 32950 22267 33258 22276
rect 33428 22234 33456 28970
rect 33416 22228 33468 22234
rect 33416 22170 33468 22176
rect 33520 22094 33548 36502
rect 33704 36417 33732 36502
rect 33690 36408 33746 36417
rect 33690 36343 33746 36352
rect 33600 35488 33652 35494
rect 33600 35430 33652 35436
rect 33612 35086 33640 35430
rect 33600 35080 33652 35086
rect 33600 35022 33652 35028
rect 33796 34474 33824 39850
rect 33888 38010 33916 40326
rect 33876 38004 33928 38010
rect 33876 37946 33928 37952
rect 34072 37806 34100 41414
rect 34164 40594 34192 41618
rect 34152 40588 34204 40594
rect 34152 40530 34204 40536
rect 34256 39522 34284 45526
rect 35084 44810 35112 53926
rect 35348 53440 35400 53446
rect 35348 53382 35400 53388
rect 35360 44946 35388 53382
rect 35348 44940 35400 44946
rect 35348 44882 35400 44888
rect 35532 44940 35584 44946
rect 35532 44882 35584 44888
rect 35072 44804 35124 44810
rect 35072 44746 35124 44752
rect 34888 44736 34940 44742
rect 34888 44678 34940 44684
rect 34796 43376 34848 43382
rect 34796 43318 34848 43324
rect 34520 43308 34572 43314
rect 34520 43250 34572 43256
rect 34532 42702 34560 43250
rect 34520 42696 34572 42702
rect 34520 42638 34572 42644
rect 34532 42362 34560 42638
rect 34520 42356 34572 42362
rect 34520 42298 34572 42304
rect 34532 41682 34560 42298
rect 34520 41676 34572 41682
rect 34520 41618 34572 41624
rect 34704 41676 34756 41682
rect 34704 41618 34756 41624
rect 34520 40112 34572 40118
rect 34520 40054 34572 40060
rect 34336 39636 34388 39642
rect 34336 39578 34388 39584
rect 34164 39494 34284 39522
rect 34060 37800 34112 37806
rect 34060 37742 34112 37748
rect 34164 37652 34192 39494
rect 34348 39438 34376 39578
rect 34336 39432 34388 39438
rect 34336 39374 34388 39380
rect 34348 38894 34376 39374
rect 34336 38888 34388 38894
rect 34336 38830 34388 38836
rect 34532 38486 34560 40054
rect 34716 40050 34744 41618
rect 34808 40934 34836 43318
rect 34796 40928 34848 40934
rect 34796 40870 34848 40876
rect 34704 40044 34756 40050
rect 34704 39986 34756 39992
rect 34716 39438 34744 39986
rect 34796 39840 34848 39846
rect 34796 39782 34848 39788
rect 34704 39432 34756 39438
rect 34704 39374 34756 39380
rect 34520 38480 34572 38486
rect 34520 38422 34572 38428
rect 34716 38418 34744 39374
rect 34808 39098 34836 39782
rect 34900 39098 34928 44678
rect 35440 44532 35492 44538
rect 35440 44474 35492 44480
rect 35072 41540 35124 41546
rect 35072 41482 35124 41488
rect 35084 40730 35112 41482
rect 35452 41414 35480 44474
rect 35544 42158 35572 44882
rect 36556 44538 36584 53926
rect 36636 53440 36688 53446
rect 36636 53382 36688 53388
rect 36648 44538 36676 53382
rect 36544 44532 36596 44538
rect 36544 44474 36596 44480
rect 36636 44532 36688 44538
rect 36636 44474 36688 44480
rect 36176 44192 36228 44198
rect 36176 44134 36228 44140
rect 36544 44192 36596 44198
rect 36544 44134 36596 44140
rect 35992 43240 36044 43246
rect 35992 43182 36044 43188
rect 36004 42294 36032 43182
rect 35992 42288 36044 42294
rect 35992 42230 36044 42236
rect 35532 42152 35584 42158
rect 35532 42094 35584 42100
rect 35544 41818 35572 42094
rect 35624 42016 35676 42022
rect 35624 41958 35676 41964
rect 35532 41812 35584 41818
rect 35532 41754 35584 41760
rect 35452 41386 35572 41414
rect 35164 40928 35216 40934
rect 35164 40870 35216 40876
rect 35072 40724 35124 40730
rect 35072 40666 35124 40672
rect 34796 39092 34848 39098
rect 34796 39034 34848 39040
rect 34888 39092 34940 39098
rect 34888 39034 34940 39040
rect 34980 38752 35032 38758
rect 34980 38694 35032 38700
rect 34704 38412 34756 38418
rect 34704 38354 34756 38360
rect 34716 37874 34744 38354
rect 34704 37868 34756 37874
rect 34704 37810 34756 37816
rect 34072 37624 34192 37652
rect 34336 37664 34388 37670
rect 33968 36712 34020 36718
rect 33968 36654 34020 36660
rect 33876 36372 33928 36378
rect 33876 36314 33928 36320
rect 33888 35290 33916 36314
rect 33980 35766 34008 36654
rect 34072 36582 34100 37624
rect 34336 37606 34388 37612
rect 34152 37460 34204 37466
rect 34152 37402 34204 37408
rect 34060 36576 34112 36582
rect 34060 36518 34112 36524
rect 33968 35760 34020 35766
rect 33968 35702 34020 35708
rect 33876 35284 33928 35290
rect 33876 35226 33928 35232
rect 33784 34468 33836 34474
rect 33784 34410 33836 34416
rect 33784 33856 33836 33862
rect 33784 33798 33836 33804
rect 33692 31884 33744 31890
rect 33692 31826 33744 31832
rect 33598 31376 33654 31385
rect 33598 31311 33600 31320
rect 33652 31311 33654 31320
rect 33600 31282 33652 31288
rect 33704 29578 33732 31826
rect 33692 29572 33744 29578
rect 33692 29514 33744 29520
rect 33796 29458 33824 33798
rect 33888 33590 33916 35226
rect 33980 34542 34008 35702
rect 33968 34536 34020 34542
rect 33968 34478 34020 34484
rect 33876 33584 33928 33590
rect 33876 33526 33928 33532
rect 33980 33522 34008 34478
rect 33968 33516 34020 33522
rect 33968 33458 34020 33464
rect 34072 31754 34100 36518
rect 33612 29430 33824 29458
rect 33888 31726 34100 31754
rect 33612 28558 33640 29430
rect 33784 29232 33836 29238
rect 33784 29174 33836 29180
rect 33690 29064 33746 29073
rect 33690 28999 33692 29008
rect 33744 28999 33746 29008
rect 33692 28970 33744 28976
rect 33600 28552 33652 28558
rect 33600 28494 33652 28500
rect 33336 22066 33548 22094
rect 33612 22094 33640 28494
rect 33692 26988 33744 26994
rect 33692 26930 33744 26936
rect 33704 26518 33732 26930
rect 33692 26512 33744 26518
rect 33692 26454 33744 26460
rect 33704 24342 33732 26454
rect 33796 25974 33824 29174
rect 33784 25968 33836 25974
rect 33784 25910 33836 25916
rect 33888 25242 33916 31726
rect 34164 31686 34192 37402
rect 34244 36848 34296 36854
rect 34244 36790 34296 36796
rect 34256 35018 34284 36790
rect 34244 35012 34296 35018
rect 34244 34954 34296 34960
rect 34244 32292 34296 32298
rect 34244 32234 34296 32240
rect 34152 31680 34204 31686
rect 34152 31622 34204 31628
rect 34256 30394 34284 32234
rect 34348 32026 34376 37606
rect 34520 37120 34572 37126
rect 34520 37062 34572 37068
rect 34428 36372 34480 36378
rect 34428 36314 34480 36320
rect 34440 34746 34468 36314
rect 34532 36038 34560 37062
rect 34992 36242 35020 38694
rect 34612 36236 34664 36242
rect 34612 36178 34664 36184
rect 34980 36236 35032 36242
rect 34980 36178 35032 36184
rect 34520 36032 34572 36038
rect 34520 35974 34572 35980
rect 34520 35692 34572 35698
rect 34520 35634 34572 35640
rect 34428 34740 34480 34746
rect 34428 34682 34480 34688
rect 34336 32020 34388 32026
rect 34336 31962 34388 31968
rect 34336 31272 34388 31278
rect 34388 31232 34468 31260
rect 34336 31214 34388 31220
rect 34440 30394 34468 31232
rect 34244 30388 34296 30394
rect 34244 30330 34296 30336
rect 34428 30388 34480 30394
rect 34428 30330 34480 30336
rect 34336 30320 34388 30326
rect 34532 30297 34560 35634
rect 34624 34746 34652 36178
rect 35176 36174 35204 40870
rect 35256 40180 35308 40186
rect 35256 40122 35308 40128
rect 35268 38894 35296 40122
rect 35256 38888 35308 38894
rect 35256 38830 35308 38836
rect 35256 38412 35308 38418
rect 35256 38354 35308 38360
rect 35268 36718 35296 38354
rect 35440 38276 35492 38282
rect 35360 38236 35440 38264
rect 35360 38010 35388 38236
rect 35440 38218 35492 38224
rect 35348 38004 35400 38010
rect 35348 37946 35400 37952
rect 35256 36712 35308 36718
rect 35256 36654 35308 36660
rect 35072 36168 35124 36174
rect 35072 36110 35124 36116
rect 35164 36168 35216 36174
rect 35164 36110 35216 36116
rect 35084 35834 35112 36110
rect 35072 35828 35124 35834
rect 35072 35770 35124 35776
rect 34612 34740 34664 34746
rect 34612 34682 34664 34688
rect 35360 34202 35388 37946
rect 35440 37120 35492 37126
rect 35440 37062 35492 37068
rect 35452 34202 35480 37062
rect 34612 34196 34664 34202
rect 34612 34138 34664 34144
rect 35348 34196 35400 34202
rect 35348 34138 35400 34144
rect 35440 34196 35492 34202
rect 35440 34138 35492 34144
rect 34624 34066 34652 34138
rect 34612 34060 34664 34066
rect 34612 34002 34664 34008
rect 34704 33448 34756 33454
rect 34704 33390 34756 33396
rect 34612 32768 34664 32774
rect 34612 32710 34664 32716
rect 34624 32434 34652 32710
rect 34716 32502 34744 33390
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 34704 32496 34756 32502
rect 34704 32438 34756 32444
rect 34612 32428 34664 32434
rect 34612 32370 34664 32376
rect 34716 31754 34744 32438
rect 34624 31726 34744 31754
rect 34624 31414 34652 31726
rect 34612 31408 34664 31414
rect 34612 31350 34664 31356
rect 34336 30262 34388 30268
rect 34518 30288 34574 30297
rect 34060 29776 34112 29782
rect 34060 29718 34112 29724
rect 33968 29096 34020 29102
rect 33968 29038 34020 29044
rect 33980 28966 34008 29038
rect 33968 28960 34020 28966
rect 33968 28902 34020 28908
rect 33980 27470 34008 28902
rect 33968 27464 34020 27470
rect 33968 27406 34020 27412
rect 34072 26926 34100 29718
rect 34152 28620 34204 28626
rect 34152 28562 34204 28568
rect 34164 28218 34192 28562
rect 34152 28212 34204 28218
rect 34152 28154 34204 28160
rect 34152 28076 34204 28082
rect 34152 28018 34204 28024
rect 34164 27062 34192 28018
rect 34152 27056 34204 27062
rect 34204 27016 34284 27044
rect 34152 26998 34204 27004
rect 34060 26920 34112 26926
rect 34060 26862 34112 26868
rect 33968 26784 34020 26790
rect 33968 26726 34020 26732
rect 33980 25362 34008 26726
rect 34072 25514 34100 26862
rect 34256 26314 34284 27016
rect 34348 26466 34376 30262
rect 34518 30223 34574 30232
rect 34520 30048 34572 30054
rect 34520 29990 34572 29996
rect 34428 26920 34480 26926
rect 34428 26862 34480 26868
rect 34440 26586 34468 26862
rect 34428 26580 34480 26586
rect 34428 26522 34480 26528
rect 34348 26438 34468 26466
rect 34244 26308 34296 26314
rect 34244 26250 34296 26256
rect 34072 25486 34192 25514
rect 34256 25498 34284 26250
rect 34336 25900 34388 25906
rect 34336 25842 34388 25848
rect 33968 25356 34020 25362
rect 33968 25298 34020 25304
rect 34060 25356 34112 25362
rect 34060 25298 34112 25304
rect 33888 25214 34008 25242
rect 33876 24812 33928 24818
rect 33876 24754 33928 24760
rect 33888 24614 33916 24754
rect 33876 24608 33928 24614
rect 33876 24550 33928 24556
rect 33692 24336 33744 24342
rect 33692 24278 33744 24284
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 33692 23724 33744 23730
rect 33692 23666 33744 23672
rect 33704 23118 33732 23666
rect 33796 23610 33824 24142
rect 33876 24064 33928 24070
rect 33876 24006 33928 24012
rect 33888 23798 33916 24006
rect 33876 23792 33928 23798
rect 33876 23734 33928 23740
rect 33796 23582 33916 23610
rect 33692 23112 33744 23118
rect 33692 23054 33744 23060
rect 33888 22098 33916 23582
rect 33612 22066 33824 22094
rect 32950 21244 33258 21253
rect 32950 21242 32956 21244
rect 33012 21242 33036 21244
rect 33092 21242 33116 21244
rect 33172 21242 33196 21244
rect 33252 21242 33258 21244
rect 33012 21190 33014 21242
rect 33194 21190 33196 21242
rect 32950 21188 32956 21190
rect 33012 21188 33036 21190
rect 33092 21188 33116 21190
rect 33172 21188 33196 21190
rect 33252 21188 33258 21190
rect 32950 21179 33258 21188
rect 32864 21004 32916 21010
rect 32864 20946 32916 20952
rect 32864 20596 32916 20602
rect 32784 20556 32864 20584
rect 32864 20538 32916 20544
rect 32496 20256 32548 20262
rect 32496 20198 32548 20204
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32324 17054 32444 17082
rect 32312 16992 32364 16998
rect 32312 16934 32364 16940
rect 32324 15638 32352 16934
rect 32312 15632 32364 15638
rect 32312 15574 32364 15580
rect 32416 15450 32444 17054
rect 32508 15502 32536 20198
rect 32950 20156 33258 20165
rect 32950 20154 32956 20156
rect 33012 20154 33036 20156
rect 33092 20154 33116 20156
rect 33172 20154 33196 20156
rect 33252 20154 33258 20156
rect 33012 20102 33014 20154
rect 33194 20102 33196 20154
rect 32950 20100 32956 20102
rect 33012 20100 33036 20102
rect 33092 20100 33116 20102
rect 33172 20100 33196 20102
rect 33252 20100 33258 20102
rect 32950 20091 33258 20100
rect 33336 19854 33364 22066
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33324 19848 33376 19854
rect 33324 19790 33376 19796
rect 33520 19378 33548 21286
rect 33796 19666 33824 22066
rect 33876 22092 33928 22098
rect 33876 22034 33928 22040
rect 33980 19854 34008 25214
rect 34072 23594 34100 25298
rect 34060 23588 34112 23594
rect 34060 23530 34112 23536
rect 34072 21486 34100 23530
rect 34164 23526 34192 25486
rect 34244 25492 34296 25498
rect 34244 25434 34296 25440
rect 34244 24880 34296 24886
rect 34244 24822 34296 24828
rect 34152 23520 34204 23526
rect 34152 23462 34204 23468
rect 34164 23322 34192 23462
rect 34256 23322 34284 24822
rect 34348 24206 34376 25842
rect 34336 24200 34388 24206
rect 34336 24142 34388 24148
rect 34336 24064 34388 24070
rect 34440 24018 34468 26438
rect 34532 25226 34560 29990
rect 34624 29306 34652 31350
rect 34704 30252 34756 30258
rect 34704 30194 34756 30200
rect 34612 29300 34664 29306
rect 34612 29242 34664 29248
rect 34624 29102 34652 29242
rect 34612 29096 34664 29102
rect 34612 29038 34664 29044
rect 34624 28762 34652 29038
rect 34612 28756 34664 28762
rect 34612 28698 34664 28704
rect 34624 28082 34652 28698
rect 34612 28076 34664 28082
rect 34612 28018 34664 28024
rect 34612 27328 34664 27334
rect 34612 27270 34664 27276
rect 34624 27033 34652 27270
rect 34610 27024 34666 27033
rect 34610 26959 34666 26968
rect 34716 26518 34744 30194
rect 34808 28558 34836 33050
rect 35440 32972 35492 32978
rect 35440 32914 35492 32920
rect 35348 32768 35400 32774
rect 35348 32710 35400 32716
rect 35164 32360 35216 32366
rect 34992 32308 35164 32314
rect 34992 32302 35216 32308
rect 34992 32298 35204 32302
rect 34980 32292 35204 32298
rect 35032 32286 35204 32292
rect 34980 32234 35032 32240
rect 34888 32224 34940 32230
rect 34888 32166 34940 32172
rect 34900 30870 34928 32166
rect 35256 31952 35308 31958
rect 35256 31894 35308 31900
rect 35164 31272 35216 31278
rect 35164 31214 35216 31220
rect 34888 30864 34940 30870
rect 34888 30806 34940 30812
rect 34980 30592 35032 30598
rect 34980 30534 35032 30540
rect 34992 28694 35020 30534
rect 35176 29306 35204 31214
rect 35164 29300 35216 29306
rect 35164 29242 35216 29248
rect 34980 28688 35032 28694
rect 34980 28630 35032 28636
rect 34796 28552 34848 28558
rect 34796 28494 34848 28500
rect 34796 28416 34848 28422
rect 34796 28358 34848 28364
rect 34980 28416 35032 28422
rect 34980 28358 35032 28364
rect 34704 26512 34756 26518
rect 34704 26454 34756 26460
rect 34716 25838 34744 26454
rect 34704 25832 34756 25838
rect 34704 25774 34756 25780
rect 34808 25226 34836 28358
rect 34992 27441 35020 28358
rect 35176 27606 35204 29242
rect 35164 27600 35216 27606
rect 35164 27542 35216 27548
rect 35268 27538 35296 31894
rect 35360 29850 35388 32710
rect 35452 30938 35480 32914
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 35544 30598 35572 41386
rect 35636 40186 35664 41958
rect 35808 41472 35860 41478
rect 35808 41414 35860 41420
rect 35820 41386 35940 41414
rect 35912 40186 35940 41386
rect 35624 40180 35676 40186
rect 35624 40122 35676 40128
rect 35900 40180 35952 40186
rect 35900 40122 35952 40128
rect 35992 39568 36044 39574
rect 35990 39536 35992 39545
rect 36044 39536 36046 39545
rect 35990 39471 36046 39480
rect 36188 39098 36216 44134
rect 36452 39976 36504 39982
rect 36452 39918 36504 39924
rect 36176 39092 36228 39098
rect 36176 39034 36228 39040
rect 36464 38894 36492 39918
rect 36452 38888 36504 38894
rect 36452 38830 36504 38836
rect 36176 38752 36228 38758
rect 35898 38720 35954 38729
rect 36228 38712 36400 38740
rect 36176 38694 36228 38700
rect 35898 38655 35954 38664
rect 35716 37120 35768 37126
rect 35716 37062 35768 37068
rect 35728 36786 35756 37062
rect 35716 36780 35768 36786
rect 35716 36722 35768 36728
rect 35624 36100 35676 36106
rect 35624 36042 35676 36048
rect 35636 32502 35664 36042
rect 35728 35086 35756 36722
rect 35808 36644 35860 36650
rect 35808 36586 35860 36592
rect 35820 36106 35848 36586
rect 35808 36100 35860 36106
rect 35808 36042 35860 36048
rect 35808 35624 35860 35630
rect 35808 35566 35860 35572
rect 35716 35080 35768 35086
rect 35716 35022 35768 35028
rect 35728 34678 35756 35022
rect 35716 34672 35768 34678
rect 35716 34614 35768 34620
rect 35728 33590 35756 34614
rect 35820 34610 35848 35566
rect 35912 35562 35940 38655
rect 36268 38548 36320 38554
rect 36268 38490 36320 38496
rect 36084 36576 36136 36582
rect 36084 36518 36136 36524
rect 35900 35556 35952 35562
rect 35900 35498 35952 35504
rect 36096 35193 36124 36518
rect 36174 35728 36230 35737
rect 36174 35663 36230 35672
rect 36188 35630 36216 35663
rect 36176 35624 36228 35630
rect 36176 35566 36228 35572
rect 36082 35184 36138 35193
rect 36082 35119 36084 35128
rect 36136 35119 36138 35128
rect 36084 35090 36136 35096
rect 35900 34944 35952 34950
rect 35900 34886 35952 34892
rect 35992 34944 36044 34950
rect 35992 34886 36044 34892
rect 35912 34746 35940 34886
rect 35900 34740 35952 34746
rect 35900 34682 35952 34688
rect 35808 34604 35860 34610
rect 35808 34546 35860 34552
rect 35808 33992 35860 33998
rect 35808 33934 35860 33940
rect 35716 33584 35768 33590
rect 35716 33526 35768 33532
rect 35716 33448 35768 33454
rect 35716 33390 35768 33396
rect 35728 32978 35756 33390
rect 35716 32972 35768 32978
rect 35716 32914 35768 32920
rect 35716 32836 35768 32842
rect 35716 32778 35768 32784
rect 35624 32496 35676 32502
rect 35624 32438 35676 32444
rect 35728 32230 35756 32778
rect 35716 32224 35768 32230
rect 35716 32166 35768 32172
rect 35820 31754 35848 33934
rect 35900 32904 35952 32910
rect 35900 32846 35952 32852
rect 35728 31726 35848 31754
rect 35728 30802 35756 31726
rect 35808 31680 35860 31686
rect 35808 31622 35860 31628
rect 35716 30796 35768 30802
rect 35716 30738 35768 30744
rect 35532 30592 35584 30598
rect 35532 30534 35584 30540
rect 35348 29844 35400 29850
rect 35348 29786 35400 29792
rect 35348 28416 35400 28422
rect 35346 28384 35348 28393
rect 35440 28416 35492 28422
rect 35400 28384 35402 28393
rect 35440 28358 35492 28364
rect 35346 28319 35402 28328
rect 35360 28150 35388 28319
rect 35348 28144 35400 28150
rect 35348 28086 35400 28092
rect 35256 27532 35308 27538
rect 35256 27474 35308 27480
rect 34978 27432 35034 27441
rect 35452 27402 35480 28358
rect 34978 27367 35034 27376
rect 35440 27396 35492 27402
rect 35440 27338 35492 27344
rect 35072 27328 35124 27334
rect 35072 27270 35124 27276
rect 34888 26784 34940 26790
rect 34888 26726 34940 26732
rect 34900 26246 34928 26726
rect 34888 26240 34940 26246
rect 34888 26182 34940 26188
rect 34900 25294 34928 26182
rect 34888 25288 34940 25294
rect 34888 25230 34940 25236
rect 34520 25220 34572 25226
rect 34520 25162 34572 25168
rect 34796 25220 34848 25226
rect 34796 25162 34848 25168
rect 34900 24614 34928 25230
rect 34888 24608 34940 24614
rect 34888 24550 34940 24556
rect 34980 24608 35032 24614
rect 34980 24550 35032 24556
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 34388 24012 34468 24018
rect 34336 24006 34468 24012
rect 34348 23990 34468 24006
rect 34152 23316 34204 23322
rect 34152 23258 34204 23264
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 34256 22574 34284 23258
rect 34244 22568 34296 22574
rect 34244 22510 34296 22516
rect 34348 22386 34376 23990
rect 34532 23866 34560 24210
rect 34900 24206 34928 24550
rect 34888 24200 34940 24206
rect 34888 24142 34940 24148
rect 34520 23860 34572 23866
rect 34520 23802 34572 23808
rect 34520 23520 34572 23526
rect 34520 23462 34572 23468
rect 34428 23112 34480 23118
rect 34428 23054 34480 23060
rect 34164 22358 34376 22386
rect 34060 21480 34112 21486
rect 34060 21422 34112 21428
rect 34164 20210 34192 22358
rect 34244 22228 34296 22234
rect 34244 22170 34296 22176
rect 34256 21690 34284 22170
rect 34336 22160 34388 22166
rect 34336 22102 34388 22108
rect 34244 21684 34296 21690
rect 34244 21626 34296 21632
rect 34256 20398 34284 21626
rect 34244 20392 34296 20398
rect 34244 20334 34296 20340
rect 34164 20182 34284 20210
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 34152 19780 34204 19786
rect 34152 19722 34204 19728
rect 33796 19638 34008 19666
rect 33508 19372 33560 19378
rect 33508 19314 33560 19320
rect 32950 19068 33258 19077
rect 32950 19066 32956 19068
rect 33012 19066 33036 19068
rect 33092 19066 33116 19068
rect 33172 19066 33196 19068
rect 33252 19066 33258 19068
rect 33012 19014 33014 19066
rect 33194 19014 33196 19066
rect 32950 19012 32956 19014
rect 33012 19012 33036 19014
rect 33092 19012 33116 19014
rect 33172 19012 33196 19014
rect 33252 19012 33258 19014
rect 32950 19003 33258 19012
rect 32864 18896 32916 18902
rect 32864 18838 32916 18844
rect 32588 18828 32640 18834
rect 32588 18770 32640 18776
rect 32600 18358 32628 18770
rect 32588 18352 32640 18358
rect 32588 18294 32640 18300
rect 32600 17882 32628 18294
rect 32588 17876 32640 17882
rect 32588 17818 32640 17824
rect 32876 17338 32904 18838
rect 33324 18216 33376 18222
rect 33324 18158 33376 18164
rect 32950 17980 33258 17989
rect 32950 17978 32956 17980
rect 33012 17978 33036 17980
rect 33092 17978 33116 17980
rect 33172 17978 33196 17980
rect 33252 17978 33258 17980
rect 33012 17926 33014 17978
rect 33194 17926 33196 17978
rect 32950 17924 32956 17926
rect 33012 17924 33036 17926
rect 33092 17924 33116 17926
rect 33172 17924 33196 17926
rect 33252 17924 33258 17926
rect 32950 17915 33258 17924
rect 33336 17678 33364 18158
rect 33324 17672 33376 17678
rect 33324 17614 33376 17620
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33324 17264 33376 17270
rect 33324 17206 33376 17212
rect 32950 16892 33258 16901
rect 32950 16890 32956 16892
rect 33012 16890 33036 16892
rect 33092 16890 33116 16892
rect 33172 16890 33196 16892
rect 33252 16890 33258 16892
rect 33012 16838 33014 16890
rect 33194 16838 33196 16890
rect 32950 16836 32956 16838
rect 33012 16836 33036 16838
rect 33092 16836 33116 16838
rect 33172 16836 33196 16838
rect 33252 16836 33258 16838
rect 32950 16827 33258 16836
rect 33336 16574 33364 17206
rect 33416 17196 33468 17202
rect 33416 17138 33468 17144
rect 33244 16546 33364 16574
rect 33140 16448 33192 16454
rect 33140 16390 33192 16396
rect 33152 16046 33180 16390
rect 33140 16040 33192 16046
rect 33140 15982 33192 15988
rect 33244 15978 33272 16546
rect 33428 16182 33456 17138
rect 33416 16176 33468 16182
rect 33416 16118 33468 16124
rect 33232 15972 33284 15978
rect 33232 15914 33284 15920
rect 33324 15972 33376 15978
rect 33324 15914 33376 15920
rect 32864 15904 32916 15910
rect 32864 15846 32916 15852
rect 32588 15632 32640 15638
rect 32588 15574 32640 15580
rect 32324 15422 32444 15450
rect 32496 15496 32548 15502
rect 32496 15438 32548 15444
rect 32220 15020 32272 15026
rect 32220 14962 32272 14968
rect 32128 14952 32180 14958
rect 32128 14894 32180 14900
rect 32140 6914 32168 14894
rect 32232 14618 32260 14962
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 32324 8566 32352 15422
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 32416 12918 32444 15302
rect 32600 13190 32628 15574
rect 32876 14958 32904 15846
rect 32950 15804 33258 15813
rect 32950 15802 32956 15804
rect 33012 15802 33036 15804
rect 33092 15802 33116 15804
rect 33172 15802 33196 15804
rect 33252 15802 33258 15804
rect 33012 15750 33014 15802
rect 33194 15750 33196 15802
rect 32950 15748 32956 15750
rect 33012 15748 33036 15750
rect 33092 15748 33116 15750
rect 33172 15748 33196 15750
rect 33252 15748 33258 15750
rect 32950 15739 33258 15748
rect 33336 15706 33364 15914
rect 33416 15904 33468 15910
rect 33416 15846 33468 15852
rect 33324 15700 33376 15706
rect 33324 15642 33376 15648
rect 33428 15502 33456 15846
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 32864 14952 32916 14958
rect 32864 14894 32916 14900
rect 32950 14716 33258 14725
rect 32950 14714 32956 14716
rect 33012 14714 33036 14716
rect 33092 14714 33116 14716
rect 33172 14714 33196 14716
rect 33252 14714 33258 14716
rect 33012 14662 33014 14714
rect 33194 14662 33196 14714
rect 32950 14660 32956 14662
rect 33012 14660 33036 14662
rect 33092 14660 33116 14662
rect 33172 14660 33196 14662
rect 33252 14660 33258 14662
rect 32950 14651 33258 14660
rect 32950 13628 33258 13637
rect 32950 13626 32956 13628
rect 33012 13626 33036 13628
rect 33092 13626 33116 13628
rect 33172 13626 33196 13628
rect 33252 13626 33258 13628
rect 33012 13574 33014 13626
rect 33194 13574 33196 13626
rect 32950 13572 32956 13574
rect 33012 13572 33036 13574
rect 33092 13572 33116 13574
rect 33172 13572 33196 13574
rect 33252 13572 33258 13574
rect 32950 13563 33258 13572
rect 33520 13326 33548 19314
rect 33692 18080 33744 18086
rect 33692 18022 33744 18028
rect 33600 17128 33652 17134
rect 33600 17070 33652 17076
rect 33612 15570 33640 17070
rect 33600 15564 33652 15570
rect 33600 15506 33652 15512
rect 33704 15502 33732 18022
rect 33784 17672 33836 17678
rect 33784 17614 33836 17620
rect 33692 15496 33744 15502
rect 33692 15438 33744 15444
rect 33796 14906 33824 17614
rect 33980 17270 34008 19638
rect 33968 17264 34020 17270
rect 33968 17206 34020 17212
rect 34058 16688 34114 16697
rect 34058 16623 34060 16632
rect 34112 16623 34114 16632
rect 34060 16594 34112 16600
rect 33704 14878 33824 14906
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33704 13258 33732 14878
rect 33784 14816 33836 14822
rect 33784 14758 33836 14764
rect 33692 13252 33744 13258
rect 33692 13194 33744 13200
rect 32588 13184 32640 13190
rect 32588 13126 32640 13132
rect 32404 12912 32456 12918
rect 32404 12854 32456 12860
rect 32312 8560 32364 8566
rect 32312 8502 32364 8508
rect 32140 6886 32260 6914
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 31668 2984 31720 2990
rect 31668 2926 31720 2932
rect 31680 800 31708 2926
rect 32232 2446 32260 6886
rect 32416 6730 32444 12854
rect 32950 12540 33258 12549
rect 32950 12538 32956 12540
rect 33012 12538 33036 12540
rect 33092 12538 33116 12540
rect 33172 12538 33196 12540
rect 33252 12538 33258 12540
rect 33012 12486 33014 12538
rect 33194 12486 33196 12538
rect 32950 12484 32956 12486
rect 33012 12484 33036 12486
rect 33092 12484 33116 12486
rect 33172 12484 33196 12486
rect 33252 12484 33258 12486
rect 32950 12475 33258 12484
rect 32950 11452 33258 11461
rect 32950 11450 32956 11452
rect 33012 11450 33036 11452
rect 33092 11450 33116 11452
rect 33172 11450 33196 11452
rect 33252 11450 33258 11452
rect 33012 11398 33014 11450
rect 33194 11398 33196 11450
rect 32950 11396 32956 11398
rect 33012 11396 33036 11398
rect 33092 11396 33116 11398
rect 33172 11396 33196 11398
rect 33252 11396 33258 11398
rect 32950 11387 33258 11396
rect 32950 10364 33258 10373
rect 32950 10362 32956 10364
rect 33012 10362 33036 10364
rect 33092 10362 33116 10364
rect 33172 10362 33196 10364
rect 33252 10362 33258 10364
rect 33012 10310 33014 10362
rect 33194 10310 33196 10362
rect 32950 10308 32956 10310
rect 33012 10308 33036 10310
rect 33092 10308 33116 10310
rect 33172 10308 33196 10310
rect 33252 10308 33258 10310
rect 32950 10299 33258 10308
rect 32950 9276 33258 9285
rect 32950 9274 32956 9276
rect 33012 9274 33036 9276
rect 33092 9274 33116 9276
rect 33172 9274 33196 9276
rect 33252 9274 33258 9276
rect 33012 9222 33014 9274
rect 33194 9222 33196 9274
rect 32950 9220 32956 9222
rect 33012 9220 33036 9222
rect 33092 9220 33116 9222
rect 33172 9220 33196 9222
rect 33252 9220 33258 9222
rect 32950 9211 33258 9220
rect 32950 8188 33258 8197
rect 32950 8186 32956 8188
rect 33012 8186 33036 8188
rect 33092 8186 33116 8188
rect 33172 8186 33196 8188
rect 33252 8186 33258 8188
rect 33012 8134 33014 8186
rect 33194 8134 33196 8186
rect 32950 8132 32956 8134
rect 33012 8132 33036 8134
rect 33092 8132 33116 8134
rect 33172 8132 33196 8134
rect 33252 8132 33258 8134
rect 32950 8123 33258 8132
rect 32950 7100 33258 7109
rect 32950 7098 32956 7100
rect 33012 7098 33036 7100
rect 33092 7098 33116 7100
rect 33172 7098 33196 7100
rect 33252 7098 33258 7100
rect 33012 7046 33014 7098
rect 33194 7046 33196 7098
rect 32950 7044 32956 7046
rect 33012 7044 33036 7046
rect 33092 7044 33116 7046
rect 33172 7044 33196 7046
rect 33252 7044 33258 7046
rect 32950 7035 33258 7044
rect 32404 6724 32456 6730
rect 32404 6666 32456 6672
rect 32950 6012 33258 6021
rect 32950 6010 32956 6012
rect 33012 6010 33036 6012
rect 33092 6010 33116 6012
rect 33172 6010 33196 6012
rect 33252 6010 33258 6012
rect 33012 5958 33014 6010
rect 33194 5958 33196 6010
rect 32950 5956 32956 5958
rect 33012 5956 33036 5958
rect 33092 5956 33116 5958
rect 33172 5956 33196 5958
rect 33252 5956 33258 5958
rect 32950 5947 33258 5956
rect 32950 4924 33258 4933
rect 32950 4922 32956 4924
rect 33012 4922 33036 4924
rect 33092 4922 33116 4924
rect 33172 4922 33196 4924
rect 33252 4922 33258 4924
rect 33012 4870 33014 4922
rect 33194 4870 33196 4922
rect 32950 4868 32956 4870
rect 33012 4868 33036 4870
rect 33092 4868 33116 4870
rect 33172 4868 33196 4870
rect 33252 4868 33258 4870
rect 32950 4859 33258 4868
rect 32950 3836 33258 3845
rect 32950 3834 32956 3836
rect 33012 3834 33036 3836
rect 33092 3834 33116 3836
rect 33172 3834 33196 3836
rect 33252 3834 33258 3836
rect 33012 3782 33014 3834
rect 33194 3782 33196 3834
rect 32950 3780 32956 3782
rect 33012 3780 33036 3782
rect 33092 3780 33116 3782
rect 33172 3780 33196 3782
rect 33252 3780 33258 3782
rect 32950 3771 33258 3780
rect 32404 2916 32456 2922
rect 32404 2858 32456 2864
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32416 800 32444 2858
rect 32950 2748 33258 2757
rect 32950 2746 32956 2748
rect 33012 2746 33036 2748
rect 33092 2746 33116 2748
rect 33172 2746 33196 2748
rect 33252 2746 33258 2748
rect 33012 2694 33014 2746
rect 33194 2694 33196 2746
rect 32950 2692 32956 2694
rect 33012 2692 33036 2694
rect 33092 2692 33116 2694
rect 33172 2692 33196 2694
rect 33252 2692 33258 2694
rect 32950 2683 33258 2692
rect 33796 2446 33824 14758
rect 33968 14476 34020 14482
rect 33968 14418 34020 14424
rect 33980 13530 34008 14418
rect 33968 13524 34020 13530
rect 33968 13466 34020 13472
rect 33980 12918 34008 13466
rect 33968 12912 34020 12918
rect 33968 12854 34020 12860
rect 33968 9444 34020 9450
rect 33968 9386 34020 9392
rect 33980 4146 34008 9386
rect 33968 4140 34020 4146
rect 33968 4082 34020 4088
rect 33876 4072 33928 4078
rect 33876 4014 33928 4020
rect 33784 2440 33836 2446
rect 33784 2382 33836 2388
rect 33140 2304 33192 2310
rect 33140 2246 33192 2252
rect 33152 800 33180 2246
rect 33888 800 33916 4014
rect 34164 3058 34192 19722
rect 34256 14414 34284 20182
rect 34348 17814 34376 22102
rect 34440 21622 34468 23054
rect 34532 22778 34560 23462
rect 34520 22772 34572 22778
rect 34520 22714 34572 22720
rect 34520 22500 34572 22506
rect 34520 22442 34572 22448
rect 34428 21616 34480 21622
rect 34428 21558 34480 21564
rect 34532 20466 34560 22442
rect 34520 20460 34572 20466
rect 34520 20402 34572 20408
rect 34428 19168 34480 19174
rect 34428 19110 34480 19116
rect 34440 18358 34468 19110
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34428 18352 34480 18358
rect 34428 18294 34480 18300
rect 34808 18222 34836 18362
rect 34796 18216 34848 18222
rect 34796 18158 34848 18164
rect 34900 18086 34928 24142
rect 34992 19854 35020 24550
rect 35084 20942 35112 27270
rect 35544 25650 35572 30534
rect 35820 30326 35848 31622
rect 35912 31142 35940 32846
rect 36004 31521 36032 34886
rect 36084 34468 36136 34474
rect 36084 34410 36136 34416
rect 36096 34066 36124 34410
rect 36084 34060 36136 34066
rect 36084 34002 36136 34008
rect 36280 32450 36308 38490
rect 36372 36530 36400 38712
rect 36452 38276 36504 38282
rect 36452 38218 36504 38224
rect 36464 37126 36492 38218
rect 36452 37120 36504 37126
rect 36452 37062 36504 37068
rect 36556 36582 36584 44134
rect 36740 43722 36768 53926
rect 37660 44402 37688 53926
rect 37844 53582 37872 55186
rect 37950 54428 38258 54437
rect 37950 54426 37956 54428
rect 38012 54426 38036 54428
rect 38092 54426 38116 54428
rect 38172 54426 38196 54428
rect 38252 54426 38258 54428
rect 38012 54374 38014 54426
rect 38194 54374 38196 54426
rect 37950 54372 37956 54374
rect 38012 54372 38036 54374
rect 38092 54372 38116 54374
rect 38172 54372 38196 54374
rect 38252 54372 38258 54374
rect 37950 54363 38258 54372
rect 38672 54194 38700 56200
rect 39408 54194 39436 56200
rect 40144 54194 40172 56200
rect 40880 54194 40908 56200
rect 38660 54188 38712 54194
rect 38660 54130 38712 54136
rect 39396 54188 39448 54194
rect 39396 54130 39448 54136
rect 40132 54188 40184 54194
rect 40132 54130 40184 54136
rect 40868 54188 40920 54194
rect 40868 54130 40920 54136
rect 40316 54052 40368 54058
rect 40316 53994 40368 54000
rect 38936 53984 38988 53990
rect 38936 53926 38988 53932
rect 37832 53576 37884 53582
rect 37832 53518 37884 53524
rect 37950 53340 38258 53349
rect 37950 53338 37956 53340
rect 38012 53338 38036 53340
rect 38092 53338 38116 53340
rect 38172 53338 38196 53340
rect 38252 53338 38258 53340
rect 38012 53286 38014 53338
rect 38194 53286 38196 53338
rect 37950 53284 37956 53286
rect 38012 53284 38036 53286
rect 38092 53284 38116 53286
rect 38172 53284 38196 53286
rect 38252 53284 38258 53286
rect 37950 53275 38258 53284
rect 37950 52252 38258 52261
rect 37950 52250 37956 52252
rect 38012 52250 38036 52252
rect 38092 52250 38116 52252
rect 38172 52250 38196 52252
rect 38252 52250 38258 52252
rect 38012 52198 38014 52250
rect 38194 52198 38196 52250
rect 37950 52196 37956 52198
rect 38012 52196 38036 52198
rect 38092 52196 38116 52198
rect 38172 52196 38196 52198
rect 38252 52196 38258 52198
rect 37950 52187 38258 52196
rect 38384 51808 38436 51814
rect 38384 51750 38436 51756
rect 37950 51164 38258 51173
rect 37950 51162 37956 51164
rect 38012 51162 38036 51164
rect 38092 51162 38116 51164
rect 38172 51162 38196 51164
rect 38252 51162 38258 51164
rect 38012 51110 38014 51162
rect 38194 51110 38196 51162
rect 37950 51108 37956 51110
rect 38012 51108 38036 51110
rect 38092 51108 38116 51110
rect 38172 51108 38196 51110
rect 38252 51108 38258 51110
rect 37950 51099 38258 51108
rect 37950 50076 38258 50085
rect 37950 50074 37956 50076
rect 38012 50074 38036 50076
rect 38092 50074 38116 50076
rect 38172 50074 38196 50076
rect 38252 50074 38258 50076
rect 38012 50022 38014 50074
rect 38194 50022 38196 50074
rect 37950 50020 37956 50022
rect 38012 50020 38036 50022
rect 38092 50020 38116 50022
rect 38172 50020 38196 50022
rect 38252 50020 38258 50022
rect 37950 50011 38258 50020
rect 37950 48988 38258 48997
rect 37950 48986 37956 48988
rect 38012 48986 38036 48988
rect 38092 48986 38116 48988
rect 38172 48986 38196 48988
rect 38252 48986 38258 48988
rect 38012 48934 38014 48986
rect 38194 48934 38196 48986
rect 37950 48932 37956 48934
rect 38012 48932 38036 48934
rect 38092 48932 38116 48934
rect 38172 48932 38196 48934
rect 38252 48932 38258 48934
rect 37950 48923 38258 48932
rect 37950 47900 38258 47909
rect 37950 47898 37956 47900
rect 38012 47898 38036 47900
rect 38092 47898 38116 47900
rect 38172 47898 38196 47900
rect 38252 47898 38258 47900
rect 38012 47846 38014 47898
rect 38194 47846 38196 47898
rect 37950 47844 37956 47846
rect 38012 47844 38036 47846
rect 38092 47844 38116 47846
rect 38172 47844 38196 47846
rect 38252 47844 38258 47846
rect 37950 47835 38258 47844
rect 37950 46812 38258 46821
rect 37950 46810 37956 46812
rect 38012 46810 38036 46812
rect 38092 46810 38116 46812
rect 38172 46810 38196 46812
rect 38252 46810 38258 46812
rect 38012 46758 38014 46810
rect 38194 46758 38196 46810
rect 37950 46756 37956 46758
rect 38012 46756 38036 46758
rect 38092 46756 38116 46758
rect 38172 46756 38196 46758
rect 38252 46756 38258 46758
rect 37950 46747 38258 46756
rect 37950 45724 38258 45733
rect 37950 45722 37956 45724
rect 38012 45722 38036 45724
rect 38092 45722 38116 45724
rect 38172 45722 38196 45724
rect 38252 45722 38258 45724
rect 38012 45670 38014 45722
rect 38194 45670 38196 45722
rect 37950 45668 37956 45670
rect 38012 45668 38036 45670
rect 38092 45668 38116 45670
rect 38172 45668 38196 45670
rect 38252 45668 38258 45670
rect 37950 45659 38258 45668
rect 37950 44636 38258 44645
rect 37950 44634 37956 44636
rect 38012 44634 38036 44636
rect 38092 44634 38116 44636
rect 38172 44634 38196 44636
rect 38252 44634 38258 44636
rect 38012 44582 38014 44634
rect 38194 44582 38196 44634
rect 37950 44580 37956 44582
rect 38012 44580 38036 44582
rect 38092 44580 38116 44582
rect 38172 44580 38196 44582
rect 38252 44580 38258 44582
rect 37950 44571 38258 44580
rect 37648 44396 37700 44402
rect 37648 44338 37700 44344
rect 36912 44328 36964 44334
rect 36912 44270 36964 44276
rect 36728 43716 36780 43722
rect 36728 43658 36780 43664
rect 36924 42770 36952 44270
rect 37660 44198 37688 44338
rect 37648 44192 37700 44198
rect 37648 44134 37700 44140
rect 38292 43852 38344 43858
rect 38292 43794 38344 43800
rect 37280 43648 37332 43654
rect 37280 43590 37332 43596
rect 36912 42764 36964 42770
rect 36912 42706 36964 42712
rect 36820 42560 36872 42566
rect 36820 42502 36872 42508
rect 36636 41540 36688 41546
rect 36636 41482 36688 41488
rect 36648 38554 36676 41482
rect 36832 41414 36860 42502
rect 36924 41818 36952 42706
rect 37004 42696 37056 42702
rect 37004 42638 37056 42644
rect 37016 42294 37044 42638
rect 37004 42288 37056 42294
rect 37004 42230 37056 42236
rect 36912 41812 36964 41818
rect 36912 41754 36964 41760
rect 37016 41478 37044 42230
rect 37004 41472 37056 41478
rect 37004 41414 37056 41420
rect 36740 41386 36860 41414
rect 36740 39982 36768 41386
rect 37016 41206 37044 41414
rect 37004 41200 37056 41206
rect 37004 41142 37056 41148
rect 36820 40180 36872 40186
rect 36820 40122 36872 40128
rect 36728 39976 36780 39982
rect 36728 39918 36780 39924
rect 36726 39536 36782 39545
rect 36726 39471 36782 39480
rect 36636 38548 36688 38554
rect 36636 38490 36688 38496
rect 36544 36576 36596 36582
rect 36372 36502 36492 36530
rect 36544 36518 36596 36524
rect 36360 36372 36412 36378
rect 36360 36314 36412 36320
rect 36372 36106 36400 36314
rect 36464 36242 36492 36502
rect 36452 36236 36504 36242
rect 36452 36178 36504 36184
rect 36360 36100 36412 36106
rect 36360 36042 36412 36048
rect 36648 35154 36676 38490
rect 36636 35148 36688 35154
rect 36636 35090 36688 35096
rect 36360 34944 36412 34950
rect 36360 34886 36412 34892
rect 36372 34134 36400 34886
rect 36360 34128 36412 34134
rect 36636 34128 36688 34134
rect 36360 34070 36412 34076
rect 36542 34096 36598 34105
rect 36636 34070 36688 34076
rect 36542 34031 36598 34040
rect 36556 33930 36584 34031
rect 36452 33924 36504 33930
rect 36452 33866 36504 33872
rect 36544 33924 36596 33930
rect 36544 33866 36596 33872
rect 36464 33386 36492 33866
rect 36648 33674 36676 34070
rect 36556 33646 36676 33674
rect 36452 33380 36504 33386
rect 36452 33322 36504 33328
rect 36556 32570 36584 33646
rect 36636 33584 36688 33590
rect 36636 33526 36688 33532
rect 36648 32842 36676 33526
rect 36636 32836 36688 32842
rect 36636 32778 36688 32784
rect 36544 32564 36596 32570
rect 36544 32506 36596 32512
rect 36636 32496 36688 32502
rect 36280 32422 36584 32450
rect 36636 32438 36688 32444
rect 36084 32292 36136 32298
rect 36084 32234 36136 32240
rect 35990 31512 36046 31521
rect 36096 31482 36124 32234
rect 36268 31952 36320 31958
rect 36268 31894 36320 31900
rect 36176 31884 36228 31890
rect 36176 31826 36228 31832
rect 35990 31447 36046 31456
rect 36084 31476 36136 31482
rect 36084 31418 36136 31424
rect 35900 31136 35952 31142
rect 35900 31078 35952 31084
rect 35808 30320 35860 30326
rect 35808 30262 35860 30268
rect 35912 30122 35940 31078
rect 35992 30184 36044 30190
rect 35992 30126 36044 30132
rect 36084 30184 36136 30190
rect 36084 30126 36136 30132
rect 35900 30116 35952 30122
rect 35900 30058 35952 30064
rect 35912 29714 35940 30058
rect 35900 29708 35952 29714
rect 35900 29650 35952 29656
rect 35900 29504 35952 29510
rect 35900 29446 35952 29452
rect 35624 28756 35676 28762
rect 35624 28698 35676 28704
rect 35636 28626 35664 28698
rect 35624 28620 35676 28626
rect 35624 28562 35676 28568
rect 35452 25622 35572 25650
rect 35348 25492 35400 25498
rect 35348 25434 35400 25440
rect 35164 25152 35216 25158
rect 35164 25094 35216 25100
rect 35176 22710 35204 25094
rect 35360 24818 35388 25434
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 35360 24274 35388 24754
rect 35348 24268 35400 24274
rect 35348 24210 35400 24216
rect 35348 24064 35400 24070
rect 35268 24012 35348 24018
rect 35268 24006 35400 24012
rect 35268 23990 35388 24006
rect 35268 23662 35296 23990
rect 35256 23656 35308 23662
rect 35256 23598 35308 23604
rect 35268 23050 35296 23598
rect 35256 23044 35308 23050
rect 35256 22986 35308 22992
rect 35164 22704 35216 22710
rect 35164 22646 35216 22652
rect 35348 21548 35400 21554
rect 35348 21490 35400 21496
rect 35360 21078 35388 21490
rect 35452 21350 35480 25622
rect 35636 25480 35664 28562
rect 35912 28218 35940 29446
rect 36004 29238 36032 30126
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 35900 28212 35952 28218
rect 35900 28154 35952 28160
rect 36096 27606 36124 30126
rect 36188 29730 36216 31826
rect 36280 30326 36308 31894
rect 36556 31346 36584 32422
rect 36648 31686 36676 32438
rect 36740 31958 36768 39471
rect 36832 36242 36860 40122
rect 37016 40118 37044 41142
rect 37004 40112 37056 40118
rect 37004 40054 37056 40060
rect 37016 39370 37044 40054
rect 37004 39364 37056 39370
rect 37004 39306 37056 39312
rect 36912 38956 36964 38962
rect 36912 38898 36964 38904
rect 36924 38350 36952 38898
rect 36912 38344 36964 38350
rect 36912 38286 36964 38292
rect 37016 38282 37044 39306
rect 37292 39098 37320 43590
rect 37950 43548 38258 43557
rect 37950 43546 37956 43548
rect 38012 43546 38036 43548
rect 38092 43546 38116 43548
rect 38172 43546 38196 43548
rect 38252 43546 38258 43548
rect 38012 43494 38014 43546
rect 38194 43494 38196 43546
rect 37950 43492 37956 43494
rect 38012 43492 38036 43494
rect 38092 43492 38116 43494
rect 38172 43492 38196 43494
rect 38252 43492 38258 43494
rect 37950 43483 38258 43492
rect 37950 42460 38258 42469
rect 37950 42458 37956 42460
rect 38012 42458 38036 42460
rect 38092 42458 38116 42460
rect 38172 42458 38196 42460
rect 38252 42458 38258 42460
rect 38012 42406 38014 42458
rect 38194 42406 38196 42458
rect 37950 42404 37956 42406
rect 38012 42404 38036 42406
rect 38092 42404 38116 42406
rect 38172 42404 38196 42406
rect 38252 42404 38258 42406
rect 37950 42395 38258 42404
rect 38304 42362 38332 43794
rect 38292 42356 38344 42362
rect 38292 42298 38344 42304
rect 37832 42152 37884 42158
rect 37832 42094 37884 42100
rect 37844 41682 37872 42094
rect 37832 41676 37884 41682
rect 37832 41618 37884 41624
rect 37844 41138 37872 41618
rect 37950 41372 38258 41381
rect 37950 41370 37956 41372
rect 38012 41370 38036 41372
rect 38092 41370 38116 41372
rect 38172 41370 38196 41372
rect 38252 41370 38258 41372
rect 38012 41318 38014 41370
rect 38194 41318 38196 41370
rect 37950 41316 37956 41318
rect 38012 41316 38036 41318
rect 38092 41316 38116 41318
rect 38172 41316 38196 41318
rect 38252 41316 38258 41318
rect 37950 41307 38258 41316
rect 37832 41132 37884 41138
rect 37832 41074 37884 41080
rect 37740 40520 37792 40526
rect 37740 40462 37792 40468
rect 37372 40384 37424 40390
rect 37372 40326 37424 40332
rect 37280 39092 37332 39098
rect 37280 39034 37332 39040
rect 37188 38888 37240 38894
rect 37188 38830 37240 38836
rect 37004 38276 37056 38282
rect 37004 38218 37056 38224
rect 37096 38276 37148 38282
rect 37096 38218 37148 38224
rect 37108 37942 37136 38218
rect 37200 38010 37228 38830
rect 37384 38418 37412 40326
rect 37556 39364 37608 39370
rect 37556 39306 37608 39312
rect 37568 39030 37596 39306
rect 37648 39296 37700 39302
rect 37648 39238 37700 39244
rect 37556 39024 37608 39030
rect 37556 38966 37608 38972
rect 37464 38752 37516 38758
rect 37464 38694 37516 38700
rect 37372 38412 37424 38418
rect 37372 38354 37424 38360
rect 37280 38208 37332 38214
rect 37280 38150 37332 38156
rect 37188 38004 37240 38010
rect 37188 37946 37240 37952
rect 37096 37936 37148 37942
rect 37096 37878 37148 37884
rect 37004 37256 37056 37262
rect 37004 37198 37056 37204
rect 36912 36576 36964 36582
rect 36912 36518 36964 36524
rect 36820 36236 36872 36242
rect 36820 36178 36872 36184
rect 36820 36032 36872 36038
rect 36820 35974 36872 35980
rect 36728 31952 36780 31958
rect 36728 31894 36780 31900
rect 36636 31680 36688 31686
rect 36636 31622 36688 31628
rect 36832 31482 36860 35974
rect 36924 31754 36952 36518
rect 37016 33658 37044 37198
rect 37292 36378 37320 38150
rect 37280 36372 37332 36378
rect 37280 36314 37332 36320
rect 37280 35488 37332 35494
rect 37280 35430 37332 35436
rect 37188 34536 37240 34542
rect 37188 34478 37240 34484
rect 37200 34066 37228 34478
rect 37188 34060 37240 34066
rect 37188 34002 37240 34008
rect 37094 33960 37150 33969
rect 37094 33895 37150 33904
rect 37108 33862 37136 33895
rect 37096 33856 37148 33862
rect 37096 33798 37148 33804
rect 37004 33652 37056 33658
rect 37004 33594 37056 33600
rect 37108 31793 37136 33798
rect 37292 33454 37320 35430
rect 37384 34626 37412 38354
rect 37476 35086 37504 38694
rect 37556 38344 37608 38350
rect 37556 38286 37608 38292
rect 37464 35080 37516 35086
rect 37464 35022 37516 35028
rect 37568 34762 37596 38286
rect 37660 34950 37688 39238
rect 37752 36922 37780 40462
rect 37844 40050 37872 41074
rect 37950 40284 38258 40293
rect 37950 40282 37956 40284
rect 38012 40282 38036 40284
rect 38092 40282 38116 40284
rect 38172 40282 38196 40284
rect 38252 40282 38258 40284
rect 38012 40230 38014 40282
rect 38194 40230 38196 40282
rect 37950 40228 37956 40230
rect 38012 40228 38036 40230
rect 38092 40228 38116 40230
rect 38172 40228 38196 40230
rect 38252 40228 38258 40230
rect 37950 40219 38258 40228
rect 37832 40044 37884 40050
rect 37832 39986 37884 39992
rect 38304 39506 38332 42298
rect 38292 39500 38344 39506
rect 38292 39442 38344 39448
rect 37832 39296 37884 39302
rect 37832 39238 37884 39244
rect 37844 39080 37872 39238
rect 37950 39196 38258 39205
rect 37950 39194 37956 39196
rect 38012 39194 38036 39196
rect 38092 39194 38116 39196
rect 38172 39194 38196 39196
rect 38252 39194 38258 39196
rect 38012 39142 38014 39194
rect 38194 39142 38196 39194
rect 37950 39140 37956 39142
rect 38012 39140 38036 39142
rect 38092 39140 38116 39142
rect 38172 39140 38196 39142
rect 38252 39140 38258 39142
rect 37950 39131 38258 39140
rect 37844 39052 37964 39080
rect 37832 38956 37884 38962
rect 37832 38898 37884 38904
rect 37844 38010 37872 38898
rect 37936 38894 37964 39052
rect 37924 38888 37976 38894
rect 37924 38830 37976 38836
rect 37950 38108 38258 38117
rect 37950 38106 37956 38108
rect 38012 38106 38036 38108
rect 38092 38106 38116 38108
rect 38172 38106 38196 38108
rect 38252 38106 38258 38108
rect 38012 38054 38014 38106
rect 38194 38054 38196 38106
rect 37950 38052 37956 38054
rect 38012 38052 38036 38054
rect 38092 38052 38116 38054
rect 38172 38052 38196 38054
rect 38252 38052 38258 38054
rect 37950 38043 38258 38052
rect 37832 38004 37884 38010
rect 37832 37946 37884 37952
rect 37832 37868 37884 37874
rect 37832 37810 37884 37816
rect 37844 37262 37872 37810
rect 38304 37806 38332 39442
rect 37924 37800 37976 37806
rect 37922 37768 37924 37777
rect 38292 37800 38344 37806
rect 37976 37768 37978 37777
rect 38292 37742 38344 37748
rect 37922 37703 37978 37712
rect 37832 37256 37884 37262
rect 37832 37198 37884 37204
rect 37950 37020 38258 37029
rect 37950 37018 37956 37020
rect 38012 37018 38036 37020
rect 38092 37018 38116 37020
rect 38172 37018 38196 37020
rect 38252 37018 38258 37020
rect 38012 36966 38014 37018
rect 38194 36966 38196 37018
rect 37950 36964 37956 36966
rect 38012 36964 38036 36966
rect 38092 36964 38116 36966
rect 38172 36964 38196 36966
rect 38252 36964 38258 36966
rect 37950 36955 38258 36964
rect 37740 36916 37792 36922
rect 37740 36858 37792 36864
rect 38014 36680 38070 36689
rect 38014 36615 38070 36624
rect 38028 36242 38056 36615
rect 38016 36236 38068 36242
rect 38016 36178 38068 36184
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 38120 36038 38148 36178
rect 38108 36032 38160 36038
rect 38108 35974 38160 35980
rect 37950 35932 38258 35941
rect 37950 35930 37956 35932
rect 38012 35930 38036 35932
rect 38092 35930 38116 35932
rect 38172 35930 38196 35932
rect 38252 35930 38258 35932
rect 38012 35878 38014 35930
rect 38194 35878 38196 35930
rect 37950 35876 37956 35878
rect 38012 35876 38036 35878
rect 38092 35876 38116 35878
rect 38172 35876 38196 35878
rect 38252 35876 38258 35878
rect 37950 35867 38258 35876
rect 38396 35578 38424 51750
rect 38844 50720 38896 50726
rect 38844 50662 38896 50668
rect 38660 49088 38712 49094
rect 38660 49030 38712 49036
rect 38568 44872 38620 44878
rect 38568 44814 38620 44820
rect 38580 40526 38608 44814
rect 38568 40520 38620 40526
rect 38672 40497 38700 49030
rect 38752 44192 38804 44198
rect 38752 44134 38804 44140
rect 38764 40594 38792 44134
rect 38752 40588 38804 40594
rect 38752 40530 38804 40536
rect 38568 40462 38620 40468
rect 38658 40488 38714 40497
rect 38658 40423 38714 40432
rect 38568 40044 38620 40050
rect 38568 39986 38620 39992
rect 38476 39568 38528 39574
rect 38476 39510 38528 39516
rect 38488 37262 38516 39510
rect 38580 39030 38608 39986
rect 38568 39024 38620 39030
rect 38568 38966 38620 38972
rect 38672 38978 38700 40423
rect 38856 39574 38884 50662
rect 38948 43314 38976 53926
rect 39304 44328 39356 44334
rect 39304 44270 39356 44276
rect 38936 43308 38988 43314
rect 38936 43250 38988 43256
rect 39316 41414 39344 44270
rect 40328 43450 40356 53994
rect 40408 53984 40460 53990
rect 40408 53926 40460 53932
rect 41328 53984 41380 53990
rect 41328 53926 41380 53932
rect 41512 53984 41564 53990
rect 41512 53926 41564 53932
rect 40316 43444 40368 43450
rect 40316 43386 40368 43392
rect 39856 43308 39908 43314
rect 39856 43250 39908 43256
rect 39672 42220 39724 42226
rect 39672 42162 39724 42168
rect 39684 41546 39712 42162
rect 39672 41540 39724 41546
rect 39672 41482 39724 41488
rect 39224 41386 39344 41414
rect 38936 41064 38988 41070
rect 38936 41006 38988 41012
rect 38844 39568 38896 39574
rect 38844 39510 38896 39516
rect 38844 39432 38896 39438
rect 38844 39374 38896 39380
rect 38856 39098 38884 39374
rect 38844 39092 38896 39098
rect 38844 39034 38896 39040
rect 38672 38950 38884 38978
rect 38660 38888 38712 38894
rect 38660 38830 38712 38836
rect 38672 38729 38700 38830
rect 38658 38720 38714 38729
rect 38658 38655 38714 38664
rect 38660 38276 38712 38282
rect 38660 38218 38712 38224
rect 38568 38208 38620 38214
rect 38568 38150 38620 38156
rect 38476 37256 38528 37262
rect 38476 37198 38528 37204
rect 38580 36825 38608 38150
rect 38672 37806 38700 38218
rect 38660 37800 38712 37806
rect 38856 37777 38884 38950
rect 38660 37742 38712 37748
rect 38842 37768 38898 37777
rect 38672 37398 38700 37742
rect 38842 37703 38898 37712
rect 38660 37392 38712 37398
rect 38660 37334 38712 37340
rect 38566 36816 38622 36825
rect 38566 36751 38622 36760
rect 38672 36718 38700 37334
rect 38476 36712 38528 36718
rect 38660 36712 38712 36718
rect 38476 36654 38528 36660
rect 38580 36660 38660 36666
rect 38580 36654 38712 36660
rect 38212 35562 38424 35578
rect 38200 35556 38424 35562
rect 38252 35550 38424 35556
rect 38200 35498 38252 35504
rect 38016 35284 38068 35290
rect 37844 35244 38016 35272
rect 37844 35154 37872 35244
rect 38016 35226 38068 35232
rect 37922 35184 37978 35193
rect 37832 35148 37884 35154
rect 37922 35119 37924 35128
rect 37832 35090 37884 35096
rect 37976 35119 37978 35128
rect 37924 35090 37976 35096
rect 37648 34944 37700 34950
rect 37648 34886 37700 34892
rect 37950 34844 38258 34853
rect 37950 34842 37956 34844
rect 38012 34842 38036 34844
rect 38092 34842 38116 34844
rect 38172 34842 38196 34844
rect 38252 34842 38258 34844
rect 38012 34790 38014 34842
rect 38194 34790 38196 34842
rect 37950 34788 37956 34790
rect 38012 34788 38036 34790
rect 38092 34788 38116 34790
rect 38172 34788 38196 34790
rect 38252 34788 38258 34790
rect 37950 34779 38258 34788
rect 37568 34734 37688 34762
rect 37384 34598 37596 34626
rect 37372 33584 37424 33590
rect 37372 33526 37424 33532
rect 37280 33448 37332 33454
rect 37280 33390 37332 33396
rect 37188 32768 37240 32774
rect 37188 32710 37240 32716
rect 37094 31784 37150 31793
rect 36924 31726 37044 31754
rect 36820 31476 36872 31482
rect 36820 31418 36872 31424
rect 37016 31385 37044 31726
rect 37094 31719 37150 31728
rect 37002 31376 37058 31385
rect 36544 31340 36596 31346
rect 37002 31311 37058 31320
rect 36544 31282 36596 31288
rect 36544 30592 36596 30598
rect 36544 30534 36596 30540
rect 36268 30320 36320 30326
rect 36268 30262 36320 30268
rect 36188 29702 36308 29730
rect 36280 29510 36308 29702
rect 36268 29504 36320 29510
rect 36268 29446 36320 29452
rect 36280 28966 36308 29446
rect 36268 28960 36320 28966
rect 36268 28902 36320 28908
rect 36360 28960 36412 28966
rect 36360 28902 36412 28908
rect 36280 28626 36308 28902
rect 36268 28620 36320 28626
rect 36268 28562 36320 28568
rect 36372 28558 36400 28902
rect 36360 28552 36412 28558
rect 36360 28494 36412 28500
rect 36450 28520 36506 28529
rect 36556 28506 36584 30534
rect 36636 29572 36688 29578
rect 36636 29514 36688 29520
rect 36648 29170 36676 29514
rect 36728 29300 36780 29306
rect 36728 29242 36780 29248
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36556 28478 36676 28506
rect 36450 28455 36506 28464
rect 36464 28218 36492 28455
rect 36544 28416 36596 28422
rect 36544 28358 36596 28364
rect 36556 28218 36584 28358
rect 36452 28212 36504 28218
rect 36452 28154 36504 28160
rect 36544 28212 36596 28218
rect 36544 28154 36596 28160
rect 36084 27600 36136 27606
rect 36084 27542 36136 27548
rect 35900 27124 35952 27130
rect 35900 27066 35952 27072
rect 35912 25838 35940 27066
rect 35900 25832 35952 25838
rect 35900 25774 35952 25780
rect 35992 25696 36044 25702
rect 35992 25638 36044 25644
rect 35544 25452 35664 25480
rect 35544 24138 35572 25452
rect 36004 25362 36032 25638
rect 35624 25356 35676 25362
rect 35624 25298 35676 25304
rect 35992 25356 36044 25362
rect 35992 25298 36044 25304
rect 35532 24132 35584 24138
rect 35532 24074 35584 24080
rect 35544 23662 35572 24074
rect 35636 24070 35664 25298
rect 35992 24948 36044 24954
rect 35992 24890 36044 24896
rect 35624 24064 35676 24070
rect 35624 24006 35676 24012
rect 35532 23656 35584 23662
rect 35532 23598 35584 23604
rect 36004 21554 36032 24890
rect 36268 24132 36320 24138
rect 36188 24092 36268 24120
rect 36188 23050 36216 24092
rect 36268 24074 36320 24080
rect 36176 23044 36228 23050
rect 36096 23004 36176 23032
rect 36096 21962 36124 23004
rect 36176 22986 36228 22992
rect 36464 22094 36492 28154
rect 36648 26858 36676 28478
rect 36636 26852 36688 26858
rect 36636 26794 36688 26800
rect 36544 25152 36596 25158
rect 36544 25094 36596 25100
rect 36556 24954 36584 25094
rect 36544 24948 36596 24954
rect 36544 24890 36596 24896
rect 36648 24410 36676 26794
rect 36636 24404 36688 24410
rect 36636 24346 36688 24352
rect 36188 22066 36492 22094
rect 36084 21956 36136 21962
rect 36084 21898 36136 21904
rect 36096 21622 36124 21898
rect 36084 21616 36136 21622
rect 36084 21558 36136 21564
rect 35992 21548 36044 21554
rect 35992 21490 36044 21496
rect 35440 21344 35492 21350
rect 35440 21286 35492 21292
rect 35348 21072 35400 21078
rect 35348 21014 35400 21020
rect 35072 20936 35124 20942
rect 35072 20878 35124 20884
rect 35162 20632 35218 20641
rect 35162 20567 35218 20576
rect 35176 20058 35204 20567
rect 35164 20052 35216 20058
rect 35164 19994 35216 20000
rect 35440 19916 35492 19922
rect 35440 19858 35492 19864
rect 34980 19848 35032 19854
rect 34980 19790 35032 19796
rect 34980 19712 35032 19718
rect 34980 19654 35032 19660
rect 34992 19417 35020 19654
rect 34978 19408 35034 19417
rect 34978 19343 35034 19352
rect 34888 18080 34940 18086
rect 34888 18022 34940 18028
rect 34336 17808 34388 17814
rect 34336 17750 34388 17756
rect 34612 17128 34664 17134
rect 34612 17070 34664 17076
rect 34624 16726 34652 17070
rect 34612 16720 34664 16726
rect 34612 16662 34664 16668
rect 34900 16658 34928 18022
rect 34888 16652 34940 16658
rect 34888 16594 34940 16600
rect 34520 16516 34572 16522
rect 34520 16458 34572 16464
rect 34336 14544 34388 14550
rect 34336 14486 34388 14492
rect 34244 14408 34296 14414
rect 34244 14350 34296 14356
rect 34244 13184 34296 13190
rect 34244 13126 34296 13132
rect 34256 3534 34284 13126
rect 34348 12782 34376 14486
rect 34532 14482 34560 16458
rect 34900 14634 34928 16594
rect 34808 14606 34928 14634
rect 34520 14476 34572 14482
rect 34520 14418 34572 14424
rect 34704 14000 34756 14006
rect 34704 13942 34756 13948
rect 34716 13190 34744 13942
rect 34704 13184 34756 13190
rect 34704 13126 34756 13132
rect 34716 12918 34744 13126
rect 34808 12986 34836 14606
rect 34888 14068 34940 14074
rect 34888 14010 34940 14016
rect 34900 13394 34928 14010
rect 34888 13388 34940 13394
rect 34888 13330 34940 13336
rect 34796 12980 34848 12986
rect 34796 12922 34848 12928
rect 34704 12912 34756 12918
rect 34704 12854 34756 12860
rect 34336 12776 34388 12782
rect 34336 12718 34388 12724
rect 34992 9654 35020 19343
rect 35452 19174 35480 19858
rect 35900 19372 35952 19378
rect 36096 19360 36124 21558
rect 36188 20874 36216 22066
rect 36176 20868 36228 20874
rect 36176 20810 36228 20816
rect 36360 20868 36412 20874
rect 36360 20810 36412 20816
rect 35952 19332 36124 19360
rect 35900 19314 35952 19320
rect 36096 19174 36124 19332
rect 35440 19168 35492 19174
rect 35440 19110 35492 19116
rect 36084 19168 36136 19174
rect 36084 19110 36136 19116
rect 36096 18358 36124 19110
rect 36084 18352 36136 18358
rect 36084 18294 36136 18300
rect 35256 18216 35308 18222
rect 35256 18158 35308 18164
rect 35268 17134 35296 18158
rect 36084 18080 36136 18086
rect 36084 18022 36136 18028
rect 35900 17740 35952 17746
rect 35900 17682 35952 17688
rect 35256 17128 35308 17134
rect 35256 17070 35308 17076
rect 35532 16652 35584 16658
rect 35532 16594 35584 16600
rect 35164 14340 35216 14346
rect 35164 14282 35216 14288
rect 34980 9648 35032 9654
rect 34980 9590 35032 9596
rect 35176 6914 35204 14282
rect 35544 13870 35572 16594
rect 35912 15570 35940 17682
rect 36096 17610 36124 18022
rect 36084 17604 36136 17610
rect 36084 17546 36136 17552
rect 36176 16788 36228 16794
rect 36176 16730 36228 16736
rect 36084 15904 36136 15910
rect 36084 15846 36136 15852
rect 35900 15564 35952 15570
rect 35900 15506 35952 15512
rect 35912 14074 35940 15506
rect 35900 14068 35952 14074
rect 35900 14010 35952 14016
rect 35532 13864 35584 13870
rect 35532 13806 35584 13812
rect 35440 13728 35492 13734
rect 35440 13670 35492 13676
rect 35452 12986 35480 13670
rect 35440 12980 35492 12986
rect 35440 12922 35492 12928
rect 36096 12714 36124 15846
rect 36188 15570 36216 16730
rect 36372 16114 36400 20810
rect 36544 20800 36596 20806
rect 36544 20742 36596 20748
rect 36452 17332 36504 17338
rect 36452 17274 36504 17280
rect 36464 16522 36492 17274
rect 36452 16516 36504 16522
rect 36452 16458 36504 16464
rect 36360 16108 36412 16114
rect 36360 16050 36412 16056
rect 36176 15564 36228 15570
rect 36176 15506 36228 15512
rect 36464 15434 36492 16458
rect 36452 15428 36504 15434
rect 36452 15370 36504 15376
rect 36556 14006 36584 20742
rect 36740 19854 36768 29242
rect 36912 25696 36964 25702
rect 36912 25638 36964 25644
rect 36924 25226 36952 25638
rect 36912 25220 36964 25226
rect 36912 25162 36964 25168
rect 36912 19916 36964 19922
rect 36912 19858 36964 19864
rect 36728 19848 36780 19854
rect 36728 19790 36780 19796
rect 36636 19236 36688 19242
rect 36636 19178 36688 19184
rect 36648 16454 36676 19178
rect 36728 18692 36780 18698
rect 36728 18634 36780 18640
rect 36636 16448 36688 16454
rect 36636 16390 36688 16396
rect 36636 15428 36688 15434
rect 36636 15370 36688 15376
rect 36544 14000 36596 14006
rect 36544 13942 36596 13948
rect 36648 13682 36676 15370
rect 36556 13654 36676 13682
rect 36556 13258 36584 13654
rect 36544 13252 36596 13258
rect 36544 13194 36596 13200
rect 36084 12708 36136 12714
rect 36084 12650 36136 12656
rect 35176 6886 35296 6914
rect 34612 3596 34664 3602
rect 34612 3538 34664 3544
rect 34244 3528 34296 3534
rect 34244 3470 34296 3476
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 34624 800 34652 3538
rect 35268 2446 35296 6886
rect 36556 4010 36584 13194
rect 36544 4004 36596 4010
rect 36544 3946 36596 3952
rect 36084 3596 36136 3602
rect 36084 3538 36136 3544
rect 35348 2508 35400 2514
rect 35348 2450 35400 2456
rect 35256 2440 35308 2446
rect 35256 2382 35308 2388
rect 35360 800 35388 2450
rect 36096 800 36124 3538
rect 36740 3534 36768 18634
rect 36820 18352 36872 18358
rect 36820 18294 36872 18300
rect 36832 17610 36860 18294
rect 36820 17604 36872 17610
rect 36820 17546 36872 17552
rect 36832 17338 36860 17546
rect 36820 17332 36872 17338
rect 36820 17274 36872 17280
rect 36820 16992 36872 16998
rect 36820 16934 36872 16940
rect 36832 15094 36860 16934
rect 36924 16640 36952 19858
rect 37016 18630 37044 31311
rect 37096 29572 37148 29578
rect 37096 29514 37148 29520
rect 37108 29102 37136 29514
rect 37200 29238 37228 32710
rect 37280 31884 37332 31890
rect 37280 31826 37332 31832
rect 37188 29232 37240 29238
rect 37188 29174 37240 29180
rect 37096 29096 37148 29102
rect 37096 29038 37148 29044
rect 37200 28506 37228 29174
rect 37108 28478 37228 28506
rect 37108 27402 37136 28478
rect 37188 28416 37240 28422
rect 37188 28358 37240 28364
rect 37096 27396 37148 27402
rect 37096 27338 37148 27344
rect 37108 27130 37136 27338
rect 37096 27124 37148 27130
rect 37096 27066 37148 27072
rect 37096 26580 37148 26586
rect 37096 26522 37148 26528
rect 37108 26353 37136 26522
rect 37094 26344 37150 26353
rect 37094 26279 37150 26288
rect 37200 24818 37228 28358
rect 37292 28121 37320 31826
rect 37384 30818 37412 33526
rect 37464 32428 37516 32434
rect 37464 32370 37516 32376
rect 37476 30938 37504 32370
rect 37568 30938 37596 34598
rect 37660 31890 37688 34734
rect 37832 34604 37884 34610
rect 37832 34546 37884 34552
rect 37740 34060 37792 34066
rect 37740 34002 37792 34008
rect 37752 33862 37780 34002
rect 37740 33856 37792 33862
rect 37740 33798 37792 33804
rect 37844 33674 37872 34546
rect 38396 34082 38424 35550
rect 38304 34054 38424 34082
rect 38488 34066 38516 36654
rect 38580 36638 38700 36654
rect 38580 35766 38608 36638
rect 38752 36032 38804 36038
rect 38752 35974 38804 35980
rect 38568 35760 38620 35766
rect 38568 35702 38620 35708
rect 38658 35048 38714 35057
rect 38658 34983 38660 34992
rect 38712 34983 38714 34992
rect 38660 34954 38712 34960
rect 38764 34354 38792 35974
rect 38948 34921 38976 41006
rect 39224 40934 39252 41386
rect 39684 41290 39712 41482
rect 39868 41414 39896 43250
rect 40040 42832 40092 42838
rect 40040 42774 40092 42780
rect 40052 41414 40080 42774
rect 40420 42566 40448 53926
rect 40684 53440 40736 53446
rect 40684 53382 40736 53388
rect 40696 44538 40724 53382
rect 40776 48544 40828 48550
rect 40776 48486 40828 48492
rect 40684 44532 40736 44538
rect 40684 44474 40736 44480
rect 40592 43240 40644 43246
rect 40592 43182 40644 43188
rect 40224 42560 40276 42566
rect 40224 42502 40276 42508
rect 40408 42560 40460 42566
rect 40408 42502 40460 42508
rect 40500 42560 40552 42566
rect 40500 42502 40552 42508
rect 39868 41386 39988 41414
rect 40052 41386 40172 41414
rect 39684 41262 39896 41290
rect 39868 41206 39896 41262
rect 39856 41200 39908 41206
rect 39856 41142 39908 41148
rect 39488 40996 39540 41002
rect 39488 40938 39540 40944
rect 39212 40928 39264 40934
rect 39212 40870 39264 40876
rect 39396 40588 39448 40594
rect 39396 40530 39448 40536
rect 39120 40384 39172 40390
rect 39120 40326 39172 40332
rect 39132 39098 39160 40326
rect 39408 39982 39436 40530
rect 39396 39976 39448 39982
rect 39396 39918 39448 39924
rect 39212 39636 39264 39642
rect 39212 39578 39264 39584
rect 39120 39092 39172 39098
rect 39120 39034 39172 39040
rect 39118 37768 39174 37777
rect 39118 37703 39174 37712
rect 39132 37126 39160 37703
rect 39120 37120 39172 37126
rect 39120 37062 39172 37068
rect 39028 36848 39080 36854
rect 39028 36790 39080 36796
rect 38934 34912 38990 34921
rect 38934 34847 38990 34856
rect 38934 34776 38990 34785
rect 38934 34711 38936 34720
rect 38988 34711 38990 34720
rect 38936 34682 38988 34688
rect 38672 34326 38792 34354
rect 38672 34218 38700 34326
rect 38626 34202 38700 34218
rect 38614 34196 38700 34202
rect 38666 34190 38700 34196
rect 38750 34232 38806 34241
rect 38750 34167 38806 34176
rect 38936 34196 38988 34202
rect 38614 34138 38666 34144
rect 38658 34096 38714 34105
rect 38476 34060 38528 34066
rect 37950 33756 38258 33765
rect 37950 33754 37956 33756
rect 38012 33754 38036 33756
rect 38092 33754 38116 33756
rect 38172 33754 38196 33756
rect 38252 33754 38258 33756
rect 38012 33702 38014 33754
rect 38194 33702 38196 33754
rect 37950 33700 37956 33702
rect 38012 33700 38036 33702
rect 38092 33700 38116 33702
rect 38172 33700 38196 33702
rect 38252 33700 38258 33702
rect 37950 33691 38258 33700
rect 37752 33646 37872 33674
rect 37752 32978 37780 33646
rect 38304 33590 38332 34054
rect 38764 34066 38792 34167
rect 38936 34138 38988 34144
rect 38658 34031 38660 34040
rect 38476 34002 38528 34008
rect 38712 34031 38714 34040
rect 38752 34060 38804 34066
rect 38660 34002 38712 34008
rect 38752 34002 38804 34008
rect 38292 33584 38344 33590
rect 37830 33552 37886 33561
rect 38292 33526 38344 33532
rect 37830 33487 37832 33496
rect 37884 33487 37886 33496
rect 37832 33458 37884 33464
rect 38384 33312 38436 33318
rect 38384 33254 38436 33260
rect 37740 32972 37792 32978
rect 37740 32914 37792 32920
rect 37832 32904 37884 32910
rect 37832 32846 37884 32852
rect 37648 31884 37700 31890
rect 37648 31826 37700 31832
rect 37844 31822 37872 32846
rect 37950 32668 38258 32677
rect 37950 32666 37956 32668
rect 38012 32666 38036 32668
rect 38092 32666 38116 32668
rect 38172 32666 38196 32668
rect 38252 32666 38258 32668
rect 38012 32614 38014 32666
rect 38194 32614 38196 32666
rect 37950 32612 37956 32614
rect 38012 32612 38036 32614
rect 38092 32612 38116 32614
rect 38172 32612 38196 32614
rect 38252 32612 38258 32614
rect 37950 32603 38258 32612
rect 38396 31872 38424 33254
rect 38488 32298 38516 34002
rect 38844 33992 38896 33998
rect 38948 33980 38976 34138
rect 38896 33952 38976 33980
rect 38844 33934 38896 33940
rect 38614 33856 38666 33862
rect 38666 33804 38976 33810
rect 38614 33798 38976 33804
rect 38626 33782 38976 33798
rect 38750 33688 38806 33697
rect 38750 33623 38806 33632
rect 38568 33040 38620 33046
rect 38568 32982 38620 32988
rect 38476 32292 38528 32298
rect 38476 32234 38528 32240
rect 38580 31929 38608 32982
rect 38764 32978 38792 33623
rect 38842 33552 38898 33561
rect 38842 33487 38898 33496
rect 38752 32972 38804 32978
rect 38752 32914 38804 32920
rect 38660 31952 38712 31958
rect 38566 31920 38622 31929
rect 38476 31884 38528 31890
rect 38396 31844 38476 31872
rect 37832 31816 37884 31822
rect 37832 31758 37884 31764
rect 37464 30932 37516 30938
rect 37464 30874 37516 30880
rect 37556 30932 37608 30938
rect 37556 30874 37608 30880
rect 37384 30790 37688 30818
rect 37556 30728 37608 30734
rect 37556 30670 37608 30676
rect 37372 30048 37424 30054
rect 37372 29990 37424 29996
rect 37464 30048 37516 30054
rect 37464 29990 37516 29996
rect 37384 28626 37412 29990
rect 37372 28620 37424 28626
rect 37372 28562 37424 28568
rect 37476 28234 37504 29990
rect 37384 28206 37504 28234
rect 37278 28112 37334 28121
rect 37278 28047 37334 28056
rect 37280 28008 37332 28014
rect 37280 27950 37332 27956
rect 37188 24812 37240 24818
rect 37188 24754 37240 24760
rect 37292 24274 37320 27950
rect 37384 25430 37412 28206
rect 37464 28076 37516 28082
rect 37464 28018 37516 28024
rect 37476 26994 37504 28018
rect 37568 27062 37596 30670
rect 37660 29714 37688 30790
rect 37740 30592 37792 30598
rect 37740 30534 37792 30540
rect 37648 29708 37700 29714
rect 37648 29650 37700 29656
rect 37556 27056 37608 27062
rect 37556 26998 37608 27004
rect 37464 26988 37516 26994
rect 37464 26930 37516 26936
rect 37476 26450 37504 26930
rect 37568 26450 37596 26998
rect 37464 26444 37516 26450
rect 37464 26386 37516 26392
rect 37556 26444 37608 26450
rect 37556 26386 37608 26392
rect 37660 26330 37688 29650
rect 37568 26302 37688 26330
rect 37752 26330 37780 30534
rect 37844 30326 37872 31758
rect 37950 31580 38258 31589
rect 37950 31578 37956 31580
rect 38012 31578 38036 31580
rect 38092 31578 38116 31580
rect 38172 31578 38196 31580
rect 38252 31578 38258 31580
rect 38012 31526 38014 31578
rect 38194 31526 38196 31578
rect 37950 31524 37956 31526
rect 38012 31524 38036 31526
rect 38092 31524 38116 31526
rect 38172 31524 38196 31526
rect 38252 31524 38258 31526
rect 37950 31515 38258 31524
rect 37924 31408 37976 31414
rect 37924 31350 37976 31356
rect 37936 30802 37964 31350
rect 38396 31346 38424 31844
rect 38660 31894 38712 31900
rect 38566 31855 38568 31864
rect 38476 31826 38528 31832
rect 38620 31855 38622 31864
rect 38568 31826 38620 31832
rect 38566 31784 38622 31793
rect 38566 31719 38622 31728
rect 38476 31680 38528 31686
rect 38476 31622 38528 31628
rect 38488 31385 38516 31622
rect 38580 31482 38608 31719
rect 38672 31482 38700 31894
rect 38568 31476 38620 31482
rect 38568 31418 38620 31424
rect 38660 31476 38712 31482
rect 38660 31418 38712 31424
rect 38474 31376 38530 31385
rect 38384 31340 38436 31346
rect 38474 31311 38530 31320
rect 38568 31340 38620 31346
rect 38384 31282 38436 31288
rect 38568 31282 38620 31288
rect 38476 31272 38528 31278
rect 38476 31214 38528 31220
rect 38488 30938 38516 31214
rect 38476 30932 38528 30938
rect 38476 30874 38528 30880
rect 37924 30796 37976 30802
rect 37924 30738 37976 30744
rect 37950 30492 38258 30501
rect 37950 30490 37956 30492
rect 38012 30490 38036 30492
rect 38092 30490 38116 30492
rect 38172 30490 38196 30492
rect 38252 30490 38258 30492
rect 38012 30438 38014 30490
rect 38194 30438 38196 30490
rect 37950 30436 37956 30438
rect 38012 30436 38036 30438
rect 38092 30436 38116 30438
rect 38172 30436 38196 30438
rect 38252 30436 38258 30438
rect 37950 30427 38258 30436
rect 37832 30320 37884 30326
rect 37924 30320 37976 30326
rect 37832 30262 37884 30268
rect 37922 30288 37924 30297
rect 37976 30288 37978 30297
rect 37922 30223 37978 30232
rect 38016 30184 38068 30190
rect 38016 30126 38068 30132
rect 38028 29850 38056 30126
rect 38384 30116 38436 30122
rect 38384 30058 38436 30064
rect 38016 29844 38068 29850
rect 38016 29786 38068 29792
rect 38292 29844 38344 29850
rect 38292 29786 38344 29792
rect 37950 29404 38258 29413
rect 37950 29402 37956 29404
rect 38012 29402 38036 29404
rect 38092 29402 38116 29404
rect 38172 29402 38196 29404
rect 38252 29402 38258 29404
rect 38012 29350 38014 29402
rect 38194 29350 38196 29402
rect 37950 29348 37956 29350
rect 38012 29348 38036 29350
rect 38092 29348 38116 29350
rect 38172 29348 38196 29350
rect 38252 29348 38258 29350
rect 37950 29339 38258 29348
rect 37832 29096 37884 29102
rect 37832 29038 37884 29044
rect 37844 27402 37872 29038
rect 37950 28316 38258 28325
rect 37950 28314 37956 28316
rect 38012 28314 38036 28316
rect 38092 28314 38116 28316
rect 38172 28314 38196 28316
rect 38252 28314 38258 28316
rect 38012 28262 38014 28314
rect 38194 28262 38196 28314
rect 37950 28260 37956 28262
rect 38012 28260 38036 28262
rect 38092 28260 38116 28262
rect 38172 28260 38196 28262
rect 38252 28260 38258 28262
rect 37950 28251 38258 28260
rect 38304 28014 38332 29786
rect 38396 29034 38424 30058
rect 38384 29028 38436 29034
rect 38384 28970 38436 28976
rect 38396 28150 38424 28970
rect 38384 28144 38436 28150
rect 38384 28086 38436 28092
rect 38292 28008 38344 28014
rect 38292 27950 38344 27956
rect 37832 27396 37884 27402
rect 37832 27338 37884 27344
rect 37950 27228 38258 27237
rect 37950 27226 37956 27228
rect 38012 27226 38036 27228
rect 38092 27226 38116 27228
rect 38172 27226 38196 27228
rect 38252 27226 38258 27228
rect 38012 27174 38014 27226
rect 38194 27174 38196 27226
rect 37950 27172 37956 27174
rect 38012 27172 38036 27174
rect 38092 27172 38116 27174
rect 38172 27172 38196 27174
rect 38252 27172 38258 27174
rect 37950 27163 38258 27172
rect 38292 26920 38344 26926
rect 38292 26862 38344 26868
rect 37752 26302 37872 26330
rect 37568 25906 37596 26302
rect 37740 26240 37792 26246
rect 37740 26182 37792 26188
rect 37752 26042 37780 26182
rect 37740 26036 37792 26042
rect 37740 25978 37792 25984
rect 37648 25968 37700 25974
rect 37648 25910 37700 25916
rect 37556 25900 37608 25906
rect 37556 25842 37608 25848
rect 37464 25764 37516 25770
rect 37464 25706 37516 25712
rect 37556 25764 37608 25770
rect 37556 25706 37608 25712
rect 37372 25424 37424 25430
rect 37372 25366 37424 25372
rect 37476 24886 37504 25706
rect 37464 24880 37516 24886
rect 37464 24822 37516 24828
rect 37280 24268 37332 24274
rect 37280 24210 37332 24216
rect 37292 23798 37320 24210
rect 37372 24064 37424 24070
rect 37372 24006 37424 24012
rect 37280 23792 37332 23798
rect 37280 23734 37332 23740
rect 37188 22976 37240 22982
rect 37188 22918 37240 22924
rect 37200 22642 37228 22918
rect 37188 22636 37240 22642
rect 37188 22578 37240 22584
rect 37292 22098 37320 23734
rect 37384 23050 37412 24006
rect 37464 23180 37516 23186
rect 37464 23122 37516 23128
rect 37372 23044 37424 23050
rect 37372 22986 37424 22992
rect 37476 22642 37504 23122
rect 37464 22636 37516 22642
rect 37464 22578 37516 22584
rect 37280 22092 37332 22098
rect 37280 22034 37332 22040
rect 37096 21344 37148 21350
rect 37096 21286 37148 21292
rect 37004 18624 37056 18630
rect 37004 18566 37056 18572
rect 37108 17814 37136 21286
rect 37476 19378 37504 22578
rect 37464 19372 37516 19378
rect 37464 19314 37516 19320
rect 37280 19304 37332 19310
rect 37280 19246 37332 19252
rect 37292 18834 37320 19246
rect 37568 19174 37596 25706
rect 37660 20874 37688 25910
rect 37740 25696 37792 25702
rect 37740 25638 37792 25644
rect 37648 20868 37700 20874
rect 37648 20810 37700 20816
rect 37556 19168 37608 19174
rect 37556 19110 37608 19116
rect 37568 18970 37596 19110
rect 37556 18964 37608 18970
rect 37556 18906 37608 18912
rect 37280 18828 37332 18834
rect 37280 18770 37332 18776
rect 37188 18692 37240 18698
rect 37188 18634 37240 18640
rect 37200 17882 37228 18634
rect 37188 17876 37240 17882
rect 37188 17818 37240 17824
rect 37096 17808 37148 17814
rect 37096 17750 37148 17756
rect 37096 17604 37148 17610
rect 37096 17546 37148 17552
rect 37108 16794 37136 17546
rect 37096 16788 37148 16794
rect 37096 16730 37148 16736
rect 37200 16658 37228 17818
rect 37292 17746 37320 18770
rect 37372 18284 37424 18290
rect 37372 18226 37424 18232
rect 37280 17740 37332 17746
rect 37280 17682 37332 17688
rect 37188 16652 37240 16658
rect 36924 16612 37136 16640
rect 36912 16448 36964 16454
rect 36912 16390 36964 16396
rect 36820 15088 36872 15094
rect 36820 15030 36872 15036
rect 36924 14958 36952 16390
rect 36912 14952 36964 14958
rect 36912 14894 36964 14900
rect 36912 14272 36964 14278
rect 36912 14214 36964 14220
rect 36924 13938 36952 14214
rect 36912 13932 36964 13938
rect 36912 13874 36964 13880
rect 37108 13326 37136 16612
rect 37188 16594 37240 16600
rect 37384 16182 37412 18226
rect 37372 16176 37424 16182
rect 37372 16118 37424 16124
rect 37568 16046 37596 18906
rect 37752 18426 37780 25638
rect 37844 25498 37872 26302
rect 37950 26140 38258 26149
rect 37950 26138 37956 26140
rect 38012 26138 38036 26140
rect 38092 26138 38116 26140
rect 38172 26138 38196 26140
rect 38252 26138 38258 26140
rect 38012 26086 38014 26138
rect 38194 26086 38196 26138
rect 37950 26084 37956 26086
rect 38012 26084 38036 26086
rect 38092 26084 38116 26086
rect 38172 26084 38196 26086
rect 38252 26084 38258 26086
rect 37950 26075 38258 26084
rect 38304 25974 38332 26862
rect 38384 26784 38436 26790
rect 38384 26726 38436 26732
rect 38292 25968 38344 25974
rect 38292 25910 38344 25916
rect 37832 25492 37884 25498
rect 37832 25434 37884 25440
rect 37844 24206 37872 25434
rect 37950 25052 38258 25061
rect 37950 25050 37956 25052
rect 38012 25050 38036 25052
rect 38092 25050 38116 25052
rect 38172 25050 38196 25052
rect 38252 25050 38258 25052
rect 38012 24998 38014 25050
rect 38194 24998 38196 25050
rect 37950 24996 37956 24998
rect 38012 24996 38036 24998
rect 38092 24996 38116 24998
rect 38172 24996 38196 24998
rect 38252 24996 38258 24998
rect 37950 24987 38258 24996
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37832 24064 37884 24070
rect 37832 24006 37884 24012
rect 37844 22982 37872 24006
rect 37950 23964 38258 23973
rect 37950 23962 37956 23964
rect 38012 23962 38036 23964
rect 38092 23962 38116 23964
rect 38172 23962 38196 23964
rect 38252 23962 38258 23964
rect 38012 23910 38014 23962
rect 38194 23910 38196 23962
rect 37950 23908 37956 23910
rect 38012 23908 38036 23910
rect 38092 23908 38116 23910
rect 38172 23908 38196 23910
rect 38252 23908 38258 23910
rect 37950 23899 38258 23908
rect 38200 23860 38252 23866
rect 38200 23802 38252 23808
rect 38212 23066 38240 23802
rect 38304 23730 38332 25910
rect 38292 23724 38344 23730
rect 38292 23666 38344 23672
rect 38396 23254 38424 26726
rect 38488 25906 38516 30874
rect 38580 30054 38608 31282
rect 38660 30796 38712 30802
rect 38660 30738 38712 30744
rect 38568 30048 38620 30054
rect 38568 29990 38620 29996
rect 38672 29050 38700 30738
rect 38752 30592 38804 30598
rect 38752 30534 38804 30540
rect 38580 29022 38700 29050
rect 38580 28762 38608 29022
rect 38660 28960 38712 28966
rect 38660 28902 38712 28908
rect 38568 28756 38620 28762
rect 38568 28698 38620 28704
rect 38568 28620 38620 28626
rect 38568 28562 38620 28568
rect 38580 27606 38608 28562
rect 38672 28558 38700 28902
rect 38660 28552 38712 28558
rect 38660 28494 38712 28500
rect 38568 27600 38620 27606
rect 38568 27542 38620 27548
rect 38476 25900 38528 25906
rect 38476 25842 38528 25848
rect 38580 25362 38608 27542
rect 38658 26344 38714 26353
rect 38658 26279 38714 26288
rect 38568 25356 38620 25362
rect 38568 25298 38620 25304
rect 38672 25242 38700 26279
rect 38580 25214 38700 25242
rect 38476 24880 38528 24886
rect 38476 24822 38528 24828
rect 38384 23248 38436 23254
rect 38384 23190 38436 23196
rect 38212 23038 38424 23066
rect 37832 22976 37884 22982
rect 37832 22918 37884 22924
rect 38292 22976 38344 22982
rect 38292 22918 38344 22924
rect 37950 22876 38258 22885
rect 37950 22874 37956 22876
rect 38012 22874 38036 22876
rect 38092 22874 38116 22876
rect 38172 22874 38196 22876
rect 38252 22874 38258 22876
rect 38012 22822 38014 22874
rect 38194 22822 38196 22874
rect 37950 22820 37956 22822
rect 38012 22820 38036 22822
rect 38092 22820 38116 22822
rect 38172 22820 38196 22822
rect 38252 22820 38258 22822
rect 37950 22811 38258 22820
rect 37832 22704 37884 22710
rect 37832 22646 37884 22652
rect 37844 21690 37872 22646
rect 37950 21788 38258 21797
rect 37950 21786 37956 21788
rect 38012 21786 38036 21788
rect 38092 21786 38116 21788
rect 38172 21786 38196 21788
rect 38252 21786 38258 21788
rect 38012 21734 38014 21786
rect 38194 21734 38196 21786
rect 37950 21732 37956 21734
rect 38012 21732 38036 21734
rect 38092 21732 38116 21734
rect 38172 21732 38196 21734
rect 38252 21732 38258 21734
rect 37950 21723 38258 21732
rect 37832 21684 37884 21690
rect 37832 21626 37884 21632
rect 37844 21010 37872 21626
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 38304 20942 38332 22918
rect 38292 20936 38344 20942
rect 38292 20878 38344 20884
rect 37950 20700 38258 20709
rect 37950 20698 37956 20700
rect 38012 20698 38036 20700
rect 38092 20698 38116 20700
rect 38172 20698 38196 20700
rect 38252 20698 38258 20700
rect 38012 20646 38014 20698
rect 38194 20646 38196 20698
rect 37950 20644 37956 20646
rect 38012 20644 38036 20646
rect 38092 20644 38116 20646
rect 38172 20644 38196 20646
rect 38252 20644 38258 20646
rect 37950 20635 38258 20644
rect 37950 19612 38258 19621
rect 37950 19610 37956 19612
rect 38012 19610 38036 19612
rect 38092 19610 38116 19612
rect 38172 19610 38196 19612
rect 38252 19610 38258 19612
rect 38012 19558 38014 19610
rect 38194 19558 38196 19610
rect 37950 19556 37956 19558
rect 38012 19556 38036 19558
rect 38092 19556 38116 19558
rect 38172 19556 38196 19558
rect 38252 19556 38258 19558
rect 37950 19547 38258 19556
rect 37950 18524 38258 18533
rect 37950 18522 37956 18524
rect 38012 18522 38036 18524
rect 38092 18522 38116 18524
rect 38172 18522 38196 18524
rect 38252 18522 38258 18524
rect 38012 18470 38014 18522
rect 38194 18470 38196 18522
rect 37950 18468 37956 18470
rect 38012 18468 38036 18470
rect 38092 18468 38116 18470
rect 38172 18468 38196 18470
rect 38252 18468 38258 18470
rect 37950 18459 38258 18468
rect 37740 18420 37792 18426
rect 37740 18362 37792 18368
rect 38016 18216 38068 18222
rect 38016 18158 38068 18164
rect 38028 17746 38056 18158
rect 38016 17740 38068 17746
rect 38016 17682 38068 17688
rect 37832 17536 37884 17542
rect 37832 17478 37884 17484
rect 37844 16590 37872 17478
rect 37950 17436 38258 17445
rect 37950 17434 37956 17436
rect 38012 17434 38036 17436
rect 38092 17434 38116 17436
rect 38172 17434 38196 17436
rect 38252 17434 38258 17436
rect 38012 17382 38014 17434
rect 38194 17382 38196 17434
rect 37950 17380 37956 17382
rect 38012 17380 38036 17382
rect 38092 17380 38116 17382
rect 38172 17380 38196 17382
rect 38252 17380 38258 17382
rect 37950 17371 38258 17380
rect 38108 16992 38160 16998
rect 38108 16934 38160 16940
rect 37832 16584 37884 16590
rect 37832 16526 37884 16532
rect 38120 16454 38148 16934
rect 38108 16448 38160 16454
rect 38108 16390 38160 16396
rect 37950 16348 38258 16357
rect 37950 16346 37956 16348
rect 38012 16346 38036 16348
rect 38092 16346 38116 16348
rect 38172 16346 38196 16348
rect 38252 16346 38258 16348
rect 38012 16294 38014 16346
rect 38194 16294 38196 16346
rect 37950 16292 37956 16294
rect 38012 16292 38036 16294
rect 38092 16292 38116 16294
rect 38172 16292 38196 16294
rect 38252 16292 38258 16294
rect 37950 16283 38258 16292
rect 37556 16040 37608 16046
rect 37556 15982 37608 15988
rect 37648 15904 37700 15910
rect 37648 15846 37700 15852
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37660 15162 37688 15846
rect 37740 15360 37792 15366
rect 37740 15302 37792 15308
rect 37648 15156 37700 15162
rect 37648 15098 37700 15104
rect 37752 14482 37780 15302
rect 37740 14476 37792 14482
rect 37660 14436 37740 14464
rect 37660 13394 37688 14436
rect 37740 14418 37792 14424
rect 37740 14340 37792 14346
rect 37740 14282 37792 14288
rect 37752 14006 37780 14282
rect 37740 14000 37792 14006
rect 37740 13942 37792 13948
rect 37648 13388 37700 13394
rect 37648 13330 37700 13336
rect 37096 13320 37148 13326
rect 37096 13262 37148 13268
rect 37280 13320 37332 13326
rect 37280 13262 37332 13268
rect 37292 12986 37320 13262
rect 37372 13252 37424 13258
rect 37372 13194 37424 13200
rect 37280 12980 37332 12986
rect 37280 12922 37332 12928
rect 36820 12708 36872 12714
rect 36820 12650 36872 12656
rect 36832 6798 36860 12650
rect 37280 9444 37332 9450
rect 37280 9386 37332 9392
rect 36820 6792 36872 6798
rect 36820 6734 36872 6740
rect 37292 3534 37320 9386
rect 36728 3528 36780 3534
rect 36728 3470 36780 3476
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 37384 3126 37412 13194
rect 37844 8566 37872 15846
rect 37950 15260 38258 15269
rect 37950 15258 37956 15260
rect 38012 15258 38036 15260
rect 38092 15258 38116 15260
rect 38172 15258 38196 15260
rect 38252 15258 38258 15260
rect 38012 15206 38014 15258
rect 38194 15206 38196 15258
rect 37950 15204 37956 15206
rect 38012 15204 38036 15206
rect 38092 15204 38116 15206
rect 38172 15204 38196 15206
rect 38252 15204 38258 15206
rect 37950 15195 38258 15204
rect 38292 14884 38344 14890
rect 38292 14826 38344 14832
rect 37950 14172 38258 14181
rect 37950 14170 37956 14172
rect 38012 14170 38036 14172
rect 38092 14170 38116 14172
rect 38172 14170 38196 14172
rect 38252 14170 38258 14172
rect 38012 14118 38014 14170
rect 38194 14118 38196 14170
rect 37950 14116 37956 14118
rect 38012 14116 38036 14118
rect 38092 14116 38116 14118
rect 38172 14116 38196 14118
rect 38252 14116 38258 14118
rect 37950 14107 38258 14116
rect 38304 13326 38332 14826
rect 38396 14006 38424 23038
rect 38488 21962 38516 24822
rect 38580 23866 38608 25214
rect 38764 25158 38792 30534
rect 38856 28082 38884 33487
rect 38948 33130 38976 33782
rect 39040 33318 39068 36790
rect 39120 35624 39172 35630
rect 39120 35566 39172 35572
rect 39028 33312 39080 33318
rect 39028 33254 39080 33260
rect 38948 33102 39068 33130
rect 38936 32972 38988 32978
rect 38936 32914 38988 32920
rect 38948 30394 38976 32914
rect 39040 32586 39068 33102
rect 39132 32774 39160 35566
rect 39224 35154 39252 39578
rect 39408 38894 39436 39918
rect 39396 38888 39448 38894
rect 39396 38830 39448 38836
rect 39500 37210 39528 40938
rect 39764 40928 39816 40934
rect 39764 40870 39816 40876
rect 39580 40724 39632 40730
rect 39580 40666 39632 40672
rect 39592 38010 39620 40666
rect 39776 39964 39804 40870
rect 39868 40186 39896 41142
rect 39960 41070 39988 41386
rect 39948 41064 40000 41070
rect 39948 41006 40000 41012
rect 39948 40928 40000 40934
rect 39948 40870 40000 40876
rect 39960 40594 39988 40870
rect 39948 40588 40000 40594
rect 39948 40530 40000 40536
rect 39948 40452 40000 40458
rect 39948 40394 40000 40400
rect 39856 40180 39908 40186
rect 39856 40122 39908 40128
rect 39776 39936 39896 39964
rect 39868 39642 39896 39936
rect 39856 39636 39908 39642
rect 39856 39578 39908 39584
rect 39672 39296 39724 39302
rect 39672 39238 39724 39244
rect 39684 38962 39712 39238
rect 39672 38956 39724 38962
rect 39672 38898 39724 38904
rect 39580 38004 39632 38010
rect 39580 37946 39632 37952
rect 39408 37182 39528 37210
rect 39302 36680 39358 36689
rect 39302 36615 39358 36624
rect 39316 35834 39344 36615
rect 39304 35828 39356 35834
rect 39304 35770 39356 35776
rect 39212 35148 39264 35154
rect 39212 35090 39264 35096
rect 39212 35012 39264 35018
rect 39212 34954 39264 34960
rect 39120 32768 39172 32774
rect 39120 32710 39172 32716
rect 39040 32558 39160 32586
rect 39028 32360 39080 32366
rect 39028 32302 39080 32308
rect 39040 31890 39068 32302
rect 39028 31884 39080 31890
rect 39028 31826 39080 31832
rect 38936 30388 38988 30394
rect 38936 30330 38988 30336
rect 39040 30326 39068 31826
rect 39028 30320 39080 30326
rect 39028 30262 39080 30268
rect 39028 30184 39080 30190
rect 39028 30126 39080 30132
rect 39040 29850 39068 30126
rect 39132 29850 39160 32558
rect 39028 29844 39080 29850
rect 39028 29786 39080 29792
rect 39120 29844 39172 29850
rect 39120 29786 39172 29792
rect 39224 29238 39252 34954
rect 39316 33697 39344 35770
rect 39408 35057 39436 37182
rect 39488 37120 39540 37126
rect 39488 37062 39540 37068
rect 39394 35048 39450 35057
rect 39394 34983 39450 34992
rect 39408 34082 39436 34983
rect 39500 34746 39528 37062
rect 39580 36848 39632 36854
rect 39580 36790 39632 36796
rect 39592 35698 39620 36790
rect 39684 36281 39712 38898
rect 39868 38894 39896 39578
rect 39856 38888 39908 38894
rect 39856 38830 39908 38836
rect 39670 36272 39726 36281
rect 39670 36207 39726 36216
rect 39580 35692 39632 35698
rect 39580 35634 39632 35640
rect 39592 35170 39620 35634
rect 39592 35142 39712 35170
rect 39580 35080 39632 35086
rect 39580 35022 39632 35028
rect 39592 34746 39620 35022
rect 39488 34740 39540 34746
rect 39488 34682 39540 34688
rect 39580 34740 39632 34746
rect 39580 34682 39632 34688
rect 39580 34128 39632 34134
rect 39578 34096 39580 34105
rect 39632 34096 39634 34105
rect 39408 34054 39528 34082
rect 39396 33924 39448 33930
rect 39396 33866 39448 33872
rect 39302 33688 39358 33697
rect 39302 33623 39358 33632
rect 39304 33584 39356 33590
rect 39304 33526 39356 33532
rect 39212 29232 39264 29238
rect 39212 29174 39264 29180
rect 39224 28218 39252 29174
rect 39212 28212 39264 28218
rect 39212 28154 39264 28160
rect 39316 28150 39344 33526
rect 39408 33454 39436 33866
rect 39396 33448 39448 33454
rect 39396 33390 39448 33396
rect 39500 30734 39528 34054
rect 39578 34031 39634 34040
rect 39580 32564 39632 32570
rect 39684 32552 39712 35142
rect 39868 34610 39896 38830
rect 39960 38654 39988 40394
rect 40040 39092 40092 39098
rect 40040 39034 40092 39040
rect 40052 38826 40080 39034
rect 40040 38820 40092 38826
rect 40040 38762 40092 38768
rect 39960 38626 40080 38654
rect 40052 36825 40080 38626
rect 40144 37806 40172 41386
rect 40132 37800 40184 37806
rect 40132 37742 40184 37748
rect 40144 37330 40172 37742
rect 40132 37324 40184 37330
rect 40132 37266 40184 37272
rect 40236 37262 40264 42502
rect 40316 42152 40368 42158
rect 40316 42094 40368 42100
rect 40328 40186 40356 42094
rect 40420 41721 40448 42502
rect 40406 41712 40462 41721
rect 40406 41647 40462 41656
rect 40316 40180 40368 40186
rect 40316 40122 40368 40128
rect 40328 37806 40356 40122
rect 40408 38412 40460 38418
rect 40408 38354 40460 38360
rect 40420 38214 40448 38354
rect 40408 38208 40460 38214
rect 40408 38150 40460 38156
rect 40408 37868 40460 37874
rect 40408 37810 40460 37816
rect 40316 37800 40368 37806
rect 40316 37742 40368 37748
rect 40316 37664 40368 37670
rect 40316 37606 40368 37612
rect 40328 37330 40356 37606
rect 40316 37324 40368 37330
rect 40316 37266 40368 37272
rect 40224 37256 40276 37262
rect 40224 37198 40276 37204
rect 40038 36816 40094 36825
rect 40038 36751 40094 36760
rect 39948 36712 40000 36718
rect 39948 36654 40000 36660
rect 39960 35834 39988 36654
rect 39948 35828 40000 35834
rect 39948 35770 40000 35776
rect 39856 34604 39908 34610
rect 39856 34546 39908 34552
rect 39960 34542 39988 35770
rect 39948 34536 40000 34542
rect 39948 34478 40000 34484
rect 39948 34400 40000 34406
rect 39948 34342 40000 34348
rect 39764 33856 39816 33862
rect 39764 33798 39816 33804
rect 39632 32524 39712 32552
rect 39580 32506 39632 32512
rect 39488 30728 39540 30734
rect 39488 30670 39540 30676
rect 39592 30326 39620 32506
rect 39672 30932 39724 30938
rect 39672 30874 39724 30880
rect 39580 30320 39632 30326
rect 39580 30262 39632 30268
rect 39684 29306 39712 30874
rect 39776 29306 39804 33798
rect 39960 32230 39988 34342
rect 40052 34241 40080 36751
rect 40224 36100 40276 36106
rect 40224 36042 40276 36048
rect 40236 35086 40264 36042
rect 40328 35494 40356 37266
rect 40420 36854 40448 37810
rect 40408 36848 40460 36854
rect 40408 36790 40460 36796
rect 40408 36576 40460 36582
rect 40408 36518 40460 36524
rect 40316 35488 40368 35494
rect 40316 35430 40368 35436
rect 40224 35080 40276 35086
rect 40224 35022 40276 35028
rect 40132 35012 40184 35018
rect 40132 34954 40184 34960
rect 40038 34232 40094 34241
rect 40038 34167 40094 34176
rect 40144 33658 40172 34954
rect 40420 34474 40448 36518
rect 40512 36242 40540 42502
rect 40604 38894 40632 43182
rect 40788 39098 40816 48486
rect 41052 47456 41104 47462
rect 41052 47398 41104 47404
rect 40960 43716 41012 43722
rect 40960 43658 41012 43664
rect 40972 39846 41000 43658
rect 40960 39840 41012 39846
rect 40960 39782 41012 39788
rect 40868 39432 40920 39438
rect 40868 39374 40920 39380
rect 40776 39092 40828 39098
rect 40776 39034 40828 39040
rect 40592 38888 40644 38894
rect 40592 38830 40644 38836
rect 40604 38418 40632 38830
rect 40592 38412 40644 38418
rect 40592 38354 40644 38360
rect 40604 36922 40632 38354
rect 40684 38208 40736 38214
rect 40684 38150 40736 38156
rect 40696 37874 40724 38150
rect 40684 37868 40736 37874
rect 40684 37810 40736 37816
rect 40684 37324 40736 37330
rect 40684 37266 40736 37272
rect 40592 36916 40644 36922
rect 40592 36858 40644 36864
rect 40604 36582 40632 36858
rect 40592 36576 40644 36582
rect 40592 36518 40644 36524
rect 40592 36304 40644 36310
rect 40592 36246 40644 36252
rect 40500 36236 40552 36242
rect 40500 36178 40552 36184
rect 40408 34468 40460 34474
rect 40408 34410 40460 34416
rect 40224 34400 40276 34406
rect 40224 34342 40276 34348
rect 40132 33652 40184 33658
rect 40132 33594 40184 33600
rect 40132 32768 40184 32774
rect 40132 32710 40184 32716
rect 40040 32496 40092 32502
rect 40040 32438 40092 32444
rect 39948 32224 40000 32230
rect 39868 32172 39948 32178
rect 39868 32166 40000 32172
rect 39868 32150 39988 32166
rect 39672 29300 39724 29306
rect 39672 29242 39724 29248
rect 39764 29300 39816 29306
rect 39764 29242 39816 29248
rect 39672 29164 39724 29170
rect 39672 29106 39724 29112
rect 39304 28144 39356 28150
rect 39304 28086 39356 28092
rect 39580 28144 39632 28150
rect 39580 28086 39632 28092
rect 38844 28076 38896 28082
rect 38844 28018 38896 28024
rect 39212 28076 39264 28082
rect 39212 28018 39264 28024
rect 38752 25152 38804 25158
rect 38752 25094 38804 25100
rect 39224 24070 39252 28018
rect 39396 27872 39448 27878
rect 39396 27814 39448 27820
rect 39408 25906 39436 27814
rect 39592 26382 39620 28086
rect 39684 28014 39712 29106
rect 39868 29102 39896 32150
rect 40052 31822 40080 32438
rect 40040 31816 40092 31822
rect 40040 31758 40092 31764
rect 40040 31476 40092 31482
rect 40040 31418 40092 31424
rect 40052 30802 40080 31418
rect 40040 30796 40092 30802
rect 40040 30738 40092 30744
rect 39948 30116 40000 30122
rect 39948 30058 40000 30064
rect 39856 29096 39908 29102
rect 39856 29038 39908 29044
rect 39672 28008 39724 28014
rect 39672 27950 39724 27956
rect 39684 27606 39712 27950
rect 39672 27600 39724 27606
rect 39672 27542 39724 27548
rect 39580 26376 39632 26382
rect 39580 26318 39632 26324
rect 39488 26308 39540 26314
rect 39488 26250 39540 26256
rect 39396 25900 39448 25906
rect 39396 25842 39448 25848
rect 39500 25498 39528 26250
rect 39960 26042 39988 30058
rect 40040 29640 40092 29646
rect 40040 29582 40092 29588
rect 40052 29034 40080 29582
rect 40040 29028 40092 29034
rect 40040 28970 40092 28976
rect 40052 27538 40080 28970
rect 40144 28490 40172 32710
rect 40236 31754 40264 34342
rect 40316 33448 40368 33454
rect 40316 33390 40368 33396
rect 40328 31890 40356 33390
rect 40512 32774 40540 36178
rect 40604 34950 40632 36246
rect 40696 36106 40724 37266
rect 40684 36100 40736 36106
rect 40684 36042 40736 36048
rect 40788 35986 40816 39034
rect 40880 39030 40908 39374
rect 40868 39024 40920 39030
rect 40868 38966 40920 38972
rect 40972 38434 41000 39782
rect 40696 35958 40816 35986
rect 40880 38406 41000 38434
rect 40696 35698 40724 35958
rect 40774 35864 40830 35873
rect 40774 35799 40830 35808
rect 40788 35766 40816 35799
rect 40776 35760 40828 35766
rect 40776 35702 40828 35708
rect 40684 35692 40736 35698
rect 40684 35634 40736 35640
rect 40684 35080 40736 35086
rect 40684 35022 40736 35028
rect 40592 34944 40644 34950
rect 40592 34886 40644 34892
rect 40604 34610 40632 34886
rect 40592 34604 40644 34610
rect 40592 34546 40644 34552
rect 40592 33448 40644 33454
rect 40592 33390 40644 33396
rect 40604 33114 40632 33390
rect 40592 33108 40644 33114
rect 40592 33050 40644 33056
rect 40590 33008 40646 33017
rect 40590 32943 40646 32952
rect 40604 32910 40632 32943
rect 40696 32910 40724 35022
rect 40880 34610 40908 38406
rect 41064 38350 41092 47398
rect 41236 43104 41288 43110
rect 41236 43046 41288 43052
rect 41144 40112 41196 40118
rect 41144 40054 41196 40060
rect 41156 38554 41184 40054
rect 41248 40050 41276 43046
rect 41340 42226 41368 53926
rect 41524 43790 41552 53926
rect 41616 53582 41644 56200
rect 41696 54324 41748 54330
rect 41696 54266 41748 54272
rect 41604 53576 41656 53582
rect 41604 53518 41656 53524
rect 41708 45554 41736 54266
rect 42352 54262 42380 56200
rect 42340 54256 42392 54262
rect 42340 54198 42392 54204
rect 43088 54194 43116 56200
rect 43824 56114 43852 56200
rect 43916 56114 43944 56222
rect 43824 56086 43944 56114
rect 44100 54194 44128 56222
rect 44546 56200 44602 57000
rect 46754 56200 46810 57000
rect 47490 56200 47546 57000
rect 48226 56200 48282 57000
rect 48962 56200 49018 57000
rect 49698 56200 49754 57000
rect 50434 56200 50490 57000
rect 44560 54194 44588 56200
rect 43076 54188 43128 54194
rect 43076 54130 43128 54136
rect 44088 54188 44140 54194
rect 44088 54130 44140 54136
rect 44548 54188 44600 54194
rect 44548 54130 44600 54136
rect 43628 54052 43680 54058
rect 43628 53994 43680 54000
rect 42950 53884 43258 53893
rect 42950 53882 42956 53884
rect 43012 53882 43036 53884
rect 43092 53882 43116 53884
rect 43172 53882 43196 53884
rect 43252 53882 43258 53884
rect 43012 53830 43014 53882
rect 43194 53830 43196 53882
rect 42950 53828 42956 53830
rect 43012 53828 43036 53830
rect 43092 53828 43116 53830
rect 43172 53828 43196 53830
rect 43252 53828 43258 53830
rect 42950 53819 43258 53828
rect 42950 52796 43258 52805
rect 42950 52794 42956 52796
rect 43012 52794 43036 52796
rect 43092 52794 43116 52796
rect 43172 52794 43196 52796
rect 43252 52794 43258 52796
rect 43012 52742 43014 52794
rect 43194 52742 43196 52794
rect 42950 52740 42956 52742
rect 43012 52740 43036 52742
rect 43092 52740 43116 52742
rect 43172 52740 43196 52742
rect 43252 52740 43258 52742
rect 42950 52731 43258 52740
rect 42950 51708 43258 51717
rect 42950 51706 42956 51708
rect 43012 51706 43036 51708
rect 43092 51706 43116 51708
rect 43172 51706 43196 51708
rect 43252 51706 43258 51708
rect 43012 51654 43014 51706
rect 43194 51654 43196 51706
rect 42950 51652 42956 51654
rect 43012 51652 43036 51654
rect 43092 51652 43116 51654
rect 43172 51652 43196 51654
rect 43252 51652 43258 51654
rect 42950 51643 43258 51652
rect 42950 50620 43258 50629
rect 42950 50618 42956 50620
rect 43012 50618 43036 50620
rect 43092 50618 43116 50620
rect 43172 50618 43196 50620
rect 43252 50618 43258 50620
rect 43012 50566 43014 50618
rect 43194 50566 43196 50618
rect 42950 50564 42956 50566
rect 43012 50564 43036 50566
rect 43092 50564 43116 50566
rect 43172 50564 43196 50566
rect 43252 50564 43258 50566
rect 42950 50555 43258 50564
rect 42950 49532 43258 49541
rect 42950 49530 42956 49532
rect 43012 49530 43036 49532
rect 43092 49530 43116 49532
rect 43172 49530 43196 49532
rect 43252 49530 43258 49532
rect 43012 49478 43014 49530
rect 43194 49478 43196 49530
rect 42950 49476 42956 49478
rect 43012 49476 43036 49478
rect 43092 49476 43116 49478
rect 43172 49476 43196 49478
rect 43252 49476 43258 49478
rect 42950 49467 43258 49476
rect 42950 48444 43258 48453
rect 42950 48442 42956 48444
rect 43012 48442 43036 48444
rect 43092 48442 43116 48444
rect 43172 48442 43196 48444
rect 43252 48442 43258 48444
rect 43012 48390 43014 48442
rect 43194 48390 43196 48442
rect 42950 48388 42956 48390
rect 43012 48388 43036 48390
rect 43092 48388 43116 48390
rect 43172 48388 43196 48390
rect 43252 48388 43258 48390
rect 42950 48379 43258 48388
rect 42950 47356 43258 47365
rect 42950 47354 42956 47356
rect 43012 47354 43036 47356
rect 43092 47354 43116 47356
rect 43172 47354 43196 47356
rect 43252 47354 43258 47356
rect 43012 47302 43014 47354
rect 43194 47302 43196 47354
rect 42950 47300 42956 47302
rect 43012 47300 43036 47302
rect 43092 47300 43116 47302
rect 43172 47300 43196 47302
rect 43252 47300 43258 47302
rect 42950 47291 43258 47300
rect 42950 46268 43258 46277
rect 42950 46266 42956 46268
rect 43012 46266 43036 46268
rect 43092 46266 43116 46268
rect 43172 46266 43196 46268
rect 43252 46266 43258 46268
rect 43012 46214 43014 46266
rect 43194 46214 43196 46266
rect 42950 46212 42956 46214
rect 43012 46212 43036 46214
rect 43092 46212 43116 46214
rect 43172 46212 43196 46214
rect 43252 46212 43258 46214
rect 42950 46203 43258 46212
rect 41616 45526 41736 45554
rect 41512 43784 41564 43790
rect 41512 43726 41564 43732
rect 41616 42362 41644 45526
rect 42950 45180 43258 45189
rect 42950 45178 42956 45180
rect 43012 45178 43036 45180
rect 43092 45178 43116 45180
rect 43172 45178 43196 45180
rect 43252 45178 43258 45180
rect 43012 45126 43014 45178
rect 43194 45126 43196 45178
rect 42950 45124 42956 45126
rect 43012 45124 43036 45126
rect 43092 45124 43116 45126
rect 43172 45124 43196 45126
rect 43252 45124 43258 45126
rect 42950 45115 43258 45124
rect 43444 44192 43496 44198
rect 43444 44134 43496 44140
rect 42950 44092 43258 44101
rect 42950 44090 42956 44092
rect 43012 44090 43036 44092
rect 43092 44090 43116 44092
rect 43172 44090 43196 44092
rect 43252 44090 43258 44092
rect 43012 44038 43014 44090
rect 43194 44038 43196 44090
rect 42950 44036 42956 44038
rect 43012 44036 43036 44038
rect 43092 44036 43116 44038
rect 43172 44036 43196 44038
rect 43252 44036 43258 44038
rect 42950 44027 43258 44036
rect 42064 43240 42116 43246
rect 42064 43182 42116 43188
rect 41604 42356 41656 42362
rect 41604 42298 41656 42304
rect 41328 42220 41380 42226
rect 41328 42162 41380 42168
rect 41340 42129 41368 42162
rect 41326 42120 41382 42129
rect 41326 42055 41382 42064
rect 41236 40044 41288 40050
rect 41236 39986 41288 39992
rect 41696 39976 41748 39982
rect 41696 39918 41748 39924
rect 41420 39364 41472 39370
rect 41420 39306 41472 39312
rect 41432 39098 41460 39306
rect 41420 39092 41472 39098
rect 41420 39034 41472 39040
rect 41708 38758 41736 39918
rect 41880 39908 41932 39914
rect 41880 39850 41932 39856
rect 41892 39030 41920 39850
rect 42076 39098 42104 43182
rect 42950 43004 43258 43013
rect 42950 43002 42956 43004
rect 43012 43002 43036 43004
rect 43092 43002 43116 43004
rect 43172 43002 43196 43004
rect 43252 43002 43258 43004
rect 43012 42950 43014 43002
rect 43194 42950 43196 43002
rect 42950 42948 42956 42950
rect 43012 42948 43036 42950
rect 43092 42948 43116 42950
rect 43172 42948 43196 42950
rect 43252 42948 43258 42950
rect 42950 42939 43258 42948
rect 42950 41916 43258 41925
rect 42950 41914 42956 41916
rect 43012 41914 43036 41916
rect 43092 41914 43116 41916
rect 43172 41914 43196 41916
rect 43252 41914 43258 41916
rect 43012 41862 43014 41914
rect 43194 41862 43196 41914
rect 42950 41860 42956 41862
rect 43012 41860 43036 41862
rect 43092 41860 43116 41862
rect 43172 41860 43196 41862
rect 43252 41860 43258 41862
rect 42950 41851 43258 41860
rect 42950 40828 43258 40837
rect 42950 40826 42956 40828
rect 43012 40826 43036 40828
rect 43092 40826 43116 40828
rect 43172 40826 43196 40828
rect 43252 40826 43258 40828
rect 43012 40774 43014 40826
rect 43194 40774 43196 40826
rect 42950 40772 42956 40774
rect 43012 40772 43036 40774
rect 43092 40772 43116 40774
rect 43172 40772 43196 40774
rect 43252 40772 43258 40774
rect 42950 40763 43258 40772
rect 42432 40180 42484 40186
rect 42432 40122 42484 40128
rect 42064 39092 42116 39098
rect 42064 39034 42116 39040
rect 41880 39024 41932 39030
rect 41880 38966 41932 38972
rect 41236 38752 41288 38758
rect 41236 38694 41288 38700
rect 41696 38752 41748 38758
rect 41696 38694 41748 38700
rect 41144 38548 41196 38554
rect 41144 38490 41196 38496
rect 41052 38344 41104 38350
rect 41052 38286 41104 38292
rect 41248 38010 41276 38694
rect 41512 38344 41564 38350
rect 41512 38286 41564 38292
rect 41236 38004 41288 38010
rect 41236 37946 41288 37952
rect 40960 37664 41012 37670
rect 40960 37606 41012 37612
rect 41420 37664 41472 37670
rect 41420 37606 41472 37612
rect 40972 36718 41000 37606
rect 41236 36780 41288 36786
rect 41236 36722 41288 36728
rect 40960 36712 41012 36718
rect 40960 36654 41012 36660
rect 41248 36378 41276 36722
rect 41236 36372 41288 36378
rect 41236 36314 41288 36320
rect 41328 36032 41380 36038
rect 41328 35974 41380 35980
rect 41142 35864 41198 35873
rect 41142 35799 41198 35808
rect 40960 35624 41012 35630
rect 40960 35566 41012 35572
rect 40868 34604 40920 34610
rect 40868 34546 40920 34552
rect 40776 34400 40828 34406
rect 40776 34342 40828 34348
rect 40592 32904 40644 32910
rect 40592 32846 40644 32852
rect 40684 32904 40736 32910
rect 40684 32846 40736 32852
rect 40500 32768 40552 32774
rect 40500 32710 40552 32716
rect 40316 31884 40368 31890
rect 40316 31826 40368 31832
rect 40224 31748 40276 31754
rect 40224 31690 40276 31696
rect 40224 31476 40276 31482
rect 40224 31418 40276 31424
rect 40236 30870 40264 31418
rect 40408 31136 40460 31142
rect 40408 31078 40460 31084
rect 40500 31136 40552 31142
rect 40500 31078 40552 31084
rect 40224 30864 40276 30870
rect 40224 30806 40276 30812
rect 40316 30864 40368 30870
rect 40316 30806 40368 30812
rect 40236 30258 40264 30806
rect 40224 30252 40276 30258
rect 40224 30194 40276 30200
rect 40328 30054 40356 30806
rect 40420 30734 40448 31078
rect 40512 30938 40540 31078
rect 40500 30932 40552 30938
rect 40500 30874 40552 30880
rect 40408 30728 40460 30734
rect 40408 30670 40460 30676
rect 40316 30048 40368 30054
rect 40316 29990 40368 29996
rect 40328 29714 40356 29990
rect 40316 29708 40368 29714
rect 40316 29650 40368 29656
rect 40328 28626 40356 29650
rect 40788 29170 40816 34342
rect 40972 33318 41000 35566
rect 41156 34785 41184 35799
rect 41142 34776 41198 34785
rect 41142 34711 41198 34720
rect 40960 33312 41012 33318
rect 40960 33254 41012 33260
rect 40868 33108 40920 33114
rect 40868 33050 40920 33056
rect 40880 33017 40908 33050
rect 40866 33008 40922 33017
rect 40866 32943 40922 32952
rect 40960 32768 41012 32774
rect 40960 32710 41012 32716
rect 40776 29164 40828 29170
rect 40776 29106 40828 29112
rect 40316 28620 40368 28626
rect 40316 28562 40368 28568
rect 40684 28620 40736 28626
rect 40684 28562 40736 28568
rect 40132 28484 40184 28490
rect 40132 28426 40184 28432
rect 40316 28416 40368 28422
rect 40316 28358 40368 28364
rect 40040 27532 40092 27538
rect 40040 27474 40092 27480
rect 40052 26994 40080 27474
rect 40040 26988 40092 26994
rect 40040 26930 40092 26936
rect 40052 26450 40080 26930
rect 40040 26444 40092 26450
rect 40040 26386 40092 26392
rect 39948 26036 40000 26042
rect 39948 25978 40000 25984
rect 39580 25832 39632 25838
rect 39580 25774 39632 25780
rect 39672 25832 39724 25838
rect 39672 25774 39724 25780
rect 39488 25492 39540 25498
rect 39488 25434 39540 25440
rect 39500 24750 39528 25434
rect 39488 24744 39540 24750
rect 39488 24686 39540 24692
rect 39212 24064 39264 24070
rect 39212 24006 39264 24012
rect 38568 23860 38620 23866
rect 38568 23802 38620 23808
rect 38568 23724 38620 23730
rect 38568 23666 38620 23672
rect 38580 22778 38608 23666
rect 39488 23656 39540 23662
rect 39488 23598 39540 23604
rect 38752 23520 38804 23526
rect 38752 23462 38804 23468
rect 38764 23186 38792 23462
rect 38752 23180 38804 23186
rect 38752 23122 38804 23128
rect 38568 22772 38620 22778
rect 38568 22714 38620 22720
rect 38476 21956 38528 21962
rect 38476 21898 38528 21904
rect 38580 21570 38608 22714
rect 38764 21622 38792 23122
rect 39028 22636 39080 22642
rect 39028 22578 39080 22584
rect 39040 21622 39068 22578
rect 39500 22574 39528 23598
rect 39592 23526 39620 25774
rect 39684 25226 39712 25774
rect 39672 25220 39724 25226
rect 39672 25162 39724 25168
rect 39684 23798 39712 25162
rect 40040 25152 40092 25158
rect 40040 25094 40092 25100
rect 40052 24206 40080 25094
rect 40328 24274 40356 28358
rect 40408 27396 40460 27402
rect 40408 27338 40460 27344
rect 40420 26042 40448 27338
rect 40696 27130 40724 28562
rect 40972 28558 41000 32710
rect 41156 30326 41184 34711
rect 41340 33998 41368 35974
rect 41432 35222 41460 37606
rect 41524 37330 41552 38286
rect 41708 38282 41736 38694
rect 41696 38276 41748 38282
rect 41696 38218 41748 38224
rect 41512 37324 41564 37330
rect 41512 37266 41564 37272
rect 41708 36242 41736 38218
rect 41786 36272 41842 36281
rect 41696 36236 41748 36242
rect 41786 36207 41788 36216
rect 41696 36178 41748 36184
rect 41840 36207 41842 36216
rect 41880 36236 41932 36242
rect 41788 36178 41840 36184
rect 41880 36178 41932 36184
rect 41604 36168 41656 36174
rect 41604 36110 41656 36116
rect 41420 35216 41472 35222
rect 41420 35158 41472 35164
rect 41420 34944 41472 34950
rect 41420 34886 41472 34892
rect 41432 34746 41460 34886
rect 41420 34740 41472 34746
rect 41420 34682 41472 34688
rect 41328 33992 41380 33998
rect 41328 33934 41380 33940
rect 41328 32836 41380 32842
rect 41328 32778 41380 32784
rect 41420 32836 41472 32842
rect 41420 32778 41472 32784
rect 41340 32570 41368 32778
rect 41328 32564 41380 32570
rect 41328 32506 41380 32512
rect 41432 32502 41460 32778
rect 41512 32564 41564 32570
rect 41512 32506 41564 32512
rect 41420 32496 41472 32502
rect 41420 32438 41472 32444
rect 41328 32292 41380 32298
rect 41328 32234 41380 32240
rect 41340 31482 41368 32234
rect 41524 31822 41552 32506
rect 41512 31816 41564 31822
rect 41512 31758 41564 31764
rect 41512 31680 41564 31686
rect 41512 31622 41564 31628
rect 41328 31476 41380 31482
rect 41328 31418 41380 31424
rect 41524 30734 41552 31622
rect 41616 30734 41644 36110
rect 41788 34944 41840 34950
rect 41788 34886 41840 34892
rect 41800 34610 41828 34886
rect 41788 34604 41840 34610
rect 41788 34546 41840 34552
rect 41892 33454 41920 36178
rect 41972 35624 42024 35630
rect 41972 35566 42024 35572
rect 41984 33658 42012 35566
rect 41972 33652 42024 33658
rect 41972 33594 42024 33600
rect 41880 33448 41932 33454
rect 41880 33390 41932 33396
rect 41984 32910 42012 33594
rect 42076 32978 42104 39034
rect 42248 37868 42300 37874
rect 42248 37810 42300 37816
rect 42156 34128 42208 34134
rect 42156 34070 42208 34076
rect 42168 33318 42196 34070
rect 42260 33998 42288 37810
rect 42444 36922 42472 40122
rect 42950 39740 43258 39749
rect 42950 39738 42956 39740
rect 43012 39738 43036 39740
rect 43092 39738 43116 39740
rect 43172 39738 43196 39740
rect 43252 39738 43258 39740
rect 43012 39686 43014 39738
rect 43194 39686 43196 39738
rect 42950 39684 42956 39686
rect 43012 39684 43036 39686
rect 43092 39684 43116 39686
rect 43172 39684 43196 39686
rect 43252 39684 43258 39686
rect 42950 39675 43258 39684
rect 42800 39500 42852 39506
rect 42800 39442 42852 39448
rect 42616 39364 42668 39370
rect 42616 39306 42668 39312
rect 42628 39030 42656 39306
rect 42616 39024 42668 39030
rect 42616 38966 42668 38972
rect 42628 38298 42656 38966
rect 42812 38554 42840 39442
rect 42950 38652 43258 38661
rect 42950 38650 42956 38652
rect 43012 38650 43036 38652
rect 43092 38650 43116 38652
rect 43172 38650 43196 38652
rect 43252 38650 43258 38652
rect 43012 38598 43014 38650
rect 43194 38598 43196 38650
rect 42950 38596 42956 38598
rect 43012 38596 43036 38598
rect 43092 38596 43116 38598
rect 43172 38596 43196 38598
rect 43252 38596 43258 38598
rect 42950 38587 43258 38596
rect 42800 38548 42852 38554
rect 42800 38490 42852 38496
rect 43352 38548 43404 38554
rect 43352 38490 43404 38496
rect 43168 38412 43220 38418
rect 43168 38354 43220 38360
rect 42800 38344 42852 38350
rect 42628 38292 42800 38298
rect 42628 38286 42852 38292
rect 42628 38270 42840 38286
rect 42800 38004 42852 38010
rect 42800 37946 42852 37952
rect 42524 37324 42576 37330
rect 42524 37266 42576 37272
rect 42432 36916 42484 36922
rect 42432 36858 42484 36864
rect 42340 36848 42392 36854
rect 42338 36816 42340 36825
rect 42392 36816 42394 36825
rect 42338 36751 42394 36760
rect 42536 35698 42564 37266
rect 42812 36174 42840 37946
rect 43180 37806 43208 38354
rect 43260 38276 43312 38282
rect 43260 38218 43312 38224
rect 43272 37942 43300 38218
rect 43260 37936 43312 37942
rect 43260 37878 43312 37884
rect 43168 37800 43220 37806
rect 43168 37742 43220 37748
rect 42950 37564 43258 37573
rect 42950 37562 42956 37564
rect 43012 37562 43036 37564
rect 43092 37562 43116 37564
rect 43172 37562 43196 37564
rect 43252 37562 43258 37564
rect 43012 37510 43014 37562
rect 43194 37510 43196 37562
rect 42950 37508 42956 37510
rect 43012 37508 43036 37510
rect 43092 37508 43116 37510
rect 43172 37508 43196 37510
rect 43252 37508 43258 37510
rect 42950 37499 43258 37508
rect 43364 36718 43392 38490
rect 43456 38010 43484 44134
rect 43536 42016 43588 42022
rect 43536 41958 43588 41964
rect 43444 38004 43496 38010
rect 43444 37946 43496 37952
rect 43444 37120 43496 37126
rect 43444 37062 43496 37068
rect 43352 36712 43404 36718
rect 43352 36654 43404 36660
rect 42950 36476 43258 36485
rect 42950 36474 42956 36476
rect 43012 36474 43036 36476
rect 43092 36474 43116 36476
rect 43172 36474 43196 36476
rect 43252 36474 43258 36476
rect 43012 36422 43014 36474
rect 43194 36422 43196 36474
rect 42950 36420 42956 36422
rect 43012 36420 43036 36422
rect 43092 36420 43116 36422
rect 43172 36420 43196 36422
rect 43252 36420 43258 36422
rect 42950 36411 43258 36420
rect 43352 36236 43404 36242
rect 43352 36178 43404 36184
rect 42800 36168 42852 36174
rect 42800 36110 42852 36116
rect 42800 36032 42852 36038
rect 42800 35974 42852 35980
rect 42892 36032 42944 36038
rect 42892 35974 42944 35980
rect 43260 36032 43312 36038
rect 43260 35974 43312 35980
rect 42524 35692 42576 35698
rect 42524 35634 42576 35640
rect 42536 35154 42564 35634
rect 42524 35148 42576 35154
rect 42524 35090 42576 35096
rect 42812 34678 42840 35974
rect 42904 35494 42932 35974
rect 43272 35894 43300 35974
rect 43180 35866 43300 35894
rect 43180 35766 43208 35866
rect 43168 35760 43220 35766
rect 43168 35702 43220 35708
rect 43364 35494 43392 36178
rect 43456 35894 43484 37062
rect 43548 36174 43576 41958
rect 43536 36168 43588 36174
rect 43536 36110 43588 36116
rect 43456 35866 43576 35894
rect 42892 35488 42944 35494
rect 42892 35430 42944 35436
rect 43352 35488 43404 35494
rect 43352 35430 43404 35436
rect 42950 35388 43258 35397
rect 42950 35386 42956 35388
rect 43012 35386 43036 35388
rect 43092 35386 43116 35388
rect 43172 35386 43196 35388
rect 43252 35386 43258 35388
rect 43012 35334 43014 35386
rect 43194 35334 43196 35386
rect 42950 35332 42956 35334
rect 43012 35332 43036 35334
rect 43092 35332 43116 35334
rect 43172 35332 43196 35334
rect 43252 35332 43258 35334
rect 42950 35323 43258 35332
rect 43364 35154 43392 35430
rect 43548 35154 43576 35866
rect 43640 35306 43668 53994
rect 44180 53984 44232 53990
rect 44180 53926 44232 53932
rect 46388 53984 46440 53990
rect 46388 53926 46440 53932
rect 44192 42702 44220 53926
rect 46112 53576 46164 53582
rect 46112 53518 46164 53524
rect 46124 53242 46152 53518
rect 46112 53236 46164 53242
rect 46112 53178 46164 53184
rect 46204 49972 46256 49978
rect 46204 49914 46256 49920
rect 44180 42696 44232 42702
rect 44180 42638 44232 42644
rect 43904 42152 43956 42158
rect 43904 42094 43956 42100
rect 43720 38208 43772 38214
rect 43720 38150 43772 38156
rect 43732 38010 43760 38150
rect 43720 38004 43772 38010
rect 43720 37946 43772 37952
rect 43812 37732 43864 37738
rect 43812 37674 43864 37680
rect 43720 37120 43772 37126
rect 43720 37062 43772 37068
rect 43732 36786 43760 37062
rect 43720 36780 43772 36786
rect 43720 36722 43772 36728
rect 43640 35278 43760 35306
rect 43352 35148 43404 35154
rect 43352 35090 43404 35096
rect 43536 35148 43588 35154
rect 43536 35090 43588 35096
rect 42800 34672 42852 34678
rect 42800 34614 42852 34620
rect 43548 34542 43576 35090
rect 43628 34944 43680 34950
rect 43628 34886 43680 34892
rect 43640 34678 43668 34886
rect 43628 34672 43680 34678
rect 43628 34614 43680 34620
rect 43352 34536 43404 34542
rect 43352 34478 43404 34484
rect 43444 34536 43496 34542
rect 43444 34478 43496 34484
rect 43536 34536 43588 34542
rect 43536 34478 43588 34484
rect 42950 34300 43258 34309
rect 42950 34298 42956 34300
rect 43012 34298 43036 34300
rect 43092 34298 43116 34300
rect 43172 34298 43196 34300
rect 43252 34298 43258 34300
rect 43012 34246 43014 34298
rect 43194 34246 43196 34298
rect 42950 34244 42956 34246
rect 43012 34244 43036 34246
rect 43092 34244 43116 34246
rect 43172 34244 43196 34246
rect 43252 34244 43258 34246
rect 42950 34235 43258 34244
rect 42248 33992 42300 33998
rect 42248 33934 42300 33940
rect 42616 33584 42668 33590
rect 42616 33526 42668 33532
rect 42156 33312 42208 33318
rect 42156 33254 42208 33260
rect 42064 32972 42116 32978
rect 42064 32914 42116 32920
rect 41972 32904 42024 32910
rect 41972 32846 42024 32852
rect 42168 32366 42196 33254
rect 42248 32972 42300 32978
rect 42248 32914 42300 32920
rect 42156 32360 42208 32366
rect 42156 32302 42208 32308
rect 42168 31346 42196 32302
rect 42156 31340 42208 31346
rect 42156 31282 42208 31288
rect 41512 30728 41564 30734
rect 41512 30670 41564 30676
rect 41604 30728 41656 30734
rect 41604 30670 41656 30676
rect 41236 30592 41288 30598
rect 41236 30534 41288 30540
rect 41144 30320 41196 30326
rect 41144 30262 41196 30268
rect 41248 29306 41276 30534
rect 41236 29300 41288 29306
rect 41236 29242 41288 29248
rect 41144 29164 41196 29170
rect 41144 29106 41196 29112
rect 41156 28762 41184 29106
rect 41144 28756 41196 28762
rect 41144 28698 41196 28704
rect 40960 28552 41012 28558
rect 40960 28494 41012 28500
rect 41604 27396 41656 27402
rect 41604 27338 41656 27344
rect 40960 27328 41012 27334
rect 40960 27270 41012 27276
rect 41052 27328 41104 27334
rect 41052 27270 41104 27276
rect 40684 27124 40736 27130
rect 40684 27066 40736 27072
rect 40500 26580 40552 26586
rect 40500 26522 40552 26528
rect 40408 26036 40460 26042
rect 40408 25978 40460 25984
rect 40512 25362 40540 26522
rect 40696 25974 40724 27066
rect 40972 26586 41000 27270
rect 41064 26790 41092 27270
rect 41616 27062 41644 27338
rect 41604 27056 41656 27062
rect 41604 26998 41656 27004
rect 41052 26784 41104 26790
rect 41052 26726 41104 26732
rect 40960 26580 41012 26586
rect 40960 26522 41012 26528
rect 41616 26314 41644 26998
rect 42260 26926 42288 32914
rect 42628 32502 42656 33526
rect 42950 33212 43258 33221
rect 42950 33210 42956 33212
rect 43012 33210 43036 33212
rect 43092 33210 43116 33212
rect 43172 33210 43196 33212
rect 43252 33210 43258 33212
rect 43012 33158 43014 33210
rect 43194 33158 43196 33210
rect 42950 33156 42956 33158
rect 43012 33156 43036 33158
rect 43092 33156 43116 33158
rect 43172 33156 43196 33158
rect 43252 33156 43258 33158
rect 42950 33147 43258 33156
rect 42616 32496 42668 32502
rect 42616 32438 42668 32444
rect 42628 31754 42656 32438
rect 42800 32224 42852 32230
rect 42800 32166 42852 32172
rect 42708 31884 42760 31890
rect 42708 31826 42760 31832
rect 42616 31748 42668 31754
rect 42616 31690 42668 31696
rect 42628 29578 42656 31690
rect 42720 29850 42748 31826
rect 42812 31482 42840 32166
rect 42950 32124 43258 32133
rect 42950 32122 42956 32124
rect 43012 32122 43036 32124
rect 43092 32122 43116 32124
rect 43172 32122 43196 32124
rect 43252 32122 43258 32124
rect 43012 32070 43014 32122
rect 43194 32070 43196 32122
rect 42950 32068 42956 32070
rect 43012 32068 43036 32070
rect 43092 32068 43116 32070
rect 43172 32068 43196 32070
rect 43252 32068 43258 32070
rect 42950 32059 43258 32068
rect 42800 31476 42852 31482
rect 42800 31418 42852 31424
rect 42950 31036 43258 31045
rect 42950 31034 42956 31036
rect 43012 31034 43036 31036
rect 43092 31034 43116 31036
rect 43172 31034 43196 31036
rect 43252 31034 43258 31036
rect 43012 30982 43014 31034
rect 43194 30982 43196 31034
rect 42950 30980 42956 30982
rect 43012 30980 43036 30982
rect 43092 30980 43116 30982
rect 43172 30980 43196 30982
rect 43252 30980 43258 30982
rect 42950 30971 43258 30980
rect 43364 30734 43392 34478
rect 43456 32178 43484 34478
rect 43732 33046 43760 35278
rect 43720 33040 43772 33046
rect 43720 32982 43772 32988
rect 43824 32910 43852 37674
rect 43916 36038 43944 42094
rect 43996 39432 44048 39438
rect 43996 39374 44048 39380
rect 44008 38350 44036 39374
rect 43996 38344 44048 38350
rect 43996 38286 44048 38292
rect 44008 37194 44036 38286
rect 46216 38282 46244 49914
rect 46400 48278 46428 53926
rect 46768 53650 46796 56200
rect 46848 55752 46900 55758
rect 46848 55694 46900 55700
rect 46860 54194 46888 55694
rect 47504 54194 47532 56200
rect 48240 54618 48268 56200
rect 48240 54590 48360 54618
rect 47950 54428 48258 54437
rect 47950 54426 47956 54428
rect 48012 54426 48036 54428
rect 48092 54426 48116 54428
rect 48172 54426 48196 54428
rect 48252 54426 48258 54428
rect 48012 54374 48014 54426
rect 48194 54374 48196 54426
rect 47950 54372 47956 54374
rect 48012 54372 48036 54374
rect 48092 54372 48116 54374
rect 48172 54372 48196 54374
rect 48252 54372 48258 54374
rect 47950 54363 48258 54372
rect 48332 54210 48360 54590
rect 46848 54188 46900 54194
rect 46848 54130 46900 54136
rect 47492 54188 47544 54194
rect 47492 54130 47544 54136
rect 47860 54188 47912 54194
rect 47860 54130 47912 54136
rect 48240 54182 48360 54210
rect 47032 53984 47084 53990
rect 47032 53926 47084 53932
rect 46756 53644 46808 53650
rect 46756 53586 46808 53592
rect 47044 53242 47072 53926
rect 47032 53236 47084 53242
rect 47032 53178 47084 53184
rect 46940 53100 46992 53106
rect 46940 53042 46992 53048
rect 46388 48272 46440 48278
rect 46388 48214 46440 48220
rect 46952 45558 46980 53042
rect 47768 48136 47820 48142
rect 47768 48078 47820 48084
rect 46940 45552 46992 45558
rect 47780 45554 47808 48078
rect 47872 47258 47900 54130
rect 48240 54126 48268 54182
rect 48228 54120 48280 54126
rect 48228 54062 48280 54068
rect 48976 53582 49004 56200
rect 48964 53576 49016 53582
rect 48964 53518 49016 53524
rect 48780 53440 48832 53446
rect 48780 53382 48832 53388
rect 47950 53340 48258 53349
rect 47950 53338 47956 53340
rect 48012 53338 48036 53340
rect 48092 53338 48116 53340
rect 48172 53338 48196 53340
rect 48252 53338 48258 53340
rect 48012 53286 48014 53338
rect 48194 53286 48196 53338
rect 47950 53284 47956 53286
rect 48012 53284 48036 53286
rect 48092 53284 48116 53286
rect 48172 53284 48196 53286
rect 48252 53284 48258 53286
rect 47950 53275 48258 53284
rect 48320 53100 48372 53106
rect 48320 53042 48372 53048
rect 47950 52252 48258 52261
rect 47950 52250 47956 52252
rect 48012 52250 48036 52252
rect 48092 52250 48116 52252
rect 48172 52250 48196 52252
rect 48252 52250 48258 52252
rect 48012 52198 48014 52250
rect 48194 52198 48196 52250
rect 47950 52196 47956 52198
rect 48012 52196 48036 52198
rect 48092 52196 48116 52198
rect 48172 52196 48196 52198
rect 48252 52196 48258 52198
rect 47950 52187 48258 52196
rect 47950 51164 48258 51173
rect 47950 51162 47956 51164
rect 48012 51162 48036 51164
rect 48092 51162 48116 51164
rect 48172 51162 48196 51164
rect 48252 51162 48258 51164
rect 48012 51110 48014 51162
rect 48194 51110 48196 51162
rect 47950 51108 47956 51110
rect 48012 51108 48036 51110
rect 48092 51108 48116 51110
rect 48172 51108 48196 51110
rect 48252 51108 48258 51110
rect 47950 51099 48258 51108
rect 47950 50076 48258 50085
rect 47950 50074 47956 50076
rect 48012 50074 48036 50076
rect 48092 50074 48116 50076
rect 48172 50074 48196 50076
rect 48252 50074 48258 50076
rect 48012 50022 48014 50074
rect 48194 50022 48196 50074
rect 47950 50020 47956 50022
rect 48012 50020 48036 50022
rect 48092 50020 48116 50022
rect 48172 50020 48196 50022
rect 48252 50020 48258 50022
rect 47950 50011 48258 50020
rect 47950 48988 48258 48997
rect 47950 48986 47956 48988
rect 48012 48986 48036 48988
rect 48092 48986 48116 48988
rect 48172 48986 48196 48988
rect 48252 48986 48258 48988
rect 48012 48934 48014 48986
rect 48194 48934 48196 48986
rect 47950 48932 47956 48934
rect 48012 48932 48036 48934
rect 48092 48932 48116 48934
rect 48172 48932 48196 48934
rect 48252 48932 48258 48934
rect 47950 48923 48258 48932
rect 48332 48278 48360 53042
rect 48320 48272 48372 48278
rect 48320 48214 48372 48220
rect 47950 47900 48258 47909
rect 47950 47898 47956 47900
rect 48012 47898 48036 47900
rect 48092 47898 48116 47900
rect 48172 47898 48196 47900
rect 48252 47898 48258 47900
rect 48012 47846 48014 47898
rect 48194 47846 48196 47898
rect 47950 47844 47956 47846
rect 48012 47844 48036 47846
rect 48092 47844 48116 47846
rect 48172 47844 48196 47846
rect 48252 47844 48258 47846
rect 47950 47835 48258 47844
rect 48792 47258 48820 53382
rect 49712 53174 49740 56200
rect 50448 55758 50476 56200
rect 50436 55752 50488 55758
rect 50436 55694 50488 55700
rect 49700 53168 49752 53174
rect 49700 53110 49752 53116
rect 49330 52592 49386 52601
rect 49330 52527 49386 52536
rect 49344 52494 49372 52527
rect 49332 52488 49384 52494
rect 49332 52430 49384 52436
rect 49148 52352 49200 52358
rect 49148 52294 49200 52300
rect 49056 52012 49108 52018
rect 49056 51954 49108 51960
rect 49068 51921 49096 51954
rect 49054 51912 49110 51921
rect 49054 51847 49110 51856
rect 49056 51400 49108 51406
rect 49056 51342 49108 51348
rect 49068 51241 49096 51342
rect 49054 51232 49110 51241
rect 49054 51167 49110 51176
rect 48964 50924 49016 50930
rect 48964 50866 49016 50872
rect 48976 50561 49004 50866
rect 48962 50552 49018 50561
rect 48962 50487 49018 50496
rect 49160 50402 49188 52294
rect 49332 51264 49384 51270
rect 49332 51206 49384 51212
rect 48976 50374 49188 50402
rect 48872 50176 48924 50182
rect 48872 50118 48924 50124
rect 47860 47252 47912 47258
rect 47860 47194 47912 47200
rect 48780 47252 48832 47258
rect 48780 47194 48832 47200
rect 48412 46980 48464 46986
rect 48412 46922 48464 46928
rect 47950 46812 48258 46821
rect 47950 46810 47956 46812
rect 48012 46810 48036 46812
rect 48092 46810 48116 46812
rect 48172 46810 48196 46812
rect 48252 46810 48258 46812
rect 48012 46758 48014 46810
rect 48194 46758 48196 46810
rect 47950 46756 47956 46758
rect 48012 46756 48036 46758
rect 48092 46756 48116 46758
rect 48172 46756 48196 46758
rect 48252 46756 48258 46758
rect 47950 46747 48258 46756
rect 47950 45724 48258 45733
rect 47950 45722 47956 45724
rect 48012 45722 48036 45724
rect 48092 45722 48116 45724
rect 48172 45722 48196 45724
rect 48252 45722 48258 45724
rect 48012 45670 48014 45722
rect 48194 45670 48196 45722
rect 47950 45668 47956 45670
rect 48012 45668 48036 45670
rect 48092 45668 48116 45670
rect 48172 45668 48196 45670
rect 48252 45668 48258 45670
rect 47950 45659 48258 45668
rect 47780 45526 47900 45554
rect 46940 45494 46992 45500
rect 46296 42220 46348 42226
rect 46296 42162 46348 42168
rect 46204 38276 46256 38282
rect 46204 38218 46256 38224
rect 43996 37188 44048 37194
rect 43996 37130 44048 37136
rect 43904 36032 43956 36038
rect 43904 35974 43956 35980
rect 43812 32904 43864 32910
rect 43812 32846 43864 32852
rect 43456 32150 43576 32178
rect 43444 32020 43496 32026
rect 43444 31962 43496 31968
rect 43352 30728 43404 30734
rect 43352 30670 43404 30676
rect 42800 30592 42852 30598
rect 42800 30534 42852 30540
rect 42708 29844 42760 29850
rect 42708 29786 42760 29792
rect 42616 29572 42668 29578
rect 42616 29514 42668 29520
rect 42628 27402 42656 29514
rect 42720 29102 42748 29786
rect 42708 29096 42760 29102
rect 42708 29038 42760 29044
rect 42616 27396 42668 27402
rect 42616 27338 42668 27344
rect 41788 26920 41840 26926
rect 41788 26862 41840 26868
rect 42248 26920 42300 26926
rect 42248 26862 42300 26868
rect 41800 26450 41828 26862
rect 41788 26444 41840 26450
rect 41788 26386 41840 26392
rect 41604 26308 41656 26314
rect 41604 26250 41656 26256
rect 40776 26036 40828 26042
rect 40776 25978 40828 25984
rect 40684 25968 40736 25974
rect 40684 25910 40736 25916
rect 40696 25362 40724 25910
rect 40500 25356 40552 25362
rect 40500 25298 40552 25304
rect 40684 25356 40736 25362
rect 40684 25298 40736 25304
rect 40408 25152 40460 25158
rect 40408 25094 40460 25100
rect 40420 24818 40448 25094
rect 40408 24812 40460 24818
rect 40408 24754 40460 24760
rect 40788 24274 40816 25978
rect 41616 25974 41644 26250
rect 42812 25974 42840 30534
rect 42950 29948 43258 29957
rect 42950 29946 42956 29948
rect 43012 29946 43036 29948
rect 43092 29946 43116 29948
rect 43172 29946 43196 29948
rect 43252 29946 43258 29948
rect 43012 29894 43014 29946
rect 43194 29894 43196 29946
rect 42950 29892 42956 29894
rect 43012 29892 43036 29894
rect 43092 29892 43116 29894
rect 43172 29892 43196 29894
rect 43252 29892 43258 29894
rect 42950 29883 43258 29892
rect 42950 28860 43258 28869
rect 42950 28858 42956 28860
rect 43012 28858 43036 28860
rect 43092 28858 43116 28860
rect 43172 28858 43196 28860
rect 43252 28858 43258 28860
rect 43012 28806 43014 28858
rect 43194 28806 43196 28858
rect 42950 28804 42956 28806
rect 43012 28804 43036 28806
rect 43092 28804 43116 28806
rect 43172 28804 43196 28806
rect 43252 28804 43258 28806
rect 42950 28795 43258 28804
rect 42950 27772 43258 27781
rect 42950 27770 42956 27772
rect 43012 27770 43036 27772
rect 43092 27770 43116 27772
rect 43172 27770 43196 27772
rect 43252 27770 43258 27772
rect 43012 27718 43014 27770
rect 43194 27718 43196 27770
rect 42950 27716 42956 27718
rect 43012 27716 43036 27718
rect 43092 27716 43116 27718
rect 43172 27716 43196 27718
rect 43252 27716 43258 27718
rect 42950 27707 43258 27716
rect 42950 26684 43258 26693
rect 42950 26682 42956 26684
rect 43012 26682 43036 26684
rect 43092 26682 43116 26684
rect 43172 26682 43196 26684
rect 43252 26682 43258 26684
rect 43012 26630 43014 26682
rect 43194 26630 43196 26682
rect 42950 26628 42956 26630
rect 43012 26628 43036 26630
rect 43092 26628 43116 26630
rect 43172 26628 43196 26630
rect 43252 26628 43258 26630
rect 42950 26619 43258 26628
rect 41604 25968 41656 25974
rect 41604 25910 41656 25916
rect 42800 25968 42852 25974
rect 42800 25910 42852 25916
rect 42950 25596 43258 25605
rect 42950 25594 42956 25596
rect 43012 25594 43036 25596
rect 43092 25594 43116 25596
rect 43172 25594 43196 25596
rect 43252 25594 43258 25596
rect 43012 25542 43014 25594
rect 43194 25542 43196 25594
rect 42950 25540 42956 25542
rect 43012 25540 43036 25542
rect 43092 25540 43116 25542
rect 43172 25540 43196 25542
rect 43252 25540 43258 25542
rect 42950 25531 43258 25540
rect 43456 25294 43484 31962
rect 43548 31414 43576 32150
rect 43916 32026 43944 35974
rect 44008 35698 44036 37130
rect 46308 36689 46336 42162
rect 46952 39438 46980 45494
rect 47872 45490 47900 45526
rect 47860 45484 47912 45490
rect 47860 45426 47912 45432
rect 46940 39432 46992 39438
rect 46940 39374 46992 39380
rect 46294 36680 46350 36689
rect 46294 36615 46350 36624
rect 44088 36576 44140 36582
rect 44088 36518 44140 36524
rect 43996 35692 44048 35698
rect 43996 35634 44048 35640
rect 44008 35018 44036 35634
rect 43996 35012 44048 35018
rect 43996 34954 44048 34960
rect 44008 33590 44036 34954
rect 43996 33584 44048 33590
rect 43996 33526 44048 33532
rect 44100 32434 44128 36518
rect 44272 34536 44324 34542
rect 44272 34478 44324 34484
rect 44088 32428 44140 32434
rect 44088 32370 44140 32376
rect 43904 32020 43956 32026
rect 43904 31962 43956 31968
rect 43536 31408 43588 31414
rect 43536 31350 43588 31356
rect 43548 30122 43576 31350
rect 44284 31346 44312 34478
rect 46388 32768 46440 32774
rect 46388 32710 46440 32716
rect 44640 32224 44692 32230
rect 44640 32166 44692 32172
rect 44272 31340 44324 31346
rect 44272 31282 44324 31288
rect 44364 31204 44416 31210
rect 44364 31146 44416 31152
rect 43536 30116 43588 30122
rect 43536 30058 43588 30064
rect 43996 29028 44048 29034
rect 43996 28970 44048 28976
rect 44008 27470 44036 28970
rect 43996 27464 44048 27470
rect 43996 27406 44048 27412
rect 43720 27328 43772 27334
rect 43720 27270 43772 27276
rect 43812 27328 43864 27334
rect 43812 27270 43864 27276
rect 43732 26450 43760 27270
rect 43720 26444 43772 26450
rect 43720 26386 43772 26392
rect 43824 26382 43852 27270
rect 43812 26376 43864 26382
rect 43812 26318 43864 26324
rect 43444 25288 43496 25294
rect 43444 25230 43496 25236
rect 44376 25226 44404 31146
rect 44652 27062 44680 32166
rect 45560 31204 45612 31210
rect 45560 31146 45612 31152
rect 45468 30592 45520 30598
rect 45468 30534 45520 30540
rect 44640 27056 44692 27062
rect 44640 26998 44692 27004
rect 45480 26994 45508 30534
rect 45468 26988 45520 26994
rect 45468 26930 45520 26936
rect 45572 25294 45600 31146
rect 46020 30660 46072 30666
rect 46020 30602 46072 30608
rect 46032 25906 46060 30602
rect 46400 27470 46428 32710
rect 47124 32564 47176 32570
rect 47124 32506 47176 32512
rect 47136 31890 47164 32506
rect 47124 31884 47176 31890
rect 47124 31826 47176 31832
rect 47872 31754 47900 45426
rect 47950 44636 48258 44645
rect 47950 44634 47956 44636
rect 48012 44634 48036 44636
rect 48092 44634 48116 44636
rect 48172 44634 48196 44636
rect 48252 44634 48258 44636
rect 48012 44582 48014 44634
rect 48194 44582 48196 44634
rect 47950 44580 47956 44582
rect 48012 44580 48036 44582
rect 48092 44580 48116 44582
rect 48172 44580 48196 44582
rect 48252 44580 48258 44582
rect 47950 44571 48258 44580
rect 47950 43548 48258 43557
rect 47950 43546 47956 43548
rect 48012 43546 48036 43548
rect 48092 43546 48116 43548
rect 48172 43546 48196 43548
rect 48252 43546 48258 43548
rect 48012 43494 48014 43546
rect 48194 43494 48196 43546
rect 47950 43492 47956 43494
rect 48012 43492 48036 43494
rect 48092 43492 48116 43494
rect 48172 43492 48196 43494
rect 48252 43492 48258 43494
rect 47950 43483 48258 43492
rect 47950 42460 48258 42469
rect 47950 42458 47956 42460
rect 48012 42458 48036 42460
rect 48092 42458 48116 42460
rect 48172 42458 48196 42460
rect 48252 42458 48258 42460
rect 48012 42406 48014 42458
rect 48194 42406 48196 42458
rect 47950 42404 47956 42406
rect 48012 42404 48036 42406
rect 48092 42404 48116 42406
rect 48172 42404 48196 42406
rect 48252 42404 48258 42406
rect 47950 42395 48258 42404
rect 48424 41614 48452 46922
rect 48688 46368 48740 46374
rect 48688 46310 48740 46316
rect 48596 45960 48648 45966
rect 48596 45902 48648 45908
rect 48608 45626 48636 45902
rect 48596 45620 48648 45626
rect 48596 45562 48648 45568
rect 48504 44872 48556 44878
rect 48504 44814 48556 44820
rect 48516 44441 48544 44814
rect 48502 44432 48558 44441
rect 48502 44367 48558 44376
rect 48504 43784 48556 43790
rect 48502 43752 48504 43761
rect 48556 43752 48558 43761
rect 48502 43687 48558 43696
rect 48504 43240 48556 43246
rect 48504 43182 48556 43188
rect 48516 43081 48544 43182
rect 48502 43072 48558 43081
rect 48502 43007 48558 43016
rect 48504 42696 48556 42702
rect 48504 42638 48556 42644
rect 48516 42401 48544 42638
rect 48502 42392 48558 42401
rect 48502 42327 48558 42336
rect 48504 42152 48556 42158
rect 48504 42094 48556 42100
rect 48516 41721 48544 42094
rect 48700 41818 48728 46310
rect 48884 45554 48912 50118
rect 48976 47002 49004 50374
rect 49056 50312 49108 50318
rect 49056 50254 49108 50260
rect 49068 49881 49096 50254
rect 49054 49872 49110 49881
rect 49054 49807 49110 49816
rect 49148 49836 49200 49842
rect 49148 49778 49200 49784
rect 49160 49201 49188 49778
rect 49240 49224 49292 49230
rect 49146 49192 49202 49201
rect 49240 49166 49292 49172
rect 49146 49127 49202 49136
rect 49056 48748 49108 48754
rect 49056 48690 49108 48696
rect 49068 47841 49096 48690
rect 49252 48521 49280 49166
rect 49238 48512 49294 48521
rect 49238 48447 49294 48456
rect 49344 48362 49372 51206
rect 49252 48334 49372 48362
rect 49054 47832 49110 47841
rect 49054 47767 49110 47776
rect 49056 47660 49108 47666
rect 49056 47602 49108 47608
rect 49068 47161 49096 47602
rect 49054 47152 49110 47161
rect 49054 47087 49110 47096
rect 48976 46974 49096 47002
rect 48884 45526 49004 45554
rect 48688 41812 48740 41818
rect 48688 41754 48740 41760
rect 48502 41712 48558 41721
rect 48502 41647 48558 41656
rect 48412 41608 48464 41614
rect 48412 41550 48464 41556
rect 47950 41372 48258 41381
rect 47950 41370 47956 41372
rect 48012 41370 48036 41372
rect 48092 41370 48116 41372
rect 48172 41370 48196 41372
rect 48252 41370 48258 41372
rect 48012 41318 48014 41370
rect 48194 41318 48196 41370
rect 47950 41316 47956 41318
rect 48012 41316 48036 41318
rect 48092 41316 48116 41318
rect 48172 41316 48196 41318
rect 48252 41316 48258 41318
rect 47950 41307 48258 41316
rect 47950 40284 48258 40293
rect 47950 40282 47956 40284
rect 48012 40282 48036 40284
rect 48092 40282 48116 40284
rect 48172 40282 48196 40284
rect 48252 40282 48258 40284
rect 48012 40230 48014 40282
rect 48194 40230 48196 40282
rect 47950 40228 47956 40230
rect 48012 40228 48036 40230
rect 48092 40228 48116 40230
rect 48172 40228 48196 40230
rect 48252 40228 48258 40230
rect 47950 40219 48258 40228
rect 47950 39196 48258 39205
rect 47950 39194 47956 39196
rect 48012 39194 48036 39196
rect 48092 39194 48116 39196
rect 48172 39194 48196 39196
rect 48252 39194 48258 39196
rect 48012 39142 48014 39194
rect 48194 39142 48196 39194
rect 47950 39140 47956 39142
rect 48012 39140 48036 39142
rect 48092 39140 48116 39142
rect 48172 39140 48196 39142
rect 48252 39140 48258 39142
rect 47950 39131 48258 39140
rect 47950 38108 48258 38117
rect 47950 38106 47956 38108
rect 48012 38106 48036 38108
rect 48092 38106 48116 38108
rect 48172 38106 48196 38108
rect 48252 38106 48258 38108
rect 48012 38054 48014 38106
rect 48194 38054 48196 38106
rect 47950 38052 47956 38054
rect 48012 38052 48036 38054
rect 48092 38052 48116 38054
rect 48172 38052 48196 38054
rect 48252 38052 48258 38054
rect 47950 38043 48258 38052
rect 47950 37020 48258 37029
rect 47950 37018 47956 37020
rect 48012 37018 48036 37020
rect 48092 37018 48116 37020
rect 48172 37018 48196 37020
rect 48252 37018 48258 37020
rect 48012 36966 48014 37018
rect 48194 36966 48196 37018
rect 47950 36964 47956 36966
rect 48012 36964 48036 36966
rect 48092 36964 48116 36966
rect 48172 36964 48196 36966
rect 48252 36964 48258 36966
rect 47950 36955 48258 36964
rect 47950 35932 48258 35941
rect 47950 35930 47956 35932
rect 48012 35930 48036 35932
rect 48092 35930 48116 35932
rect 48172 35930 48196 35932
rect 48252 35930 48258 35932
rect 48012 35878 48014 35930
rect 48194 35878 48196 35930
rect 47950 35876 47956 35878
rect 48012 35876 48036 35878
rect 48092 35876 48116 35878
rect 48172 35876 48196 35878
rect 48252 35876 48258 35878
rect 47950 35867 48258 35876
rect 47950 34844 48258 34853
rect 47950 34842 47956 34844
rect 48012 34842 48036 34844
rect 48092 34842 48116 34844
rect 48172 34842 48196 34844
rect 48252 34842 48258 34844
rect 48012 34790 48014 34842
rect 48194 34790 48196 34842
rect 47950 34788 47956 34790
rect 48012 34788 48036 34790
rect 48092 34788 48116 34790
rect 48172 34788 48196 34790
rect 48252 34788 48258 34790
rect 47950 34779 48258 34788
rect 48320 33924 48372 33930
rect 48320 33866 48372 33872
rect 47950 33756 48258 33765
rect 47950 33754 47956 33756
rect 48012 33754 48036 33756
rect 48092 33754 48116 33756
rect 48172 33754 48196 33756
rect 48252 33754 48258 33756
rect 48012 33702 48014 33754
rect 48194 33702 48196 33754
rect 47950 33700 47956 33702
rect 48012 33700 48036 33702
rect 48092 33700 48116 33702
rect 48172 33700 48196 33702
rect 48252 33700 48258 33702
rect 47950 33691 48258 33700
rect 47950 32668 48258 32677
rect 47950 32666 47956 32668
rect 48012 32666 48036 32668
rect 48092 32666 48116 32668
rect 48172 32666 48196 32668
rect 48252 32666 48258 32668
rect 48012 32614 48014 32666
rect 48194 32614 48196 32666
rect 47950 32612 47956 32614
rect 48012 32612 48036 32614
rect 48092 32612 48116 32614
rect 48172 32612 48196 32614
rect 48252 32612 48258 32614
rect 47950 32603 48258 32612
rect 47780 31726 47900 31754
rect 46388 27464 46440 27470
rect 46388 27406 46440 27412
rect 47584 27396 47636 27402
rect 47584 27338 47636 27344
rect 46848 26784 46900 26790
rect 46848 26726 46900 26732
rect 46020 25900 46072 25906
rect 46020 25842 46072 25848
rect 46204 25764 46256 25770
rect 46204 25706 46256 25712
rect 45560 25288 45612 25294
rect 45560 25230 45612 25236
rect 44364 25220 44416 25226
rect 44364 25162 44416 25168
rect 45468 25220 45520 25226
rect 45468 25162 45520 25168
rect 44456 25152 44508 25158
rect 44456 25094 44508 25100
rect 42950 24508 43258 24517
rect 42950 24506 42956 24508
rect 43012 24506 43036 24508
rect 43092 24506 43116 24508
rect 43172 24506 43196 24508
rect 43252 24506 43258 24508
rect 43012 24454 43014 24506
rect 43194 24454 43196 24506
rect 42950 24452 42956 24454
rect 43012 24452 43036 24454
rect 43092 24452 43116 24454
rect 43172 24452 43196 24454
rect 43252 24452 43258 24454
rect 42950 24443 43258 24452
rect 40316 24268 40368 24274
rect 40316 24210 40368 24216
rect 40776 24268 40828 24274
rect 40776 24210 40828 24216
rect 40040 24200 40092 24206
rect 40040 24142 40092 24148
rect 40040 24064 40092 24070
rect 40040 24006 40092 24012
rect 39672 23792 39724 23798
rect 39672 23734 39724 23740
rect 39580 23520 39632 23526
rect 39580 23462 39632 23468
rect 39684 22778 39712 23734
rect 39672 22772 39724 22778
rect 39672 22714 39724 22720
rect 39488 22568 39540 22574
rect 39488 22510 39540 22516
rect 38488 21554 38608 21570
rect 38752 21616 38804 21622
rect 38752 21558 38804 21564
rect 39028 21616 39080 21622
rect 39028 21558 39080 21564
rect 38476 21548 38608 21554
rect 38528 21542 38608 21548
rect 38476 21490 38528 21496
rect 38568 21344 38620 21350
rect 38568 21286 38620 21292
rect 38476 19508 38528 19514
rect 38476 19450 38528 19456
rect 38488 18222 38516 19450
rect 38476 18216 38528 18222
rect 38476 18158 38528 18164
rect 38580 17746 38608 21286
rect 39040 19446 39068 21558
rect 39948 20256 40000 20262
rect 39948 20198 40000 20204
rect 39028 19440 39080 19446
rect 39028 19382 39080 19388
rect 38660 18692 38712 18698
rect 38660 18634 38712 18640
rect 38568 17740 38620 17746
rect 38568 17682 38620 17688
rect 38672 17610 38700 18634
rect 38660 17604 38712 17610
rect 38660 17546 38712 17552
rect 38672 17338 38700 17546
rect 39960 17542 39988 20198
rect 39948 17536 40000 17542
rect 39948 17478 40000 17484
rect 38660 17332 38712 17338
rect 38660 17274 38712 17280
rect 40052 16114 40080 24006
rect 42950 23420 43258 23429
rect 42950 23418 42956 23420
rect 43012 23418 43036 23420
rect 43092 23418 43116 23420
rect 43172 23418 43196 23420
rect 43252 23418 43258 23420
rect 43012 23366 43014 23418
rect 43194 23366 43196 23418
rect 42950 23364 42956 23366
rect 43012 23364 43036 23366
rect 43092 23364 43116 23366
rect 43172 23364 43196 23366
rect 43252 23364 43258 23366
rect 42950 23355 43258 23364
rect 41236 23316 41288 23322
rect 41236 23258 41288 23264
rect 41248 19854 41276 23258
rect 42950 22332 43258 22341
rect 42950 22330 42956 22332
rect 43012 22330 43036 22332
rect 43092 22330 43116 22332
rect 43172 22330 43196 22332
rect 43252 22330 43258 22332
rect 43012 22278 43014 22330
rect 43194 22278 43196 22330
rect 42950 22276 42956 22278
rect 43012 22276 43036 22278
rect 43092 22276 43116 22278
rect 43172 22276 43196 22278
rect 43252 22276 43258 22278
rect 42950 22267 43258 22276
rect 43812 21956 43864 21962
rect 43812 21898 43864 21904
rect 41328 21888 41380 21894
rect 41328 21830 41380 21836
rect 41236 19848 41288 19854
rect 41236 19790 41288 19796
rect 41340 18766 41368 21830
rect 43824 21622 43852 21898
rect 43812 21616 43864 21622
rect 43812 21558 43864 21564
rect 42950 21244 43258 21253
rect 42950 21242 42956 21244
rect 43012 21242 43036 21244
rect 43092 21242 43116 21244
rect 43172 21242 43196 21244
rect 43252 21242 43258 21244
rect 43012 21190 43014 21242
rect 43194 21190 43196 21242
rect 42950 21188 42956 21190
rect 43012 21188 43036 21190
rect 43092 21188 43116 21190
rect 43172 21188 43196 21190
rect 43252 21188 43258 21190
rect 42950 21179 43258 21188
rect 43720 21072 43772 21078
rect 43720 21014 43772 21020
rect 42950 20156 43258 20165
rect 42950 20154 42956 20156
rect 43012 20154 43036 20156
rect 43092 20154 43116 20156
rect 43172 20154 43196 20156
rect 43252 20154 43258 20156
rect 43012 20102 43014 20154
rect 43194 20102 43196 20154
rect 42950 20100 42956 20102
rect 43012 20100 43036 20102
rect 43092 20100 43116 20102
rect 43172 20100 43196 20102
rect 43252 20100 43258 20102
rect 42950 20091 43258 20100
rect 42950 19068 43258 19077
rect 42950 19066 42956 19068
rect 43012 19066 43036 19068
rect 43092 19066 43116 19068
rect 43172 19066 43196 19068
rect 43252 19066 43258 19068
rect 43012 19014 43014 19066
rect 43194 19014 43196 19066
rect 42950 19012 42956 19014
rect 43012 19012 43036 19014
rect 43092 19012 43116 19014
rect 43172 19012 43196 19014
rect 43252 19012 43258 19014
rect 42950 19003 43258 19012
rect 41328 18760 41380 18766
rect 41328 18702 41380 18708
rect 41788 18080 41840 18086
rect 41788 18022 41840 18028
rect 40224 17060 40276 17066
rect 40224 17002 40276 17008
rect 40132 16516 40184 16522
rect 40132 16458 40184 16464
rect 40040 16108 40092 16114
rect 40040 16050 40092 16056
rect 39120 15972 39172 15978
rect 39120 15914 39172 15920
rect 38384 14000 38436 14006
rect 38384 13942 38436 13948
rect 38936 14000 38988 14006
rect 38936 13942 38988 13948
rect 38476 13864 38528 13870
rect 38476 13806 38528 13812
rect 38292 13320 38344 13326
rect 38292 13262 38344 13268
rect 37950 13084 38258 13093
rect 37950 13082 37956 13084
rect 38012 13082 38036 13084
rect 38092 13082 38116 13084
rect 38172 13082 38196 13084
rect 38252 13082 38258 13084
rect 38012 13030 38014 13082
rect 38194 13030 38196 13082
rect 37950 13028 37956 13030
rect 38012 13028 38036 13030
rect 38092 13028 38116 13030
rect 38172 13028 38196 13030
rect 38252 13028 38258 13030
rect 37950 13019 38258 13028
rect 37950 11996 38258 12005
rect 37950 11994 37956 11996
rect 38012 11994 38036 11996
rect 38092 11994 38116 11996
rect 38172 11994 38196 11996
rect 38252 11994 38258 11996
rect 38012 11942 38014 11994
rect 38194 11942 38196 11994
rect 37950 11940 37956 11942
rect 38012 11940 38036 11942
rect 38092 11940 38116 11942
rect 38172 11940 38196 11942
rect 38252 11940 38258 11942
rect 37950 11931 38258 11940
rect 37950 10908 38258 10917
rect 37950 10906 37956 10908
rect 38012 10906 38036 10908
rect 38092 10906 38116 10908
rect 38172 10906 38196 10908
rect 38252 10906 38258 10908
rect 38012 10854 38014 10906
rect 38194 10854 38196 10906
rect 37950 10852 37956 10854
rect 38012 10852 38036 10854
rect 38092 10852 38116 10854
rect 38172 10852 38196 10854
rect 38252 10852 38258 10854
rect 37950 10843 38258 10852
rect 37950 9820 38258 9829
rect 37950 9818 37956 9820
rect 38012 9818 38036 9820
rect 38092 9818 38116 9820
rect 38172 9818 38196 9820
rect 38252 9818 38258 9820
rect 38012 9766 38014 9818
rect 38194 9766 38196 9818
rect 37950 9764 37956 9766
rect 38012 9764 38036 9766
rect 38092 9764 38116 9766
rect 38172 9764 38196 9766
rect 38252 9764 38258 9766
rect 37950 9755 38258 9764
rect 37950 8732 38258 8741
rect 37950 8730 37956 8732
rect 38012 8730 38036 8732
rect 38092 8730 38116 8732
rect 38172 8730 38196 8732
rect 38252 8730 38258 8732
rect 38012 8678 38014 8730
rect 38194 8678 38196 8730
rect 37950 8676 37956 8678
rect 38012 8676 38036 8678
rect 38092 8676 38116 8678
rect 38172 8676 38196 8678
rect 38252 8676 38258 8678
rect 37950 8667 38258 8676
rect 37832 8560 37884 8566
rect 37832 8502 37884 8508
rect 37648 8356 37700 8362
rect 37648 8298 37700 8304
rect 37372 3120 37424 3126
rect 37372 3062 37424 3068
rect 37660 3058 37688 8298
rect 37950 7644 38258 7653
rect 37950 7642 37956 7644
rect 38012 7642 38036 7644
rect 38092 7642 38116 7644
rect 38172 7642 38196 7644
rect 38252 7642 38258 7644
rect 38012 7590 38014 7642
rect 38194 7590 38196 7642
rect 37950 7588 37956 7590
rect 38012 7588 38036 7590
rect 38092 7588 38116 7590
rect 38172 7588 38196 7590
rect 38252 7588 38258 7590
rect 37950 7579 38258 7588
rect 37950 6556 38258 6565
rect 37950 6554 37956 6556
rect 38012 6554 38036 6556
rect 38092 6554 38116 6556
rect 38172 6554 38196 6556
rect 38252 6554 38258 6556
rect 38012 6502 38014 6554
rect 38194 6502 38196 6554
rect 37950 6500 37956 6502
rect 38012 6500 38036 6502
rect 38092 6500 38116 6502
rect 38172 6500 38196 6502
rect 38252 6500 38258 6502
rect 37950 6491 38258 6500
rect 37950 5468 38258 5477
rect 37950 5466 37956 5468
rect 38012 5466 38036 5468
rect 38092 5466 38116 5468
rect 38172 5466 38196 5468
rect 38252 5466 38258 5468
rect 38012 5414 38014 5466
rect 38194 5414 38196 5466
rect 37950 5412 37956 5414
rect 38012 5412 38036 5414
rect 38092 5412 38116 5414
rect 38172 5412 38196 5414
rect 38252 5412 38258 5414
rect 37950 5403 38258 5412
rect 37950 4380 38258 4389
rect 37950 4378 37956 4380
rect 38012 4378 38036 4380
rect 38092 4378 38116 4380
rect 38172 4378 38196 4380
rect 38252 4378 38258 4380
rect 38012 4326 38014 4378
rect 38194 4326 38196 4378
rect 37950 4324 37956 4326
rect 38012 4324 38036 4326
rect 38092 4324 38116 4326
rect 38172 4324 38196 4326
rect 38252 4324 38258 4326
rect 37950 4315 38258 4324
rect 38488 4146 38516 13806
rect 38948 13802 38976 13942
rect 39132 13938 39160 15914
rect 40040 14408 40092 14414
rect 40040 14350 40092 14356
rect 39120 13932 39172 13938
rect 39120 13874 39172 13880
rect 38936 13796 38988 13802
rect 38936 13738 38988 13744
rect 39856 13184 39908 13190
rect 39856 13126 39908 13132
rect 38934 12336 38990 12345
rect 39868 12306 39896 13126
rect 39948 12640 40000 12646
rect 39948 12582 40000 12588
rect 38934 12271 38990 12280
rect 39856 12300 39908 12306
rect 38948 12238 38976 12271
rect 39856 12242 39908 12248
rect 38936 12232 38988 12238
rect 38936 12174 38988 12180
rect 39960 10674 39988 12582
rect 39948 10668 40000 10674
rect 39948 10610 40000 10616
rect 38476 4140 38528 4146
rect 38476 4082 38528 4088
rect 39028 4072 39080 4078
rect 39028 4014 39080 4020
rect 37950 3292 38258 3301
rect 37950 3290 37956 3292
rect 38012 3290 38036 3292
rect 38092 3290 38116 3292
rect 38172 3290 38196 3292
rect 38252 3290 38258 3292
rect 38012 3238 38014 3290
rect 38194 3238 38196 3290
rect 37950 3236 37956 3238
rect 38012 3236 38036 3238
rect 38092 3236 38116 3238
rect 38172 3236 38196 3238
rect 38252 3236 38258 3238
rect 37950 3227 38258 3236
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 36820 2984 36872 2990
rect 36820 2926 36872 2932
rect 36832 800 36860 2926
rect 37556 2916 37608 2922
rect 37556 2858 37608 2864
rect 37568 800 37596 2858
rect 38292 2508 38344 2514
rect 38292 2450 38344 2456
rect 37950 2204 38258 2213
rect 37950 2202 37956 2204
rect 38012 2202 38036 2204
rect 38092 2202 38116 2204
rect 38172 2202 38196 2204
rect 38252 2202 38258 2204
rect 38012 2150 38014 2202
rect 38194 2150 38196 2202
rect 37950 2148 37956 2150
rect 38012 2148 38036 2150
rect 38092 2148 38116 2150
rect 38172 2148 38196 2150
rect 38252 2148 38258 2150
rect 37950 2139 38258 2148
rect 38304 800 38332 2450
rect 39040 800 39068 4014
rect 39764 3596 39816 3602
rect 39764 3538 39816 3544
rect 39776 800 39804 3538
rect 40052 2446 40080 14350
rect 40144 13938 40172 16458
rect 40236 14414 40264 17002
rect 41800 15026 41828 18022
rect 42950 17980 43258 17989
rect 42950 17978 42956 17980
rect 43012 17978 43036 17980
rect 43092 17978 43116 17980
rect 43172 17978 43196 17980
rect 43252 17978 43258 17980
rect 43012 17926 43014 17978
rect 43194 17926 43196 17978
rect 42950 17924 42956 17926
rect 43012 17924 43036 17926
rect 43092 17924 43116 17926
rect 43172 17924 43196 17926
rect 43252 17924 43258 17926
rect 42950 17915 43258 17924
rect 43732 17270 43760 21014
rect 44468 18766 44496 25094
rect 45100 21412 45152 21418
rect 45100 21354 45152 21360
rect 44456 18760 44508 18766
rect 44456 18702 44508 18708
rect 44824 17808 44876 17814
rect 44824 17750 44876 17756
rect 43720 17264 43772 17270
rect 43720 17206 43772 17212
rect 42950 16892 43258 16901
rect 42950 16890 42956 16892
rect 43012 16890 43036 16892
rect 43092 16890 43116 16892
rect 43172 16890 43196 16892
rect 43252 16890 43258 16892
rect 43012 16838 43014 16890
rect 43194 16838 43196 16890
rect 42950 16836 42956 16838
rect 43012 16836 43036 16838
rect 43092 16836 43116 16838
rect 43172 16836 43196 16838
rect 43252 16836 43258 16838
rect 42950 16827 43258 16836
rect 42950 15804 43258 15813
rect 42950 15802 42956 15804
rect 43012 15802 43036 15804
rect 43092 15802 43116 15804
rect 43172 15802 43196 15804
rect 43252 15802 43258 15804
rect 43012 15750 43014 15802
rect 43194 15750 43196 15802
rect 42950 15748 42956 15750
rect 43012 15748 43036 15750
rect 43092 15748 43116 15750
rect 43172 15748 43196 15750
rect 43252 15748 43258 15750
rect 42950 15739 43258 15748
rect 41788 15020 41840 15026
rect 41788 14962 41840 14968
rect 41236 14816 41288 14822
rect 41236 14758 41288 14764
rect 44180 14816 44232 14822
rect 44180 14758 44232 14764
rect 40224 14408 40276 14414
rect 40224 14350 40276 14356
rect 40132 13932 40184 13938
rect 40132 13874 40184 13880
rect 40592 13864 40644 13870
rect 40592 13806 40644 13812
rect 40604 13326 40632 13806
rect 40592 13320 40644 13326
rect 40592 13262 40644 13268
rect 41248 12238 41276 14758
rect 42950 14716 43258 14725
rect 42950 14714 42956 14716
rect 43012 14714 43036 14716
rect 43092 14714 43116 14716
rect 43172 14714 43196 14716
rect 43252 14714 43258 14716
rect 43012 14662 43014 14714
rect 43194 14662 43196 14714
rect 42950 14660 42956 14662
rect 43012 14660 43036 14662
rect 43092 14660 43116 14662
rect 43172 14660 43196 14662
rect 43252 14660 43258 14662
rect 42950 14651 43258 14660
rect 41328 14544 41380 14550
rect 41328 14486 41380 14492
rect 41236 12232 41288 12238
rect 41236 12174 41288 12180
rect 41340 11762 41368 14486
rect 42800 14272 42852 14278
rect 42800 14214 42852 14220
rect 42708 14000 42760 14006
rect 42708 13942 42760 13948
rect 41880 12164 41932 12170
rect 41880 12106 41932 12112
rect 41328 11756 41380 11762
rect 41328 11698 41380 11704
rect 41420 7336 41472 7342
rect 41420 7278 41472 7284
rect 40132 6792 40184 6798
rect 40132 6734 40184 6740
rect 40144 4146 40172 6734
rect 40132 4140 40184 4146
rect 40132 4082 40184 4088
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 40592 2508 40644 2514
rect 40512 2468 40592 2496
rect 40040 2440 40092 2446
rect 40040 2382 40092 2388
rect 40512 800 40540 2468
rect 40592 2450 40644 2456
rect 41248 800 41276 3538
rect 41432 2446 41460 7278
rect 41892 3534 41920 12106
rect 42720 11762 42748 13942
rect 42708 11756 42760 11762
rect 42708 11698 42760 11704
rect 42812 11694 42840 14214
rect 43720 14068 43772 14074
rect 43720 14010 43772 14016
rect 42950 13628 43258 13637
rect 42950 13626 42956 13628
rect 43012 13626 43036 13628
rect 43092 13626 43116 13628
rect 43172 13626 43196 13628
rect 43252 13626 43258 13628
rect 43012 13574 43014 13626
rect 43194 13574 43196 13626
rect 42950 13572 42956 13574
rect 43012 13572 43036 13574
rect 43092 13572 43116 13574
rect 43172 13572 43196 13574
rect 43252 13572 43258 13574
rect 42950 13563 43258 13572
rect 43732 12918 43760 14010
rect 43720 12912 43772 12918
rect 43720 12854 43772 12860
rect 42950 12540 43258 12549
rect 42950 12538 42956 12540
rect 43012 12538 43036 12540
rect 43092 12538 43116 12540
rect 43172 12538 43196 12540
rect 43252 12538 43258 12540
rect 43012 12486 43014 12538
rect 43194 12486 43196 12538
rect 42950 12484 42956 12486
rect 43012 12484 43036 12486
rect 43092 12484 43116 12486
rect 43172 12484 43196 12486
rect 43252 12484 43258 12486
rect 42950 12475 43258 12484
rect 43352 12096 43404 12102
rect 43352 12038 43404 12044
rect 42800 11688 42852 11694
rect 42800 11630 42852 11636
rect 42950 11452 43258 11461
rect 42950 11450 42956 11452
rect 43012 11450 43036 11452
rect 43092 11450 43116 11452
rect 43172 11450 43196 11452
rect 43252 11450 43258 11452
rect 43012 11398 43014 11450
rect 43194 11398 43196 11450
rect 42950 11396 42956 11398
rect 43012 11396 43036 11398
rect 43092 11396 43116 11398
rect 43172 11396 43196 11398
rect 43252 11396 43258 11398
rect 42950 11387 43258 11396
rect 42708 10464 42760 10470
rect 42708 10406 42760 10412
rect 42720 8566 42748 10406
rect 42950 10364 43258 10373
rect 42950 10362 42956 10364
rect 43012 10362 43036 10364
rect 43092 10362 43116 10364
rect 43172 10362 43196 10364
rect 43252 10362 43258 10364
rect 43012 10310 43014 10362
rect 43194 10310 43196 10362
rect 42950 10308 42956 10310
rect 43012 10308 43036 10310
rect 43092 10308 43116 10310
rect 43172 10308 43196 10310
rect 43252 10308 43258 10310
rect 42950 10299 43258 10308
rect 42950 9276 43258 9285
rect 42950 9274 42956 9276
rect 43012 9274 43036 9276
rect 43092 9274 43116 9276
rect 43172 9274 43196 9276
rect 43252 9274 43258 9276
rect 43012 9222 43014 9274
rect 43194 9222 43196 9274
rect 42950 9220 42956 9222
rect 43012 9220 43036 9222
rect 43092 9220 43116 9222
rect 43172 9220 43196 9222
rect 43252 9220 43258 9222
rect 42950 9211 43258 9220
rect 43364 8974 43392 12038
rect 44192 11830 44220 14758
rect 44364 13864 44416 13870
rect 44364 13806 44416 13812
rect 44272 12096 44324 12102
rect 44272 12038 44324 12044
rect 44180 11824 44232 11830
rect 44180 11766 44232 11772
rect 44180 11552 44232 11558
rect 44180 11494 44232 11500
rect 44192 9586 44220 11494
rect 44284 11150 44312 12038
rect 44272 11144 44324 11150
rect 44272 11086 44324 11092
rect 44376 11082 44404 13806
rect 44836 13326 44864 17750
rect 45112 17678 45140 21354
rect 45480 19378 45508 25162
rect 46216 21554 46244 25706
rect 46860 23730 46888 26726
rect 47216 26240 47268 26246
rect 47216 26182 47268 26188
rect 46940 25764 46992 25770
rect 46940 25706 46992 25712
rect 46848 23724 46900 23730
rect 46848 23666 46900 23672
rect 46664 23044 46716 23050
rect 46664 22986 46716 22992
rect 46204 21548 46256 21554
rect 46204 21490 46256 21496
rect 46204 19780 46256 19786
rect 46204 19722 46256 19728
rect 45468 19372 45520 19378
rect 45468 19314 45520 19320
rect 45100 17672 45152 17678
rect 45100 17614 45152 17620
rect 46216 16590 46244 19722
rect 46676 18290 46704 22986
rect 46952 20942 46980 25706
rect 47228 24818 47256 26182
rect 47492 25220 47544 25226
rect 47492 25162 47544 25168
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 47504 23662 47532 25162
rect 47492 23656 47544 23662
rect 47492 23598 47544 23604
rect 47596 22030 47624 27338
rect 47676 26784 47728 26790
rect 47676 26726 47728 26732
rect 47688 23118 47716 26726
rect 47676 23112 47728 23118
rect 47676 23054 47728 23060
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 46940 20936 46992 20942
rect 46940 20878 46992 20884
rect 46664 18284 46716 18290
rect 46664 18226 46716 18232
rect 46848 17604 46900 17610
rect 46848 17546 46900 17552
rect 46664 17536 46716 17542
rect 46664 17478 46716 17484
rect 46204 16584 46256 16590
rect 46204 16526 46256 16532
rect 46676 13938 46704 17478
rect 46756 17060 46808 17066
rect 46756 17002 46808 17008
rect 46768 15026 46796 17002
rect 46860 15502 46888 17546
rect 46848 15496 46900 15502
rect 46848 15438 46900 15444
rect 46756 15020 46808 15026
rect 46756 14962 46808 14968
rect 46664 13932 46716 13938
rect 46664 13874 46716 13880
rect 44824 13320 44876 13326
rect 44824 13262 44876 13268
rect 46756 13184 46808 13190
rect 46756 13126 46808 13132
rect 46768 12850 46796 13126
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 44732 12708 44784 12714
rect 44732 12650 44784 12656
rect 44744 12238 44772 12650
rect 44732 12232 44784 12238
rect 44732 12174 44784 12180
rect 45652 11620 45704 11626
rect 45652 11562 45704 11568
rect 46848 11620 46900 11626
rect 46848 11562 46900 11568
rect 44364 11076 44416 11082
rect 44364 11018 44416 11024
rect 45664 10062 45692 11562
rect 46388 11552 46440 11558
rect 46388 11494 46440 11500
rect 45652 10056 45704 10062
rect 45652 9998 45704 10004
rect 44180 9580 44232 9586
rect 44180 9522 44232 9528
rect 43352 8968 43404 8974
rect 43352 8910 43404 8916
rect 46204 8900 46256 8906
rect 46204 8842 46256 8848
rect 42708 8560 42760 8566
rect 42708 8502 42760 8508
rect 42616 8424 42668 8430
rect 42616 8366 42668 8372
rect 41880 3528 41932 3534
rect 41880 3470 41932 3476
rect 42628 3058 42656 8366
rect 45928 8356 45980 8362
rect 45928 8298 45980 8304
rect 42950 8188 43258 8197
rect 42950 8186 42956 8188
rect 43012 8186 43036 8188
rect 43092 8186 43116 8188
rect 43172 8186 43196 8188
rect 43252 8186 43258 8188
rect 43012 8134 43014 8186
rect 43194 8134 43196 8186
rect 42950 8132 42956 8134
rect 43012 8132 43036 8134
rect 43092 8132 43116 8134
rect 43172 8132 43196 8134
rect 43252 8132 43258 8134
rect 42950 8123 43258 8132
rect 45192 7268 45244 7274
rect 45192 7210 45244 7216
rect 42950 7100 43258 7109
rect 42950 7098 42956 7100
rect 43012 7098 43036 7100
rect 43092 7098 43116 7100
rect 43172 7098 43196 7100
rect 43252 7098 43258 7100
rect 43012 7046 43014 7098
rect 43194 7046 43196 7098
rect 42950 7044 42956 7046
rect 43012 7044 43036 7046
rect 43092 7044 43116 7046
rect 43172 7044 43196 7046
rect 43252 7044 43258 7046
rect 42950 7035 43258 7044
rect 44456 6724 44508 6730
rect 44456 6666 44508 6672
rect 42950 6012 43258 6021
rect 42950 6010 42956 6012
rect 43012 6010 43036 6012
rect 43092 6010 43116 6012
rect 43172 6010 43196 6012
rect 43252 6010 43258 6012
rect 43012 5958 43014 6010
rect 43194 5958 43196 6010
rect 42950 5956 42956 5958
rect 43012 5956 43036 5958
rect 43092 5956 43116 5958
rect 43172 5956 43196 5958
rect 43252 5956 43258 5958
rect 42950 5947 43258 5956
rect 42950 4924 43258 4933
rect 42950 4922 42956 4924
rect 43012 4922 43036 4924
rect 43092 4922 43116 4924
rect 43172 4922 43196 4924
rect 43252 4922 43258 4924
rect 43012 4870 43014 4922
rect 43194 4870 43196 4922
rect 42950 4868 42956 4870
rect 43012 4868 43036 4870
rect 43092 4868 43116 4870
rect 43172 4868 43196 4870
rect 43252 4868 43258 4870
rect 42950 4859 43258 4868
rect 43444 4072 43496 4078
rect 43444 4014 43496 4020
rect 42950 3836 43258 3845
rect 42950 3834 42956 3836
rect 43012 3834 43036 3836
rect 43092 3834 43116 3836
rect 43172 3834 43196 3836
rect 43252 3834 43258 3836
rect 43012 3782 43014 3834
rect 43194 3782 43196 3834
rect 42950 3780 42956 3782
rect 43012 3780 43036 3782
rect 43092 3780 43116 3782
rect 43172 3780 43196 3782
rect 43252 3780 43258 3782
rect 42950 3771 43258 3780
rect 42616 3052 42668 3058
rect 42616 2994 42668 3000
rect 41972 2984 42024 2990
rect 41972 2926 42024 2932
rect 41420 2440 41472 2446
rect 41420 2382 41472 2388
rect 41984 800 42012 2926
rect 42708 2916 42760 2922
rect 42708 2858 42760 2864
rect 42720 800 42748 2858
rect 42950 2748 43258 2757
rect 42950 2746 42956 2748
rect 43012 2746 43036 2748
rect 43092 2746 43116 2748
rect 43172 2746 43196 2748
rect 43252 2746 43258 2748
rect 43012 2694 43014 2746
rect 43194 2694 43196 2746
rect 42950 2692 42956 2694
rect 43012 2692 43036 2694
rect 43092 2692 43116 2694
rect 43172 2692 43196 2694
rect 43252 2692 43258 2694
rect 42950 2683 43258 2692
rect 43456 800 43484 4014
rect 44180 3596 44232 3602
rect 44180 3538 44232 3544
rect 44192 800 44220 3538
rect 44468 3058 44496 6666
rect 45204 3534 45232 7210
rect 45940 6798 45968 8298
rect 45928 6792 45980 6798
rect 45928 6734 45980 6740
rect 46216 5710 46244 8842
rect 46400 7886 46428 11494
rect 46480 11076 46532 11082
rect 46480 11018 46532 11024
rect 46492 8498 46520 11018
rect 46860 9586 46888 11562
rect 47584 10668 47636 10674
rect 47584 10610 47636 10616
rect 46848 9580 46900 9586
rect 46848 9522 46900 9528
rect 47124 8900 47176 8906
rect 47124 8842 47176 8848
rect 46480 8492 46532 8498
rect 46480 8434 46532 8440
rect 46388 7880 46440 7886
rect 46388 7822 46440 7828
rect 46204 5704 46256 5710
rect 46204 5646 46256 5652
rect 46020 4140 46072 4146
rect 46020 4082 46072 4088
rect 46032 4010 46060 4082
rect 46020 4004 46072 4010
rect 46020 3946 46072 3952
rect 45192 3528 45244 3534
rect 44914 3496 44970 3505
rect 45192 3470 45244 3476
rect 44914 3431 44970 3440
rect 44456 3052 44508 3058
rect 44456 2994 44508 3000
rect 44928 800 44956 3431
rect 46032 2650 46060 3946
rect 47136 3194 47164 8842
rect 47596 7274 47624 10610
rect 47780 9518 47808 31726
rect 47950 31580 48258 31589
rect 47950 31578 47956 31580
rect 48012 31578 48036 31580
rect 48092 31578 48116 31580
rect 48172 31578 48196 31580
rect 48252 31578 48258 31580
rect 48012 31526 48014 31578
rect 48194 31526 48196 31578
rect 47950 31524 47956 31526
rect 48012 31524 48036 31526
rect 48092 31524 48116 31526
rect 48172 31524 48196 31526
rect 48252 31524 48258 31526
rect 47950 31515 48258 31524
rect 48332 31346 48360 33866
rect 48320 31340 48372 31346
rect 48320 31282 48372 31288
rect 47860 31136 47912 31142
rect 47860 31078 47912 31084
rect 47872 28082 47900 31078
rect 47950 30492 48258 30501
rect 47950 30490 47956 30492
rect 48012 30490 48036 30492
rect 48092 30490 48116 30492
rect 48172 30490 48196 30492
rect 48252 30490 48258 30492
rect 48012 30438 48014 30490
rect 48194 30438 48196 30490
rect 47950 30436 47956 30438
rect 48012 30436 48036 30438
rect 48092 30436 48116 30438
rect 48172 30436 48196 30438
rect 48252 30436 48258 30438
rect 47950 30427 48258 30436
rect 47950 29404 48258 29413
rect 47950 29402 47956 29404
rect 48012 29402 48036 29404
rect 48092 29402 48116 29404
rect 48172 29402 48196 29404
rect 48252 29402 48258 29404
rect 48012 29350 48014 29402
rect 48194 29350 48196 29402
rect 47950 29348 47956 29350
rect 48012 29348 48036 29350
rect 48092 29348 48116 29350
rect 48172 29348 48196 29350
rect 48252 29348 48258 29350
rect 47950 29339 48258 29348
rect 47950 28316 48258 28325
rect 47950 28314 47956 28316
rect 48012 28314 48036 28316
rect 48092 28314 48116 28316
rect 48172 28314 48196 28316
rect 48252 28314 48258 28316
rect 48012 28262 48014 28314
rect 48194 28262 48196 28314
rect 47950 28260 47956 28262
rect 48012 28260 48036 28262
rect 48092 28260 48116 28262
rect 48172 28260 48196 28262
rect 48252 28260 48258 28262
rect 47950 28251 48258 28260
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 47860 27872 47912 27878
rect 47860 27814 47912 27820
rect 47872 24206 47900 27814
rect 47950 27228 48258 27237
rect 47950 27226 47956 27228
rect 48012 27226 48036 27228
rect 48092 27226 48116 27228
rect 48172 27226 48196 27228
rect 48252 27226 48258 27228
rect 48012 27174 48014 27226
rect 48194 27174 48196 27226
rect 47950 27172 47956 27174
rect 48012 27172 48036 27174
rect 48092 27172 48116 27174
rect 48172 27172 48196 27174
rect 48252 27172 48258 27174
rect 47950 27163 48258 27172
rect 47950 26140 48258 26149
rect 47950 26138 47956 26140
rect 48012 26138 48036 26140
rect 48092 26138 48116 26140
rect 48172 26138 48196 26140
rect 48252 26138 48258 26140
rect 48012 26086 48014 26138
rect 48194 26086 48196 26138
rect 47950 26084 47956 26086
rect 48012 26084 48036 26086
rect 48092 26084 48116 26086
rect 48172 26084 48196 26086
rect 48252 26084 48258 26086
rect 47950 26075 48258 26084
rect 47950 25052 48258 25061
rect 47950 25050 47956 25052
rect 48012 25050 48036 25052
rect 48092 25050 48116 25052
rect 48172 25050 48196 25052
rect 48252 25050 48258 25052
rect 48012 24998 48014 25050
rect 48194 24998 48196 25050
rect 47950 24996 47956 24998
rect 48012 24996 48036 24998
rect 48092 24996 48116 24998
rect 48172 24996 48196 24998
rect 48252 24996 48258 24998
rect 47950 24987 48258 24996
rect 47860 24200 47912 24206
rect 47860 24142 47912 24148
rect 47950 23964 48258 23973
rect 47950 23962 47956 23964
rect 48012 23962 48036 23964
rect 48092 23962 48116 23964
rect 48172 23962 48196 23964
rect 48252 23962 48258 23964
rect 48012 23910 48014 23962
rect 48194 23910 48196 23962
rect 47950 23908 47956 23910
rect 48012 23908 48036 23910
rect 48092 23908 48116 23910
rect 48172 23908 48196 23910
rect 48252 23908 48258 23910
rect 47950 23899 48258 23908
rect 47860 23656 47912 23662
rect 47860 23598 47912 23604
rect 47872 20466 47900 23598
rect 47950 22876 48258 22885
rect 47950 22874 47956 22876
rect 48012 22874 48036 22876
rect 48092 22874 48116 22876
rect 48172 22874 48196 22876
rect 48252 22874 48258 22876
rect 48012 22822 48014 22874
rect 48194 22822 48196 22874
rect 47950 22820 47956 22822
rect 48012 22820 48036 22822
rect 48092 22820 48116 22822
rect 48172 22820 48196 22822
rect 48252 22820 48258 22822
rect 47950 22811 48258 22820
rect 47950 21788 48258 21797
rect 47950 21786 47956 21788
rect 48012 21786 48036 21788
rect 48092 21786 48116 21788
rect 48172 21786 48196 21788
rect 48252 21786 48258 21788
rect 48012 21734 48014 21786
rect 48194 21734 48196 21786
rect 47950 21732 47956 21734
rect 48012 21732 48036 21734
rect 48092 21732 48116 21734
rect 48172 21732 48196 21734
rect 48252 21732 48258 21734
rect 47950 21723 48258 21732
rect 47950 20700 48258 20709
rect 47950 20698 47956 20700
rect 48012 20698 48036 20700
rect 48092 20698 48116 20700
rect 48172 20698 48196 20700
rect 48252 20698 48258 20700
rect 48012 20646 48014 20698
rect 48194 20646 48196 20698
rect 47950 20644 47956 20646
rect 48012 20644 48036 20646
rect 48092 20644 48116 20646
rect 48172 20644 48196 20646
rect 48252 20644 48258 20646
rect 47950 20635 48258 20644
rect 47860 20460 47912 20466
rect 47860 20402 47912 20408
rect 47950 19612 48258 19621
rect 47950 19610 47956 19612
rect 48012 19610 48036 19612
rect 48092 19610 48116 19612
rect 48172 19610 48196 19612
rect 48252 19610 48258 19612
rect 48012 19558 48014 19610
rect 48194 19558 48196 19610
rect 47950 19556 47956 19558
rect 48012 19556 48036 19558
rect 48092 19556 48116 19558
rect 48172 19556 48196 19558
rect 48252 19556 48258 19558
rect 47950 19547 48258 19556
rect 47860 18692 47912 18698
rect 47860 18634 47912 18640
rect 47872 16114 47900 18634
rect 47950 18524 48258 18533
rect 47950 18522 47956 18524
rect 48012 18522 48036 18524
rect 48092 18522 48116 18524
rect 48172 18522 48196 18524
rect 48252 18522 48258 18524
rect 48012 18470 48014 18522
rect 48194 18470 48196 18522
rect 47950 18468 47956 18470
rect 48012 18468 48036 18470
rect 48092 18468 48116 18470
rect 48172 18468 48196 18470
rect 48252 18468 48258 18470
rect 47950 18459 48258 18468
rect 47950 17436 48258 17445
rect 47950 17434 47956 17436
rect 48012 17434 48036 17436
rect 48092 17434 48116 17436
rect 48172 17434 48196 17436
rect 48252 17434 48258 17436
rect 48012 17382 48014 17434
rect 48194 17382 48196 17434
rect 47950 17380 47956 17382
rect 48012 17380 48036 17382
rect 48092 17380 48116 17382
rect 48172 17380 48196 17382
rect 48252 17380 48258 17382
rect 47950 17371 48258 17380
rect 47950 16348 48258 16357
rect 47950 16346 47956 16348
rect 48012 16346 48036 16348
rect 48092 16346 48116 16348
rect 48172 16346 48196 16348
rect 48252 16346 48258 16348
rect 48012 16294 48014 16346
rect 48194 16294 48196 16346
rect 47950 16292 47956 16294
rect 48012 16292 48036 16294
rect 48092 16292 48116 16294
rect 48172 16292 48196 16294
rect 48252 16292 48258 16294
rect 47950 16283 48258 16292
rect 47860 16108 47912 16114
rect 47860 16050 47912 16056
rect 47950 15260 48258 15269
rect 47950 15258 47956 15260
rect 48012 15258 48036 15260
rect 48092 15258 48116 15260
rect 48172 15258 48196 15260
rect 48252 15258 48258 15260
rect 48012 15206 48014 15258
rect 48194 15206 48196 15258
rect 47950 15204 47956 15206
rect 48012 15204 48036 15206
rect 48092 15204 48116 15206
rect 48172 15204 48196 15206
rect 48252 15204 48258 15206
rect 47950 15195 48258 15204
rect 47950 14172 48258 14181
rect 47950 14170 47956 14172
rect 48012 14170 48036 14172
rect 48092 14170 48116 14172
rect 48172 14170 48196 14172
rect 48252 14170 48258 14172
rect 48012 14118 48014 14170
rect 48194 14118 48196 14170
rect 47950 14116 47956 14118
rect 48012 14116 48036 14118
rect 48092 14116 48116 14118
rect 48172 14116 48196 14118
rect 48252 14116 48258 14118
rect 47950 14107 48258 14116
rect 47950 13084 48258 13093
rect 47950 13082 47956 13084
rect 48012 13082 48036 13084
rect 48092 13082 48116 13084
rect 48172 13082 48196 13084
rect 48252 13082 48258 13084
rect 48012 13030 48014 13082
rect 48194 13030 48196 13082
rect 47950 13028 47956 13030
rect 48012 13028 48036 13030
rect 48092 13028 48116 13030
rect 48172 13028 48196 13030
rect 48252 13028 48258 13030
rect 47950 13019 48258 13028
rect 47950 11996 48258 12005
rect 47950 11994 47956 11996
rect 48012 11994 48036 11996
rect 48092 11994 48116 11996
rect 48172 11994 48196 11996
rect 48252 11994 48258 11996
rect 48012 11942 48014 11994
rect 48194 11942 48196 11994
rect 47950 11940 47956 11942
rect 48012 11940 48036 11942
rect 48092 11940 48116 11942
rect 48172 11940 48196 11942
rect 48252 11940 48258 11942
rect 47950 11931 48258 11940
rect 47950 10908 48258 10917
rect 47950 10906 47956 10908
rect 48012 10906 48036 10908
rect 48092 10906 48116 10908
rect 48172 10906 48196 10908
rect 48252 10906 48258 10908
rect 48012 10854 48014 10906
rect 48194 10854 48196 10906
rect 47950 10852 47956 10854
rect 48012 10852 48036 10854
rect 48092 10852 48116 10854
rect 48172 10852 48196 10854
rect 48252 10852 48258 10854
rect 47950 10843 48258 10852
rect 47950 9820 48258 9829
rect 47950 9818 47956 9820
rect 48012 9818 48036 9820
rect 48092 9818 48116 9820
rect 48172 9818 48196 9820
rect 48252 9818 48258 9820
rect 48012 9766 48014 9818
rect 48194 9766 48196 9818
rect 47950 9764 47956 9766
rect 48012 9764 48036 9766
rect 48092 9764 48116 9766
rect 48172 9764 48196 9766
rect 48252 9764 48258 9766
rect 47950 9755 48258 9764
rect 47768 9512 47820 9518
rect 47768 9454 47820 9460
rect 47768 9376 47820 9382
rect 47768 9318 47820 9324
rect 47676 8968 47728 8974
rect 47676 8910 47728 8916
rect 47584 7268 47636 7274
rect 47584 7210 47636 7216
rect 47688 3534 47716 8910
rect 47780 7410 47808 9318
rect 48424 8906 48452 41550
rect 48504 41064 48556 41070
rect 48502 41032 48504 41041
rect 48556 41032 48558 41041
rect 48502 40967 48558 40976
rect 48778 40624 48834 40633
rect 48778 40559 48780 40568
rect 48832 40559 48834 40568
rect 48780 40530 48832 40536
rect 48504 40520 48556 40526
rect 48504 40462 48556 40468
rect 48516 40361 48544 40462
rect 48502 40352 48558 40361
rect 48502 40287 48558 40296
rect 48504 39976 48556 39982
rect 48504 39918 48556 39924
rect 48596 39976 48648 39982
rect 48596 39918 48648 39924
rect 48516 39681 48544 39918
rect 48502 39672 48558 39681
rect 48502 39607 48558 39616
rect 48504 39432 48556 39438
rect 48504 39374 48556 39380
rect 48516 39001 48544 39374
rect 48502 38992 48558 39001
rect 48502 38927 48558 38936
rect 48608 38010 48636 39918
rect 48976 39574 49004 45526
rect 49068 45354 49096 46974
rect 49148 45892 49200 45898
rect 49148 45834 49200 45840
rect 49160 45801 49188 45834
rect 49146 45792 49202 45801
rect 49146 45727 49202 45736
rect 49056 45348 49108 45354
rect 49056 45290 49108 45296
rect 48964 39568 49016 39574
rect 48778 39536 48834 39545
rect 48964 39510 49016 39516
rect 48778 39471 48780 39480
rect 48832 39471 48834 39480
rect 48780 39442 48832 39448
rect 49148 38208 49200 38214
rect 49148 38150 49200 38156
rect 48596 38004 48648 38010
rect 48596 37946 48648 37952
rect 49160 37466 49188 38150
rect 49148 37460 49200 37466
rect 49148 37402 49200 37408
rect 48504 37324 48556 37330
rect 48504 37266 48556 37272
rect 48516 36961 48544 37266
rect 48780 37256 48832 37262
rect 48780 37198 48832 37204
rect 48502 36952 48558 36961
rect 48502 36887 48558 36896
rect 48792 36854 48820 37198
rect 48780 36848 48832 36854
rect 48780 36790 48832 36796
rect 49148 36576 49200 36582
rect 49148 36518 49200 36524
rect 49160 36310 49188 36518
rect 49148 36304 49200 36310
rect 49148 36246 49200 36252
rect 49056 35828 49108 35834
rect 49056 35770 49108 35776
rect 49068 34542 49096 35770
rect 49148 34944 49200 34950
rect 49148 34886 49200 34892
rect 49160 34678 49188 34886
rect 49148 34672 49200 34678
rect 49148 34614 49200 34620
rect 49056 34536 49108 34542
rect 49056 34478 49108 34484
rect 49252 33969 49280 48334
rect 49332 46572 49384 46578
rect 49332 46514 49384 46520
rect 49344 46481 49372 46514
rect 49330 46472 49386 46481
rect 49330 46407 49386 46416
rect 49330 45112 49386 45121
rect 49330 45047 49386 45056
rect 49344 44402 49372 45047
rect 49332 44396 49384 44402
rect 49332 44338 49384 44344
rect 49332 38344 49384 38350
rect 49330 38312 49332 38321
rect 49384 38312 49386 38321
rect 49330 38247 49386 38256
rect 49332 37868 49384 37874
rect 49332 37810 49384 37816
rect 49344 37641 49372 37810
rect 49330 37632 49386 37641
rect 49330 37567 49386 37576
rect 49332 36780 49384 36786
rect 49332 36722 49384 36728
rect 49344 36281 49372 36722
rect 49330 36272 49386 36281
rect 49330 36207 49386 36216
rect 49332 35692 49384 35698
rect 49332 35634 49384 35640
rect 49344 35601 49372 35634
rect 49330 35592 49386 35601
rect 49330 35527 49386 35536
rect 49332 35080 49384 35086
rect 49332 35022 49384 35028
rect 49344 34921 49372 35022
rect 49330 34912 49386 34921
rect 49330 34847 49386 34856
rect 49332 34604 49384 34610
rect 49332 34546 49384 34552
rect 49344 34241 49372 34546
rect 49330 34232 49386 34241
rect 49330 34167 49386 34176
rect 49332 33992 49384 33998
rect 49238 33960 49294 33969
rect 49332 33934 49384 33940
rect 49238 33895 49294 33904
rect 48596 33856 48648 33862
rect 48596 33798 48648 33804
rect 48504 32360 48556 32366
rect 48504 32302 48556 32308
rect 48516 32201 48544 32302
rect 48502 32192 48558 32201
rect 48502 32127 48558 32136
rect 48504 31816 48556 31822
rect 48504 31758 48556 31764
rect 48516 31521 48544 31758
rect 48502 31512 48558 31521
rect 48502 31447 48558 31456
rect 48504 31272 48556 31278
rect 48504 31214 48556 31220
rect 48516 30841 48544 31214
rect 48502 30832 48558 30841
rect 48608 30802 48636 33798
rect 49344 33561 49372 33934
rect 49330 33552 49386 33561
rect 49330 33487 49386 33496
rect 48780 33108 48832 33114
rect 48780 33050 48832 33056
rect 48792 32434 48820 33050
rect 49332 32904 49384 32910
rect 49330 32872 49332 32881
rect 49384 32872 49386 32881
rect 49330 32807 49386 32816
rect 49148 32768 49200 32774
rect 49148 32710 49200 32716
rect 48780 32428 48832 32434
rect 48780 32370 48832 32376
rect 49160 32298 49188 32710
rect 49148 32292 49200 32298
rect 49148 32234 49200 32240
rect 48502 30767 48558 30776
rect 48596 30796 48648 30802
rect 48596 30738 48648 30744
rect 49332 30252 49384 30258
rect 49332 30194 49384 30200
rect 49344 30161 49372 30194
rect 49330 30152 49386 30161
rect 49330 30087 49386 30096
rect 48504 29640 48556 29646
rect 48504 29582 48556 29588
rect 48516 29481 48544 29582
rect 48502 29472 48558 29481
rect 48502 29407 48558 29416
rect 49332 29164 49384 29170
rect 49332 29106 49384 29112
rect 49344 28801 49372 29106
rect 49330 28792 49386 28801
rect 49330 28727 49386 28736
rect 49332 28552 49384 28558
rect 49332 28494 49384 28500
rect 49148 28416 49200 28422
rect 49148 28358 49200 28364
rect 49160 28150 49188 28358
rect 49148 28144 49200 28150
rect 49344 28121 49372 28494
rect 49148 28086 49200 28092
rect 49330 28112 49386 28121
rect 49330 28047 49386 28056
rect 48504 27464 48556 27470
rect 48502 27432 48504 27441
rect 48596 27464 48648 27470
rect 48556 27432 48558 27441
rect 48596 27406 48648 27412
rect 48502 27367 48558 27376
rect 48504 26920 48556 26926
rect 48504 26862 48556 26868
rect 48516 26761 48544 26862
rect 48502 26752 48558 26761
rect 48502 26687 48558 26696
rect 48608 26518 48636 27406
rect 48780 26920 48832 26926
rect 48780 26862 48832 26868
rect 48792 26586 48820 26862
rect 48780 26580 48832 26586
rect 48780 26522 48832 26528
rect 48596 26512 48648 26518
rect 48596 26454 48648 26460
rect 48504 26376 48556 26382
rect 48504 26318 48556 26324
rect 48516 26081 48544 26318
rect 48502 26072 48558 26081
rect 48502 26007 48558 26016
rect 49332 25900 49384 25906
rect 49332 25842 49384 25848
rect 49148 25696 49200 25702
rect 49148 25638 49200 25644
rect 49160 25430 49188 25638
rect 49148 25424 49200 25430
rect 49344 25401 49372 25842
rect 49148 25366 49200 25372
rect 49330 25392 49386 25401
rect 49330 25327 49386 25336
rect 49148 24744 49200 24750
rect 49146 24712 49148 24721
rect 49200 24712 49202 24721
rect 49146 24647 49202 24656
rect 49148 24132 49200 24138
rect 49148 24074 49200 24080
rect 49160 24041 49188 24074
rect 49146 24032 49202 24041
rect 49146 23967 49202 23976
rect 49148 23656 49200 23662
rect 49148 23598 49200 23604
rect 49160 23361 49188 23598
rect 49146 23352 49202 23361
rect 49146 23287 49202 23296
rect 49148 23044 49200 23050
rect 49148 22986 49200 22992
rect 49160 22681 49188 22986
rect 49146 22672 49202 22681
rect 49146 22607 49202 22616
rect 49148 22024 49200 22030
rect 49146 21992 49148 22001
rect 49200 21992 49202 22001
rect 49146 21927 49202 21936
rect 49148 21480 49200 21486
rect 49148 21422 49200 21428
rect 49160 21321 49188 21422
rect 49146 21312 49202 21321
rect 49146 21247 49202 21256
rect 49148 20868 49200 20874
rect 49148 20810 49200 20816
rect 49160 20641 49188 20810
rect 49146 20632 49202 20641
rect 49146 20567 49202 20576
rect 49148 20392 49200 20398
rect 49148 20334 49200 20340
rect 49160 19961 49188 20334
rect 49146 19952 49202 19961
rect 49146 19887 49202 19896
rect 49148 19372 49200 19378
rect 49148 19314 49200 19320
rect 49160 19281 49188 19314
rect 49146 19272 49202 19281
rect 49146 19207 49202 19216
rect 49148 18692 49200 18698
rect 49148 18634 49200 18640
rect 49160 18601 49188 18634
rect 49146 18592 49202 18601
rect 49146 18527 49202 18536
rect 49148 18216 49200 18222
rect 49148 18158 49200 18164
rect 49160 17921 49188 18158
rect 49146 17912 49202 17921
rect 49146 17847 49202 17856
rect 49148 17604 49200 17610
rect 49148 17546 49200 17552
rect 49160 17241 49188 17546
rect 49146 17232 49202 17241
rect 49146 17167 49202 17176
rect 49146 16552 49202 16561
rect 49146 16487 49148 16496
rect 49200 16487 49202 16496
rect 49148 16458 49200 16464
rect 49148 16040 49200 16046
rect 49148 15982 49200 15988
rect 49160 15881 49188 15982
rect 49146 15872 49202 15881
rect 49146 15807 49202 15816
rect 49148 15428 49200 15434
rect 49148 15370 49200 15376
rect 49160 15201 49188 15370
rect 49146 15192 49202 15201
rect 49146 15127 49202 15136
rect 49148 14952 49200 14958
rect 49148 14894 49200 14900
rect 49160 14521 49188 14894
rect 49146 14512 49202 14521
rect 49146 14447 49202 14456
rect 49148 13864 49200 13870
rect 49146 13832 49148 13841
rect 49200 13832 49202 13841
rect 49146 13767 49202 13776
rect 49148 13252 49200 13258
rect 49148 13194 49200 13200
rect 49160 13161 49188 13194
rect 49146 13152 49202 13161
rect 49146 13087 49202 13096
rect 49148 12776 49200 12782
rect 49148 12718 49200 12724
rect 49160 12481 49188 12718
rect 49146 12472 49202 12481
rect 49146 12407 49202 12416
rect 49148 12164 49200 12170
rect 49148 12106 49200 12112
rect 49160 11801 49188 12106
rect 49146 11792 49202 11801
rect 49146 11727 49202 11736
rect 49148 11144 49200 11150
rect 49146 11112 49148 11121
rect 49200 11112 49202 11121
rect 49146 11047 49202 11056
rect 49148 10600 49200 10606
rect 49148 10542 49200 10548
rect 49160 10441 49188 10542
rect 49146 10432 49202 10441
rect 49146 10367 49202 10376
rect 49148 9988 49200 9994
rect 49148 9930 49200 9936
rect 49160 9761 49188 9930
rect 49146 9752 49202 9761
rect 49146 9687 49202 9696
rect 48688 9512 48740 9518
rect 48688 9454 48740 9460
rect 49148 9512 49200 9518
rect 49148 9454 49200 9460
rect 48700 8906 48728 9454
rect 49160 9081 49188 9454
rect 49146 9072 49202 9081
rect 49146 9007 49202 9016
rect 48412 8900 48464 8906
rect 48412 8842 48464 8848
rect 48688 8900 48740 8906
rect 48688 8842 48740 8848
rect 47860 8832 47912 8838
rect 47860 8774 47912 8780
rect 47768 7404 47820 7410
rect 47768 7346 47820 7352
rect 47768 7268 47820 7274
rect 47768 7210 47820 7216
rect 47780 5030 47808 7210
rect 47768 5024 47820 5030
rect 47768 4966 47820 4972
rect 47768 3936 47820 3942
rect 47768 3878 47820 3884
rect 47676 3528 47728 3534
rect 47676 3470 47728 3476
rect 47124 3188 47176 3194
rect 47124 3130 47176 3136
rect 47124 3052 47176 3058
rect 47124 2994 47176 3000
rect 46388 2848 46440 2854
rect 46388 2790 46440 2796
rect 46020 2644 46072 2650
rect 46020 2586 46072 2592
rect 45652 2372 45704 2378
rect 45652 2314 45704 2320
rect 45664 800 45692 2314
rect 46400 800 46428 2790
rect 47136 800 47164 2994
rect 47780 2446 47808 3878
rect 47872 3126 47900 8774
rect 47950 8732 48258 8741
rect 47950 8730 47956 8732
rect 48012 8730 48036 8732
rect 48092 8730 48116 8732
rect 48172 8730 48196 8732
rect 48252 8730 48258 8732
rect 48012 8678 48014 8730
rect 48194 8678 48196 8730
rect 47950 8676 47956 8678
rect 48012 8676 48036 8678
rect 48092 8676 48116 8678
rect 48172 8676 48196 8678
rect 48252 8676 48258 8678
rect 47950 8667 48258 8676
rect 47950 7644 48258 7653
rect 47950 7642 47956 7644
rect 48012 7642 48036 7644
rect 48092 7642 48116 7644
rect 48172 7642 48196 7644
rect 48252 7642 48258 7644
rect 48012 7590 48014 7642
rect 48194 7590 48196 7642
rect 47950 7588 47956 7590
rect 48012 7588 48036 7590
rect 48092 7588 48116 7590
rect 48172 7588 48196 7590
rect 48252 7588 48258 7590
rect 47950 7579 48258 7588
rect 48700 6914 48728 8842
rect 49148 8424 49200 8430
rect 49146 8392 49148 8401
rect 49200 8392 49202 8401
rect 49146 8327 49202 8336
rect 49148 7812 49200 7818
rect 49148 7754 49200 7760
rect 49160 7721 49188 7754
rect 49146 7712 49202 7721
rect 49146 7647 49202 7656
rect 49148 7336 49200 7342
rect 49148 7278 49200 7284
rect 49160 7041 49188 7278
rect 49146 7032 49202 7041
rect 49146 6967 49202 6976
rect 48700 6886 48912 6914
rect 47950 6556 48258 6565
rect 47950 6554 47956 6556
rect 48012 6554 48036 6556
rect 48092 6554 48116 6556
rect 48172 6554 48196 6556
rect 48252 6554 48258 6556
rect 48012 6502 48014 6554
rect 48194 6502 48196 6554
rect 47950 6500 47956 6502
rect 48012 6500 48036 6502
rect 48092 6500 48116 6502
rect 48172 6500 48196 6502
rect 48252 6500 48258 6502
rect 47950 6491 48258 6500
rect 47950 5468 48258 5477
rect 47950 5466 47956 5468
rect 48012 5466 48036 5468
rect 48092 5466 48116 5468
rect 48172 5466 48196 5468
rect 48252 5466 48258 5468
rect 48012 5414 48014 5466
rect 48194 5414 48196 5466
rect 47950 5412 47956 5414
rect 48012 5412 48036 5414
rect 48092 5412 48116 5414
rect 48172 5412 48196 5414
rect 48252 5412 48258 5414
rect 47950 5403 48258 5412
rect 47950 4380 48258 4389
rect 47950 4378 47956 4380
rect 48012 4378 48036 4380
rect 48092 4378 48116 4380
rect 48172 4378 48196 4380
rect 48252 4378 48258 4380
rect 48012 4326 48014 4378
rect 48194 4326 48196 4378
rect 47950 4324 47956 4326
rect 48012 4324 48036 4326
rect 48092 4324 48116 4326
rect 48172 4324 48196 4326
rect 48252 4324 48258 4326
rect 47950 4315 48258 4324
rect 48596 4140 48648 4146
rect 48596 4082 48648 4088
rect 47950 3292 48258 3301
rect 47950 3290 47956 3292
rect 48012 3290 48036 3292
rect 48092 3290 48116 3292
rect 48172 3290 48196 3292
rect 48252 3290 48258 3292
rect 48012 3238 48014 3290
rect 48194 3238 48196 3290
rect 47950 3236 47956 3238
rect 48012 3236 48036 3238
rect 48092 3236 48116 3238
rect 48172 3236 48196 3238
rect 48252 3236 48258 3238
rect 47950 3227 48258 3236
rect 47860 3120 47912 3126
rect 47860 3062 47912 3068
rect 47860 2984 47912 2990
rect 47860 2926 47912 2932
rect 47768 2440 47820 2446
rect 47768 2382 47820 2388
rect 47872 800 47900 2926
rect 48320 2848 48372 2854
rect 48320 2790 48372 2796
rect 48332 2514 48360 2790
rect 48320 2508 48372 2514
rect 48320 2450 48372 2456
rect 47950 2204 48258 2213
rect 47950 2202 47956 2204
rect 48012 2202 48036 2204
rect 48092 2202 48116 2204
rect 48172 2202 48196 2204
rect 48252 2202 48258 2204
rect 48012 2150 48014 2202
rect 48194 2150 48196 2202
rect 47950 2148 47956 2150
rect 48012 2148 48036 2150
rect 48092 2148 48116 2150
rect 48172 2148 48196 2150
rect 48252 2148 48258 2150
rect 47950 2139 48258 2148
rect 48608 800 48636 4082
rect 48884 4010 48912 6886
rect 49148 6724 49200 6730
rect 49148 6666 49200 6672
rect 49160 6361 49188 6666
rect 49146 6352 49202 6361
rect 49146 6287 49202 6296
rect 49148 5704 49200 5710
rect 49146 5672 49148 5681
rect 49200 5672 49202 5681
rect 49146 5607 49202 5616
rect 49332 5024 49384 5030
rect 49330 4992 49332 5001
rect 49384 4992 49386 5001
rect 49330 4927 49386 4936
rect 49148 4548 49200 4554
rect 49148 4490 49200 4496
rect 49160 4321 49188 4490
rect 49146 4312 49202 4321
rect 49146 4247 49202 4256
rect 48872 4004 48924 4010
rect 48872 3946 48924 3952
rect 49332 3460 49384 3466
rect 49332 3402 49384 3408
rect 49344 800 49372 3402
rect 28092 734 28396 762
rect 28722 0 28778 800
rect 29458 0 29514 800
rect 30194 0 30250 800
rect 30930 0 30986 800
rect 31666 0 31722 800
rect 32402 0 32458 800
rect 33138 0 33194 800
rect 33874 0 33930 800
rect 34610 0 34666 800
rect 35346 0 35402 800
rect 36082 0 36138 800
rect 36818 0 36874 800
rect 37554 0 37610 800
rect 38290 0 38346 800
rect 39026 0 39082 800
rect 39762 0 39818 800
rect 40498 0 40554 800
rect 41234 0 41290 800
rect 41970 0 42026 800
rect 42706 0 42762 800
rect 43442 0 43498 800
rect 44178 0 44234 800
rect 44914 0 44970 800
rect 45650 0 45706 800
rect 46386 0 46442 800
rect 47122 0 47178 800
rect 47858 0 47914 800
rect 48594 0 48650 800
rect 49330 0 49386 800
<< via2 >>
rect 938 52672 994 52728
rect 2778 54984 2834 55040
rect 938 50360 994 50416
rect 938 48068 994 48104
rect 938 48048 940 48068
rect 940 48048 992 48068
rect 992 48048 994 48068
rect 938 45736 994 45792
rect 938 43424 994 43480
rect 2956 53882 3012 53884
rect 3036 53882 3092 53884
rect 3116 53882 3172 53884
rect 3196 53882 3252 53884
rect 2956 53830 3002 53882
rect 3002 53830 3012 53882
rect 3036 53830 3066 53882
rect 3066 53830 3078 53882
rect 3078 53830 3092 53882
rect 3116 53830 3130 53882
rect 3130 53830 3142 53882
rect 3142 53830 3172 53882
rect 3196 53830 3206 53882
rect 3206 53830 3252 53882
rect 2956 53828 3012 53830
rect 3036 53828 3092 53830
rect 3116 53828 3172 53830
rect 3196 53828 3252 53830
rect 2956 52794 3012 52796
rect 3036 52794 3092 52796
rect 3116 52794 3172 52796
rect 3196 52794 3252 52796
rect 2956 52742 3002 52794
rect 3002 52742 3012 52794
rect 3036 52742 3066 52794
rect 3066 52742 3078 52794
rect 3078 52742 3092 52794
rect 3116 52742 3130 52794
rect 3130 52742 3142 52794
rect 3142 52742 3172 52794
rect 3196 52742 3206 52794
rect 3206 52742 3252 52794
rect 2956 52740 3012 52742
rect 3036 52740 3092 52742
rect 3116 52740 3172 52742
rect 3196 52740 3252 52742
rect 2956 51706 3012 51708
rect 3036 51706 3092 51708
rect 3116 51706 3172 51708
rect 3196 51706 3252 51708
rect 2956 51654 3002 51706
rect 3002 51654 3012 51706
rect 3036 51654 3066 51706
rect 3066 51654 3078 51706
rect 3078 51654 3092 51706
rect 3116 51654 3130 51706
rect 3130 51654 3142 51706
rect 3142 51654 3172 51706
rect 3196 51654 3206 51706
rect 3206 51654 3252 51706
rect 2956 51652 3012 51654
rect 3036 51652 3092 51654
rect 3116 51652 3172 51654
rect 3196 51652 3252 51654
rect 1674 41112 1730 41168
rect 2956 50618 3012 50620
rect 3036 50618 3092 50620
rect 3116 50618 3172 50620
rect 3196 50618 3252 50620
rect 2956 50566 3002 50618
rect 3002 50566 3012 50618
rect 3036 50566 3066 50618
rect 3066 50566 3078 50618
rect 3078 50566 3092 50618
rect 3116 50566 3130 50618
rect 3130 50566 3142 50618
rect 3142 50566 3172 50618
rect 3196 50566 3206 50618
rect 3206 50566 3252 50618
rect 2956 50564 3012 50566
rect 3036 50564 3092 50566
rect 3116 50564 3172 50566
rect 3196 50564 3252 50566
rect 2956 49530 3012 49532
rect 3036 49530 3092 49532
rect 3116 49530 3172 49532
rect 3196 49530 3252 49532
rect 2956 49478 3002 49530
rect 3002 49478 3012 49530
rect 3036 49478 3066 49530
rect 3066 49478 3078 49530
rect 3078 49478 3092 49530
rect 3116 49478 3130 49530
rect 3130 49478 3142 49530
rect 3142 49478 3172 49530
rect 3196 49478 3206 49530
rect 3206 49478 3252 49530
rect 2956 49476 3012 49478
rect 3036 49476 3092 49478
rect 3116 49476 3172 49478
rect 3196 49476 3252 49478
rect 2956 48442 3012 48444
rect 3036 48442 3092 48444
rect 3116 48442 3172 48444
rect 3196 48442 3252 48444
rect 2956 48390 3002 48442
rect 3002 48390 3012 48442
rect 3036 48390 3066 48442
rect 3066 48390 3078 48442
rect 3078 48390 3092 48442
rect 3116 48390 3130 48442
rect 3130 48390 3142 48442
rect 3142 48390 3172 48442
rect 3196 48390 3206 48442
rect 3206 48390 3252 48442
rect 2956 48388 3012 48390
rect 3036 48388 3092 48390
rect 3116 48388 3172 48390
rect 3196 48388 3252 48390
rect 2956 47354 3012 47356
rect 3036 47354 3092 47356
rect 3116 47354 3172 47356
rect 3196 47354 3252 47356
rect 2956 47302 3002 47354
rect 3002 47302 3012 47354
rect 3036 47302 3066 47354
rect 3066 47302 3078 47354
rect 3078 47302 3092 47354
rect 3116 47302 3130 47354
rect 3130 47302 3142 47354
rect 3142 47302 3172 47354
rect 3196 47302 3206 47354
rect 3206 47302 3252 47354
rect 2956 47300 3012 47302
rect 3036 47300 3092 47302
rect 3116 47300 3172 47302
rect 3196 47300 3252 47302
rect 2956 46266 3012 46268
rect 3036 46266 3092 46268
rect 3116 46266 3172 46268
rect 3196 46266 3252 46268
rect 2956 46214 3002 46266
rect 3002 46214 3012 46266
rect 3036 46214 3066 46266
rect 3066 46214 3078 46266
rect 3078 46214 3092 46266
rect 3116 46214 3130 46266
rect 3130 46214 3142 46266
rect 3142 46214 3172 46266
rect 3196 46214 3206 46266
rect 3206 46214 3252 46266
rect 2956 46212 3012 46214
rect 3036 46212 3092 46214
rect 3116 46212 3172 46214
rect 3196 46212 3252 46214
rect 2956 45178 3012 45180
rect 3036 45178 3092 45180
rect 3116 45178 3172 45180
rect 3196 45178 3252 45180
rect 2956 45126 3002 45178
rect 3002 45126 3012 45178
rect 3036 45126 3066 45178
rect 3066 45126 3078 45178
rect 3078 45126 3092 45178
rect 3116 45126 3130 45178
rect 3130 45126 3142 45178
rect 3142 45126 3172 45178
rect 3196 45126 3206 45178
rect 3206 45126 3252 45178
rect 2956 45124 3012 45126
rect 3036 45124 3092 45126
rect 3116 45124 3172 45126
rect 3196 45124 3252 45126
rect 2956 44090 3012 44092
rect 3036 44090 3092 44092
rect 3116 44090 3172 44092
rect 3196 44090 3252 44092
rect 2956 44038 3002 44090
rect 3002 44038 3012 44090
rect 3036 44038 3066 44090
rect 3066 44038 3078 44090
rect 3078 44038 3092 44090
rect 3116 44038 3130 44090
rect 3130 44038 3142 44090
rect 3142 44038 3172 44090
rect 3196 44038 3206 44090
rect 3206 44038 3252 44090
rect 2956 44036 3012 44038
rect 3036 44036 3092 44038
rect 3116 44036 3172 44038
rect 3196 44036 3252 44038
rect 2956 43002 3012 43004
rect 3036 43002 3092 43004
rect 3116 43002 3172 43004
rect 3196 43002 3252 43004
rect 2956 42950 3002 43002
rect 3002 42950 3012 43002
rect 3036 42950 3066 43002
rect 3066 42950 3078 43002
rect 3078 42950 3092 43002
rect 3116 42950 3130 43002
rect 3130 42950 3142 43002
rect 3142 42950 3172 43002
rect 3196 42950 3206 43002
rect 3206 42950 3252 43002
rect 2956 42948 3012 42950
rect 3036 42948 3092 42950
rect 3116 42948 3172 42950
rect 3196 42948 3252 42950
rect 2956 41914 3012 41916
rect 3036 41914 3092 41916
rect 3116 41914 3172 41916
rect 3196 41914 3252 41916
rect 2956 41862 3002 41914
rect 3002 41862 3012 41914
rect 3036 41862 3066 41914
rect 3066 41862 3078 41914
rect 3078 41862 3092 41914
rect 3116 41862 3130 41914
rect 3130 41862 3142 41914
rect 3142 41862 3172 41914
rect 3196 41862 3206 41914
rect 3206 41862 3252 41914
rect 2956 41860 3012 41862
rect 3036 41860 3092 41862
rect 3116 41860 3172 41862
rect 3196 41860 3252 41862
rect 7956 54426 8012 54428
rect 8036 54426 8092 54428
rect 8116 54426 8172 54428
rect 8196 54426 8252 54428
rect 7956 54374 8002 54426
rect 8002 54374 8012 54426
rect 8036 54374 8066 54426
rect 8066 54374 8078 54426
rect 8078 54374 8092 54426
rect 8116 54374 8130 54426
rect 8130 54374 8142 54426
rect 8142 54374 8172 54426
rect 8196 54374 8206 54426
rect 8206 54374 8252 54426
rect 7956 54372 8012 54374
rect 8036 54372 8092 54374
rect 8116 54372 8172 54374
rect 8196 54372 8252 54374
rect 7956 53338 8012 53340
rect 8036 53338 8092 53340
rect 8116 53338 8172 53340
rect 8196 53338 8252 53340
rect 7956 53286 8002 53338
rect 8002 53286 8012 53338
rect 8036 53286 8066 53338
rect 8066 53286 8078 53338
rect 8078 53286 8092 53338
rect 8116 53286 8130 53338
rect 8130 53286 8142 53338
rect 8142 53286 8172 53338
rect 8196 53286 8206 53338
rect 8206 53286 8252 53338
rect 7956 53284 8012 53286
rect 8036 53284 8092 53286
rect 8116 53284 8172 53286
rect 8196 53284 8252 53286
rect 7956 52250 8012 52252
rect 8036 52250 8092 52252
rect 8116 52250 8172 52252
rect 8196 52250 8252 52252
rect 7956 52198 8002 52250
rect 8002 52198 8012 52250
rect 8036 52198 8066 52250
rect 8066 52198 8078 52250
rect 8078 52198 8092 52250
rect 8116 52198 8130 52250
rect 8130 52198 8142 52250
rect 8142 52198 8172 52250
rect 8196 52198 8206 52250
rect 8206 52198 8252 52250
rect 7956 52196 8012 52198
rect 8036 52196 8092 52198
rect 8116 52196 8172 52198
rect 8196 52196 8252 52198
rect 7956 51162 8012 51164
rect 8036 51162 8092 51164
rect 8116 51162 8172 51164
rect 8196 51162 8252 51164
rect 7956 51110 8002 51162
rect 8002 51110 8012 51162
rect 8036 51110 8066 51162
rect 8066 51110 8078 51162
rect 8078 51110 8092 51162
rect 8116 51110 8130 51162
rect 8130 51110 8142 51162
rect 8142 51110 8172 51162
rect 8196 51110 8206 51162
rect 8206 51110 8252 51162
rect 7956 51108 8012 51110
rect 8036 51108 8092 51110
rect 8116 51108 8172 51110
rect 8196 51108 8252 51110
rect 7956 50074 8012 50076
rect 8036 50074 8092 50076
rect 8116 50074 8172 50076
rect 8196 50074 8252 50076
rect 7956 50022 8002 50074
rect 8002 50022 8012 50074
rect 8036 50022 8066 50074
rect 8066 50022 8078 50074
rect 8078 50022 8092 50074
rect 8116 50022 8130 50074
rect 8130 50022 8142 50074
rect 8142 50022 8172 50074
rect 8196 50022 8206 50074
rect 8206 50022 8252 50074
rect 7956 50020 8012 50022
rect 8036 50020 8092 50022
rect 8116 50020 8172 50022
rect 8196 50020 8252 50022
rect 7956 48986 8012 48988
rect 8036 48986 8092 48988
rect 8116 48986 8172 48988
rect 8196 48986 8252 48988
rect 7956 48934 8002 48986
rect 8002 48934 8012 48986
rect 8036 48934 8066 48986
rect 8066 48934 8078 48986
rect 8078 48934 8092 48986
rect 8116 48934 8130 48986
rect 8130 48934 8142 48986
rect 8142 48934 8172 48986
rect 8196 48934 8206 48986
rect 8206 48934 8252 48986
rect 7956 48932 8012 48934
rect 8036 48932 8092 48934
rect 8116 48932 8172 48934
rect 8196 48932 8252 48934
rect 7956 47898 8012 47900
rect 8036 47898 8092 47900
rect 8116 47898 8172 47900
rect 8196 47898 8252 47900
rect 7956 47846 8002 47898
rect 8002 47846 8012 47898
rect 8036 47846 8066 47898
rect 8066 47846 8078 47898
rect 8078 47846 8092 47898
rect 8116 47846 8130 47898
rect 8130 47846 8142 47898
rect 8142 47846 8172 47898
rect 8196 47846 8206 47898
rect 8206 47846 8252 47898
rect 7956 47844 8012 47846
rect 8036 47844 8092 47846
rect 8116 47844 8172 47846
rect 8196 47844 8252 47846
rect 7956 46810 8012 46812
rect 8036 46810 8092 46812
rect 8116 46810 8172 46812
rect 8196 46810 8252 46812
rect 7956 46758 8002 46810
rect 8002 46758 8012 46810
rect 8036 46758 8066 46810
rect 8066 46758 8078 46810
rect 8078 46758 8092 46810
rect 8116 46758 8130 46810
rect 8130 46758 8142 46810
rect 8142 46758 8172 46810
rect 8196 46758 8206 46810
rect 8206 46758 8252 46810
rect 7956 46756 8012 46758
rect 8036 46756 8092 46758
rect 8116 46756 8172 46758
rect 8196 46756 8252 46758
rect 7956 45722 8012 45724
rect 8036 45722 8092 45724
rect 8116 45722 8172 45724
rect 8196 45722 8252 45724
rect 7956 45670 8002 45722
rect 8002 45670 8012 45722
rect 8036 45670 8066 45722
rect 8066 45670 8078 45722
rect 8078 45670 8092 45722
rect 8116 45670 8130 45722
rect 8130 45670 8142 45722
rect 8142 45670 8172 45722
rect 8196 45670 8206 45722
rect 8206 45670 8252 45722
rect 7956 45668 8012 45670
rect 8036 45668 8092 45670
rect 8116 45668 8172 45670
rect 8196 45668 8252 45670
rect 7956 44634 8012 44636
rect 8036 44634 8092 44636
rect 8116 44634 8172 44636
rect 8196 44634 8252 44636
rect 7956 44582 8002 44634
rect 8002 44582 8012 44634
rect 8036 44582 8066 44634
rect 8066 44582 8078 44634
rect 8078 44582 8092 44634
rect 8116 44582 8130 44634
rect 8130 44582 8142 44634
rect 8142 44582 8172 44634
rect 8196 44582 8206 44634
rect 8206 44582 8252 44634
rect 7956 44580 8012 44582
rect 8036 44580 8092 44582
rect 8116 44580 8172 44582
rect 8196 44580 8252 44582
rect 7956 43546 8012 43548
rect 8036 43546 8092 43548
rect 8116 43546 8172 43548
rect 8196 43546 8252 43548
rect 7956 43494 8002 43546
rect 8002 43494 8012 43546
rect 8036 43494 8066 43546
rect 8066 43494 8078 43546
rect 8078 43494 8092 43546
rect 8116 43494 8130 43546
rect 8130 43494 8142 43546
rect 8142 43494 8172 43546
rect 8196 43494 8206 43546
rect 8206 43494 8252 43546
rect 7956 43492 8012 43494
rect 8036 43492 8092 43494
rect 8116 43492 8172 43494
rect 8196 43492 8252 43494
rect 7956 42458 8012 42460
rect 8036 42458 8092 42460
rect 8116 42458 8172 42460
rect 8196 42458 8252 42460
rect 7956 42406 8002 42458
rect 8002 42406 8012 42458
rect 8036 42406 8066 42458
rect 8066 42406 8078 42458
rect 8078 42406 8092 42458
rect 8116 42406 8130 42458
rect 8130 42406 8142 42458
rect 8142 42406 8172 42458
rect 8196 42406 8206 42458
rect 8206 42406 8252 42458
rect 7956 42404 8012 42406
rect 8036 42404 8092 42406
rect 8116 42404 8172 42406
rect 8196 42404 8252 42406
rect 2956 40826 3012 40828
rect 3036 40826 3092 40828
rect 3116 40826 3172 40828
rect 3196 40826 3252 40828
rect 2956 40774 3002 40826
rect 3002 40774 3012 40826
rect 3036 40774 3066 40826
rect 3066 40774 3078 40826
rect 3078 40774 3092 40826
rect 3116 40774 3130 40826
rect 3130 40774 3142 40826
rect 3142 40774 3172 40826
rect 3196 40774 3206 40826
rect 3206 40774 3252 40826
rect 2956 40772 3012 40774
rect 3036 40772 3092 40774
rect 3116 40772 3172 40774
rect 3196 40772 3252 40774
rect 2956 39738 3012 39740
rect 3036 39738 3092 39740
rect 3116 39738 3172 39740
rect 3196 39738 3252 39740
rect 2956 39686 3002 39738
rect 3002 39686 3012 39738
rect 3036 39686 3066 39738
rect 3066 39686 3078 39738
rect 3078 39686 3092 39738
rect 3116 39686 3130 39738
rect 3130 39686 3142 39738
rect 3142 39686 3172 39738
rect 3196 39686 3206 39738
rect 3206 39686 3252 39738
rect 2956 39684 3012 39686
rect 3036 39684 3092 39686
rect 3116 39684 3172 39686
rect 3196 39684 3252 39686
rect 938 38800 994 38856
rect 2956 38650 3012 38652
rect 3036 38650 3092 38652
rect 3116 38650 3172 38652
rect 3196 38650 3252 38652
rect 2956 38598 3002 38650
rect 3002 38598 3012 38650
rect 3036 38598 3066 38650
rect 3066 38598 3078 38650
rect 3078 38598 3092 38650
rect 3116 38598 3130 38650
rect 3130 38598 3142 38650
rect 3142 38598 3172 38650
rect 3196 38598 3206 38650
rect 3206 38598 3252 38650
rect 2956 38596 3012 38598
rect 3036 38596 3092 38598
rect 3116 38596 3172 38598
rect 3196 38596 3252 38598
rect 2956 37562 3012 37564
rect 3036 37562 3092 37564
rect 3116 37562 3172 37564
rect 3196 37562 3252 37564
rect 2956 37510 3002 37562
rect 3002 37510 3012 37562
rect 3036 37510 3066 37562
rect 3066 37510 3078 37562
rect 3078 37510 3092 37562
rect 3116 37510 3130 37562
rect 3130 37510 3142 37562
rect 3142 37510 3172 37562
rect 3196 37510 3206 37562
rect 3206 37510 3252 37562
rect 2956 37508 3012 37510
rect 3036 37508 3092 37510
rect 3116 37508 3172 37510
rect 3196 37508 3252 37510
rect 938 36488 994 36544
rect 2956 36474 3012 36476
rect 3036 36474 3092 36476
rect 3116 36474 3172 36476
rect 3196 36474 3252 36476
rect 2956 36422 3002 36474
rect 3002 36422 3012 36474
rect 3036 36422 3066 36474
rect 3066 36422 3078 36474
rect 3078 36422 3092 36474
rect 3116 36422 3130 36474
rect 3130 36422 3142 36474
rect 3142 36422 3172 36474
rect 3196 36422 3206 36474
rect 3206 36422 3252 36474
rect 2956 36420 3012 36422
rect 3036 36420 3092 36422
rect 3116 36420 3172 36422
rect 3196 36420 3252 36422
rect 2956 35386 3012 35388
rect 3036 35386 3092 35388
rect 3116 35386 3172 35388
rect 3196 35386 3252 35388
rect 2956 35334 3002 35386
rect 3002 35334 3012 35386
rect 3036 35334 3066 35386
rect 3066 35334 3078 35386
rect 3078 35334 3092 35386
rect 3116 35334 3130 35386
rect 3130 35334 3142 35386
rect 3142 35334 3172 35386
rect 3196 35334 3206 35386
rect 3206 35334 3252 35386
rect 2956 35332 3012 35334
rect 3036 35332 3092 35334
rect 3116 35332 3172 35334
rect 3196 35332 3252 35334
rect 2956 34298 3012 34300
rect 3036 34298 3092 34300
rect 3116 34298 3172 34300
rect 3196 34298 3252 34300
rect 2956 34246 3002 34298
rect 3002 34246 3012 34298
rect 3036 34246 3066 34298
rect 3066 34246 3078 34298
rect 3078 34246 3092 34298
rect 3116 34246 3130 34298
rect 3130 34246 3142 34298
rect 3142 34246 3172 34298
rect 3196 34246 3206 34298
rect 3206 34246 3252 34298
rect 2956 34244 3012 34246
rect 3036 34244 3092 34246
rect 3116 34244 3172 34246
rect 3196 34244 3252 34246
rect 1766 34176 1822 34232
rect 2956 33210 3012 33212
rect 3036 33210 3092 33212
rect 3116 33210 3172 33212
rect 3196 33210 3252 33212
rect 2956 33158 3002 33210
rect 3002 33158 3012 33210
rect 3036 33158 3066 33210
rect 3066 33158 3078 33210
rect 3078 33158 3092 33210
rect 3116 33158 3130 33210
rect 3130 33158 3142 33210
rect 3142 33158 3172 33210
rect 3196 33158 3206 33210
rect 3206 33158 3252 33210
rect 2956 33156 3012 33158
rect 3036 33156 3092 33158
rect 3116 33156 3172 33158
rect 3196 33156 3252 33158
rect 2956 32122 3012 32124
rect 3036 32122 3092 32124
rect 3116 32122 3172 32124
rect 3196 32122 3252 32124
rect 2956 32070 3002 32122
rect 3002 32070 3012 32122
rect 3036 32070 3066 32122
rect 3066 32070 3078 32122
rect 3078 32070 3092 32122
rect 3116 32070 3130 32122
rect 3130 32070 3142 32122
rect 3142 32070 3172 32122
rect 3196 32070 3206 32122
rect 3206 32070 3252 32122
rect 2956 32068 3012 32070
rect 3036 32068 3092 32070
rect 3116 32068 3172 32070
rect 3196 32068 3252 32070
rect 938 31864 994 31920
rect 2956 31034 3012 31036
rect 3036 31034 3092 31036
rect 3116 31034 3172 31036
rect 3196 31034 3252 31036
rect 2956 30982 3002 31034
rect 3002 30982 3012 31034
rect 3036 30982 3066 31034
rect 3066 30982 3078 31034
rect 3078 30982 3092 31034
rect 3116 30982 3130 31034
rect 3130 30982 3142 31034
rect 3142 30982 3172 31034
rect 3196 30982 3206 31034
rect 3206 30982 3252 31034
rect 2956 30980 3012 30982
rect 3036 30980 3092 30982
rect 3116 30980 3172 30982
rect 3196 30980 3252 30982
rect 2956 29946 3012 29948
rect 3036 29946 3092 29948
rect 3116 29946 3172 29948
rect 3196 29946 3252 29948
rect 2956 29894 3002 29946
rect 3002 29894 3012 29946
rect 3036 29894 3066 29946
rect 3066 29894 3078 29946
rect 3078 29894 3092 29946
rect 3116 29894 3130 29946
rect 3130 29894 3142 29946
rect 3142 29894 3172 29946
rect 3196 29894 3206 29946
rect 3206 29894 3252 29946
rect 2956 29892 3012 29894
rect 3036 29892 3092 29894
rect 3116 29892 3172 29894
rect 3196 29892 3252 29894
rect 1306 29552 1362 29608
rect 2956 28858 3012 28860
rect 3036 28858 3092 28860
rect 3116 28858 3172 28860
rect 3196 28858 3252 28860
rect 2956 28806 3002 28858
rect 3002 28806 3012 28858
rect 3036 28806 3066 28858
rect 3066 28806 3078 28858
rect 3078 28806 3092 28858
rect 3116 28806 3130 28858
rect 3130 28806 3142 28858
rect 3142 28806 3172 28858
rect 3196 28806 3206 28858
rect 3206 28806 3252 28858
rect 2956 28804 3012 28806
rect 3036 28804 3092 28806
rect 3116 28804 3172 28806
rect 3196 28804 3252 28806
rect 7956 41370 8012 41372
rect 8036 41370 8092 41372
rect 8116 41370 8172 41372
rect 8196 41370 8252 41372
rect 7956 41318 8002 41370
rect 8002 41318 8012 41370
rect 8036 41318 8066 41370
rect 8066 41318 8078 41370
rect 8078 41318 8092 41370
rect 8116 41318 8130 41370
rect 8130 41318 8142 41370
rect 8142 41318 8172 41370
rect 8196 41318 8206 41370
rect 8206 41318 8252 41370
rect 7956 41316 8012 41318
rect 8036 41316 8092 41318
rect 8116 41316 8172 41318
rect 8196 41316 8252 41318
rect 7956 40282 8012 40284
rect 8036 40282 8092 40284
rect 8116 40282 8172 40284
rect 8196 40282 8252 40284
rect 7956 40230 8002 40282
rect 8002 40230 8012 40282
rect 8036 40230 8066 40282
rect 8066 40230 8078 40282
rect 8078 40230 8092 40282
rect 8116 40230 8130 40282
rect 8130 40230 8142 40282
rect 8142 40230 8172 40282
rect 8196 40230 8206 40282
rect 8206 40230 8252 40282
rect 7956 40228 8012 40230
rect 8036 40228 8092 40230
rect 8116 40228 8172 40230
rect 8196 40228 8252 40230
rect 7956 39194 8012 39196
rect 8036 39194 8092 39196
rect 8116 39194 8172 39196
rect 8196 39194 8252 39196
rect 7956 39142 8002 39194
rect 8002 39142 8012 39194
rect 8036 39142 8066 39194
rect 8066 39142 8078 39194
rect 8078 39142 8092 39194
rect 8116 39142 8130 39194
rect 8130 39142 8142 39194
rect 8142 39142 8172 39194
rect 8196 39142 8206 39194
rect 8206 39142 8252 39194
rect 7956 39140 8012 39142
rect 8036 39140 8092 39142
rect 8116 39140 8172 39142
rect 8196 39140 8252 39142
rect 7956 38106 8012 38108
rect 8036 38106 8092 38108
rect 8116 38106 8172 38108
rect 8196 38106 8252 38108
rect 7956 38054 8002 38106
rect 8002 38054 8012 38106
rect 8036 38054 8066 38106
rect 8066 38054 8078 38106
rect 8078 38054 8092 38106
rect 8116 38054 8130 38106
rect 8130 38054 8142 38106
rect 8142 38054 8172 38106
rect 8196 38054 8206 38106
rect 8206 38054 8252 38106
rect 7956 38052 8012 38054
rect 8036 38052 8092 38054
rect 8116 38052 8172 38054
rect 8196 38052 8252 38054
rect 7956 37018 8012 37020
rect 8036 37018 8092 37020
rect 8116 37018 8172 37020
rect 8196 37018 8252 37020
rect 7956 36966 8002 37018
rect 8002 36966 8012 37018
rect 8036 36966 8066 37018
rect 8066 36966 8078 37018
rect 8078 36966 8092 37018
rect 8116 36966 8130 37018
rect 8130 36966 8142 37018
rect 8142 36966 8172 37018
rect 8196 36966 8206 37018
rect 8206 36966 8252 37018
rect 7956 36964 8012 36966
rect 8036 36964 8092 36966
rect 8116 36964 8172 36966
rect 8196 36964 8252 36966
rect 2956 27770 3012 27772
rect 3036 27770 3092 27772
rect 3116 27770 3172 27772
rect 3196 27770 3252 27772
rect 2956 27718 3002 27770
rect 3002 27718 3012 27770
rect 3036 27718 3066 27770
rect 3066 27718 3078 27770
rect 3078 27718 3092 27770
rect 3116 27718 3130 27770
rect 3130 27718 3142 27770
rect 3142 27718 3172 27770
rect 3196 27718 3206 27770
rect 3206 27718 3252 27770
rect 2956 27716 3012 27718
rect 3036 27716 3092 27718
rect 3116 27716 3172 27718
rect 3196 27716 3252 27718
rect 1306 27240 1362 27296
rect 2956 26682 3012 26684
rect 3036 26682 3092 26684
rect 3116 26682 3172 26684
rect 3196 26682 3252 26684
rect 2956 26630 3002 26682
rect 3002 26630 3012 26682
rect 3036 26630 3066 26682
rect 3066 26630 3078 26682
rect 3078 26630 3092 26682
rect 3116 26630 3130 26682
rect 3130 26630 3142 26682
rect 3142 26630 3172 26682
rect 3196 26630 3206 26682
rect 3206 26630 3252 26682
rect 2956 26628 3012 26630
rect 3036 26628 3092 26630
rect 3116 26628 3172 26630
rect 3196 26628 3252 26630
rect 2956 25594 3012 25596
rect 3036 25594 3092 25596
rect 3116 25594 3172 25596
rect 3196 25594 3252 25596
rect 2956 25542 3002 25594
rect 3002 25542 3012 25594
rect 3036 25542 3066 25594
rect 3066 25542 3078 25594
rect 3078 25542 3092 25594
rect 3116 25542 3130 25594
rect 3130 25542 3142 25594
rect 3142 25542 3172 25594
rect 3196 25542 3206 25594
rect 3206 25542 3252 25594
rect 2956 25540 3012 25542
rect 3036 25540 3092 25542
rect 3116 25540 3172 25542
rect 3196 25540 3252 25542
rect 1306 24928 1362 24984
rect 2956 24506 3012 24508
rect 3036 24506 3092 24508
rect 3116 24506 3172 24508
rect 3196 24506 3252 24508
rect 2956 24454 3002 24506
rect 3002 24454 3012 24506
rect 3036 24454 3066 24506
rect 3066 24454 3078 24506
rect 3078 24454 3092 24506
rect 3116 24454 3130 24506
rect 3130 24454 3142 24506
rect 3142 24454 3172 24506
rect 3196 24454 3206 24506
rect 3206 24454 3252 24506
rect 2956 24452 3012 24454
rect 3036 24452 3092 24454
rect 3116 24452 3172 24454
rect 3196 24452 3252 24454
rect 2956 23418 3012 23420
rect 3036 23418 3092 23420
rect 3116 23418 3172 23420
rect 3196 23418 3252 23420
rect 2956 23366 3002 23418
rect 3002 23366 3012 23418
rect 3036 23366 3066 23418
rect 3066 23366 3078 23418
rect 3078 23366 3092 23418
rect 3116 23366 3130 23418
rect 3130 23366 3142 23418
rect 3142 23366 3172 23418
rect 3196 23366 3206 23418
rect 3206 23366 3252 23418
rect 2956 23364 3012 23366
rect 3036 23364 3092 23366
rect 3116 23364 3172 23366
rect 3196 23364 3252 23366
rect 7956 35930 8012 35932
rect 8036 35930 8092 35932
rect 8116 35930 8172 35932
rect 8196 35930 8252 35932
rect 7956 35878 8002 35930
rect 8002 35878 8012 35930
rect 8036 35878 8066 35930
rect 8066 35878 8078 35930
rect 8078 35878 8092 35930
rect 8116 35878 8130 35930
rect 8130 35878 8142 35930
rect 8142 35878 8172 35930
rect 8196 35878 8206 35930
rect 8206 35878 8252 35930
rect 7956 35876 8012 35878
rect 8036 35876 8092 35878
rect 8116 35876 8172 35878
rect 8196 35876 8252 35878
rect 7956 34842 8012 34844
rect 8036 34842 8092 34844
rect 8116 34842 8172 34844
rect 8196 34842 8252 34844
rect 7956 34790 8002 34842
rect 8002 34790 8012 34842
rect 8036 34790 8066 34842
rect 8066 34790 8078 34842
rect 8078 34790 8092 34842
rect 8116 34790 8130 34842
rect 8130 34790 8142 34842
rect 8142 34790 8172 34842
rect 8196 34790 8206 34842
rect 8206 34790 8252 34842
rect 7956 34788 8012 34790
rect 8036 34788 8092 34790
rect 8116 34788 8172 34790
rect 8196 34788 8252 34790
rect 7956 33754 8012 33756
rect 8036 33754 8092 33756
rect 8116 33754 8172 33756
rect 8196 33754 8252 33756
rect 7956 33702 8002 33754
rect 8002 33702 8012 33754
rect 8036 33702 8066 33754
rect 8066 33702 8078 33754
rect 8078 33702 8092 33754
rect 8116 33702 8130 33754
rect 8130 33702 8142 33754
rect 8142 33702 8172 33754
rect 8196 33702 8206 33754
rect 8206 33702 8252 33754
rect 7956 33700 8012 33702
rect 8036 33700 8092 33702
rect 8116 33700 8172 33702
rect 8196 33700 8252 33702
rect 7956 32666 8012 32668
rect 8036 32666 8092 32668
rect 8116 32666 8172 32668
rect 8196 32666 8252 32668
rect 7956 32614 8002 32666
rect 8002 32614 8012 32666
rect 8036 32614 8066 32666
rect 8066 32614 8078 32666
rect 8078 32614 8092 32666
rect 8116 32614 8130 32666
rect 8130 32614 8142 32666
rect 8142 32614 8172 32666
rect 8196 32614 8206 32666
rect 8206 32614 8252 32666
rect 7956 32612 8012 32614
rect 8036 32612 8092 32614
rect 8116 32612 8172 32614
rect 8196 32612 8252 32614
rect 7956 31578 8012 31580
rect 8036 31578 8092 31580
rect 8116 31578 8172 31580
rect 8196 31578 8252 31580
rect 7956 31526 8002 31578
rect 8002 31526 8012 31578
rect 8036 31526 8066 31578
rect 8066 31526 8078 31578
rect 8078 31526 8092 31578
rect 8116 31526 8130 31578
rect 8130 31526 8142 31578
rect 8142 31526 8172 31578
rect 8196 31526 8206 31578
rect 8206 31526 8252 31578
rect 7956 31524 8012 31526
rect 8036 31524 8092 31526
rect 8116 31524 8172 31526
rect 8196 31524 8252 31526
rect 9770 31184 9826 31240
rect 7956 30490 8012 30492
rect 8036 30490 8092 30492
rect 8116 30490 8172 30492
rect 8196 30490 8252 30492
rect 7956 30438 8002 30490
rect 8002 30438 8012 30490
rect 8036 30438 8066 30490
rect 8066 30438 8078 30490
rect 8078 30438 8092 30490
rect 8116 30438 8130 30490
rect 8130 30438 8142 30490
rect 8142 30438 8172 30490
rect 8196 30438 8206 30490
rect 8206 30438 8252 30490
rect 7956 30436 8012 30438
rect 8036 30436 8092 30438
rect 8116 30436 8172 30438
rect 8196 30436 8252 30438
rect 7956 29402 8012 29404
rect 8036 29402 8092 29404
rect 8116 29402 8172 29404
rect 8196 29402 8252 29404
rect 7956 29350 8002 29402
rect 8002 29350 8012 29402
rect 8036 29350 8066 29402
rect 8066 29350 8078 29402
rect 8078 29350 8092 29402
rect 8116 29350 8130 29402
rect 8130 29350 8142 29402
rect 8142 29350 8172 29402
rect 8196 29350 8206 29402
rect 8206 29350 8252 29402
rect 7956 29348 8012 29350
rect 8036 29348 8092 29350
rect 8116 29348 8172 29350
rect 8196 29348 8252 29350
rect 7956 28314 8012 28316
rect 8036 28314 8092 28316
rect 8116 28314 8172 28316
rect 8196 28314 8252 28316
rect 7956 28262 8002 28314
rect 8002 28262 8012 28314
rect 8036 28262 8066 28314
rect 8066 28262 8078 28314
rect 8078 28262 8092 28314
rect 8116 28262 8130 28314
rect 8130 28262 8142 28314
rect 8142 28262 8172 28314
rect 8196 28262 8206 28314
rect 8206 28262 8252 28314
rect 7956 28260 8012 28262
rect 8036 28260 8092 28262
rect 8116 28260 8172 28262
rect 8196 28260 8252 28262
rect 7956 27226 8012 27228
rect 8036 27226 8092 27228
rect 8116 27226 8172 27228
rect 8196 27226 8252 27228
rect 7956 27174 8002 27226
rect 8002 27174 8012 27226
rect 8036 27174 8066 27226
rect 8066 27174 8078 27226
rect 8078 27174 8092 27226
rect 8116 27174 8130 27226
rect 8130 27174 8142 27226
rect 8142 27174 8172 27226
rect 8196 27174 8206 27226
rect 8206 27174 8252 27226
rect 7956 27172 8012 27174
rect 8036 27172 8092 27174
rect 8116 27172 8172 27174
rect 8196 27172 8252 27174
rect 7956 26138 8012 26140
rect 8036 26138 8092 26140
rect 8116 26138 8172 26140
rect 8196 26138 8252 26140
rect 7956 26086 8002 26138
rect 8002 26086 8012 26138
rect 8036 26086 8066 26138
rect 8066 26086 8078 26138
rect 8078 26086 8092 26138
rect 8116 26086 8130 26138
rect 8130 26086 8142 26138
rect 8142 26086 8172 26138
rect 8196 26086 8206 26138
rect 8206 26086 8252 26138
rect 7956 26084 8012 26086
rect 8036 26084 8092 26086
rect 8116 26084 8172 26086
rect 8196 26084 8252 26086
rect 7956 25050 8012 25052
rect 8036 25050 8092 25052
rect 8116 25050 8172 25052
rect 8196 25050 8252 25052
rect 7956 24998 8002 25050
rect 8002 24998 8012 25050
rect 8036 24998 8066 25050
rect 8066 24998 8078 25050
rect 8078 24998 8092 25050
rect 8116 24998 8130 25050
rect 8130 24998 8142 25050
rect 8142 24998 8172 25050
rect 8196 24998 8206 25050
rect 8206 24998 8252 25050
rect 7956 24996 8012 24998
rect 8036 24996 8092 24998
rect 8116 24996 8172 24998
rect 8196 24996 8252 24998
rect 8850 24928 8906 24984
rect 7956 23962 8012 23964
rect 8036 23962 8092 23964
rect 8116 23962 8172 23964
rect 8196 23962 8252 23964
rect 7956 23910 8002 23962
rect 8002 23910 8012 23962
rect 8036 23910 8066 23962
rect 8066 23910 8078 23962
rect 8078 23910 8092 23962
rect 8116 23910 8130 23962
rect 8130 23910 8142 23962
rect 8142 23910 8172 23962
rect 8196 23910 8206 23962
rect 8206 23910 8252 23962
rect 7956 23908 8012 23910
rect 8036 23908 8092 23910
rect 8116 23908 8172 23910
rect 8196 23908 8252 23910
rect 1306 22616 1362 22672
rect 2956 22330 3012 22332
rect 3036 22330 3092 22332
rect 3116 22330 3172 22332
rect 3196 22330 3252 22332
rect 2956 22278 3002 22330
rect 3002 22278 3012 22330
rect 3036 22278 3066 22330
rect 3066 22278 3078 22330
rect 3078 22278 3092 22330
rect 3116 22278 3130 22330
rect 3130 22278 3142 22330
rect 3142 22278 3172 22330
rect 3196 22278 3206 22330
rect 3206 22278 3252 22330
rect 2956 22276 3012 22278
rect 3036 22276 3092 22278
rect 3116 22276 3172 22278
rect 3196 22276 3252 22278
rect 2956 21242 3012 21244
rect 3036 21242 3092 21244
rect 3116 21242 3172 21244
rect 3196 21242 3252 21244
rect 2956 21190 3002 21242
rect 3002 21190 3012 21242
rect 3036 21190 3066 21242
rect 3066 21190 3078 21242
rect 3078 21190 3092 21242
rect 3116 21190 3130 21242
rect 3130 21190 3142 21242
rect 3142 21190 3172 21242
rect 3196 21190 3206 21242
rect 3206 21190 3252 21242
rect 2956 21188 3012 21190
rect 3036 21188 3092 21190
rect 3116 21188 3172 21190
rect 3196 21188 3252 21190
rect 7956 22874 8012 22876
rect 8036 22874 8092 22876
rect 8116 22874 8172 22876
rect 8196 22874 8252 22876
rect 7956 22822 8002 22874
rect 8002 22822 8012 22874
rect 8036 22822 8066 22874
rect 8066 22822 8078 22874
rect 8078 22822 8092 22874
rect 8116 22822 8130 22874
rect 8130 22822 8142 22874
rect 8142 22822 8172 22874
rect 8196 22822 8206 22874
rect 8206 22822 8252 22874
rect 7956 22820 8012 22822
rect 8036 22820 8092 22822
rect 8116 22820 8172 22822
rect 8196 22820 8252 22822
rect 7956 21786 8012 21788
rect 8036 21786 8092 21788
rect 8116 21786 8172 21788
rect 8196 21786 8252 21788
rect 7956 21734 8002 21786
rect 8002 21734 8012 21786
rect 8036 21734 8066 21786
rect 8066 21734 8078 21786
rect 8078 21734 8092 21786
rect 8116 21734 8130 21786
rect 8130 21734 8142 21786
rect 8142 21734 8172 21786
rect 8196 21734 8206 21786
rect 8206 21734 8252 21786
rect 7956 21732 8012 21734
rect 8036 21732 8092 21734
rect 8116 21732 8172 21734
rect 8196 21732 8252 21734
rect 1306 20340 1308 20360
rect 1308 20340 1360 20360
rect 1360 20340 1362 20360
rect 1306 20304 1362 20340
rect 1306 17992 1362 18048
rect 7956 20698 8012 20700
rect 8036 20698 8092 20700
rect 8116 20698 8172 20700
rect 8196 20698 8252 20700
rect 7956 20646 8002 20698
rect 8002 20646 8012 20698
rect 8036 20646 8066 20698
rect 8066 20646 8078 20698
rect 8078 20646 8092 20698
rect 8116 20646 8130 20698
rect 8130 20646 8142 20698
rect 8142 20646 8172 20698
rect 8196 20646 8206 20698
rect 8206 20646 8252 20698
rect 7956 20644 8012 20646
rect 8036 20644 8092 20646
rect 8116 20644 8172 20646
rect 8196 20644 8252 20646
rect 2956 20154 3012 20156
rect 3036 20154 3092 20156
rect 3116 20154 3172 20156
rect 3196 20154 3252 20156
rect 2956 20102 3002 20154
rect 3002 20102 3012 20154
rect 3036 20102 3066 20154
rect 3066 20102 3078 20154
rect 3078 20102 3092 20154
rect 3116 20102 3130 20154
rect 3130 20102 3142 20154
rect 3142 20102 3172 20154
rect 3196 20102 3206 20154
rect 3206 20102 3252 20154
rect 2956 20100 3012 20102
rect 3036 20100 3092 20102
rect 3116 20100 3172 20102
rect 3196 20100 3252 20102
rect 7956 19610 8012 19612
rect 8036 19610 8092 19612
rect 8116 19610 8172 19612
rect 8196 19610 8252 19612
rect 7956 19558 8002 19610
rect 8002 19558 8012 19610
rect 8036 19558 8066 19610
rect 8066 19558 8078 19610
rect 8078 19558 8092 19610
rect 8116 19558 8130 19610
rect 8130 19558 8142 19610
rect 8142 19558 8172 19610
rect 8196 19558 8206 19610
rect 8206 19558 8252 19610
rect 7956 19556 8012 19558
rect 8036 19556 8092 19558
rect 8116 19556 8172 19558
rect 8196 19556 8252 19558
rect 2956 19066 3012 19068
rect 3036 19066 3092 19068
rect 3116 19066 3172 19068
rect 3196 19066 3252 19068
rect 2956 19014 3002 19066
rect 3002 19014 3012 19066
rect 3036 19014 3066 19066
rect 3066 19014 3078 19066
rect 3078 19014 3092 19066
rect 3116 19014 3130 19066
rect 3130 19014 3142 19066
rect 3142 19014 3172 19066
rect 3196 19014 3206 19066
rect 3206 19014 3252 19066
rect 2956 19012 3012 19014
rect 3036 19012 3092 19014
rect 3116 19012 3172 19014
rect 3196 19012 3252 19014
rect 7956 18522 8012 18524
rect 8036 18522 8092 18524
rect 8116 18522 8172 18524
rect 8196 18522 8252 18524
rect 7956 18470 8002 18522
rect 8002 18470 8012 18522
rect 8036 18470 8066 18522
rect 8066 18470 8078 18522
rect 8078 18470 8092 18522
rect 8116 18470 8130 18522
rect 8130 18470 8142 18522
rect 8142 18470 8172 18522
rect 8196 18470 8206 18522
rect 8206 18470 8252 18522
rect 7956 18468 8012 18470
rect 8036 18468 8092 18470
rect 8116 18468 8172 18470
rect 8196 18468 8252 18470
rect 2956 17978 3012 17980
rect 3036 17978 3092 17980
rect 3116 17978 3172 17980
rect 3196 17978 3252 17980
rect 2956 17926 3002 17978
rect 3002 17926 3012 17978
rect 3036 17926 3066 17978
rect 3066 17926 3078 17978
rect 3078 17926 3092 17978
rect 3116 17926 3130 17978
rect 3130 17926 3142 17978
rect 3142 17926 3172 17978
rect 3196 17926 3206 17978
rect 3206 17926 3252 17978
rect 2956 17924 3012 17926
rect 3036 17924 3092 17926
rect 3116 17924 3172 17926
rect 3196 17924 3252 17926
rect 7956 17434 8012 17436
rect 8036 17434 8092 17436
rect 8116 17434 8172 17436
rect 8196 17434 8252 17436
rect 7956 17382 8002 17434
rect 8002 17382 8012 17434
rect 8036 17382 8066 17434
rect 8066 17382 8078 17434
rect 8078 17382 8092 17434
rect 8116 17382 8130 17434
rect 8130 17382 8142 17434
rect 8142 17382 8172 17434
rect 8196 17382 8206 17434
rect 8206 17382 8252 17434
rect 7956 17380 8012 17382
rect 8036 17380 8092 17382
rect 8116 17380 8172 17382
rect 8196 17380 8252 17382
rect 2956 16890 3012 16892
rect 3036 16890 3092 16892
rect 3116 16890 3172 16892
rect 3196 16890 3252 16892
rect 2956 16838 3002 16890
rect 3002 16838 3012 16890
rect 3036 16838 3066 16890
rect 3066 16838 3078 16890
rect 3078 16838 3092 16890
rect 3116 16838 3130 16890
rect 3130 16838 3142 16890
rect 3142 16838 3172 16890
rect 3196 16838 3206 16890
rect 3206 16838 3252 16890
rect 2956 16836 3012 16838
rect 3036 16836 3092 16838
rect 3116 16836 3172 16838
rect 3196 16836 3252 16838
rect 8942 22616 8998 22672
rect 8942 22072 8998 22128
rect 2956 15802 3012 15804
rect 3036 15802 3092 15804
rect 3116 15802 3172 15804
rect 3196 15802 3252 15804
rect 2956 15750 3002 15802
rect 3002 15750 3012 15802
rect 3036 15750 3066 15802
rect 3066 15750 3078 15802
rect 3078 15750 3092 15802
rect 3116 15750 3130 15802
rect 3130 15750 3142 15802
rect 3142 15750 3172 15802
rect 3196 15750 3206 15802
rect 3206 15750 3252 15802
rect 2956 15748 3012 15750
rect 3036 15748 3092 15750
rect 3116 15748 3172 15750
rect 3196 15748 3252 15750
rect 1306 15680 1362 15736
rect 2956 14714 3012 14716
rect 3036 14714 3092 14716
rect 3116 14714 3172 14716
rect 3196 14714 3252 14716
rect 2956 14662 3002 14714
rect 3002 14662 3012 14714
rect 3036 14662 3066 14714
rect 3066 14662 3078 14714
rect 3078 14662 3092 14714
rect 3116 14662 3130 14714
rect 3130 14662 3142 14714
rect 3142 14662 3172 14714
rect 3196 14662 3206 14714
rect 3206 14662 3252 14714
rect 2956 14660 3012 14662
rect 3036 14660 3092 14662
rect 3116 14660 3172 14662
rect 3196 14660 3252 14662
rect 7956 16346 8012 16348
rect 8036 16346 8092 16348
rect 8116 16346 8172 16348
rect 8196 16346 8252 16348
rect 7956 16294 8002 16346
rect 8002 16294 8012 16346
rect 8036 16294 8066 16346
rect 8066 16294 8078 16346
rect 8078 16294 8092 16346
rect 8116 16294 8130 16346
rect 8130 16294 8142 16346
rect 8142 16294 8172 16346
rect 8196 16294 8206 16346
rect 8206 16294 8252 16346
rect 7956 16292 8012 16294
rect 8036 16292 8092 16294
rect 8116 16292 8172 16294
rect 8196 16292 8252 16294
rect 7956 15258 8012 15260
rect 8036 15258 8092 15260
rect 8116 15258 8172 15260
rect 8196 15258 8252 15260
rect 7956 15206 8002 15258
rect 8002 15206 8012 15258
rect 8036 15206 8066 15258
rect 8066 15206 8078 15258
rect 8078 15206 8092 15258
rect 8116 15206 8130 15258
rect 8130 15206 8142 15258
rect 8142 15206 8172 15258
rect 8196 15206 8206 15258
rect 8206 15206 8252 15258
rect 7956 15204 8012 15206
rect 8036 15204 8092 15206
rect 8116 15204 8172 15206
rect 8196 15204 8252 15206
rect 7956 14170 8012 14172
rect 8036 14170 8092 14172
rect 8116 14170 8172 14172
rect 8196 14170 8252 14172
rect 7956 14118 8002 14170
rect 8002 14118 8012 14170
rect 8036 14118 8066 14170
rect 8066 14118 8078 14170
rect 8078 14118 8092 14170
rect 8116 14118 8130 14170
rect 8130 14118 8142 14170
rect 8142 14118 8172 14170
rect 8196 14118 8206 14170
rect 8206 14118 8252 14170
rect 7956 14116 8012 14118
rect 8036 14116 8092 14118
rect 8116 14116 8172 14118
rect 8196 14116 8252 14118
rect 2956 13626 3012 13628
rect 3036 13626 3092 13628
rect 3116 13626 3172 13628
rect 3196 13626 3252 13628
rect 2956 13574 3002 13626
rect 3002 13574 3012 13626
rect 3036 13574 3066 13626
rect 3066 13574 3078 13626
rect 3078 13574 3092 13626
rect 3116 13574 3130 13626
rect 3130 13574 3142 13626
rect 3142 13574 3172 13626
rect 3196 13574 3206 13626
rect 3206 13574 3252 13626
rect 2956 13572 3012 13574
rect 3036 13572 3092 13574
rect 3116 13572 3172 13574
rect 3196 13572 3252 13574
rect 2778 13368 2834 13424
rect 7956 13082 8012 13084
rect 8036 13082 8092 13084
rect 8116 13082 8172 13084
rect 8196 13082 8252 13084
rect 7956 13030 8002 13082
rect 8002 13030 8012 13082
rect 8036 13030 8066 13082
rect 8066 13030 8078 13082
rect 8078 13030 8092 13082
rect 8116 13030 8130 13082
rect 8130 13030 8142 13082
rect 8142 13030 8172 13082
rect 8196 13030 8206 13082
rect 8206 13030 8252 13082
rect 7956 13028 8012 13030
rect 8036 13028 8092 13030
rect 8116 13028 8172 13030
rect 8196 13028 8252 13030
rect 2956 12538 3012 12540
rect 3036 12538 3092 12540
rect 3116 12538 3172 12540
rect 3196 12538 3252 12540
rect 2956 12486 3002 12538
rect 3002 12486 3012 12538
rect 3036 12486 3066 12538
rect 3066 12486 3078 12538
rect 3078 12486 3092 12538
rect 3116 12486 3130 12538
rect 3130 12486 3142 12538
rect 3142 12486 3172 12538
rect 3196 12486 3206 12538
rect 3206 12486 3252 12538
rect 2956 12484 3012 12486
rect 3036 12484 3092 12486
rect 3116 12484 3172 12486
rect 3196 12484 3252 12486
rect 2956 11450 3012 11452
rect 3036 11450 3092 11452
rect 3116 11450 3172 11452
rect 3196 11450 3252 11452
rect 2956 11398 3002 11450
rect 3002 11398 3012 11450
rect 3036 11398 3066 11450
rect 3066 11398 3078 11450
rect 3078 11398 3092 11450
rect 3116 11398 3130 11450
rect 3130 11398 3142 11450
rect 3142 11398 3172 11450
rect 3196 11398 3206 11450
rect 3206 11398 3252 11450
rect 2956 11396 3012 11398
rect 3036 11396 3092 11398
rect 3116 11396 3172 11398
rect 3196 11396 3252 11398
rect 7956 11994 8012 11996
rect 8036 11994 8092 11996
rect 8116 11994 8172 11996
rect 8196 11994 8252 11996
rect 7956 11942 8002 11994
rect 8002 11942 8012 11994
rect 8036 11942 8066 11994
rect 8066 11942 8078 11994
rect 8078 11942 8092 11994
rect 8116 11942 8130 11994
rect 8130 11942 8142 11994
rect 8142 11942 8172 11994
rect 8196 11942 8206 11994
rect 8206 11942 8252 11994
rect 7956 11940 8012 11942
rect 8036 11940 8092 11942
rect 8116 11940 8172 11942
rect 8196 11940 8252 11942
rect 3330 11056 3386 11112
rect 2956 10362 3012 10364
rect 3036 10362 3092 10364
rect 3116 10362 3172 10364
rect 3196 10362 3252 10364
rect 2956 10310 3002 10362
rect 3002 10310 3012 10362
rect 3036 10310 3066 10362
rect 3066 10310 3078 10362
rect 3078 10310 3092 10362
rect 3116 10310 3130 10362
rect 3130 10310 3142 10362
rect 3142 10310 3172 10362
rect 3196 10310 3206 10362
rect 3206 10310 3252 10362
rect 2956 10308 3012 10310
rect 3036 10308 3092 10310
rect 3116 10308 3172 10310
rect 3196 10308 3252 10310
rect 2956 9274 3012 9276
rect 3036 9274 3092 9276
rect 3116 9274 3172 9276
rect 3196 9274 3252 9276
rect 2956 9222 3002 9274
rect 3002 9222 3012 9274
rect 3036 9222 3066 9274
rect 3066 9222 3078 9274
rect 3078 9222 3092 9274
rect 3116 9222 3130 9274
rect 3130 9222 3142 9274
rect 3142 9222 3172 9274
rect 3196 9222 3206 9274
rect 3206 9222 3252 9274
rect 2956 9220 3012 9222
rect 3036 9220 3092 9222
rect 3116 9220 3172 9222
rect 3196 9220 3252 9222
rect 3330 8744 3386 8800
rect 2956 8186 3012 8188
rect 3036 8186 3092 8188
rect 3116 8186 3172 8188
rect 3196 8186 3252 8188
rect 2956 8134 3002 8186
rect 3002 8134 3012 8186
rect 3036 8134 3066 8186
rect 3066 8134 3078 8186
rect 3078 8134 3092 8186
rect 3116 8134 3130 8186
rect 3130 8134 3142 8186
rect 3142 8134 3172 8186
rect 3196 8134 3206 8186
rect 3206 8134 3252 8186
rect 2956 8132 3012 8134
rect 3036 8132 3092 8134
rect 3116 8132 3172 8134
rect 3196 8132 3252 8134
rect 2956 7098 3012 7100
rect 3036 7098 3092 7100
rect 3116 7098 3172 7100
rect 3196 7098 3252 7100
rect 2956 7046 3002 7098
rect 3002 7046 3012 7098
rect 3036 7046 3066 7098
rect 3066 7046 3078 7098
rect 3078 7046 3092 7098
rect 3116 7046 3130 7098
rect 3130 7046 3142 7098
rect 3142 7046 3172 7098
rect 3196 7046 3206 7098
rect 3206 7046 3252 7098
rect 2956 7044 3012 7046
rect 3036 7044 3092 7046
rect 3116 7044 3172 7046
rect 3196 7044 3252 7046
rect 3422 6432 3478 6488
rect 2956 6010 3012 6012
rect 3036 6010 3092 6012
rect 3116 6010 3172 6012
rect 3196 6010 3252 6012
rect 2956 5958 3002 6010
rect 3002 5958 3012 6010
rect 3036 5958 3066 6010
rect 3066 5958 3078 6010
rect 3078 5958 3092 6010
rect 3116 5958 3130 6010
rect 3130 5958 3142 6010
rect 3142 5958 3172 6010
rect 3196 5958 3206 6010
rect 3206 5958 3252 6010
rect 2956 5956 3012 5958
rect 3036 5956 3092 5958
rect 3116 5956 3172 5958
rect 3196 5956 3252 5958
rect 2956 4922 3012 4924
rect 3036 4922 3092 4924
rect 3116 4922 3172 4924
rect 3196 4922 3252 4924
rect 2956 4870 3002 4922
rect 3002 4870 3012 4922
rect 3036 4870 3066 4922
rect 3066 4870 3078 4922
rect 3078 4870 3092 4922
rect 3116 4870 3130 4922
rect 3130 4870 3142 4922
rect 3142 4870 3172 4922
rect 3196 4870 3206 4922
rect 3206 4870 3252 4922
rect 2956 4868 3012 4870
rect 3036 4868 3092 4870
rect 3116 4868 3172 4870
rect 3196 4868 3252 4870
rect 3422 4120 3478 4176
rect 2956 3834 3012 3836
rect 3036 3834 3092 3836
rect 3116 3834 3172 3836
rect 3196 3834 3252 3836
rect 2956 3782 3002 3834
rect 3002 3782 3012 3834
rect 3036 3782 3066 3834
rect 3066 3782 3078 3834
rect 3078 3782 3092 3834
rect 3116 3782 3130 3834
rect 3130 3782 3142 3834
rect 3142 3782 3172 3834
rect 3196 3782 3206 3834
rect 3206 3782 3252 3834
rect 2956 3780 3012 3782
rect 3036 3780 3092 3782
rect 3116 3780 3172 3782
rect 3196 3780 3252 3782
rect 7956 10906 8012 10908
rect 8036 10906 8092 10908
rect 8116 10906 8172 10908
rect 8196 10906 8252 10908
rect 7956 10854 8002 10906
rect 8002 10854 8012 10906
rect 8036 10854 8066 10906
rect 8066 10854 8078 10906
rect 8078 10854 8092 10906
rect 8116 10854 8130 10906
rect 8130 10854 8142 10906
rect 8142 10854 8172 10906
rect 8196 10854 8206 10906
rect 8206 10854 8252 10906
rect 7956 10852 8012 10854
rect 8036 10852 8092 10854
rect 8116 10852 8172 10854
rect 8196 10852 8252 10854
rect 7956 9818 8012 9820
rect 8036 9818 8092 9820
rect 8116 9818 8172 9820
rect 8196 9818 8252 9820
rect 7956 9766 8002 9818
rect 8002 9766 8012 9818
rect 8036 9766 8066 9818
rect 8066 9766 8078 9818
rect 8078 9766 8092 9818
rect 8116 9766 8130 9818
rect 8130 9766 8142 9818
rect 8142 9766 8172 9818
rect 8196 9766 8206 9818
rect 8206 9766 8252 9818
rect 7956 9764 8012 9766
rect 8036 9764 8092 9766
rect 8116 9764 8172 9766
rect 8196 9764 8252 9766
rect 7956 8730 8012 8732
rect 8036 8730 8092 8732
rect 8116 8730 8172 8732
rect 8196 8730 8252 8732
rect 7956 8678 8002 8730
rect 8002 8678 8012 8730
rect 8036 8678 8066 8730
rect 8066 8678 8078 8730
rect 8078 8678 8092 8730
rect 8116 8678 8130 8730
rect 8130 8678 8142 8730
rect 8142 8678 8172 8730
rect 8196 8678 8206 8730
rect 8206 8678 8252 8730
rect 7956 8676 8012 8678
rect 8036 8676 8092 8678
rect 8116 8676 8172 8678
rect 8196 8676 8252 8678
rect 7956 7642 8012 7644
rect 8036 7642 8092 7644
rect 8116 7642 8172 7644
rect 8196 7642 8252 7644
rect 7956 7590 8002 7642
rect 8002 7590 8012 7642
rect 8036 7590 8066 7642
rect 8066 7590 8078 7642
rect 8078 7590 8092 7642
rect 8116 7590 8130 7642
rect 8130 7590 8142 7642
rect 8142 7590 8172 7642
rect 8196 7590 8206 7642
rect 8206 7590 8252 7642
rect 7956 7588 8012 7590
rect 8036 7588 8092 7590
rect 8116 7588 8172 7590
rect 8196 7588 8252 7590
rect 9402 22072 9458 22128
rect 12956 53882 13012 53884
rect 13036 53882 13092 53884
rect 13116 53882 13172 53884
rect 13196 53882 13252 53884
rect 12956 53830 13002 53882
rect 13002 53830 13012 53882
rect 13036 53830 13066 53882
rect 13066 53830 13078 53882
rect 13078 53830 13092 53882
rect 13116 53830 13130 53882
rect 13130 53830 13142 53882
rect 13142 53830 13172 53882
rect 13196 53830 13206 53882
rect 13206 53830 13252 53882
rect 12956 53828 13012 53830
rect 13036 53828 13092 53830
rect 13116 53828 13172 53830
rect 13196 53828 13252 53830
rect 12956 52794 13012 52796
rect 13036 52794 13092 52796
rect 13116 52794 13172 52796
rect 13196 52794 13252 52796
rect 12956 52742 13002 52794
rect 13002 52742 13012 52794
rect 13036 52742 13066 52794
rect 13066 52742 13078 52794
rect 13078 52742 13092 52794
rect 13116 52742 13130 52794
rect 13130 52742 13142 52794
rect 13142 52742 13172 52794
rect 13196 52742 13206 52794
rect 13206 52742 13252 52794
rect 12956 52740 13012 52742
rect 13036 52740 13092 52742
rect 13116 52740 13172 52742
rect 13196 52740 13252 52742
rect 12956 51706 13012 51708
rect 13036 51706 13092 51708
rect 13116 51706 13172 51708
rect 13196 51706 13252 51708
rect 12956 51654 13002 51706
rect 13002 51654 13012 51706
rect 13036 51654 13066 51706
rect 13066 51654 13078 51706
rect 13078 51654 13092 51706
rect 13116 51654 13130 51706
rect 13130 51654 13142 51706
rect 13142 51654 13172 51706
rect 13196 51654 13206 51706
rect 13206 51654 13252 51706
rect 12956 51652 13012 51654
rect 13036 51652 13092 51654
rect 13116 51652 13172 51654
rect 13196 51652 13252 51654
rect 12956 50618 13012 50620
rect 13036 50618 13092 50620
rect 13116 50618 13172 50620
rect 13196 50618 13252 50620
rect 12956 50566 13002 50618
rect 13002 50566 13012 50618
rect 13036 50566 13066 50618
rect 13066 50566 13078 50618
rect 13078 50566 13092 50618
rect 13116 50566 13130 50618
rect 13130 50566 13142 50618
rect 13142 50566 13172 50618
rect 13196 50566 13206 50618
rect 13206 50566 13252 50618
rect 12956 50564 13012 50566
rect 13036 50564 13092 50566
rect 13116 50564 13172 50566
rect 13196 50564 13252 50566
rect 12956 49530 13012 49532
rect 13036 49530 13092 49532
rect 13116 49530 13172 49532
rect 13196 49530 13252 49532
rect 12956 49478 13002 49530
rect 13002 49478 13012 49530
rect 13036 49478 13066 49530
rect 13066 49478 13078 49530
rect 13078 49478 13092 49530
rect 13116 49478 13130 49530
rect 13130 49478 13142 49530
rect 13142 49478 13172 49530
rect 13196 49478 13206 49530
rect 13206 49478 13252 49530
rect 12956 49476 13012 49478
rect 13036 49476 13092 49478
rect 13116 49476 13172 49478
rect 13196 49476 13252 49478
rect 12956 48442 13012 48444
rect 13036 48442 13092 48444
rect 13116 48442 13172 48444
rect 13196 48442 13252 48444
rect 12956 48390 13002 48442
rect 13002 48390 13012 48442
rect 13036 48390 13066 48442
rect 13066 48390 13078 48442
rect 13078 48390 13092 48442
rect 13116 48390 13130 48442
rect 13130 48390 13142 48442
rect 13142 48390 13172 48442
rect 13196 48390 13206 48442
rect 13206 48390 13252 48442
rect 12956 48388 13012 48390
rect 13036 48388 13092 48390
rect 13116 48388 13172 48390
rect 13196 48388 13252 48390
rect 12956 47354 13012 47356
rect 13036 47354 13092 47356
rect 13116 47354 13172 47356
rect 13196 47354 13252 47356
rect 12956 47302 13002 47354
rect 13002 47302 13012 47354
rect 13036 47302 13066 47354
rect 13066 47302 13078 47354
rect 13078 47302 13092 47354
rect 13116 47302 13130 47354
rect 13130 47302 13142 47354
rect 13142 47302 13172 47354
rect 13196 47302 13206 47354
rect 13206 47302 13252 47354
rect 12956 47300 13012 47302
rect 13036 47300 13092 47302
rect 13116 47300 13172 47302
rect 13196 47300 13252 47302
rect 12956 46266 13012 46268
rect 13036 46266 13092 46268
rect 13116 46266 13172 46268
rect 13196 46266 13252 46268
rect 12956 46214 13002 46266
rect 13002 46214 13012 46266
rect 13036 46214 13066 46266
rect 13066 46214 13078 46266
rect 13078 46214 13092 46266
rect 13116 46214 13130 46266
rect 13130 46214 13142 46266
rect 13142 46214 13172 46266
rect 13196 46214 13206 46266
rect 13206 46214 13252 46266
rect 12956 46212 13012 46214
rect 13036 46212 13092 46214
rect 13116 46212 13172 46214
rect 13196 46212 13252 46214
rect 12956 45178 13012 45180
rect 13036 45178 13092 45180
rect 13116 45178 13172 45180
rect 13196 45178 13252 45180
rect 12956 45126 13002 45178
rect 13002 45126 13012 45178
rect 13036 45126 13066 45178
rect 13066 45126 13078 45178
rect 13078 45126 13092 45178
rect 13116 45126 13130 45178
rect 13130 45126 13142 45178
rect 13142 45126 13172 45178
rect 13196 45126 13206 45178
rect 13206 45126 13252 45178
rect 12956 45124 13012 45126
rect 13036 45124 13092 45126
rect 13116 45124 13172 45126
rect 13196 45124 13252 45126
rect 12956 44090 13012 44092
rect 13036 44090 13092 44092
rect 13116 44090 13172 44092
rect 13196 44090 13252 44092
rect 12956 44038 13002 44090
rect 13002 44038 13012 44090
rect 13036 44038 13066 44090
rect 13066 44038 13078 44090
rect 13078 44038 13092 44090
rect 13116 44038 13130 44090
rect 13130 44038 13142 44090
rect 13142 44038 13172 44090
rect 13196 44038 13206 44090
rect 13206 44038 13252 44090
rect 12956 44036 13012 44038
rect 13036 44036 13092 44038
rect 13116 44036 13172 44038
rect 13196 44036 13252 44038
rect 12956 43002 13012 43004
rect 13036 43002 13092 43004
rect 13116 43002 13172 43004
rect 13196 43002 13252 43004
rect 12956 42950 13002 43002
rect 13002 42950 13012 43002
rect 13036 42950 13066 43002
rect 13066 42950 13078 43002
rect 13078 42950 13092 43002
rect 13116 42950 13130 43002
rect 13130 42950 13142 43002
rect 13142 42950 13172 43002
rect 13196 42950 13206 43002
rect 13206 42950 13252 43002
rect 12956 42948 13012 42950
rect 13036 42948 13092 42950
rect 13116 42948 13172 42950
rect 13196 42948 13252 42950
rect 12956 41914 13012 41916
rect 13036 41914 13092 41916
rect 13116 41914 13172 41916
rect 13196 41914 13252 41916
rect 12956 41862 13002 41914
rect 13002 41862 13012 41914
rect 13036 41862 13066 41914
rect 13066 41862 13078 41914
rect 13078 41862 13092 41914
rect 13116 41862 13130 41914
rect 13130 41862 13142 41914
rect 13142 41862 13172 41914
rect 13196 41862 13206 41914
rect 13206 41862 13252 41914
rect 12956 41860 13012 41862
rect 13036 41860 13092 41862
rect 13116 41860 13172 41862
rect 13196 41860 13252 41862
rect 12956 40826 13012 40828
rect 13036 40826 13092 40828
rect 13116 40826 13172 40828
rect 13196 40826 13252 40828
rect 12956 40774 13002 40826
rect 13002 40774 13012 40826
rect 13036 40774 13066 40826
rect 13066 40774 13078 40826
rect 13078 40774 13092 40826
rect 13116 40774 13130 40826
rect 13130 40774 13142 40826
rect 13142 40774 13172 40826
rect 13196 40774 13206 40826
rect 13206 40774 13252 40826
rect 12956 40772 13012 40774
rect 13036 40772 13092 40774
rect 13116 40772 13172 40774
rect 13196 40772 13252 40774
rect 12956 39738 13012 39740
rect 13036 39738 13092 39740
rect 13116 39738 13172 39740
rect 13196 39738 13252 39740
rect 12956 39686 13002 39738
rect 13002 39686 13012 39738
rect 13036 39686 13066 39738
rect 13066 39686 13078 39738
rect 13078 39686 13092 39738
rect 13116 39686 13130 39738
rect 13130 39686 13142 39738
rect 13142 39686 13172 39738
rect 13196 39686 13206 39738
rect 13206 39686 13252 39738
rect 12956 39684 13012 39686
rect 13036 39684 13092 39686
rect 13116 39684 13172 39686
rect 13196 39684 13252 39686
rect 12956 38650 13012 38652
rect 13036 38650 13092 38652
rect 13116 38650 13172 38652
rect 13196 38650 13252 38652
rect 12956 38598 13002 38650
rect 13002 38598 13012 38650
rect 13036 38598 13066 38650
rect 13066 38598 13078 38650
rect 13078 38598 13092 38650
rect 13116 38598 13130 38650
rect 13130 38598 13142 38650
rect 13142 38598 13172 38650
rect 13196 38598 13206 38650
rect 13206 38598 13252 38650
rect 12956 38596 13012 38598
rect 13036 38596 13092 38598
rect 13116 38596 13172 38598
rect 13196 38596 13252 38598
rect 12956 37562 13012 37564
rect 13036 37562 13092 37564
rect 13116 37562 13172 37564
rect 13196 37562 13252 37564
rect 12956 37510 13002 37562
rect 13002 37510 13012 37562
rect 13036 37510 13066 37562
rect 13066 37510 13078 37562
rect 13078 37510 13092 37562
rect 13116 37510 13130 37562
rect 13130 37510 13142 37562
rect 13142 37510 13172 37562
rect 13196 37510 13206 37562
rect 13206 37510 13252 37562
rect 12956 37508 13012 37510
rect 13036 37508 13092 37510
rect 13116 37508 13172 37510
rect 13196 37508 13252 37510
rect 12956 36474 13012 36476
rect 13036 36474 13092 36476
rect 13116 36474 13172 36476
rect 13196 36474 13252 36476
rect 12956 36422 13002 36474
rect 13002 36422 13012 36474
rect 13036 36422 13066 36474
rect 13066 36422 13078 36474
rect 13078 36422 13092 36474
rect 13116 36422 13130 36474
rect 13130 36422 13142 36474
rect 13142 36422 13172 36474
rect 13196 36422 13206 36474
rect 13206 36422 13252 36474
rect 12956 36420 13012 36422
rect 13036 36420 13092 36422
rect 13116 36420 13172 36422
rect 13196 36420 13252 36422
rect 12956 35386 13012 35388
rect 13036 35386 13092 35388
rect 13116 35386 13172 35388
rect 13196 35386 13252 35388
rect 12956 35334 13002 35386
rect 13002 35334 13012 35386
rect 13036 35334 13066 35386
rect 13066 35334 13078 35386
rect 13078 35334 13092 35386
rect 13116 35334 13130 35386
rect 13130 35334 13142 35386
rect 13142 35334 13172 35386
rect 13196 35334 13206 35386
rect 13206 35334 13252 35386
rect 12956 35332 13012 35334
rect 13036 35332 13092 35334
rect 13116 35332 13172 35334
rect 13196 35332 13252 35334
rect 12956 34298 13012 34300
rect 13036 34298 13092 34300
rect 13116 34298 13172 34300
rect 13196 34298 13252 34300
rect 12956 34246 13002 34298
rect 13002 34246 13012 34298
rect 13036 34246 13066 34298
rect 13066 34246 13078 34298
rect 13078 34246 13092 34298
rect 13116 34246 13130 34298
rect 13130 34246 13142 34298
rect 13142 34246 13172 34298
rect 13196 34246 13206 34298
rect 13206 34246 13252 34298
rect 12956 34244 13012 34246
rect 13036 34244 13092 34246
rect 13116 34244 13172 34246
rect 13196 34244 13252 34246
rect 12956 33210 13012 33212
rect 13036 33210 13092 33212
rect 13116 33210 13172 33212
rect 13196 33210 13252 33212
rect 12956 33158 13002 33210
rect 13002 33158 13012 33210
rect 13036 33158 13066 33210
rect 13066 33158 13078 33210
rect 13078 33158 13092 33210
rect 13116 33158 13130 33210
rect 13130 33158 13142 33210
rect 13142 33158 13172 33210
rect 13196 33158 13206 33210
rect 13206 33158 13252 33210
rect 12956 33156 13012 33158
rect 13036 33156 13092 33158
rect 13116 33156 13172 33158
rect 13196 33156 13252 33158
rect 12956 32122 13012 32124
rect 13036 32122 13092 32124
rect 13116 32122 13172 32124
rect 13196 32122 13252 32124
rect 12956 32070 13002 32122
rect 13002 32070 13012 32122
rect 13036 32070 13066 32122
rect 13066 32070 13078 32122
rect 13078 32070 13092 32122
rect 13116 32070 13130 32122
rect 13130 32070 13142 32122
rect 13142 32070 13172 32122
rect 13196 32070 13206 32122
rect 13206 32070 13252 32122
rect 12956 32068 13012 32070
rect 13036 32068 13092 32070
rect 13116 32068 13172 32070
rect 13196 32068 13252 32070
rect 12956 31034 13012 31036
rect 13036 31034 13092 31036
rect 13116 31034 13172 31036
rect 13196 31034 13252 31036
rect 12956 30982 13002 31034
rect 13002 30982 13012 31034
rect 13036 30982 13066 31034
rect 13066 30982 13078 31034
rect 13078 30982 13092 31034
rect 13116 30982 13130 31034
rect 13130 30982 13142 31034
rect 13142 30982 13172 31034
rect 13196 30982 13206 31034
rect 13206 30982 13252 31034
rect 12956 30980 13012 30982
rect 13036 30980 13092 30982
rect 13116 30980 13172 30982
rect 13196 30980 13252 30982
rect 12956 29946 13012 29948
rect 13036 29946 13092 29948
rect 13116 29946 13172 29948
rect 13196 29946 13252 29948
rect 12956 29894 13002 29946
rect 13002 29894 13012 29946
rect 13036 29894 13066 29946
rect 13066 29894 13078 29946
rect 13078 29894 13092 29946
rect 13116 29894 13130 29946
rect 13130 29894 13142 29946
rect 13142 29894 13172 29946
rect 13196 29894 13206 29946
rect 13206 29894 13252 29946
rect 12956 29892 13012 29894
rect 13036 29892 13092 29894
rect 13116 29892 13172 29894
rect 13196 29892 13252 29894
rect 12956 28858 13012 28860
rect 13036 28858 13092 28860
rect 13116 28858 13172 28860
rect 13196 28858 13252 28860
rect 12956 28806 13002 28858
rect 13002 28806 13012 28858
rect 13036 28806 13066 28858
rect 13066 28806 13078 28858
rect 13078 28806 13092 28858
rect 13116 28806 13130 28858
rect 13130 28806 13142 28858
rect 13142 28806 13172 28858
rect 13196 28806 13206 28858
rect 13206 28806 13252 28858
rect 12956 28804 13012 28806
rect 13036 28804 13092 28806
rect 13116 28804 13172 28806
rect 13196 28804 13252 28806
rect 12956 27770 13012 27772
rect 13036 27770 13092 27772
rect 13116 27770 13172 27772
rect 13196 27770 13252 27772
rect 12956 27718 13002 27770
rect 13002 27718 13012 27770
rect 13036 27718 13066 27770
rect 13066 27718 13078 27770
rect 13078 27718 13092 27770
rect 13116 27718 13130 27770
rect 13130 27718 13142 27770
rect 13142 27718 13172 27770
rect 13196 27718 13206 27770
rect 13206 27718 13252 27770
rect 12956 27716 13012 27718
rect 13036 27716 13092 27718
rect 13116 27716 13172 27718
rect 13196 27716 13252 27718
rect 12956 26682 13012 26684
rect 13036 26682 13092 26684
rect 13116 26682 13172 26684
rect 13196 26682 13252 26684
rect 12956 26630 13002 26682
rect 13002 26630 13012 26682
rect 13036 26630 13066 26682
rect 13066 26630 13078 26682
rect 13078 26630 13092 26682
rect 13116 26630 13130 26682
rect 13130 26630 13142 26682
rect 13142 26630 13172 26682
rect 13196 26630 13206 26682
rect 13206 26630 13252 26682
rect 12956 26628 13012 26630
rect 13036 26628 13092 26630
rect 13116 26628 13172 26630
rect 13196 26628 13252 26630
rect 12956 25594 13012 25596
rect 13036 25594 13092 25596
rect 13116 25594 13172 25596
rect 13196 25594 13252 25596
rect 12956 25542 13002 25594
rect 13002 25542 13012 25594
rect 13036 25542 13066 25594
rect 13066 25542 13078 25594
rect 13078 25542 13092 25594
rect 13116 25542 13130 25594
rect 13130 25542 13142 25594
rect 13142 25542 13172 25594
rect 13196 25542 13206 25594
rect 13206 25542 13252 25594
rect 12956 25540 13012 25542
rect 13036 25540 13092 25542
rect 13116 25540 13172 25542
rect 13196 25540 13252 25542
rect 9586 25200 9642 25256
rect 9586 24928 9642 24984
rect 12956 24506 13012 24508
rect 13036 24506 13092 24508
rect 13116 24506 13172 24508
rect 13196 24506 13252 24508
rect 12956 24454 13002 24506
rect 13002 24454 13012 24506
rect 13036 24454 13066 24506
rect 13066 24454 13078 24506
rect 13078 24454 13092 24506
rect 13116 24454 13130 24506
rect 13130 24454 13142 24506
rect 13142 24454 13172 24506
rect 13196 24454 13206 24506
rect 13206 24454 13252 24506
rect 12956 24452 13012 24454
rect 13036 24452 13092 24454
rect 13116 24452 13172 24454
rect 13196 24452 13252 24454
rect 7956 6554 8012 6556
rect 8036 6554 8092 6556
rect 8116 6554 8172 6556
rect 8196 6554 8252 6556
rect 7956 6502 8002 6554
rect 8002 6502 8012 6554
rect 8036 6502 8066 6554
rect 8066 6502 8078 6554
rect 8078 6502 8092 6554
rect 8116 6502 8130 6554
rect 8130 6502 8142 6554
rect 8142 6502 8172 6554
rect 8196 6502 8206 6554
rect 8206 6502 8252 6554
rect 7956 6500 8012 6502
rect 8036 6500 8092 6502
rect 8116 6500 8172 6502
rect 8196 6500 8252 6502
rect 7956 5466 8012 5468
rect 8036 5466 8092 5468
rect 8116 5466 8172 5468
rect 8196 5466 8252 5468
rect 7956 5414 8002 5466
rect 8002 5414 8012 5466
rect 8036 5414 8066 5466
rect 8066 5414 8078 5466
rect 8078 5414 8092 5466
rect 8116 5414 8130 5466
rect 8130 5414 8142 5466
rect 8142 5414 8172 5466
rect 8196 5414 8206 5466
rect 8206 5414 8252 5466
rect 7956 5412 8012 5414
rect 8036 5412 8092 5414
rect 8116 5412 8172 5414
rect 8196 5412 8252 5414
rect 7956 4378 8012 4380
rect 8036 4378 8092 4380
rect 8116 4378 8172 4380
rect 8196 4378 8252 4380
rect 7956 4326 8002 4378
rect 8002 4326 8012 4378
rect 8036 4326 8066 4378
rect 8066 4326 8078 4378
rect 8078 4326 8092 4378
rect 8116 4326 8130 4378
rect 8130 4326 8142 4378
rect 8142 4326 8172 4378
rect 8196 4326 8206 4378
rect 8206 4326 8252 4378
rect 7956 4324 8012 4326
rect 8036 4324 8092 4326
rect 8116 4324 8172 4326
rect 8196 4324 8252 4326
rect 7956 3290 8012 3292
rect 8036 3290 8092 3292
rect 8116 3290 8172 3292
rect 8196 3290 8252 3292
rect 7956 3238 8002 3290
rect 8002 3238 8012 3290
rect 8036 3238 8066 3290
rect 8066 3238 8078 3290
rect 8078 3238 8092 3290
rect 8116 3238 8130 3290
rect 8130 3238 8142 3290
rect 8142 3238 8172 3290
rect 8196 3238 8206 3290
rect 8206 3238 8252 3290
rect 7956 3236 8012 3238
rect 8036 3236 8092 3238
rect 8116 3236 8172 3238
rect 8196 3236 8252 3238
rect 2956 2746 3012 2748
rect 3036 2746 3092 2748
rect 3116 2746 3172 2748
rect 3196 2746 3252 2748
rect 2956 2694 3002 2746
rect 3002 2694 3012 2746
rect 3036 2694 3066 2746
rect 3066 2694 3078 2746
rect 3078 2694 3092 2746
rect 3116 2694 3130 2746
rect 3130 2694 3142 2746
rect 3142 2694 3172 2746
rect 3196 2694 3206 2746
rect 3206 2694 3252 2746
rect 2956 2692 3012 2694
rect 3036 2692 3092 2694
rect 3116 2692 3172 2694
rect 3196 2692 3252 2694
rect 2778 1808 2834 1864
rect 4986 2372 5042 2408
rect 4986 2352 4988 2372
rect 4988 2352 5040 2372
rect 5040 2352 5042 2372
rect 5722 2896 5778 2952
rect 9494 2508 9550 2544
rect 9494 2488 9496 2508
rect 9496 2488 9548 2508
rect 9548 2488 9550 2508
rect 7956 2202 8012 2204
rect 8036 2202 8092 2204
rect 8116 2202 8172 2204
rect 8196 2202 8252 2204
rect 7956 2150 8002 2202
rect 8002 2150 8012 2202
rect 8036 2150 8066 2202
rect 8066 2150 8078 2202
rect 8078 2150 8092 2202
rect 8116 2150 8130 2202
rect 8130 2150 8142 2202
rect 8142 2150 8172 2202
rect 8196 2150 8206 2202
rect 8206 2150 8252 2202
rect 7956 2148 8012 2150
rect 8036 2148 8092 2150
rect 8116 2148 8172 2150
rect 8196 2148 8252 2150
rect 12956 23418 13012 23420
rect 13036 23418 13092 23420
rect 13116 23418 13172 23420
rect 13196 23418 13252 23420
rect 12956 23366 13002 23418
rect 13002 23366 13012 23418
rect 13036 23366 13066 23418
rect 13066 23366 13078 23418
rect 13078 23366 13092 23418
rect 13116 23366 13130 23418
rect 13130 23366 13142 23418
rect 13142 23366 13172 23418
rect 13196 23366 13206 23418
rect 13206 23366 13252 23418
rect 12956 23364 13012 23366
rect 13036 23364 13092 23366
rect 13116 23364 13172 23366
rect 13196 23364 13252 23366
rect 12956 22330 13012 22332
rect 13036 22330 13092 22332
rect 13116 22330 13172 22332
rect 13196 22330 13252 22332
rect 12956 22278 13002 22330
rect 13002 22278 13012 22330
rect 13036 22278 13066 22330
rect 13066 22278 13078 22330
rect 13078 22278 13092 22330
rect 13116 22278 13130 22330
rect 13130 22278 13142 22330
rect 13142 22278 13172 22330
rect 13196 22278 13206 22330
rect 13206 22278 13252 22330
rect 12956 22276 13012 22278
rect 13036 22276 13092 22278
rect 13116 22276 13172 22278
rect 13196 22276 13252 22278
rect 12956 21242 13012 21244
rect 13036 21242 13092 21244
rect 13116 21242 13172 21244
rect 13196 21242 13252 21244
rect 12956 21190 13002 21242
rect 13002 21190 13012 21242
rect 13036 21190 13066 21242
rect 13066 21190 13078 21242
rect 13078 21190 13092 21242
rect 13116 21190 13130 21242
rect 13130 21190 13142 21242
rect 13142 21190 13172 21242
rect 13196 21190 13206 21242
rect 13206 21190 13252 21242
rect 12956 21188 13012 21190
rect 13036 21188 13092 21190
rect 13116 21188 13172 21190
rect 13196 21188 13252 21190
rect 12956 20154 13012 20156
rect 13036 20154 13092 20156
rect 13116 20154 13172 20156
rect 13196 20154 13252 20156
rect 12956 20102 13002 20154
rect 13002 20102 13012 20154
rect 13036 20102 13066 20154
rect 13066 20102 13078 20154
rect 13078 20102 13092 20154
rect 13116 20102 13130 20154
rect 13130 20102 13142 20154
rect 13142 20102 13172 20154
rect 13196 20102 13206 20154
rect 13206 20102 13252 20154
rect 12956 20100 13012 20102
rect 13036 20100 13092 20102
rect 13116 20100 13172 20102
rect 13196 20100 13252 20102
rect 12956 19066 13012 19068
rect 13036 19066 13092 19068
rect 13116 19066 13172 19068
rect 13196 19066 13252 19068
rect 12956 19014 13002 19066
rect 13002 19014 13012 19066
rect 13036 19014 13066 19066
rect 13066 19014 13078 19066
rect 13078 19014 13092 19066
rect 13116 19014 13130 19066
rect 13130 19014 13142 19066
rect 13142 19014 13172 19066
rect 13196 19014 13206 19066
rect 13206 19014 13252 19066
rect 12956 19012 13012 19014
rect 13036 19012 13092 19014
rect 13116 19012 13172 19014
rect 13196 19012 13252 19014
rect 12956 17978 13012 17980
rect 13036 17978 13092 17980
rect 13116 17978 13172 17980
rect 13196 17978 13252 17980
rect 12956 17926 13002 17978
rect 13002 17926 13012 17978
rect 13036 17926 13066 17978
rect 13066 17926 13078 17978
rect 13078 17926 13092 17978
rect 13116 17926 13130 17978
rect 13130 17926 13142 17978
rect 13142 17926 13172 17978
rect 13196 17926 13206 17978
rect 13206 17926 13252 17978
rect 12956 17924 13012 17926
rect 13036 17924 13092 17926
rect 13116 17924 13172 17926
rect 13196 17924 13252 17926
rect 12956 16890 13012 16892
rect 13036 16890 13092 16892
rect 13116 16890 13172 16892
rect 13196 16890 13252 16892
rect 12956 16838 13002 16890
rect 13002 16838 13012 16890
rect 13036 16838 13066 16890
rect 13066 16838 13078 16890
rect 13078 16838 13092 16890
rect 13116 16838 13130 16890
rect 13130 16838 13142 16890
rect 13142 16838 13172 16890
rect 13196 16838 13206 16890
rect 13206 16838 13252 16890
rect 12956 16836 13012 16838
rect 13036 16836 13092 16838
rect 13116 16836 13172 16838
rect 13196 16836 13252 16838
rect 12956 15802 13012 15804
rect 13036 15802 13092 15804
rect 13116 15802 13172 15804
rect 13196 15802 13252 15804
rect 12956 15750 13002 15802
rect 13002 15750 13012 15802
rect 13036 15750 13066 15802
rect 13066 15750 13078 15802
rect 13078 15750 13092 15802
rect 13116 15750 13130 15802
rect 13130 15750 13142 15802
rect 13142 15750 13172 15802
rect 13196 15750 13206 15802
rect 13206 15750 13252 15802
rect 12956 15748 13012 15750
rect 13036 15748 13092 15750
rect 13116 15748 13172 15750
rect 13196 15748 13252 15750
rect 12956 14714 13012 14716
rect 13036 14714 13092 14716
rect 13116 14714 13172 14716
rect 13196 14714 13252 14716
rect 12956 14662 13002 14714
rect 13002 14662 13012 14714
rect 13036 14662 13066 14714
rect 13066 14662 13078 14714
rect 13078 14662 13092 14714
rect 13116 14662 13130 14714
rect 13130 14662 13142 14714
rect 13142 14662 13172 14714
rect 13196 14662 13206 14714
rect 13206 14662 13252 14714
rect 12956 14660 13012 14662
rect 13036 14660 13092 14662
rect 13116 14660 13172 14662
rect 13196 14660 13252 14662
rect 12956 13626 13012 13628
rect 13036 13626 13092 13628
rect 13116 13626 13172 13628
rect 13196 13626 13252 13628
rect 12956 13574 13002 13626
rect 13002 13574 13012 13626
rect 13036 13574 13066 13626
rect 13066 13574 13078 13626
rect 13078 13574 13092 13626
rect 13116 13574 13130 13626
rect 13130 13574 13142 13626
rect 13142 13574 13172 13626
rect 13196 13574 13206 13626
rect 13206 13574 13252 13626
rect 12956 13572 13012 13574
rect 13036 13572 13092 13574
rect 13116 13572 13172 13574
rect 13196 13572 13252 13574
rect 12956 12538 13012 12540
rect 13036 12538 13092 12540
rect 13116 12538 13172 12540
rect 13196 12538 13252 12540
rect 12956 12486 13002 12538
rect 13002 12486 13012 12538
rect 13036 12486 13066 12538
rect 13066 12486 13078 12538
rect 13078 12486 13092 12538
rect 13116 12486 13130 12538
rect 13130 12486 13142 12538
rect 13142 12486 13172 12538
rect 13196 12486 13206 12538
rect 13206 12486 13252 12538
rect 12956 12484 13012 12486
rect 13036 12484 13092 12486
rect 13116 12484 13172 12486
rect 13196 12484 13252 12486
rect 12956 11450 13012 11452
rect 13036 11450 13092 11452
rect 13116 11450 13172 11452
rect 13196 11450 13252 11452
rect 12956 11398 13002 11450
rect 13002 11398 13012 11450
rect 13036 11398 13066 11450
rect 13066 11398 13078 11450
rect 13078 11398 13092 11450
rect 13116 11398 13130 11450
rect 13130 11398 13142 11450
rect 13142 11398 13172 11450
rect 13196 11398 13206 11450
rect 13206 11398 13252 11450
rect 12956 11396 13012 11398
rect 13036 11396 13092 11398
rect 13116 11396 13172 11398
rect 13196 11396 13252 11398
rect 12956 10362 13012 10364
rect 13036 10362 13092 10364
rect 13116 10362 13172 10364
rect 13196 10362 13252 10364
rect 12956 10310 13002 10362
rect 13002 10310 13012 10362
rect 13036 10310 13066 10362
rect 13066 10310 13078 10362
rect 13078 10310 13092 10362
rect 13116 10310 13130 10362
rect 13130 10310 13142 10362
rect 13142 10310 13172 10362
rect 13196 10310 13206 10362
rect 13206 10310 13252 10362
rect 12956 10308 13012 10310
rect 13036 10308 13092 10310
rect 13116 10308 13172 10310
rect 13196 10308 13252 10310
rect 12956 9274 13012 9276
rect 13036 9274 13092 9276
rect 13116 9274 13172 9276
rect 13196 9274 13252 9276
rect 12956 9222 13002 9274
rect 13002 9222 13012 9274
rect 13036 9222 13066 9274
rect 13066 9222 13078 9274
rect 13078 9222 13092 9274
rect 13116 9222 13130 9274
rect 13130 9222 13142 9274
rect 13142 9222 13172 9274
rect 13196 9222 13206 9274
rect 13206 9222 13252 9274
rect 12956 9220 13012 9222
rect 13036 9220 13092 9222
rect 13116 9220 13172 9222
rect 13196 9220 13252 9222
rect 12956 8186 13012 8188
rect 13036 8186 13092 8188
rect 13116 8186 13172 8188
rect 13196 8186 13252 8188
rect 12956 8134 13002 8186
rect 13002 8134 13012 8186
rect 13036 8134 13066 8186
rect 13066 8134 13078 8186
rect 13078 8134 13092 8186
rect 13116 8134 13130 8186
rect 13130 8134 13142 8186
rect 13142 8134 13172 8186
rect 13196 8134 13206 8186
rect 13206 8134 13252 8186
rect 12956 8132 13012 8134
rect 13036 8132 13092 8134
rect 13116 8132 13172 8134
rect 13196 8132 13252 8134
rect 12956 7098 13012 7100
rect 13036 7098 13092 7100
rect 13116 7098 13172 7100
rect 13196 7098 13252 7100
rect 12956 7046 13002 7098
rect 13002 7046 13012 7098
rect 13036 7046 13066 7098
rect 13066 7046 13078 7098
rect 13078 7046 13092 7098
rect 13116 7046 13130 7098
rect 13130 7046 13142 7098
rect 13142 7046 13172 7098
rect 13196 7046 13206 7098
rect 13206 7046 13252 7098
rect 12956 7044 13012 7046
rect 13036 7044 13092 7046
rect 13116 7044 13172 7046
rect 13196 7044 13252 7046
rect 12956 6010 13012 6012
rect 13036 6010 13092 6012
rect 13116 6010 13172 6012
rect 13196 6010 13252 6012
rect 12956 5958 13002 6010
rect 13002 5958 13012 6010
rect 13036 5958 13066 6010
rect 13066 5958 13078 6010
rect 13078 5958 13092 6010
rect 13116 5958 13130 6010
rect 13130 5958 13142 6010
rect 13142 5958 13172 6010
rect 13196 5958 13206 6010
rect 13206 5958 13252 6010
rect 12956 5956 13012 5958
rect 13036 5956 13092 5958
rect 13116 5956 13172 5958
rect 13196 5956 13252 5958
rect 12956 4922 13012 4924
rect 13036 4922 13092 4924
rect 13116 4922 13172 4924
rect 13196 4922 13252 4924
rect 12956 4870 13002 4922
rect 13002 4870 13012 4922
rect 13036 4870 13066 4922
rect 13066 4870 13078 4922
rect 13078 4870 13092 4922
rect 13116 4870 13130 4922
rect 13130 4870 13142 4922
rect 13142 4870 13172 4922
rect 13196 4870 13206 4922
rect 13206 4870 13252 4922
rect 12956 4868 13012 4870
rect 13036 4868 13092 4870
rect 13116 4868 13172 4870
rect 13196 4868 13252 4870
rect 12956 3834 13012 3836
rect 13036 3834 13092 3836
rect 13116 3834 13172 3836
rect 13196 3834 13252 3836
rect 12956 3782 13002 3834
rect 13002 3782 13012 3834
rect 13036 3782 13066 3834
rect 13066 3782 13078 3834
rect 13078 3782 13092 3834
rect 13116 3782 13130 3834
rect 13130 3782 13142 3834
rect 13142 3782 13172 3834
rect 13196 3782 13206 3834
rect 13206 3782 13252 3834
rect 12956 3780 13012 3782
rect 13036 3780 13092 3782
rect 13116 3780 13172 3782
rect 13196 3780 13252 3782
rect 17956 54426 18012 54428
rect 18036 54426 18092 54428
rect 18116 54426 18172 54428
rect 18196 54426 18252 54428
rect 17956 54374 18002 54426
rect 18002 54374 18012 54426
rect 18036 54374 18066 54426
rect 18066 54374 18078 54426
rect 18078 54374 18092 54426
rect 18116 54374 18130 54426
rect 18130 54374 18142 54426
rect 18142 54374 18172 54426
rect 18196 54374 18206 54426
rect 18206 54374 18252 54426
rect 17956 54372 18012 54374
rect 18036 54372 18092 54374
rect 18116 54372 18172 54374
rect 18196 54372 18252 54374
rect 17956 53338 18012 53340
rect 18036 53338 18092 53340
rect 18116 53338 18172 53340
rect 18196 53338 18252 53340
rect 17956 53286 18002 53338
rect 18002 53286 18012 53338
rect 18036 53286 18066 53338
rect 18066 53286 18078 53338
rect 18078 53286 18092 53338
rect 18116 53286 18130 53338
rect 18130 53286 18142 53338
rect 18142 53286 18172 53338
rect 18196 53286 18206 53338
rect 18206 53286 18252 53338
rect 17956 53284 18012 53286
rect 18036 53284 18092 53286
rect 18116 53284 18172 53286
rect 18196 53284 18252 53286
rect 17956 52250 18012 52252
rect 18036 52250 18092 52252
rect 18116 52250 18172 52252
rect 18196 52250 18252 52252
rect 17956 52198 18002 52250
rect 18002 52198 18012 52250
rect 18036 52198 18066 52250
rect 18066 52198 18078 52250
rect 18078 52198 18092 52250
rect 18116 52198 18130 52250
rect 18130 52198 18142 52250
rect 18142 52198 18172 52250
rect 18196 52198 18206 52250
rect 18206 52198 18252 52250
rect 17956 52196 18012 52198
rect 18036 52196 18092 52198
rect 18116 52196 18172 52198
rect 18196 52196 18252 52198
rect 17956 51162 18012 51164
rect 18036 51162 18092 51164
rect 18116 51162 18172 51164
rect 18196 51162 18252 51164
rect 17956 51110 18002 51162
rect 18002 51110 18012 51162
rect 18036 51110 18066 51162
rect 18066 51110 18078 51162
rect 18078 51110 18092 51162
rect 18116 51110 18130 51162
rect 18130 51110 18142 51162
rect 18142 51110 18172 51162
rect 18196 51110 18206 51162
rect 18206 51110 18252 51162
rect 17956 51108 18012 51110
rect 18036 51108 18092 51110
rect 18116 51108 18172 51110
rect 18196 51108 18252 51110
rect 17956 50074 18012 50076
rect 18036 50074 18092 50076
rect 18116 50074 18172 50076
rect 18196 50074 18252 50076
rect 17956 50022 18002 50074
rect 18002 50022 18012 50074
rect 18036 50022 18066 50074
rect 18066 50022 18078 50074
rect 18078 50022 18092 50074
rect 18116 50022 18130 50074
rect 18130 50022 18142 50074
rect 18142 50022 18172 50074
rect 18196 50022 18206 50074
rect 18206 50022 18252 50074
rect 17956 50020 18012 50022
rect 18036 50020 18092 50022
rect 18116 50020 18172 50022
rect 18196 50020 18252 50022
rect 17956 48986 18012 48988
rect 18036 48986 18092 48988
rect 18116 48986 18172 48988
rect 18196 48986 18252 48988
rect 17956 48934 18002 48986
rect 18002 48934 18012 48986
rect 18036 48934 18066 48986
rect 18066 48934 18078 48986
rect 18078 48934 18092 48986
rect 18116 48934 18130 48986
rect 18130 48934 18142 48986
rect 18142 48934 18172 48986
rect 18196 48934 18206 48986
rect 18206 48934 18252 48986
rect 17956 48932 18012 48934
rect 18036 48932 18092 48934
rect 18116 48932 18172 48934
rect 18196 48932 18252 48934
rect 17956 47898 18012 47900
rect 18036 47898 18092 47900
rect 18116 47898 18172 47900
rect 18196 47898 18252 47900
rect 17956 47846 18002 47898
rect 18002 47846 18012 47898
rect 18036 47846 18066 47898
rect 18066 47846 18078 47898
rect 18078 47846 18092 47898
rect 18116 47846 18130 47898
rect 18130 47846 18142 47898
rect 18142 47846 18172 47898
rect 18196 47846 18206 47898
rect 18206 47846 18252 47898
rect 17956 47844 18012 47846
rect 18036 47844 18092 47846
rect 18116 47844 18172 47846
rect 18196 47844 18252 47846
rect 17956 46810 18012 46812
rect 18036 46810 18092 46812
rect 18116 46810 18172 46812
rect 18196 46810 18252 46812
rect 17956 46758 18002 46810
rect 18002 46758 18012 46810
rect 18036 46758 18066 46810
rect 18066 46758 18078 46810
rect 18078 46758 18092 46810
rect 18116 46758 18130 46810
rect 18130 46758 18142 46810
rect 18142 46758 18172 46810
rect 18196 46758 18206 46810
rect 18206 46758 18252 46810
rect 17956 46756 18012 46758
rect 18036 46756 18092 46758
rect 18116 46756 18172 46758
rect 18196 46756 18252 46758
rect 17956 45722 18012 45724
rect 18036 45722 18092 45724
rect 18116 45722 18172 45724
rect 18196 45722 18252 45724
rect 17956 45670 18002 45722
rect 18002 45670 18012 45722
rect 18036 45670 18066 45722
rect 18066 45670 18078 45722
rect 18078 45670 18092 45722
rect 18116 45670 18130 45722
rect 18130 45670 18142 45722
rect 18142 45670 18172 45722
rect 18196 45670 18206 45722
rect 18206 45670 18252 45722
rect 17956 45668 18012 45670
rect 18036 45668 18092 45670
rect 18116 45668 18172 45670
rect 18196 45668 18252 45670
rect 17956 44634 18012 44636
rect 18036 44634 18092 44636
rect 18116 44634 18172 44636
rect 18196 44634 18252 44636
rect 17956 44582 18002 44634
rect 18002 44582 18012 44634
rect 18036 44582 18066 44634
rect 18066 44582 18078 44634
rect 18078 44582 18092 44634
rect 18116 44582 18130 44634
rect 18130 44582 18142 44634
rect 18142 44582 18172 44634
rect 18196 44582 18206 44634
rect 18206 44582 18252 44634
rect 17956 44580 18012 44582
rect 18036 44580 18092 44582
rect 18116 44580 18172 44582
rect 18196 44580 18252 44582
rect 17956 43546 18012 43548
rect 18036 43546 18092 43548
rect 18116 43546 18172 43548
rect 18196 43546 18252 43548
rect 17956 43494 18002 43546
rect 18002 43494 18012 43546
rect 18036 43494 18066 43546
rect 18066 43494 18078 43546
rect 18078 43494 18092 43546
rect 18116 43494 18130 43546
rect 18130 43494 18142 43546
rect 18142 43494 18172 43546
rect 18196 43494 18206 43546
rect 18206 43494 18252 43546
rect 17956 43492 18012 43494
rect 18036 43492 18092 43494
rect 18116 43492 18172 43494
rect 18196 43492 18252 43494
rect 17956 42458 18012 42460
rect 18036 42458 18092 42460
rect 18116 42458 18172 42460
rect 18196 42458 18252 42460
rect 17956 42406 18002 42458
rect 18002 42406 18012 42458
rect 18036 42406 18066 42458
rect 18066 42406 18078 42458
rect 18078 42406 18092 42458
rect 18116 42406 18130 42458
rect 18130 42406 18142 42458
rect 18142 42406 18172 42458
rect 18196 42406 18206 42458
rect 18206 42406 18252 42458
rect 17956 42404 18012 42406
rect 18036 42404 18092 42406
rect 18116 42404 18172 42406
rect 18196 42404 18252 42406
rect 17956 41370 18012 41372
rect 18036 41370 18092 41372
rect 18116 41370 18172 41372
rect 18196 41370 18252 41372
rect 17956 41318 18002 41370
rect 18002 41318 18012 41370
rect 18036 41318 18066 41370
rect 18066 41318 18078 41370
rect 18078 41318 18092 41370
rect 18116 41318 18130 41370
rect 18130 41318 18142 41370
rect 18142 41318 18172 41370
rect 18196 41318 18206 41370
rect 18206 41318 18252 41370
rect 17956 41316 18012 41318
rect 18036 41316 18092 41318
rect 18116 41316 18172 41318
rect 18196 41316 18252 41318
rect 17956 40282 18012 40284
rect 18036 40282 18092 40284
rect 18116 40282 18172 40284
rect 18196 40282 18252 40284
rect 17956 40230 18002 40282
rect 18002 40230 18012 40282
rect 18036 40230 18066 40282
rect 18066 40230 18078 40282
rect 18078 40230 18092 40282
rect 18116 40230 18130 40282
rect 18130 40230 18142 40282
rect 18142 40230 18172 40282
rect 18196 40230 18206 40282
rect 18206 40230 18252 40282
rect 17956 40228 18012 40230
rect 18036 40228 18092 40230
rect 18116 40228 18172 40230
rect 18196 40228 18252 40230
rect 17956 39194 18012 39196
rect 18036 39194 18092 39196
rect 18116 39194 18172 39196
rect 18196 39194 18252 39196
rect 17956 39142 18002 39194
rect 18002 39142 18012 39194
rect 18036 39142 18066 39194
rect 18066 39142 18078 39194
rect 18078 39142 18092 39194
rect 18116 39142 18130 39194
rect 18130 39142 18142 39194
rect 18142 39142 18172 39194
rect 18196 39142 18206 39194
rect 18206 39142 18252 39194
rect 17956 39140 18012 39142
rect 18036 39140 18092 39142
rect 18116 39140 18172 39142
rect 18196 39140 18252 39142
rect 17956 38106 18012 38108
rect 18036 38106 18092 38108
rect 18116 38106 18172 38108
rect 18196 38106 18252 38108
rect 17956 38054 18002 38106
rect 18002 38054 18012 38106
rect 18036 38054 18066 38106
rect 18066 38054 18078 38106
rect 18078 38054 18092 38106
rect 18116 38054 18130 38106
rect 18130 38054 18142 38106
rect 18142 38054 18172 38106
rect 18196 38054 18206 38106
rect 18206 38054 18252 38106
rect 17956 38052 18012 38054
rect 18036 38052 18092 38054
rect 18116 38052 18172 38054
rect 18196 38052 18252 38054
rect 17956 37018 18012 37020
rect 18036 37018 18092 37020
rect 18116 37018 18172 37020
rect 18196 37018 18252 37020
rect 17956 36966 18002 37018
rect 18002 36966 18012 37018
rect 18036 36966 18066 37018
rect 18066 36966 18078 37018
rect 18078 36966 18092 37018
rect 18116 36966 18130 37018
rect 18130 36966 18142 37018
rect 18142 36966 18172 37018
rect 18196 36966 18206 37018
rect 18206 36966 18252 37018
rect 17956 36964 18012 36966
rect 18036 36964 18092 36966
rect 18116 36964 18172 36966
rect 18196 36964 18252 36966
rect 17956 35930 18012 35932
rect 18036 35930 18092 35932
rect 18116 35930 18172 35932
rect 18196 35930 18252 35932
rect 17956 35878 18002 35930
rect 18002 35878 18012 35930
rect 18036 35878 18066 35930
rect 18066 35878 18078 35930
rect 18078 35878 18092 35930
rect 18116 35878 18130 35930
rect 18130 35878 18142 35930
rect 18142 35878 18172 35930
rect 18196 35878 18206 35930
rect 18206 35878 18252 35930
rect 17956 35876 18012 35878
rect 18036 35876 18092 35878
rect 18116 35876 18172 35878
rect 18196 35876 18252 35878
rect 17956 34842 18012 34844
rect 18036 34842 18092 34844
rect 18116 34842 18172 34844
rect 18196 34842 18252 34844
rect 17956 34790 18002 34842
rect 18002 34790 18012 34842
rect 18036 34790 18066 34842
rect 18066 34790 18078 34842
rect 18078 34790 18092 34842
rect 18116 34790 18130 34842
rect 18130 34790 18142 34842
rect 18142 34790 18172 34842
rect 18196 34790 18206 34842
rect 18206 34790 18252 34842
rect 17956 34788 18012 34790
rect 18036 34788 18092 34790
rect 18116 34788 18172 34790
rect 18196 34788 18252 34790
rect 17956 33754 18012 33756
rect 18036 33754 18092 33756
rect 18116 33754 18172 33756
rect 18196 33754 18252 33756
rect 17956 33702 18002 33754
rect 18002 33702 18012 33754
rect 18036 33702 18066 33754
rect 18066 33702 18078 33754
rect 18078 33702 18092 33754
rect 18116 33702 18130 33754
rect 18130 33702 18142 33754
rect 18142 33702 18172 33754
rect 18196 33702 18206 33754
rect 18206 33702 18252 33754
rect 17956 33700 18012 33702
rect 18036 33700 18092 33702
rect 18116 33700 18172 33702
rect 18196 33700 18252 33702
rect 17956 32666 18012 32668
rect 18036 32666 18092 32668
rect 18116 32666 18172 32668
rect 18196 32666 18252 32668
rect 17956 32614 18002 32666
rect 18002 32614 18012 32666
rect 18036 32614 18066 32666
rect 18066 32614 18078 32666
rect 18078 32614 18092 32666
rect 18116 32614 18130 32666
rect 18130 32614 18142 32666
rect 18142 32614 18172 32666
rect 18196 32614 18206 32666
rect 18206 32614 18252 32666
rect 17956 32612 18012 32614
rect 18036 32612 18092 32614
rect 18116 32612 18172 32614
rect 18196 32612 18252 32614
rect 17956 31578 18012 31580
rect 18036 31578 18092 31580
rect 18116 31578 18172 31580
rect 18196 31578 18252 31580
rect 17956 31526 18002 31578
rect 18002 31526 18012 31578
rect 18036 31526 18066 31578
rect 18066 31526 18078 31578
rect 18078 31526 18092 31578
rect 18116 31526 18130 31578
rect 18130 31526 18142 31578
rect 18142 31526 18172 31578
rect 18196 31526 18206 31578
rect 18206 31526 18252 31578
rect 17956 31524 18012 31526
rect 18036 31524 18092 31526
rect 18116 31524 18172 31526
rect 18196 31524 18252 31526
rect 17956 30490 18012 30492
rect 18036 30490 18092 30492
rect 18116 30490 18172 30492
rect 18196 30490 18252 30492
rect 17956 30438 18002 30490
rect 18002 30438 18012 30490
rect 18036 30438 18066 30490
rect 18066 30438 18078 30490
rect 18078 30438 18092 30490
rect 18116 30438 18130 30490
rect 18130 30438 18142 30490
rect 18142 30438 18172 30490
rect 18196 30438 18206 30490
rect 18206 30438 18252 30490
rect 17956 30436 18012 30438
rect 18036 30436 18092 30438
rect 18116 30436 18172 30438
rect 18196 30436 18252 30438
rect 17956 29402 18012 29404
rect 18036 29402 18092 29404
rect 18116 29402 18172 29404
rect 18196 29402 18252 29404
rect 17956 29350 18002 29402
rect 18002 29350 18012 29402
rect 18036 29350 18066 29402
rect 18066 29350 18078 29402
rect 18078 29350 18092 29402
rect 18116 29350 18130 29402
rect 18130 29350 18142 29402
rect 18142 29350 18172 29402
rect 18196 29350 18206 29402
rect 18206 29350 18252 29402
rect 17956 29348 18012 29350
rect 18036 29348 18092 29350
rect 18116 29348 18172 29350
rect 18196 29348 18252 29350
rect 12956 2746 13012 2748
rect 13036 2746 13092 2748
rect 13116 2746 13172 2748
rect 13196 2746 13252 2748
rect 12956 2694 13002 2746
rect 13002 2694 13012 2746
rect 13036 2694 13066 2746
rect 13066 2694 13078 2746
rect 13078 2694 13092 2746
rect 13116 2694 13130 2746
rect 13130 2694 13142 2746
rect 13142 2694 13172 2746
rect 13196 2694 13206 2746
rect 13206 2694 13252 2746
rect 12956 2692 13012 2694
rect 13036 2692 13092 2694
rect 13116 2692 13172 2694
rect 13196 2692 13252 2694
rect 13634 2644 13690 2680
rect 13634 2624 13636 2644
rect 13636 2624 13688 2644
rect 13688 2624 13690 2644
rect 17956 28314 18012 28316
rect 18036 28314 18092 28316
rect 18116 28314 18172 28316
rect 18196 28314 18252 28316
rect 17956 28262 18002 28314
rect 18002 28262 18012 28314
rect 18036 28262 18066 28314
rect 18066 28262 18078 28314
rect 18078 28262 18092 28314
rect 18116 28262 18130 28314
rect 18130 28262 18142 28314
rect 18142 28262 18172 28314
rect 18196 28262 18206 28314
rect 18206 28262 18252 28314
rect 17956 28260 18012 28262
rect 18036 28260 18092 28262
rect 18116 28260 18172 28262
rect 18196 28260 18252 28262
rect 17956 27226 18012 27228
rect 18036 27226 18092 27228
rect 18116 27226 18172 27228
rect 18196 27226 18252 27228
rect 17956 27174 18002 27226
rect 18002 27174 18012 27226
rect 18036 27174 18066 27226
rect 18066 27174 18078 27226
rect 18078 27174 18092 27226
rect 18116 27174 18130 27226
rect 18130 27174 18142 27226
rect 18142 27174 18172 27226
rect 18196 27174 18206 27226
rect 18206 27174 18252 27226
rect 17956 27172 18012 27174
rect 18036 27172 18092 27174
rect 18116 27172 18172 27174
rect 18196 27172 18252 27174
rect 17956 26138 18012 26140
rect 18036 26138 18092 26140
rect 18116 26138 18172 26140
rect 18196 26138 18252 26140
rect 17956 26086 18002 26138
rect 18002 26086 18012 26138
rect 18036 26086 18066 26138
rect 18066 26086 18078 26138
rect 18078 26086 18092 26138
rect 18116 26086 18130 26138
rect 18130 26086 18142 26138
rect 18142 26086 18172 26138
rect 18196 26086 18206 26138
rect 18206 26086 18252 26138
rect 17956 26084 18012 26086
rect 18036 26084 18092 26086
rect 18116 26084 18172 26086
rect 18196 26084 18252 26086
rect 17956 25050 18012 25052
rect 18036 25050 18092 25052
rect 18116 25050 18172 25052
rect 18196 25050 18252 25052
rect 17956 24998 18002 25050
rect 18002 24998 18012 25050
rect 18036 24998 18066 25050
rect 18066 24998 18078 25050
rect 18078 24998 18092 25050
rect 18116 24998 18130 25050
rect 18130 24998 18142 25050
rect 18142 24998 18172 25050
rect 18196 24998 18206 25050
rect 18206 24998 18252 25050
rect 17956 24996 18012 24998
rect 18036 24996 18092 24998
rect 18116 24996 18172 24998
rect 18196 24996 18252 24998
rect 17956 23962 18012 23964
rect 18036 23962 18092 23964
rect 18116 23962 18172 23964
rect 18196 23962 18252 23964
rect 17956 23910 18002 23962
rect 18002 23910 18012 23962
rect 18036 23910 18066 23962
rect 18066 23910 18078 23962
rect 18078 23910 18092 23962
rect 18116 23910 18130 23962
rect 18130 23910 18142 23962
rect 18142 23910 18172 23962
rect 18196 23910 18206 23962
rect 18206 23910 18252 23962
rect 17956 23908 18012 23910
rect 18036 23908 18092 23910
rect 18116 23908 18172 23910
rect 18196 23908 18252 23910
rect 17956 22874 18012 22876
rect 18036 22874 18092 22876
rect 18116 22874 18172 22876
rect 18196 22874 18252 22876
rect 17956 22822 18002 22874
rect 18002 22822 18012 22874
rect 18036 22822 18066 22874
rect 18066 22822 18078 22874
rect 18078 22822 18092 22874
rect 18116 22822 18130 22874
rect 18130 22822 18142 22874
rect 18142 22822 18172 22874
rect 18196 22822 18206 22874
rect 18206 22822 18252 22874
rect 17956 22820 18012 22822
rect 18036 22820 18092 22822
rect 18116 22820 18172 22822
rect 18196 22820 18252 22822
rect 22956 53882 23012 53884
rect 23036 53882 23092 53884
rect 23116 53882 23172 53884
rect 23196 53882 23252 53884
rect 22956 53830 23002 53882
rect 23002 53830 23012 53882
rect 23036 53830 23066 53882
rect 23066 53830 23078 53882
rect 23078 53830 23092 53882
rect 23116 53830 23130 53882
rect 23130 53830 23142 53882
rect 23142 53830 23172 53882
rect 23196 53830 23206 53882
rect 23206 53830 23252 53882
rect 22956 53828 23012 53830
rect 23036 53828 23092 53830
rect 23116 53828 23172 53830
rect 23196 53828 23252 53830
rect 27956 54426 28012 54428
rect 28036 54426 28092 54428
rect 28116 54426 28172 54428
rect 28196 54426 28252 54428
rect 27956 54374 28002 54426
rect 28002 54374 28012 54426
rect 28036 54374 28066 54426
rect 28066 54374 28078 54426
rect 28078 54374 28092 54426
rect 28116 54374 28130 54426
rect 28130 54374 28142 54426
rect 28142 54374 28172 54426
rect 28196 54374 28206 54426
rect 28206 54374 28252 54426
rect 27956 54372 28012 54374
rect 28036 54372 28092 54374
rect 28116 54372 28172 54374
rect 28196 54372 28252 54374
rect 24950 53932 24952 53952
rect 24952 53932 25004 53952
rect 25004 53932 25006 53952
rect 24950 53896 25006 53932
rect 22956 52794 23012 52796
rect 23036 52794 23092 52796
rect 23116 52794 23172 52796
rect 23196 52794 23252 52796
rect 22956 52742 23002 52794
rect 23002 52742 23012 52794
rect 23036 52742 23066 52794
rect 23066 52742 23078 52794
rect 23078 52742 23092 52794
rect 23116 52742 23130 52794
rect 23130 52742 23142 52794
rect 23142 52742 23172 52794
rect 23196 52742 23206 52794
rect 23206 52742 23252 52794
rect 22956 52740 23012 52742
rect 23036 52740 23092 52742
rect 23116 52740 23172 52742
rect 23196 52740 23252 52742
rect 22956 51706 23012 51708
rect 23036 51706 23092 51708
rect 23116 51706 23172 51708
rect 23196 51706 23252 51708
rect 22956 51654 23002 51706
rect 23002 51654 23012 51706
rect 23036 51654 23066 51706
rect 23066 51654 23078 51706
rect 23078 51654 23092 51706
rect 23116 51654 23130 51706
rect 23130 51654 23142 51706
rect 23142 51654 23172 51706
rect 23196 51654 23206 51706
rect 23206 51654 23252 51706
rect 22956 51652 23012 51654
rect 23036 51652 23092 51654
rect 23116 51652 23172 51654
rect 23196 51652 23252 51654
rect 22956 50618 23012 50620
rect 23036 50618 23092 50620
rect 23116 50618 23172 50620
rect 23196 50618 23252 50620
rect 22956 50566 23002 50618
rect 23002 50566 23012 50618
rect 23036 50566 23066 50618
rect 23066 50566 23078 50618
rect 23078 50566 23092 50618
rect 23116 50566 23130 50618
rect 23130 50566 23142 50618
rect 23142 50566 23172 50618
rect 23196 50566 23206 50618
rect 23206 50566 23252 50618
rect 22956 50564 23012 50566
rect 23036 50564 23092 50566
rect 23116 50564 23172 50566
rect 23196 50564 23252 50566
rect 22956 49530 23012 49532
rect 23036 49530 23092 49532
rect 23116 49530 23172 49532
rect 23196 49530 23252 49532
rect 22956 49478 23002 49530
rect 23002 49478 23012 49530
rect 23036 49478 23066 49530
rect 23066 49478 23078 49530
rect 23078 49478 23092 49530
rect 23116 49478 23130 49530
rect 23130 49478 23142 49530
rect 23142 49478 23172 49530
rect 23196 49478 23206 49530
rect 23206 49478 23252 49530
rect 22956 49476 23012 49478
rect 23036 49476 23092 49478
rect 23116 49476 23172 49478
rect 23196 49476 23252 49478
rect 22956 48442 23012 48444
rect 23036 48442 23092 48444
rect 23116 48442 23172 48444
rect 23196 48442 23252 48444
rect 22956 48390 23002 48442
rect 23002 48390 23012 48442
rect 23036 48390 23066 48442
rect 23066 48390 23078 48442
rect 23078 48390 23092 48442
rect 23116 48390 23130 48442
rect 23130 48390 23142 48442
rect 23142 48390 23172 48442
rect 23196 48390 23206 48442
rect 23206 48390 23252 48442
rect 22956 48388 23012 48390
rect 23036 48388 23092 48390
rect 23116 48388 23172 48390
rect 23196 48388 23252 48390
rect 22956 47354 23012 47356
rect 23036 47354 23092 47356
rect 23116 47354 23172 47356
rect 23196 47354 23252 47356
rect 22956 47302 23002 47354
rect 23002 47302 23012 47354
rect 23036 47302 23066 47354
rect 23066 47302 23078 47354
rect 23078 47302 23092 47354
rect 23116 47302 23130 47354
rect 23130 47302 23142 47354
rect 23142 47302 23172 47354
rect 23196 47302 23206 47354
rect 23206 47302 23252 47354
rect 22956 47300 23012 47302
rect 23036 47300 23092 47302
rect 23116 47300 23172 47302
rect 23196 47300 23252 47302
rect 22956 46266 23012 46268
rect 23036 46266 23092 46268
rect 23116 46266 23172 46268
rect 23196 46266 23252 46268
rect 22956 46214 23002 46266
rect 23002 46214 23012 46266
rect 23036 46214 23066 46266
rect 23066 46214 23078 46266
rect 23078 46214 23092 46266
rect 23116 46214 23130 46266
rect 23130 46214 23142 46266
rect 23142 46214 23172 46266
rect 23196 46214 23206 46266
rect 23206 46214 23252 46266
rect 22956 46212 23012 46214
rect 23036 46212 23092 46214
rect 23116 46212 23172 46214
rect 23196 46212 23252 46214
rect 22956 45178 23012 45180
rect 23036 45178 23092 45180
rect 23116 45178 23172 45180
rect 23196 45178 23252 45180
rect 22956 45126 23002 45178
rect 23002 45126 23012 45178
rect 23036 45126 23066 45178
rect 23066 45126 23078 45178
rect 23078 45126 23092 45178
rect 23116 45126 23130 45178
rect 23130 45126 23142 45178
rect 23142 45126 23172 45178
rect 23196 45126 23206 45178
rect 23206 45126 23252 45178
rect 22956 45124 23012 45126
rect 23036 45124 23092 45126
rect 23116 45124 23172 45126
rect 23196 45124 23252 45126
rect 22956 44090 23012 44092
rect 23036 44090 23092 44092
rect 23116 44090 23172 44092
rect 23196 44090 23252 44092
rect 22956 44038 23002 44090
rect 23002 44038 23012 44090
rect 23036 44038 23066 44090
rect 23066 44038 23078 44090
rect 23078 44038 23092 44090
rect 23116 44038 23130 44090
rect 23130 44038 23142 44090
rect 23142 44038 23172 44090
rect 23196 44038 23206 44090
rect 23206 44038 23252 44090
rect 22956 44036 23012 44038
rect 23036 44036 23092 44038
rect 23116 44036 23172 44038
rect 23196 44036 23252 44038
rect 22956 43002 23012 43004
rect 23036 43002 23092 43004
rect 23116 43002 23172 43004
rect 23196 43002 23252 43004
rect 22956 42950 23002 43002
rect 23002 42950 23012 43002
rect 23036 42950 23066 43002
rect 23066 42950 23078 43002
rect 23078 42950 23092 43002
rect 23116 42950 23130 43002
rect 23130 42950 23142 43002
rect 23142 42950 23172 43002
rect 23196 42950 23206 43002
rect 23206 42950 23252 43002
rect 22956 42948 23012 42950
rect 23036 42948 23092 42950
rect 23116 42948 23172 42950
rect 23196 42948 23252 42950
rect 22956 41914 23012 41916
rect 23036 41914 23092 41916
rect 23116 41914 23172 41916
rect 23196 41914 23252 41916
rect 22956 41862 23002 41914
rect 23002 41862 23012 41914
rect 23036 41862 23066 41914
rect 23066 41862 23078 41914
rect 23078 41862 23092 41914
rect 23116 41862 23130 41914
rect 23130 41862 23142 41914
rect 23142 41862 23172 41914
rect 23196 41862 23206 41914
rect 23206 41862 23252 41914
rect 22956 41860 23012 41862
rect 23036 41860 23092 41862
rect 23116 41860 23172 41862
rect 23196 41860 23252 41862
rect 17956 21786 18012 21788
rect 18036 21786 18092 21788
rect 18116 21786 18172 21788
rect 18196 21786 18252 21788
rect 17956 21734 18002 21786
rect 18002 21734 18012 21786
rect 18036 21734 18066 21786
rect 18066 21734 18078 21786
rect 18078 21734 18092 21786
rect 18116 21734 18130 21786
rect 18130 21734 18142 21786
rect 18142 21734 18172 21786
rect 18196 21734 18206 21786
rect 18206 21734 18252 21786
rect 17956 21732 18012 21734
rect 18036 21732 18092 21734
rect 18116 21732 18172 21734
rect 18196 21732 18252 21734
rect 17956 20698 18012 20700
rect 18036 20698 18092 20700
rect 18116 20698 18172 20700
rect 18196 20698 18252 20700
rect 17956 20646 18002 20698
rect 18002 20646 18012 20698
rect 18036 20646 18066 20698
rect 18066 20646 18078 20698
rect 18078 20646 18092 20698
rect 18116 20646 18130 20698
rect 18130 20646 18142 20698
rect 18142 20646 18172 20698
rect 18196 20646 18206 20698
rect 18206 20646 18252 20698
rect 17956 20644 18012 20646
rect 18036 20644 18092 20646
rect 18116 20644 18172 20646
rect 18196 20644 18252 20646
rect 17956 19610 18012 19612
rect 18036 19610 18092 19612
rect 18116 19610 18172 19612
rect 18196 19610 18252 19612
rect 17956 19558 18002 19610
rect 18002 19558 18012 19610
rect 18036 19558 18066 19610
rect 18066 19558 18078 19610
rect 18078 19558 18092 19610
rect 18116 19558 18130 19610
rect 18130 19558 18142 19610
rect 18142 19558 18172 19610
rect 18196 19558 18206 19610
rect 18206 19558 18252 19610
rect 17956 19556 18012 19558
rect 18036 19556 18092 19558
rect 18116 19556 18172 19558
rect 18196 19556 18252 19558
rect 17956 18522 18012 18524
rect 18036 18522 18092 18524
rect 18116 18522 18172 18524
rect 18196 18522 18252 18524
rect 17956 18470 18002 18522
rect 18002 18470 18012 18522
rect 18036 18470 18066 18522
rect 18066 18470 18078 18522
rect 18078 18470 18092 18522
rect 18116 18470 18130 18522
rect 18130 18470 18142 18522
rect 18142 18470 18172 18522
rect 18196 18470 18206 18522
rect 18206 18470 18252 18522
rect 17956 18468 18012 18470
rect 18036 18468 18092 18470
rect 18116 18468 18172 18470
rect 18196 18468 18252 18470
rect 17956 17434 18012 17436
rect 18036 17434 18092 17436
rect 18116 17434 18172 17436
rect 18196 17434 18252 17436
rect 17956 17382 18002 17434
rect 18002 17382 18012 17434
rect 18036 17382 18066 17434
rect 18066 17382 18078 17434
rect 18078 17382 18092 17434
rect 18116 17382 18130 17434
rect 18130 17382 18142 17434
rect 18142 17382 18172 17434
rect 18196 17382 18206 17434
rect 18206 17382 18252 17434
rect 17956 17380 18012 17382
rect 18036 17380 18092 17382
rect 18116 17380 18172 17382
rect 18196 17380 18252 17382
rect 17956 16346 18012 16348
rect 18036 16346 18092 16348
rect 18116 16346 18172 16348
rect 18196 16346 18252 16348
rect 17956 16294 18002 16346
rect 18002 16294 18012 16346
rect 18036 16294 18066 16346
rect 18066 16294 18078 16346
rect 18078 16294 18092 16346
rect 18116 16294 18130 16346
rect 18130 16294 18142 16346
rect 18142 16294 18172 16346
rect 18196 16294 18206 16346
rect 18206 16294 18252 16346
rect 17956 16292 18012 16294
rect 18036 16292 18092 16294
rect 18116 16292 18172 16294
rect 18196 16292 18252 16294
rect 17956 15258 18012 15260
rect 18036 15258 18092 15260
rect 18116 15258 18172 15260
rect 18196 15258 18252 15260
rect 17956 15206 18002 15258
rect 18002 15206 18012 15258
rect 18036 15206 18066 15258
rect 18066 15206 18078 15258
rect 18078 15206 18092 15258
rect 18116 15206 18130 15258
rect 18130 15206 18142 15258
rect 18142 15206 18172 15258
rect 18196 15206 18206 15258
rect 18206 15206 18252 15258
rect 17956 15204 18012 15206
rect 18036 15204 18092 15206
rect 18116 15204 18172 15206
rect 18196 15204 18252 15206
rect 17956 14170 18012 14172
rect 18036 14170 18092 14172
rect 18116 14170 18172 14172
rect 18196 14170 18252 14172
rect 17956 14118 18002 14170
rect 18002 14118 18012 14170
rect 18036 14118 18066 14170
rect 18066 14118 18078 14170
rect 18078 14118 18092 14170
rect 18116 14118 18130 14170
rect 18130 14118 18142 14170
rect 18142 14118 18172 14170
rect 18196 14118 18206 14170
rect 18206 14118 18252 14170
rect 17956 14116 18012 14118
rect 18036 14116 18092 14118
rect 18116 14116 18172 14118
rect 18196 14116 18252 14118
rect 17956 13082 18012 13084
rect 18036 13082 18092 13084
rect 18116 13082 18172 13084
rect 18196 13082 18252 13084
rect 17956 13030 18002 13082
rect 18002 13030 18012 13082
rect 18036 13030 18066 13082
rect 18066 13030 18078 13082
rect 18078 13030 18092 13082
rect 18116 13030 18130 13082
rect 18130 13030 18142 13082
rect 18142 13030 18172 13082
rect 18196 13030 18206 13082
rect 18206 13030 18252 13082
rect 17956 13028 18012 13030
rect 18036 13028 18092 13030
rect 18116 13028 18172 13030
rect 18196 13028 18252 13030
rect 17956 11994 18012 11996
rect 18036 11994 18092 11996
rect 18116 11994 18172 11996
rect 18196 11994 18252 11996
rect 17956 11942 18002 11994
rect 18002 11942 18012 11994
rect 18036 11942 18066 11994
rect 18066 11942 18078 11994
rect 18078 11942 18092 11994
rect 18116 11942 18130 11994
rect 18130 11942 18142 11994
rect 18142 11942 18172 11994
rect 18196 11942 18206 11994
rect 18206 11942 18252 11994
rect 17956 11940 18012 11942
rect 18036 11940 18092 11942
rect 18116 11940 18172 11942
rect 18196 11940 18252 11942
rect 17956 10906 18012 10908
rect 18036 10906 18092 10908
rect 18116 10906 18172 10908
rect 18196 10906 18252 10908
rect 17956 10854 18002 10906
rect 18002 10854 18012 10906
rect 18036 10854 18066 10906
rect 18066 10854 18078 10906
rect 18078 10854 18092 10906
rect 18116 10854 18130 10906
rect 18130 10854 18142 10906
rect 18142 10854 18172 10906
rect 18196 10854 18206 10906
rect 18206 10854 18252 10906
rect 17956 10852 18012 10854
rect 18036 10852 18092 10854
rect 18116 10852 18172 10854
rect 18196 10852 18252 10854
rect 17956 9818 18012 9820
rect 18036 9818 18092 9820
rect 18116 9818 18172 9820
rect 18196 9818 18252 9820
rect 17956 9766 18002 9818
rect 18002 9766 18012 9818
rect 18036 9766 18066 9818
rect 18066 9766 18078 9818
rect 18078 9766 18092 9818
rect 18116 9766 18130 9818
rect 18130 9766 18142 9818
rect 18142 9766 18172 9818
rect 18196 9766 18206 9818
rect 18206 9766 18252 9818
rect 17956 9764 18012 9766
rect 18036 9764 18092 9766
rect 18116 9764 18172 9766
rect 18196 9764 18252 9766
rect 17956 8730 18012 8732
rect 18036 8730 18092 8732
rect 18116 8730 18172 8732
rect 18196 8730 18252 8732
rect 17956 8678 18002 8730
rect 18002 8678 18012 8730
rect 18036 8678 18066 8730
rect 18066 8678 18078 8730
rect 18078 8678 18092 8730
rect 18116 8678 18130 8730
rect 18130 8678 18142 8730
rect 18142 8678 18172 8730
rect 18196 8678 18206 8730
rect 18206 8678 18252 8730
rect 17956 8676 18012 8678
rect 18036 8676 18092 8678
rect 18116 8676 18172 8678
rect 18196 8676 18252 8678
rect 17956 7642 18012 7644
rect 18036 7642 18092 7644
rect 18116 7642 18172 7644
rect 18196 7642 18252 7644
rect 17956 7590 18002 7642
rect 18002 7590 18012 7642
rect 18036 7590 18066 7642
rect 18066 7590 18078 7642
rect 18078 7590 18092 7642
rect 18116 7590 18130 7642
rect 18130 7590 18142 7642
rect 18142 7590 18172 7642
rect 18196 7590 18206 7642
rect 18206 7590 18252 7642
rect 17956 7588 18012 7590
rect 18036 7588 18092 7590
rect 18116 7588 18172 7590
rect 18196 7588 18252 7590
rect 17956 6554 18012 6556
rect 18036 6554 18092 6556
rect 18116 6554 18172 6556
rect 18196 6554 18252 6556
rect 17956 6502 18002 6554
rect 18002 6502 18012 6554
rect 18036 6502 18066 6554
rect 18066 6502 18078 6554
rect 18078 6502 18092 6554
rect 18116 6502 18130 6554
rect 18130 6502 18142 6554
rect 18142 6502 18172 6554
rect 18196 6502 18206 6554
rect 18206 6502 18252 6554
rect 17956 6500 18012 6502
rect 18036 6500 18092 6502
rect 18116 6500 18172 6502
rect 18196 6500 18252 6502
rect 17956 5466 18012 5468
rect 18036 5466 18092 5468
rect 18116 5466 18172 5468
rect 18196 5466 18252 5468
rect 17956 5414 18002 5466
rect 18002 5414 18012 5466
rect 18036 5414 18066 5466
rect 18066 5414 18078 5466
rect 18078 5414 18092 5466
rect 18116 5414 18130 5466
rect 18130 5414 18142 5466
rect 18142 5414 18172 5466
rect 18196 5414 18206 5466
rect 18206 5414 18252 5466
rect 17956 5412 18012 5414
rect 18036 5412 18092 5414
rect 18116 5412 18172 5414
rect 18196 5412 18252 5414
rect 17956 4378 18012 4380
rect 18036 4378 18092 4380
rect 18116 4378 18172 4380
rect 18196 4378 18252 4380
rect 17956 4326 18002 4378
rect 18002 4326 18012 4378
rect 18036 4326 18066 4378
rect 18066 4326 18078 4378
rect 18078 4326 18092 4378
rect 18116 4326 18130 4378
rect 18130 4326 18142 4378
rect 18142 4326 18172 4378
rect 18196 4326 18206 4378
rect 18206 4326 18252 4378
rect 17956 4324 18012 4326
rect 18036 4324 18092 4326
rect 18116 4324 18172 4326
rect 18196 4324 18252 4326
rect 17956 3290 18012 3292
rect 18036 3290 18092 3292
rect 18116 3290 18172 3292
rect 18196 3290 18252 3292
rect 17956 3238 18002 3290
rect 18002 3238 18012 3290
rect 18036 3238 18066 3290
rect 18066 3238 18078 3290
rect 18078 3238 18092 3290
rect 18116 3238 18130 3290
rect 18130 3238 18142 3290
rect 18142 3238 18172 3290
rect 18196 3238 18206 3290
rect 18206 3238 18252 3290
rect 17956 3236 18012 3238
rect 18036 3236 18092 3238
rect 18116 3236 18172 3238
rect 18196 3236 18252 3238
rect 22098 30096 22154 30152
rect 17956 2202 18012 2204
rect 18036 2202 18092 2204
rect 18116 2202 18172 2204
rect 18196 2202 18252 2204
rect 17956 2150 18002 2202
rect 18002 2150 18012 2202
rect 18036 2150 18066 2202
rect 18066 2150 18078 2202
rect 18078 2150 18092 2202
rect 18116 2150 18130 2202
rect 18130 2150 18142 2202
rect 18142 2150 18172 2202
rect 18196 2150 18206 2202
rect 18206 2150 18252 2202
rect 17956 2148 18012 2150
rect 18036 2148 18092 2150
rect 18116 2148 18172 2150
rect 18196 2148 18252 2150
rect 22374 38936 22430 38992
rect 22956 40826 23012 40828
rect 23036 40826 23092 40828
rect 23116 40826 23172 40828
rect 23196 40826 23252 40828
rect 22956 40774 23002 40826
rect 23002 40774 23012 40826
rect 23036 40774 23066 40826
rect 23066 40774 23078 40826
rect 23078 40774 23092 40826
rect 23116 40774 23130 40826
rect 23130 40774 23142 40826
rect 23142 40774 23172 40826
rect 23196 40774 23206 40826
rect 23206 40774 23252 40826
rect 22956 40772 23012 40774
rect 23036 40772 23092 40774
rect 23116 40772 23172 40774
rect 23196 40772 23252 40774
rect 22956 39738 23012 39740
rect 23036 39738 23092 39740
rect 23116 39738 23172 39740
rect 23196 39738 23252 39740
rect 22956 39686 23002 39738
rect 23002 39686 23012 39738
rect 23036 39686 23066 39738
rect 23066 39686 23078 39738
rect 23078 39686 23092 39738
rect 23116 39686 23130 39738
rect 23130 39686 23142 39738
rect 23142 39686 23172 39738
rect 23196 39686 23206 39738
rect 23206 39686 23252 39738
rect 22956 39684 23012 39686
rect 23036 39684 23092 39686
rect 23116 39684 23172 39686
rect 23196 39684 23252 39686
rect 22956 38650 23012 38652
rect 23036 38650 23092 38652
rect 23116 38650 23172 38652
rect 23196 38650 23252 38652
rect 22956 38598 23002 38650
rect 23002 38598 23012 38650
rect 23036 38598 23066 38650
rect 23066 38598 23078 38650
rect 23078 38598 23092 38650
rect 23116 38598 23130 38650
rect 23130 38598 23142 38650
rect 23142 38598 23172 38650
rect 23196 38598 23206 38650
rect 23206 38598 23252 38650
rect 22956 38596 23012 38598
rect 23036 38596 23092 38598
rect 23116 38596 23172 38598
rect 23196 38596 23252 38598
rect 22956 37562 23012 37564
rect 23036 37562 23092 37564
rect 23116 37562 23172 37564
rect 23196 37562 23252 37564
rect 22956 37510 23002 37562
rect 23002 37510 23012 37562
rect 23036 37510 23066 37562
rect 23066 37510 23078 37562
rect 23078 37510 23092 37562
rect 23116 37510 23130 37562
rect 23130 37510 23142 37562
rect 23142 37510 23172 37562
rect 23196 37510 23206 37562
rect 23206 37510 23252 37562
rect 22956 37508 23012 37510
rect 23036 37508 23092 37510
rect 23116 37508 23172 37510
rect 23196 37508 23252 37510
rect 22956 36474 23012 36476
rect 23036 36474 23092 36476
rect 23116 36474 23172 36476
rect 23196 36474 23252 36476
rect 22956 36422 23002 36474
rect 23002 36422 23012 36474
rect 23036 36422 23066 36474
rect 23066 36422 23078 36474
rect 23078 36422 23092 36474
rect 23116 36422 23130 36474
rect 23130 36422 23142 36474
rect 23142 36422 23172 36474
rect 23196 36422 23206 36474
rect 23206 36422 23252 36474
rect 22956 36420 23012 36422
rect 23036 36420 23092 36422
rect 23116 36420 23172 36422
rect 23196 36420 23252 36422
rect 22466 31220 22468 31240
rect 22468 31220 22520 31240
rect 22520 31220 22522 31240
rect 22466 31184 22522 31220
rect 22956 35386 23012 35388
rect 23036 35386 23092 35388
rect 23116 35386 23172 35388
rect 23196 35386 23252 35388
rect 22956 35334 23002 35386
rect 23002 35334 23012 35386
rect 23036 35334 23066 35386
rect 23066 35334 23078 35386
rect 23078 35334 23092 35386
rect 23116 35334 23130 35386
rect 23130 35334 23142 35386
rect 23142 35334 23172 35386
rect 23196 35334 23206 35386
rect 23206 35334 23252 35386
rect 22956 35332 23012 35334
rect 23036 35332 23092 35334
rect 23116 35332 23172 35334
rect 23196 35332 23252 35334
rect 22956 34298 23012 34300
rect 23036 34298 23092 34300
rect 23116 34298 23172 34300
rect 23196 34298 23252 34300
rect 22956 34246 23002 34298
rect 23002 34246 23012 34298
rect 23036 34246 23066 34298
rect 23066 34246 23078 34298
rect 23078 34246 23092 34298
rect 23116 34246 23130 34298
rect 23130 34246 23142 34298
rect 23142 34246 23172 34298
rect 23196 34246 23206 34298
rect 23206 34246 23252 34298
rect 22956 34244 23012 34246
rect 23036 34244 23092 34246
rect 23116 34244 23172 34246
rect 23196 34244 23252 34246
rect 22956 33210 23012 33212
rect 23036 33210 23092 33212
rect 23116 33210 23172 33212
rect 23196 33210 23252 33212
rect 22956 33158 23002 33210
rect 23002 33158 23012 33210
rect 23036 33158 23066 33210
rect 23066 33158 23078 33210
rect 23078 33158 23092 33210
rect 23116 33158 23130 33210
rect 23130 33158 23142 33210
rect 23142 33158 23172 33210
rect 23196 33158 23206 33210
rect 23206 33158 23252 33210
rect 22956 33156 23012 33158
rect 23036 33156 23092 33158
rect 23116 33156 23172 33158
rect 23196 33156 23252 33158
rect 22956 32122 23012 32124
rect 23036 32122 23092 32124
rect 23116 32122 23172 32124
rect 23196 32122 23252 32124
rect 22956 32070 23002 32122
rect 23002 32070 23012 32122
rect 23036 32070 23066 32122
rect 23066 32070 23078 32122
rect 23078 32070 23092 32122
rect 23116 32070 23130 32122
rect 23130 32070 23142 32122
rect 23142 32070 23172 32122
rect 23196 32070 23206 32122
rect 23206 32070 23252 32122
rect 22956 32068 23012 32070
rect 23036 32068 23092 32070
rect 23116 32068 23172 32070
rect 23196 32068 23252 32070
rect 22956 31034 23012 31036
rect 23036 31034 23092 31036
rect 23116 31034 23172 31036
rect 23196 31034 23252 31036
rect 22956 30982 23002 31034
rect 23002 30982 23012 31034
rect 23036 30982 23066 31034
rect 23066 30982 23078 31034
rect 23078 30982 23092 31034
rect 23116 30982 23130 31034
rect 23130 30982 23142 31034
rect 23142 30982 23172 31034
rect 23196 30982 23206 31034
rect 23206 30982 23252 31034
rect 22956 30980 23012 30982
rect 23036 30980 23092 30982
rect 23116 30980 23172 30982
rect 23196 30980 23252 30982
rect 24398 35264 24454 35320
rect 24214 32816 24270 32872
rect 22956 29946 23012 29948
rect 23036 29946 23092 29948
rect 23116 29946 23172 29948
rect 23196 29946 23252 29948
rect 22956 29894 23002 29946
rect 23002 29894 23012 29946
rect 23036 29894 23066 29946
rect 23066 29894 23078 29946
rect 23078 29894 23092 29946
rect 23116 29894 23130 29946
rect 23130 29894 23142 29946
rect 23142 29894 23172 29946
rect 23196 29894 23206 29946
rect 23206 29894 23252 29946
rect 22956 29892 23012 29894
rect 23036 29892 23092 29894
rect 23116 29892 23172 29894
rect 23196 29892 23252 29894
rect 22956 28858 23012 28860
rect 23036 28858 23092 28860
rect 23116 28858 23172 28860
rect 23196 28858 23252 28860
rect 22956 28806 23002 28858
rect 23002 28806 23012 28858
rect 23036 28806 23066 28858
rect 23066 28806 23078 28858
rect 23078 28806 23092 28858
rect 23116 28806 23130 28858
rect 23130 28806 23142 28858
rect 23142 28806 23172 28858
rect 23196 28806 23206 28858
rect 23206 28806 23252 28858
rect 22956 28804 23012 28806
rect 23036 28804 23092 28806
rect 23116 28804 23172 28806
rect 23196 28804 23252 28806
rect 22956 27770 23012 27772
rect 23036 27770 23092 27772
rect 23116 27770 23172 27772
rect 23196 27770 23252 27772
rect 22956 27718 23002 27770
rect 23002 27718 23012 27770
rect 23036 27718 23066 27770
rect 23066 27718 23078 27770
rect 23078 27718 23092 27770
rect 23116 27718 23130 27770
rect 23130 27718 23142 27770
rect 23142 27718 23172 27770
rect 23196 27718 23206 27770
rect 23206 27718 23252 27770
rect 22956 27716 23012 27718
rect 23036 27716 23092 27718
rect 23116 27716 23172 27718
rect 23196 27716 23252 27718
rect 22956 26682 23012 26684
rect 23036 26682 23092 26684
rect 23116 26682 23172 26684
rect 23196 26682 23252 26684
rect 22956 26630 23002 26682
rect 23002 26630 23012 26682
rect 23036 26630 23066 26682
rect 23066 26630 23078 26682
rect 23078 26630 23092 26682
rect 23116 26630 23130 26682
rect 23130 26630 23142 26682
rect 23142 26630 23172 26682
rect 23196 26630 23206 26682
rect 23206 26630 23252 26682
rect 22956 26628 23012 26630
rect 23036 26628 23092 26630
rect 23116 26628 23172 26630
rect 23196 26628 23252 26630
rect 22466 23568 22522 23624
rect 22956 25594 23012 25596
rect 23036 25594 23092 25596
rect 23116 25594 23172 25596
rect 23196 25594 23252 25596
rect 22956 25542 23002 25594
rect 23002 25542 23012 25594
rect 23036 25542 23066 25594
rect 23066 25542 23078 25594
rect 23078 25542 23092 25594
rect 23116 25542 23130 25594
rect 23130 25542 23142 25594
rect 23142 25542 23172 25594
rect 23196 25542 23206 25594
rect 23206 25542 23252 25594
rect 22956 25540 23012 25542
rect 23036 25540 23092 25542
rect 23116 25540 23172 25542
rect 23196 25540 23252 25542
rect 22956 24506 23012 24508
rect 23036 24506 23092 24508
rect 23116 24506 23172 24508
rect 23196 24506 23252 24508
rect 22956 24454 23002 24506
rect 23002 24454 23012 24506
rect 23036 24454 23066 24506
rect 23066 24454 23078 24506
rect 23078 24454 23092 24506
rect 23116 24454 23130 24506
rect 23130 24454 23142 24506
rect 23142 24454 23172 24506
rect 23196 24454 23206 24506
rect 23206 24454 23252 24506
rect 22956 24452 23012 24454
rect 23036 24452 23092 24454
rect 23116 24452 23172 24454
rect 23196 24452 23252 24454
rect 22558 20440 22614 20496
rect 23386 23588 23442 23624
rect 23386 23568 23388 23588
rect 23388 23568 23440 23588
rect 23440 23568 23442 23588
rect 23386 23432 23442 23488
rect 22956 23418 23012 23420
rect 23036 23418 23092 23420
rect 23116 23418 23172 23420
rect 23196 23418 23252 23420
rect 22956 23366 23002 23418
rect 23002 23366 23012 23418
rect 23036 23366 23066 23418
rect 23066 23366 23078 23418
rect 23078 23366 23092 23418
rect 23116 23366 23130 23418
rect 23130 23366 23142 23418
rect 23142 23366 23172 23418
rect 23196 23366 23206 23418
rect 23206 23366 23252 23418
rect 22956 23364 23012 23366
rect 23036 23364 23092 23366
rect 23116 23364 23172 23366
rect 23196 23364 23252 23366
rect 22956 22330 23012 22332
rect 23036 22330 23092 22332
rect 23116 22330 23172 22332
rect 23196 22330 23252 22332
rect 22956 22278 23002 22330
rect 23002 22278 23012 22330
rect 23036 22278 23066 22330
rect 23066 22278 23078 22330
rect 23078 22278 23092 22330
rect 23116 22278 23130 22330
rect 23130 22278 23142 22330
rect 23142 22278 23172 22330
rect 23196 22278 23206 22330
rect 23206 22278 23252 22330
rect 22956 22276 23012 22278
rect 23036 22276 23092 22278
rect 23116 22276 23172 22278
rect 23196 22276 23252 22278
rect 22956 21242 23012 21244
rect 23036 21242 23092 21244
rect 23116 21242 23172 21244
rect 23196 21242 23252 21244
rect 22956 21190 23002 21242
rect 23002 21190 23012 21242
rect 23036 21190 23066 21242
rect 23066 21190 23078 21242
rect 23078 21190 23092 21242
rect 23116 21190 23130 21242
rect 23130 21190 23142 21242
rect 23142 21190 23172 21242
rect 23196 21190 23206 21242
rect 23206 21190 23252 21242
rect 22956 21188 23012 21190
rect 23036 21188 23092 21190
rect 23116 21188 23172 21190
rect 23196 21188 23252 21190
rect 23294 20476 23296 20496
rect 23296 20476 23348 20496
rect 23348 20476 23350 20496
rect 23294 20440 23350 20476
rect 22956 20154 23012 20156
rect 23036 20154 23092 20156
rect 23116 20154 23172 20156
rect 23196 20154 23252 20156
rect 22956 20102 23002 20154
rect 23002 20102 23012 20154
rect 23036 20102 23066 20154
rect 23066 20102 23078 20154
rect 23078 20102 23092 20154
rect 23116 20102 23130 20154
rect 23130 20102 23142 20154
rect 23142 20102 23172 20154
rect 23196 20102 23206 20154
rect 23206 20102 23252 20154
rect 22956 20100 23012 20102
rect 23036 20100 23092 20102
rect 23116 20100 23172 20102
rect 23196 20100 23252 20102
rect 22956 19066 23012 19068
rect 23036 19066 23092 19068
rect 23116 19066 23172 19068
rect 23196 19066 23252 19068
rect 22956 19014 23002 19066
rect 23002 19014 23012 19066
rect 23036 19014 23066 19066
rect 23066 19014 23078 19066
rect 23078 19014 23092 19066
rect 23116 19014 23130 19066
rect 23130 19014 23142 19066
rect 23142 19014 23172 19066
rect 23196 19014 23206 19066
rect 23206 19014 23252 19066
rect 22956 19012 23012 19014
rect 23036 19012 23092 19014
rect 23116 19012 23172 19014
rect 23196 19012 23252 19014
rect 22834 18808 22890 18864
rect 22956 17978 23012 17980
rect 23036 17978 23092 17980
rect 23116 17978 23172 17980
rect 23196 17978 23252 17980
rect 22956 17926 23002 17978
rect 23002 17926 23012 17978
rect 23036 17926 23066 17978
rect 23066 17926 23078 17978
rect 23078 17926 23092 17978
rect 23116 17926 23130 17978
rect 23130 17926 23142 17978
rect 23142 17926 23172 17978
rect 23196 17926 23206 17978
rect 23206 17926 23252 17978
rect 22956 17924 23012 17926
rect 23036 17924 23092 17926
rect 23116 17924 23172 17926
rect 23196 17924 23252 17926
rect 22956 16890 23012 16892
rect 23036 16890 23092 16892
rect 23116 16890 23172 16892
rect 23196 16890 23252 16892
rect 22956 16838 23002 16890
rect 23002 16838 23012 16890
rect 23036 16838 23066 16890
rect 23066 16838 23078 16890
rect 23078 16838 23092 16890
rect 23116 16838 23130 16890
rect 23130 16838 23142 16890
rect 23142 16838 23172 16890
rect 23196 16838 23206 16890
rect 23206 16838 23252 16890
rect 22956 16836 23012 16838
rect 23036 16836 23092 16838
rect 23116 16836 23172 16838
rect 23196 16836 23252 16838
rect 22956 15802 23012 15804
rect 23036 15802 23092 15804
rect 23116 15802 23172 15804
rect 23196 15802 23252 15804
rect 22956 15750 23002 15802
rect 23002 15750 23012 15802
rect 23036 15750 23066 15802
rect 23066 15750 23078 15802
rect 23078 15750 23092 15802
rect 23116 15750 23130 15802
rect 23130 15750 23142 15802
rect 23142 15750 23172 15802
rect 23196 15750 23206 15802
rect 23206 15750 23252 15802
rect 22956 15748 23012 15750
rect 23036 15748 23092 15750
rect 23116 15748 23172 15750
rect 23196 15748 23252 15750
rect 21086 2352 21142 2408
rect 22956 14714 23012 14716
rect 23036 14714 23092 14716
rect 23116 14714 23172 14716
rect 23196 14714 23252 14716
rect 22956 14662 23002 14714
rect 23002 14662 23012 14714
rect 23036 14662 23066 14714
rect 23066 14662 23078 14714
rect 23078 14662 23092 14714
rect 23116 14662 23130 14714
rect 23130 14662 23142 14714
rect 23142 14662 23172 14714
rect 23196 14662 23206 14714
rect 23206 14662 23252 14714
rect 22956 14660 23012 14662
rect 23036 14660 23092 14662
rect 23116 14660 23172 14662
rect 23196 14660 23252 14662
rect 22956 13626 23012 13628
rect 23036 13626 23092 13628
rect 23116 13626 23172 13628
rect 23196 13626 23252 13628
rect 22956 13574 23002 13626
rect 23002 13574 23012 13626
rect 23036 13574 23066 13626
rect 23066 13574 23078 13626
rect 23078 13574 23092 13626
rect 23116 13574 23130 13626
rect 23130 13574 23142 13626
rect 23142 13574 23172 13626
rect 23196 13574 23206 13626
rect 23206 13574 23252 13626
rect 22956 13572 23012 13574
rect 23036 13572 23092 13574
rect 23116 13572 23172 13574
rect 23196 13572 23252 13574
rect 22956 12538 23012 12540
rect 23036 12538 23092 12540
rect 23116 12538 23172 12540
rect 23196 12538 23252 12540
rect 22956 12486 23002 12538
rect 23002 12486 23012 12538
rect 23036 12486 23066 12538
rect 23066 12486 23078 12538
rect 23078 12486 23092 12538
rect 23116 12486 23130 12538
rect 23130 12486 23142 12538
rect 23142 12486 23172 12538
rect 23196 12486 23206 12538
rect 23206 12486 23252 12538
rect 22956 12484 23012 12486
rect 23036 12484 23092 12486
rect 23116 12484 23172 12486
rect 23196 12484 23252 12486
rect 22956 11450 23012 11452
rect 23036 11450 23092 11452
rect 23116 11450 23172 11452
rect 23196 11450 23252 11452
rect 22956 11398 23002 11450
rect 23002 11398 23012 11450
rect 23036 11398 23066 11450
rect 23066 11398 23078 11450
rect 23078 11398 23092 11450
rect 23116 11398 23130 11450
rect 23130 11398 23142 11450
rect 23142 11398 23172 11450
rect 23196 11398 23206 11450
rect 23206 11398 23252 11450
rect 22956 11396 23012 11398
rect 23036 11396 23092 11398
rect 23116 11396 23172 11398
rect 23196 11396 23252 11398
rect 22956 10362 23012 10364
rect 23036 10362 23092 10364
rect 23116 10362 23172 10364
rect 23196 10362 23252 10364
rect 22956 10310 23002 10362
rect 23002 10310 23012 10362
rect 23036 10310 23066 10362
rect 23066 10310 23078 10362
rect 23078 10310 23092 10362
rect 23116 10310 23130 10362
rect 23130 10310 23142 10362
rect 23142 10310 23172 10362
rect 23196 10310 23206 10362
rect 23206 10310 23252 10362
rect 22956 10308 23012 10310
rect 23036 10308 23092 10310
rect 23116 10308 23172 10310
rect 23196 10308 23252 10310
rect 22956 9274 23012 9276
rect 23036 9274 23092 9276
rect 23116 9274 23172 9276
rect 23196 9274 23252 9276
rect 22956 9222 23002 9274
rect 23002 9222 23012 9274
rect 23036 9222 23066 9274
rect 23066 9222 23078 9274
rect 23078 9222 23092 9274
rect 23116 9222 23130 9274
rect 23130 9222 23142 9274
rect 23142 9222 23172 9274
rect 23196 9222 23206 9274
rect 23206 9222 23252 9274
rect 22956 9220 23012 9222
rect 23036 9220 23092 9222
rect 23116 9220 23172 9222
rect 23196 9220 23252 9222
rect 22956 8186 23012 8188
rect 23036 8186 23092 8188
rect 23116 8186 23172 8188
rect 23196 8186 23252 8188
rect 22956 8134 23002 8186
rect 23002 8134 23012 8186
rect 23036 8134 23066 8186
rect 23066 8134 23078 8186
rect 23078 8134 23092 8186
rect 23116 8134 23130 8186
rect 23130 8134 23142 8186
rect 23142 8134 23172 8186
rect 23196 8134 23206 8186
rect 23206 8134 23252 8186
rect 22956 8132 23012 8134
rect 23036 8132 23092 8134
rect 23116 8132 23172 8134
rect 23196 8132 23252 8134
rect 22956 7098 23012 7100
rect 23036 7098 23092 7100
rect 23116 7098 23172 7100
rect 23196 7098 23252 7100
rect 22956 7046 23002 7098
rect 23002 7046 23012 7098
rect 23036 7046 23066 7098
rect 23066 7046 23078 7098
rect 23078 7046 23092 7098
rect 23116 7046 23130 7098
rect 23130 7046 23142 7098
rect 23142 7046 23172 7098
rect 23196 7046 23206 7098
rect 23206 7046 23252 7098
rect 22956 7044 23012 7046
rect 23036 7044 23092 7046
rect 23116 7044 23172 7046
rect 23196 7044 23252 7046
rect 22956 6010 23012 6012
rect 23036 6010 23092 6012
rect 23116 6010 23172 6012
rect 23196 6010 23252 6012
rect 22956 5958 23002 6010
rect 23002 5958 23012 6010
rect 23036 5958 23066 6010
rect 23066 5958 23078 6010
rect 23078 5958 23092 6010
rect 23116 5958 23130 6010
rect 23130 5958 23142 6010
rect 23142 5958 23172 6010
rect 23196 5958 23206 6010
rect 23206 5958 23252 6010
rect 22956 5956 23012 5958
rect 23036 5956 23092 5958
rect 23116 5956 23172 5958
rect 23196 5956 23252 5958
rect 22956 4922 23012 4924
rect 23036 4922 23092 4924
rect 23116 4922 23172 4924
rect 23196 4922 23252 4924
rect 22956 4870 23002 4922
rect 23002 4870 23012 4922
rect 23036 4870 23066 4922
rect 23066 4870 23078 4922
rect 23078 4870 23092 4922
rect 23116 4870 23130 4922
rect 23130 4870 23142 4922
rect 23142 4870 23172 4922
rect 23196 4870 23206 4922
rect 23206 4870 23252 4922
rect 22956 4868 23012 4870
rect 23036 4868 23092 4870
rect 23116 4868 23172 4870
rect 23196 4868 23252 4870
rect 22956 3834 23012 3836
rect 23036 3834 23092 3836
rect 23116 3834 23172 3836
rect 23196 3834 23252 3836
rect 22956 3782 23002 3834
rect 23002 3782 23012 3834
rect 23036 3782 23066 3834
rect 23066 3782 23078 3834
rect 23078 3782 23092 3834
rect 23116 3782 23130 3834
rect 23130 3782 23142 3834
rect 23142 3782 23172 3834
rect 23196 3782 23206 3834
rect 23206 3782 23252 3834
rect 22956 3780 23012 3782
rect 23036 3780 23092 3782
rect 23116 3780 23172 3782
rect 23196 3780 23252 3782
rect 22956 2746 23012 2748
rect 23036 2746 23092 2748
rect 23116 2746 23172 2748
rect 23196 2746 23252 2748
rect 22956 2694 23002 2746
rect 23002 2694 23012 2746
rect 23036 2694 23066 2746
rect 23066 2694 23078 2746
rect 23078 2694 23092 2746
rect 23116 2694 23130 2746
rect 23130 2694 23142 2746
rect 23142 2694 23172 2746
rect 23196 2694 23206 2746
rect 23206 2694 23252 2746
rect 22956 2692 23012 2694
rect 23036 2692 23092 2694
rect 23116 2692 23172 2694
rect 23196 2692 23252 2694
rect 25594 35944 25650 36000
rect 25042 22924 25044 22944
rect 25044 22924 25096 22944
rect 25096 22924 25098 22944
rect 25042 22888 25098 22924
rect 25778 35672 25834 35728
rect 27066 40024 27122 40080
rect 27342 36896 27398 36952
rect 27956 53338 28012 53340
rect 28036 53338 28092 53340
rect 28116 53338 28172 53340
rect 28196 53338 28252 53340
rect 27956 53286 28002 53338
rect 28002 53286 28012 53338
rect 28036 53286 28066 53338
rect 28066 53286 28078 53338
rect 28078 53286 28092 53338
rect 28116 53286 28130 53338
rect 28130 53286 28142 53338
rect 28142 53286 28172 53338
rect 28196 53286 28206 53338
rect 28206 53286 28252 53338
rect 27956 53284 28012 53286
rect 28036 53284 28092 53286
rect 28116 53284 28172 53286
rect 28196 53284 28252 53286
rect 27956 52250 28012 52252
rect 28036 52250 28092 52252
rect 28116 52250 28172 52252
rect 28196 52250 28252 52252
rect 27956 52198 28002 52250
rect 28002 52198 28012 52250
rect 28036 52198 28066 52250
rect 28066 52198 28078 52250
rect 28078 52198 28092 52250
rect 28116 52198 28130 52250
rect 28130 52198 28142 52250
rect 28142 52198 28172 52250
rect 28196 52198 28206 52250
rect 28206 52198 28252 52250
rect 27956 52196 28012 52198
rect 28036 52196 28092 52198
rect 28116 52196 28172 52198
rect 28196 52196 28252 52198
rect 27956 51162 28012 51164
rect 28036 51162 28092 51164
rect 28116 51162 28172 51164
rect 28196 51162 28252 51164
rect 27956 51110 28002 51162
rect 28002 51110 28012 51162
rect 28036 51110 28066 51162
rect 28066 51110 28078 51162
rect 28078 51110 28092 51162
rect 28116 51110 28130 51162
rect 28130 51110 28142 51162
rect 28142 51110 28172 51162
rect 28196 51110 28206 51162
rect 28206 51110 28252 51162
rect 27956 51108 28012 51110
rect 28036 51108 28092 51110
rect 28116 51108 28172 51110
rect 28196 51108 28252 51110
rect 27956 50074 28012 50076
rect 28036 50074 28092 50076
rect 28116 50074 28172 50076
rect 28196 50074 28252 50076
rect 27956 50022 28002 50074
rect 28002 50022 28012 50074
rect 28036 50022 28066 50074
rect 28066 50022 28078 50074
rect 28078 50022 28092 50074
rect 28116 50022 28130 50074
rect 28130 50022 28142 50074
rect 28142 50022 28172 50074
rect 28196 50022 28206 50074
rect 28206 50022 28252 50074
rect 27956 50020 28012 50022
rect 28036 50020 28092 50022
rect 28116 50020 28172 50022
rect 28196 50020 28252 50022
rect 27956 48986 28012 48988
rect 28036 48986 28092 48988
rect 28116 48986 28172 48988
rect 28196 48986 28252 48988
rect 27956 48934 28002 48986
rect 28002 48934 28012 48986
rect 28036 48934 28066 48986
rect 28066 48934 28078 48986
rect 28078 48934 28092 48986
rect 28116 48934 28130 48986
rect 28130 48934 28142 48986
rect 28142 48934 28172 48986
rect 28196 48934 28206 48986
rect 28206 48934 28252 48986
rect 27956 48932 28012 48934
rect 28036 48932 28092 48934
rect 28116 48932 28172 48934
rect 28196 48932 28252 48934
rect 27956 47898 28012 47900
rect 28036 47898 28092 47900
rect 28116 47898 28172 47900
rect 28196 47898 28252 47900
rect 27956 47846 28002 47898
rect 28002 47846 28012 47898
rect 28036 47846 28066 47898
rect 28066 47846 28078 47898
rect 28078 47846 28092 47898
rect 28116 47846 28130 47898
rect 28130 47846 28142 47898
rect 28142 47846 28172 47898
rect 28196 47846 28206 47898
rect 28206 47846 28252 47898
rect 27956 47844 28012 47846
rect 28036 47844 28092 47846
rect 28116 47844 28172 47846
rect 28196 47844 28252 47846
rect 27956 46810 28012 46812
rect 28036 46810 28092 46812
rect 28116 46810 28172 46812
rect 28196 46810 28252 46812
rect 27956 46758 28002 46810
rect 28002 46758 28012 46810
rect 28036 46758 28066 46810
rect 28066 46758 28078 46810
rect 28078 46758 28092 46810
rect 28116 46758 28130 46810
rect 28130 46758 28142 46810
rect 28142 46758 28172 46810
rect 28196 46758 28206 46810
rect 28206 46758 28252 46810
rect 27956 46756 28012 46758
rect 28036 46756 28092 46758
rect 28116 46756 28172 46758
rect 28196 46756 28252 46758
rect 27956 45722 28012 45724
rect 28036 45722 28092 45724
rect 28116 45722 28172 45724
rect 28196 45722 28252 45724
rect 27956 45670 28002 45722
rect 28002 45670 28012 45722
rect 28036 45670 28066 45722
rect 28066 45670 28078 45722
rect 28078 45670 28092 45722
rect 28116 45670 28130 45722
rect 28130 45670 28142 45722
rect 28142 45670 28172 45722
rect 28196 45670 28206 45722
rect 28206 45670 28252 45722
rect 27956 45668 28012 45670
rect 28036 45668 28092 45670
rect 28116 45668 28172 45670
rect 28196 45668 28252 45670
rect 27956 44634 28012 44636
rect 28036 44634 28092 44636
rect 28116 44634 28172 44636
rect 28196 44634 28252 44636
rect 27956 44582 28002 44634
rect 28002 44582 28012 44634
rect 28036 44582 28066 44634
rect 28066 44582 28078 44634
rect 28078 44582 28092 44634
rect 28116 44582 28130 44634
rect 28130 44582 28142 44634
rect 28142 44582 28172 44634
rect 28196 44582 28206 44634
rect 28206 44582 28252 44634
rect 27956 44580 28012 44582
rect 28036 44580 28092 44582
rect 28116 44580 28172 44582
rect 28196 44580 28252 44582
rect 27956 43546 28012 43548
rect 28036 43546 28092 43548
rect 28116 43546 28172 43548
rect 28196 43546 28252 43548
rect 27956 43494 28002 43546
rect 28002 43494 28012 43546
rect 28036 43494 28066 43546
rect 28066 43494 28078 43546
rect 28078 43494 28092 43546
rect 28116 43494 28130 43546
rect 28130 43494 28142 43546
rect 28142 43494 28172 43546
rect 28196 43494 28206 43546
rect 28206 43494 28252 43546
rect 27956 43492 28012 43494
rect 28036 43492 28092 43494
rect 28116 43492 28172 43494
rect 28196 43492 28252 43494
rect 27956 42458 28012 42460
rect 28036 42458 28092 42460
rect 28116 42458 28172 42460
rect 28196 42458 28252 42460
rect 27956 42406 28002 42458
rect 28002 42406 28012 42458
rect 28036 42406 28066 42458
rect 28066 42406 28078 42458
rect 28078 42406 28092 42458
rect 28116 42406 28130 42458
rect 28130 42406 28142 42458
rect 28142 42406 28172 42458
rect 28196 42406 28206 42458
rect 28206 42406 28252 42458
rect 27956 42404 28012 42406
rect 28036 42404 28092 42406
rect 28116 42404 28172 42406
rect 28196 42404 28252 42406
rect 27956 41370 28012 41372
rect 28036 41370 28092 41372
rect 28116 41370 28172 41372
rect 28196 41370 28252 41372
rect 27956 41318 28002 41370
rect 28002 41318 28012 41370
rect 28036 41318 28066 41370
rect 28066 41318 28078 41370
rect 28078 41318 28092 41370
rect 28116 41318 28130 41370
rect 28130 41318 28142 41370
rect 28142 41318 28172 41370
rect 28196 41318 28206 41370
rect 28206 41318 28252 41370
rect 27956 41316 28012 41318
rect 28036 41316 28092 41318
rect 28116 41316 28172 41318
rect 28196 41316 28252 41318
rect 27956 40282 28012 40284
rect 28036 40282 28092 40284
rect 28116 40282 28172 40284
rect 28196 40282 28252 40284
rect 27956 40230 28002 40282
rect 28002 40230 28012 40282
rect 28036 40230 28066 40282
rect 28066 40230 28078 40282
rect 28078 40230 28092 40282
rect 28116 40230 28130 40282
rect 28130 40230 28142 40282
rect 28142 40230 28172 40282
rect 28196 40230 28206 40282
rect 28206 40230 28252 40282
rect 27956 40228 28012 40230
rect 28036 40228 28092 40230
rect 28116 40228 28172 40230
rect 28196 40228 28252 40230
rect 27956 39194 28012 39196
rect 28036 39194 28092 39196
rect 28116 39194 28172 39196
rect 28196 39194 28252 39196
rect 27956 39142 28002 39194
rect 28002 39142 28012 39194
rect 28036 39142 28066 39194
rect 28066 39142 28078 39194
rect 28078 39142 28092 39194
rect 28116 39142 28130 39194
rect 28130 39142 28142 39194
rect 28142 39142 28172 39194
rect 28196 39142 28206 39194
rect 28206 39142 28252 39194
rect 27956 39140 28012 39142
rect 28036 39140 28092 39142
rect 28116 39140 28172 39142
rect 28196 39140 28252 39142
rect 27986 38936 28042 38992
rect 27956 38106 28012 38108
rect 28036 38106 28092 38108
rect 28116 38106 28172 38108
rect 28196 38106 28252 38108
rect 27956 38054 28002 38106
rect 28002 38054 28012 38106
rect 28036 38054 28066 38106
rect 28066 38054 28078 38106
rect 28078 38054 28092 38106
rect 28116 38054 28130 38106
rect 28130 38054 28142 38106
rect 28142 38054 28172 38106
rect 28196 38054 28206 38106
rect 28206 38054 28252 38106
rect 27956 38052 28012 38054
rect 28036 38052 28092 38054
rect 28116 38052 28172 38054
rect 28196 38052 28252 38054
rect 27956 37018 28012 37020
rect 28036 37018 28092 37020
rect 28116 37018 28172 37020
rect 28196 37018 28252 37020
rect 27956 36966 28002 37018
rect 28002 36966 28012 37018
rect 28036 36966 28066 37018
rect 28066 36966 28078 37018
rect 28078 36966 28092 37018
rect 28116 36966 28130 37018
rect 28130 36966 28142 37018
rect 28142 36966 28172 37018
rect 28196 36966 28206 37018
rect 28206 36966 28252 37018
rect 27956 36964 28012 36966
rect 28036 36964 28092 36966
rect 28116 36964 28172 36966
rect 28196 36964 28252 36966
rect 27802 36896 27858 36952
rect 28170 36116 28172 36136
rect 28172 36116 28224 36136
rect 28224 36116 28226 36136
rect 28170 36080 28226 36116
rect 27956 35930 28012 35932
rect 28036 35930 28092 35932
rect 28116 35930 28172 35932
rect 28196 35930 28252 35932
rect 27956 35878 28002 35930
rect 28002 35878 28012 35930
rect 28036 35878 28066 35930
rect 28066 35878 28078 35930
rect 28078 35878 28092 35930
rect 28116 35878 28130 35930
rect 28130 35878 28142 35930
rect 28142 35878 28172 35930
rect 28196 35878 28206 35930
rect 28206 35878 28252 35930
rect 27956 35876 28012 35878
rect 28036 35876 28092 35878
rect 28116 35876 28172 35878
rect 28196 35876 28252 35878
rect 27710 35264 27766 35320
rect 26974 33224 27030 33280
rect 26698 32816 26754 32872
rect 26054 30368 26110 30424
rect 25502 24248 25558 24304
rect 25962 22480 26018 22536
rect 26146 24792 26202 24848
rect 26238 23568 26294 23624
rect 27342 33768 27398 33824
rect 27066 27648 27122 27704
rect 27956 34842 28012 34844
rect 28036 34842 28092 34844
rect 28116 34842 28172 34844
rect 28196 34842 28252 34844
rect 27956 34790 28002 34842
rect 28002 34790 28012 34842
rect 28036 34790 28066 34842
rect 28066 34790 28078 34842
rect 28078 34790 28092 34842
rect 28116 34790 28130 34842
rect 28130 34790 28142 34842
rect 28142 34790 28172 34842
rect 28196 34790 28206 34842
rect 28206 34790 28252 34842
rect 27956 34788 28012 34790
rect 28036 34788 28092 34790
rect 28116 34788 28172 34790
rect 28196 34788 28252 34790
rect 27986 33904 28042 33960
rect 27956 33754 28012 33756
rect 28036 33754 28092 33756
rect 28116 33754 28172 33756
rect 28196 33754 28252 33756
rect 27956 33702 28002 33754
rect 28002 33702 28012 33754
rect 28036 33702 28066 33754
rect 28066 33702 28078 33754
rect 28078 33702 28092 33754
rect 28116 33702 28130 33754
rect 28130 33702 28142 33754
rect 28142 33702 28172 33754
rect 28196 33702 28206 33754
rect 28206 33702 28252 33754
rect 27956 33700 28012 33702
rect 28036 33700 28092 33702
rect 28116 33700 28172 33702
rect 28196 33700 28252 33702
rect 27956 32666 28012 32668
rect 28036 32666 28092 32668
rect 28116 32666 28172 32668
rect 28196 32666 28252 32668
rect 27956 32614 28002 32666
rect 28002 32614 28012 32666
rect 28036 32614 28066 32666
rect 28066 32614 28078 32666
rect 28078 32614 28092 32666
rect 28116 32614 28130 32666
rect 28130 32614 28142 32666
rect 28142 32614 28172 32666
rect 28196 32614 28206 32666
rect 28206 32614 28252 32666
rect 27956 32612 28012 32614
rect 28036 32612 28092 32614
rect 28116 32612 28172 32614
rect 28196 32612 28252 32614
rect 26698 24928 26754 24984
rect 27956 31578 28012 31580
rect 28036 31578 28092 31580
rect 28116 31578 28172 31580
rect 28196 31578 28252 31580
rect 27956 31526 28002 31578
rect 28002 31526 28012 31578
rect 28036 31526 28066 31578
rect 28066 31526 28078 31578
rect 28078 31526 28092 31578
rect 28116 31526 28130 31578
rect 28130 31526 28142 31578
rect 28142 31526 28172 31578
rect 28196 31526 28206 31578
rect 28206 31526 28252 31578
rect 27956 31524 28012 31526
rect 28036 31524 28092 31526
rect 28116 31524 28172 31526
rect 28196 31524 28252 31526
rect 27956 30490 28012 30492
rect 28036 30490 28092 30492
rect 28116 30490 28172 30492
rect 28196 30490 28252 30492
rect 27956 30438 28002 30490
rect 28002 30438 28012 30490
rect 28036 30438 28066 30490
rect 28066 30438 28078 30490
rect 28078 30438 28092 30490
rect 28116 30438 28130 30490
rect 28130 30438 28142 30490
rect 28142 30438 28172 30490
rect 28196 30438 28206 30490
rect 28206 30438 28252 30490
rect 27956 30436 28012 30438
rect 28036 30436 28092 30438
rect 28116 30436 28172 30438
rect 28196 30436 28252 30438
rect 28262 30232 28318 30288
rect 27956 29402 28012 29404
rect 28036 29402 28092 29404
rect 28116 29402 28172 29404
rect 28196 29402 28252 29404
rect 27956 29350 28002 29402
rect 28002 29350 28012 29402
rect 28036 29350 28066 29402
rect 28066 29350 28078 29402
rect 28078 29350 28092 29402
rect 28116 29350 28130 29402
rect 28130 29350 28142 29402
rect 28142 29350 28172 29402
rect 28196 29350 28206 29402
rect 28206 29350 28252 29402
rect 27956 29348 28012 29350
rect 28036 29348 28092 29350
rect 28116 29348 28172 29350
rect 28196 29348 28252 29350
rect 27956 28314 28012 28316
rect 28036 28314 28092 28316
rect 28116 28314 28172 28316
rect 28196 28314 28252 28316
rect 27956 28262 28002 28314
rect 28002 28262 28012 28314
rect 28036 28262 28066 28314
rect 28066 28262 28078 28314
rect 28078 28262 28092 28314
rect 28116 28262 28130 28314
rect 28130 28262 28142 28314
rect 28142 28262 28172 28314
rect 28196 28262 28206 28314
rect 28206 28262 28252 28314
rect 27956 28260 28012 28262
rect 28036 28260 28092 28262
rect 28116 28260 28172 28262
rect 28196 28260 28252 28262
rect 27710 28192 27766 28248
rect 27956 27226 28012 27228
rect 28036 27226 28092 27228
rect 28116 27226 28172 27228
rect 28196 27226 28252 27228
rect 27956 27174 28002 27226
rect 28002 27174 28012 27226
rect 28036 27174 28066 27226
rect 28066 27174 28078 27226
rect 28078 27174 28092 27226
rect 28116 27174 28130 27226
rect 28130 27174 28142 27226
rect 28142 27174 28172 27226
rect 28196 27174 28206 27226
rect 28206 27174 28252 27226
rect 27956 27172 28012 27174
rect 28036 27172 28092 27174
rect 28116 27172 28172 27174
rect 28196 27172 28252 27174
rect 28906 34992 28962 35048
rect 28722 32952 28778 33008
rect 28538 32136 28594 32192
rect 27956 26138 28012 26140
rect 28036 26138 28092 26140
rect 28116 26138 28172 26140
rect 28196 26138 28252 26140
rect 27956 26086 28002 26138
rect 28002 26086 28012 26138
rect 28036 26086 28066 26138
rect 28066 26086 28078 26138
rect 28078 26086 28092 26138
rect 28116 26086 28130 26138
rect 28130 26086 28142 26138
rect 28142 26086 28172 26138
rect 28196 26086 28206 26138
rect 28206 26086 28252 26138
rect 27956 26084 28012 26086
rect 28036 26084 28092 26086
rect 28116 26084 28172 26086
rect 28196 26084 28252 26086
rect 27066 19236 27122 19272
rect 27066 19216 27068 19236
rect 27068 19216 27120 19236
rect 27120 19216 27122 19236
rect 27710 24928 27766 24984
rect 27618 24792 27674 24848
rect 27710 24112 27766 24168
rect 27956 25050 28012 25052
rect 28036 25050 28092 25052
rect 28116 25050 28172 25052
rect 28196 25050 28252 25052
rect 27956 24998 28002 25050
rect 28002 24998 28012 25050
rect 28036 24998 28066 25050
rect 28066 24998 28078 25050
rect 28078 24998 28092 25050
rect 28116 24998 28130 25050
rect 28130 24998 28142 25050
rect 28142 24998 28172 25050
rect 28196 24998 28206 25050
rect 28206 24998 28252 25050
rect 27956 24996 28012 24998
rect 28036 24996 28092 24998
rect 28116 24996 28172 24998
rect 28196 24996 28252 24998
rect 28722 32852 28724 32872
rect 28724 32852 28776 32872
rect 28776 32852 28778 32872
rect 28722 32816 28778 32852
rect 28906 32836 28962 32872
rect 28906 32816 28908 32836
rect 28908 32816 28960 32836
rect 28960 32816 28962 32836
rect 28906 30132 28908 30152
rect 28908 30132 28960 30152
rect 28960 30132 28962 30152
rect 28906 30096 28962 30132
rect 27956 23962 28012 23964
rect 28036 23962 28092 23964
rect 28116 23962 28172 23964
rect 28196 23962 28252 23964
rect 27956 23910 28002 23962
rect 28002 23910 28012 23962
rect 28036 23910 28066 23962
rect 28066 23910 28078 23962
rect 28078 23910 28092 23962
rect 28116 23910 28130 23962
rect 28130 23910 28142 23962
rect 28142 23910 28172 23962
rect 28196 23910 28206 23962
rect 28206 23910 28252 23962
rect 27956 23908 28012 23910
rect 28036 23908 28092 23910
rect 28116 23908 28172 23910
rect 28196 23908 28252 23910
rect 28538 23432 28594 23488
rect 29642 37712 29698 37768
rect 29458 36624 29514 36680
rect 28906 25064 28962 25120
rect 28814 24928 28870 24984
rect 28814 24656 28870 24712
rect 29458 27240 29514 27296
rect 27956 22874 28012 22876
rect 28036 22874 28092 22876
rect 28116 22874 28172 22876
rect 28196 22874 28252 22876
rect 27956 22822 28002 22874
rect 28002 22822 28012 22874
rect 28036 22822 28066 22874
rect 28066 22822 28078 22874
rect 28078 22822 28092 22874
rect 28116 22822 28130 22874
rect 28130 22822 28142 22874
rect 28142 22822 28172 22874
rect 28196 22822 28206 22874
rect 28206 22822 28252 22874
rect 27956 22820 28012 22822
rect 28036 22820 28092 22822
rect 28116 22820 28172 22822
rect 28196 22820 28252 22822
rect 27802 22480 27858 22536
rect 27956 21786 28012 21788
rect 28036 21786 28092 21788
rect 28116 21786 28172 21788
rect 28196 21786 28252 21788
rect 27956 21734 28002 21786
rect 28002 21734 28012 21786
rect 28036 21734 28066 21786
rect 28066 21734 28078 21786
rect 28078 21734 28092 21786
rect 28116 21734 28130 21786
rect 28130 21734 28142 21786
rect 28142 21734 28172 21786
rect 28196 21734 28206 21786
rect 28206 21734 28252 21786
rect 27956 21732 28012 21734
rect 28036 21732 28092 21734
rect 28116 21732 28172 21734
rect 28196 21732 28252 21734
rect 27956 20698 28012 20700
rect 28036 20698 28092 20700
rect 28116 20698 28172 20700
rect 28196 20698 28252 20700
rect 27956 20646 28002 20698
rect 28002 20646 28012 20698
rect 28036 20646 28066 20698
rect 28066 20646 28078 20698
rect 28078 20646 28092 20698
rect 28116 20646 28130 20698
rect 28130 20646 28142 20698
rect 28142 20646 28172 20698
rect 28196 20646 28206 20698
rect 28206 20646 28252 20698
rect 27956 20644 28012 20646
rect 28036 20644 28092 20646
rect 28116 20644 28172 20646
rect 28196 20644 28252 20646
rect 27956 19610 28012 19612
rect 28036 19610 28092 19612
rect 28116 19610 28172 19612
rect 28196 19610 28252 19612
rect 27956 19558 28002 19610
rect 28002 19558 28012 19610
rect 28036 19558 28066 19610
rect 28066 19558 28078 19610
rect 28078 19558 28092 19610
rect 28116 19558 28130 19610
rect 28130 19558 28142 19610
rect 28142 19558 28172 19610
rect 28196 19558 28206 19610
rect 28206 19558 28252 19610
rect 27956 19556 28012 19558
rect 28036 19556 28092 19558
rect 28116 19556 28172 19558
rect 28196 19556 28252 19558
rect 27956 18522 28012 18524
rect 28036 18522 28092 18524
rect 28116 18522 28172 18524
rect 28196 18522 28252 18524
rect 27956 18470 28002 18522
rect 28002 18470 28012 18522
rect 28036 18470 28066 18522
rect 28066 18470 28078 18522
rect 28078 18470 28092 18522
rect 28116 18470 28130 18522
rect 28130 18470 28142 18522
rect 28142 18470 28172 18522
rect 28196 18470 28206 18522
rect 28206 18470 28252 18522
rect 27956 18468 28012 18470
rect 28036 18468 28092 18470
rect 28116 18468 28172 18470
rect 28196 18468 28252 18470
rect 27956 17434 28012 17436
rect 28036 17434 28092 17436
rect 28116 17434 28172 17436
rect 28196 17434 28252 17436
rect 27956 17382 28002 17434
rect 28002 17382 28012 17434
rect 28036 17382 28066 17434
rect 28066 17382 28078 17434
rect 28078 17382 28092 17434
rect 28116 17382 28130 17434
rect 28130 17382 28142 17434
rect 28142 17382 28172 17434
rect 28196 17382 28206 17434
rect 28206 17382 28252 17434
rect 27956 17380 28012 17382
rect 28036 17380 28092 17382
rect 28116 17380 28172 17382
rect 28196 17380 28252 17382
rect 27956 16346 28012 16348
rect 28036 16346 28092 16348
rect 28116 16346 28172 16348
rect 28196 16346 28252 16348
rect 27956 16294 28002 16346
rect 28002 16294 28012 16346
rect 28036 16294 28066 16346
rect 28066 16294 28078 16346
rect 28078 16294 28092 16346
rect 28116 16294 28130 16346
rect 28130 16294 28142 16346
rect 28142 16294 28172 16346
rect 28196 16294 28206 16346
rect 28206 16294 28252 16346
rect 27956 16292 28012 16294
rect 28036 16292 28092 16294
rect 28116 16292 28172 16294
rect 28196 16292 28252 16294
rect 27956 15258 28012 15260
rect 28036 15258 28092 15260
rect 28116 15258 28172 15260
rect 28196 15258 28252 15260
rect 27956 15206 28002 15258
rect 28002 15206 28012 15258
rect 28036 15206 28066 15258
rect 28066 15206 28078 15258
rect 28078 15206 28092 15258
rect 28116 15206 28130 15258
rect 28130 15206 28142 15258
rect 28142 15206 28172 15258
rect 28196 15206 28206 15258
rect 28206 15206 28252 15258
rect 27956 15204 28012 15206
rect 28036 15204 28092 15206
rect 28116 15204 28172 15206
rect 28196 15204 28252 15206
rect 27956 14170 28012 14172
rect 28036 14170 28092 14172
rect 28116 14170 28172 14172
rect 28196 14170 28252 14172
rect 27956 14118 28002 14170
rect 28002 14118 28012 14170
rect 28036 14118 28066 14170
rect 28066 14118 28078 14170
rect 28078 14118 28092 14170
rect 28116 14118 28130 14170
rect 28130 14118 28142 14170
rect 28142 14118 28172 14170
rect 28196 14118 28206 14170
rect 28206 14118 28252 14170
rect 27956 14116 28012 14118
rect 28036 14116 28092 14118
rect 28116 14116 28172 14118
rect 28196 14116 28252 14118
rect 27956 13082 28012 13084
rect 28036 13082 28092 13084
rect 28116 13082 28172 13084
rect 28196 13082 28252 13084
rect 27956 13030 28002 13082
rect 28002 13030 28012 13082
rect 28036 13030 28066 13082
rect 28066 13030 28078 13082
rect 28078 13030 28092 13082
rect 28116 13030 28130 13082
rect 28130 13030 28142 13082
rect 28142 13030 28172 13082
rect 28196 13030 28206 13082
rect 28206 13030 28252 13082
rect 27956 13028 28012 13030
rect 28036 13028 28092 13030
rect 28116 13028 28172 13030
rect 28196 13028 28252 13030
rect 28906 23588 28962 23624
rect 28906 23568 28908 23588
rect 28908 23568 28960 23588
rect 28960 23568 28962 23588
rect 28538 21936 28594 21992
rect 28538 19236 28594 19272
rect 28538 19216 28540 19236
rect 28540 19216 28592 19236
rect 28592 19216 28594 19236
rect 27956 11994 28012 11996
rect 28036 11994 28092 11996
rect 28116 11994 28172 11996
rect 28196 11994 28252 11996
rect 27956 11942 28002 11994
rect 28002 11942 28012 11994
rect 28036 11942 28066 11994
rect 28066 11942 28078 11994
rect 28078 11942 28092 11994
rect 28116 11942 28130 11994
rect 28130 11942 28142 11994
rect 28142 11942 28172 11994
rect 28196 11942 28206 11994
rect 28206 11942 28252 11994
rect 27956 11940 28012 11942
rect 28036 11940 28092 11942
rect 28116 11940 28172 11942
rect 28196 11940 28252 11942
rect 27956 10906 28012 10908
rect 28036 10906 28092 10908
rect 28116 10906 28172 10908
rect 28196 10906 28252 10908
rect 27956 10854 28002 10906
rect 28002 10854 28012 10906
rect 28036 10854 28066 10906
rect 28066 10854 28078 10906
rect 28078 10854 28092 10906
rect 28116 10854 28130 10906
rect 28130 10854 28142 10906
rect 28142 10854 28172 10906
rect 28196 10854 28206 10906
rect 28206 10854 28252 10906
rect 27956 10852 28012 10854
rect 28036 10852 28092 10854
rect 28116 10852 28172 10854
rect 28196 10852 28252 10854
rect 27956 9818 28012 9820
rect 28036 9818 28092 9820
rect 28116 9818 28172 9820
rect 28196 9818 28252 9820
rect 27956 9766 28002 9818
rect 28002 9766 28012 9818
rect 28036 9766 28066 9818
rect 28066 9766 28078 9818
rect 28078 9766 28092 9818
rect 28116 9766 28130 9818
rect 28130 9766 28142 9818
rect 28142 9766 28172 9818
rect 28196 9766 28206 9818
rect 28206 9766 28252 9818
rect 27956 9764 28012 9766
rect 28036 9764 28092 9766
rect 28116 9764 28172 9766
rect 28196 9764 28252 9766
rect 27956 8730 28012 8732
rect 28036 8730 28092 8732
rect 28116 8730 28172 8732
rect 28196 8730 28252 8732
rect 27956 8678 28002 8730
rect 28002 8678 28012 8730
rect 28036 8678 28066 8730
rect 28066 8678 28078 8730
rect 28078 8678 28092 8730
rect 28116 8678 28130 8730
rect 28130 8678 28142 8730
rect 28142 8678 28172 8730
rect 28196 8678 28206 8730
rect 28206 8678 28252 8730
rect 27956 8676 28012 8678
rect 28036 8676 28092 8678
rect 28116 8676 28172 8678
rect 28196 8676 28252 8678
rect 27956 7642 28012 7644
rect 28036 7642 28092 7644
rect 28116 7642 28172 7644
rect 28196 7642 28252 7644
rect 27956 7590 28002 7642
rect 28002 7590 28012 7642
rect 28036 7590 28066 7642
rect 28066 7590 28078 7642
rect 28078 7590 28092 7642
rect 28116 7590 28130 7642
rect 28130 7590 28142 7642
rect 28142 7590 28172 7642
rect 28196 7590 28206 7642
rect 28206 7590 28252 7642
rect 27956 7588 28012 7590
rect 28036 7588 28092 7590
rect 28116 7588 28172 7590
rect 28196 7588 28252 7590
rect 27956 6554 28012 6556
rect 28036 6554 28092 6556
rect 28116 6554 28172 6556
rect 28196 6554 28252 6556
rect 27956 6502 28002 6554
rect 28002 6502 28012 6554
rect 28036 6502 28066 6554
rect 28066 6502 28078 6554
rect 28078 6502 28092 6554
rect 28116 6502 28130 6554
rect 28130 6502 28142 6554
rect 28142 6502 28172 6554
rect 28196 6502 28206 6554
rect 28206 6502 28252 6554
rect 27956 6500 28012 6502
rect 28036 6500 28092 6502
rect 28116 6500 28172 6502
rect 28196 6500 28252 6502
rect 27956 5466 28012 5468
rect 28036 5466 28092 5468
rect 28116 5466 28172 5468
rect 28196 5466 28252 5468
rect 27956 5414 28002 5466
rect 28002 5414 28012 5466
rect 28036 5414 28066 5466
rect 28066 5414 28078 5466
rect 28078 5414 28092 5466
rect 28116 5414 28130 5466
rect 28130 5414 28142 5466
rect 28142 5414 28172 5466
rect 28196 5414 28206 5466
rect 28206 5414 28252 5466
rect 27956 5412 28012 5414
rect 28036 5412 28092 5414
rect 28116 5412 28172 5414
rect 28196 5412 28252 5414
rect 27956 4378 28012 4380
rect 28036 4378 28092 4380
rect 28116 4378 28172 4380
rect 28196 4378 28252 4380
rect 27956 4326 28002 4378
rect 28002 4326 28012 4378
rect 28036 4326 28066 4378
rect 28066 4326 28078 4378
rect 28078 4326 28092 4378
rect 28116 4326 28130 4378
rect 28130 4326 28142 4378
rect 28142 4326 28172 4378
rect 28196 4326 28206 4378
rect 28206 4326 28252 4378
rect 27956 4324 28012 4326
rect 28036 4324 28092 4326
rect 28116 4324 28172 4326
rect 28196 4324 28252 4326
rect 27956 3290 28012 3292
rect 28036 3290 28092 3292
rect 28116 3290 28172 3292
rect 28196 3290 28252 3292
rect 27956 3238 28002 3290
rect 28002 3238 28012 3290
rect 28036 3238 28066 3290
rect 28066 3238 28078 3290
rect 28078 3238 28092 3290
rect 28116 3238 28130 3290
rect 28130 3238 28142 3290
rect 28142 3238 28172 3290
rect 28196 3238 28206 3290
rect 28206 3238 28252 3290
rect 27956 3236 28012 3238
rect 28036 3236 28092 3238
rect 28116 3236 28172 3238
rect 28196 3236 28252 3238
rect 27956 2202 28012 2204
rect 28036 2202 28092 2204
rect 28116 2202 28172 2204
rect 28196 2202 28252 2204
rect 27956 2150 28002 2202
rect 28002 2150 28012 2202
rect 28036 2150 28066 2202
rect 28066 2150 28078 2202
rect 28078 2150 28092 2202
rect 28116 2150 28130 2202
rect 28130 2150 28142 2202
rect 28142 2150 28172 2202
rect 28196 2150 28206 2202
rect 28206 2150 28252 2202
rect 27956 2148 28012 2150
rect 28036 2148 28092 2150
rect 28116 2148 28172 2150
rect 28196 2148 28252 2150
rect 28538 12416 28594 12472
rect 28814 17332 28870 17368
rect 28814 17312 28816 17332
rect 28816 17312 28868 17332
rect 28868 17312 28870 17332
rect 29090 19372 29146 19408
rect 29090 19352 29092 19372
rect 29092 19352 29144 19372
rect 29144 19352 29146 19372
rect 29090 18028 29092 18048
rect 29092 18028 29144 18048
rect 29144 18028 29146 18048
rect 29090 17992 29146 18028
rect 30194 30640 30250 30696
rect 32956 53882 33012 53884
rect 33036 53882 33092 53884
rect 33116 53882 33172 53884
rect 33196 53882 33252 53884
rect 32956 53830 33002 53882
rect 33002 53830 33012 53882
rect 33036 53830 33066 53882
rect 33066 53830 33078 53882
rect 33078 53830 33092 53882
rect 33116 53830 33130 53882
rect 33130 53830 33142 53882
rect 33142 53830 33172 53882
rect 33196 53830 33206 53882
rect 33206 53830 33252 53882
rect 32956 53828 33012 53830
rect 33036 53828 33092 53830
rect 33116 53828 33172 53830
rect 33196 53828 33252 53830
rect 32956 52794 33012 52796
rect 33036 52794 33092 52796
rect 33116 52794 33172 52796
rect 33196 52794 33252 52796
rect 32956 52742 33002 52794
rect 33002 52742 33012 52794
rect 33036 52742 33066 52794
rect 33066 52742 33078 52794
rect 33078 52742 33092 52794
rect 33116 52742 33130 52794
rect 33130 52742 33142 52794
rect 33142 52742 33172 52794
rect 33196 52742 33206 52794
rect 33206 52742 33252 52794
rect 32956 52740 33012 52742
rect 33036 52740 33092 52742
rect 33116 52740 33172 52742
rect 33196 52740 33252 52742
rect 32956 51706 33012 51708
rect 33036 51706 33092 51708
rect 33116 51706 33172 51708
rect 33196 51706 33252 51708
rect 32956 51654 33002 51706
rect 33002 51654 33012 51706
rect 33036 51654 33066 51706
rect 33066 51654 33078 51706
rect 33078 51654 33092 51706
rect 33116 51654 33130 51706
rect 33130 51654 33142 51706
rect 33142 51654 33172 51706
rect 33196 51654 33206 51706
rect 33206 51654 33252 51706
rect 32956 51652 33012 51654
rect 33036 51652 33092 51654
rect 33116 51652 33172 51654
rect 33196 51652 33252 51654
rect 32956 50618 33012 50620
rect 33036 50618 33092 50620
rect 33116 50618 33172 50620
rect 33196 50618 33252 50620
rect 32956 50566 33002 50618
rect 33002 50566 33012 50618
rect 33036 50566 33066 50618
rect 33066 50566 33078 50618
rect 33078 50566 33092 50618
rect 33116 50566 33130 50618
rect 33130 50566 33142 50618
rect 33142 50566 33172 50618
rect 33196 50566 33206 50618
rect 33206 50566 33252 50618
rect 32956 50564 33012 50566
rect 33036 50564 33092 50566
rect 33116 50564 33172 50566
rect 33196 50564 33252 50566
rect 32956 49530 33012 49532
rect 33036 49530 33092 49532
rect 33116 49530 33172 49532
rect 33196 49530 33252 49532
rect 32956 49478 33002 49530
rect 33002 49478 33012 49530
rect 33036 49478 33066 49530
rect 33066 49478 33078 49530
rect 33078 49478 33092 49530
rect 33116 49478 33130 49530
rect 33130 49478 33142 49530
rect 33142 49478 33172 49530
rect 33196 49478 33206 49530
rect 33206 49478 33252 49530
rect 32956 49476 33012 49478
rect 33036 49476 33092 49478
rect 33116 49476 33172 49478
rect 33196 49476 33252 49478
rect 32956 48442 33012 48444
rect 33036 48442 33092 48444
rect 33116 48442 33172 48444
rect 33196 48442 33252 48444
rect 32956 48390 33002 48442
rect 33002 48390 33012 48442
rect 33036 48390 33066 48442
rect 33066 48390 33078 48442
rect 33078 48390 33092 48442
rect 33116 48390 33130 48442
rect 33130 48390 33142 48442
rect 33142 48390 33172 48442
rect 33196 48390 33206 48442
rect 33206 48390 33252 48442
rect 32956 48388 33012 48390
rect 33036 48388 33092 48390
rect 33116 48388 33172 48390
rect 33196 48388 33252 48390
rect 32956 47354 33012 47356
rect 33036 47354 33092 47356
rect 33116 47354 33172 47356
rect 33196 47354 33252 47356
rect 32956 47302 33002 47354
rect 33002 47302 33012 47354
rect 33036 47302 33066 47354
rect 33066 47302 33078 47354
rect 33078 47302 33092 47354
rect 33116 47302 33130 47354
rect 33130 47302 33142 47354
rect 33142 47302 33172 47354
rect 33196 47302 33206 47354
rect 33206 47302 33252 47354
rect 32956 47300 33012 47302
rect 33036 47300 33092 47302
rect 33116 47300 33172 47302
rect 33196 47300 33252 47302
rect 32956 46266 33012 46268
rect 33036 46266 33092 46268
rect 33116 46266 33172 46268
rect 33196 46266 33252 46268
rect 32956 46214 33002 46266
rect 33002 46214 33012 46266
rect 33036 46214 33066 46266
rect 33066 46214 33078 46266
rect 33078 46214 33092 46266
rect 33116 46214 33130 46266
rect 33130 46214 33142 46266
rect 33142 46214 33172 46266
rect 33196 46214 33206 46266
rect 33206 46214 33252 46266
rect 32956 46212 33012 46214
rect 33036 46212 33092 46214
rect 33116 46212 33172 46214
rect 33196 46212 33252 46214
rect 30746 40024 30802 40080
rect 31022 36624 31078 36680
rect 30654 30096 30710 30152
rect 31574 34040 31630 34096
rect 32956 45178 33012 45180
rect 33036 45178 33092 45180
rect 33116 45178 33172 45180
rect 33196 45178 33252 45180
rect 32956 45126 33002 45178
rect 33002 45126 33012 45178
rect 33036 45126 33066 45178
rect 33066 45126 33078 45178
rect 33078 45126 33092 45178
rect 33116 45126 33130 45178
rect 33130 45126 33142 45178
rect 33142 45126 33172 45178
rect 33196 45126 33206 45178
rect 33206 45126 33252 45178
rect 32956 45124 33012 45126
rect 33036 45124 33092 45126
rect 33116 45124 33172 45126
rect 33196 45124 33252 45126
rect 32956 44090 33012 44092
rect 33036 44090 33092 44092
rect 33116 44090 33172 44092
rect 33196 44090 33252 44092
rect 32956 44038 33002 44090
rect 33002 44038 33012 44090
rect 33036 44038 33066 44090
rect 33066 44038 33078 44090
rect 33078 44038 33092 44090
rect 33116 44038 33130 44090
rect 33130 44038 33142 44090
rect 33142 44038 33172 44090
rect 33196 44038 33206 44090
rect 33206 44038 33252 44090
rect 32956 44036 33012 44038
rect 33036 44036 33092 44038
rect 33116 44036 33172 44038
rect 33196 44036 33252 44038
rect 32956 43002 33012 43004
rect 33036 43002 33092 43004
rect 33116 43002 33172 43004
rect 33196 43002 33252 43004
rect 32956 42950 33002 43002
rect 33002 42950 33012 43002
rect 33036 42950 33066 43002
rect 33066 42950 33078 43002
rect 33078 42950 33092 43002
rect 33116 42950 33130 43002
rect 33130 42950 33142 43002
rect 33142 42950 33172 43002
rect 33196 42950 33206 43002
rect 33206 42950 33252 43002
rect 32956 42948 33012 42950
rect 33036 42948 33092 42950
rect 33116 42948 33172 42950
rect 33196 42948 33252 42950
rect 32956 41914 33012 41916
rect 33036 41914 33092 41916
rect 33116 41914 33172 41916
rect 33196 41914 33252 41916
rect 32956 41862 33002 41914
rect 33002 41862 33012 41914
rect 33036 41862 33066 41914
rect 33066 41862 33078 41914
rect 33078 41862 33092 41914
rect 33116 41862 33130 41914
rect 33130 41862 33142 41914
rect 33142 41862 33172 41914
rect 33196 41862 33206 41914
rect 33206 41862 33252 41914
rect 32956 41860 33012 41862
rect 33036 41860 33092 41862
rect 33116 41860 33172 41862
rect 33196 41860 33252 41862
rect 32956 40826 33012 40828
rect 33036 40826 33092 40828
rect 33116 40826 33172 40828
rect 33196 40826 33252 40828
rect 32956 40774 33002 40826
rect 33002 40774 33012 40826
rect 33036 40774 33066 40826
rect 33066 40774 33078 40826
rect 33078 40774 33092 40826
rect 33116 40774 33130 40826
rect 33130 40774 33142 40826
rect 33142 40774 33172 40826
rect 33196 40774 33206 40826
rect 33206 40774 33252 40826
rect 32956 40772 33012 40774
rect 33036 40772 33092 40774
rect 33116 40772 33172 40774
rect 33196 40772 33252 40774
rect 32494 36216 32550 36272
rect 29918 23432 29974 23488
rect 28814 12552 28870 12608
rect 31206 28056 31262 28112
rect 30930 27240 30986 27296
rect 31298 27004 31300 27024
rect 31300 27004 31352 27024
rect 31352 27004 31354 27024
rect 31022 26288 31078 26344
rect 30378 22652 30380 22672
rect 30380 22652 30432 22672
rect 30432 22652 30434 22672
rect 30378 22616 30434 22652
rect 30470 20596 30526 20632
rect 30470 20576 30472 20596
rect 30472 20576 30524 20596
rect 30524 20576 30526 20596
rect 31298 26968 31354 27004
rect 31574 27376 31630 27432
rect 32956 39738 33012 39740
rect 33036 39738 33092 39740
rect 33116 39738 33172 39740
rect 33196 39738 33252 39740
rect 32956 39686 33002 39738
rect 33002 39686 33012 39738
rect 33036 39686 33066 39738
rect 33066 39686 33078 39738
rect 33078 39686 33092 39738
rect 33116 39686 33130 39738
rect 33130 39686 33142 39738
rect 33142 39686 33172 39738
rect 33196 39686 33206 39738
rect 33206 39686 33252 39738
rect 32956 39684 33012 39686
rect 33036 39684 33092 39686
rect 33116 39684 33172 39686
rect 33196 39684 33252 39686
rect 32956 38650 33012 38652
rect 33036 38650 33092 38652
rect 33116 38650 33172 38652
rect 33196 38650 33252 38652
rect 32956 38598 33002 38650
rect 33002 38598 33012 38650
rect 33036 38598 33066 38650
rect 33066 38598 33078 38650
rect 33078 38598 33092 38650
rect 33116 38598 33130 38650
rect 33130 38598 33142 38650
rect 33142 38598 33172 38650
rect 33196 38598 33206 38650
rect 33206 38598 33252 38650
rect 32956 38596 33012 38598
rect 33036 38596 33092 38598
rect 33116 38596 33172 38598
rect 33196 38596 33252 38598
rect 33230 37712 33286 37768
rect 32956 37562 33012 37564
rect 33036 37562 33092 37564
rect 33116 37562 33172 37564
rect 33196 37562 33252 37564
rect 32956 37510 33002 37562
rect 33002 37510 33012 37562
rect 33036 37510 33066 37562
rect 33066 37510 33078 37562
rect 33078 37510 33092 37562
rect 33116 37510 33130 37562
rect 33130 37510 33142 37562
rect 33142 37510 33172 37562
rect 33196 37510 33206 37562
rect 33206 37510 33252 37562
rect 32956 37508 33012 37510
rect 33036 37508 33092 37510
rect 33116 37508 33172 37510
rect 33196 37508 33252 37510
rect 32956 36474 33012 36476
rect 33036 36474 33092 36476
rect 33116 36474 33172 36476
rect 33196 36474 33252 36476
rect 32956 36422 33002 36474
rect 33002 36422 33012 36474
rect 33036 36422 33066 36474
rect 33066 36422 33078 36474
rect 33078 36422 33092 36474
rect 33116 36422 33130 36474
rect 33130 36422 33142 36474
rect 33142 36422 33172 36474
rect 33196 36422 33206 36474
rect 33206 36422 33252 36474
rect 32956 36420 33012 36422
rect 33036 36420 33092 36422
rect 33116 36420 33172 36422
rect 33196 36420 33252 36422
rect 32770 35572 32772 35592
rect 32772 35572 32824 35592
rect 32824 35572 32826 35592
rect 32770 35536 32826 35572
rect 32956 35386 33012 35388
rect 33036 35386 33092 35388
rect 33116 35386 33172 35388
rect 33196 35386 33252 35388
rect 32956 35334 33002 35386
rect 33002 35334 33012 35386
rect 33036 35334 33066 35386
rect 33066 35334 33078 35386
rect 33078 35334 33092 35386
rect 33116 35334 33130 35386
rect 33130 35334 33142 35386
rect 33142 35334 33172 35386
rect 33196 35334 33206 35386
rect 33206 35334 33252 35386
rect 32956 35332 33012 35334
rect 33036 35332 33092 35334
rect 33116 35332 33172 35334
rect 33196 35332 33252 35334
rect 32956 34298 33012 34300
rect 33036 34298 33092 34300
rect 33116 34298 33172 34300
rect 33196 34298 33252 34300
rect 32956 34246 33002 34298
rect 33002 34246 33012 34298
rect 33036 34246 33066 34298
rect 33066 34246 33078 34298
rect 33078 34246 33092 34298
rect 33116 34246 33130 34298
rect 33130 34246 33142 34298
rect 33142 34246 33172 34298
rect 33196 34246 33206 34298
rect 33206 34246 33252 34298
rect 32956 34244 33012 34246
rect 33036 34244 33092 34246
rect 33116 34244 33172 34246
rect 33196 34244 33252 34246
rect 32956 33210 33012 33212
rect 33036 33210 33092 33212
rect 33116 33210 33172 33212
rect 33196 33210 33252 33212
rect 32956 33158 33002 33210
rect 33002 33158 33012 33210
rect 33036 33158 33066 33210
rect 33066 33158 33078 33210
rect 33078 33158 33092 33210
rect 33116 33158 33130 33210
rect 33130 33158 33142 33210
rect 33142 33158 33172 33210
rect 33196 33158 33206 33210
rect 33206 33158 33252 33210
rect 32956 33156 33012 33158
rect 33036 33156 33092 33158
rect 33116 33156 33172 33158
rect 33196 33156 33252 33158
rect 32956 32122 33012 32124
rect 33036 32122 33092 32124
rect 33116 32122 33172 32124
rect 33196 32122 33252 32124
rect 32956 32070 33002 32122
rect 33002 32070 33012 32122
rect 33036 32070 33066 32122
rect 33066 32070 33078 32122
rect 33078 32070 33092 32122
rect 33116 32070 33130 32122
rect 33130 32070 33142 32122
rect 33142 32070 33172 32122
rect 33196 32070 33206 32122
rect 33206 32070 33252 32122
rect 32956 32068 33012 32070
rect 33036 32068 33092 32070
rect 33116 32068 33172 32070
rect 33196 32068 33252 32070
rect 32126 26288 32182 26344
rect 32956 31034 33012 31036
rect 33036 31034 33092 31036
rect 33116 31034 33172 31036
rect 33196 31034 33252 31036
rect 32956 30982 33002 31034
rect 33002 30982 33012 31034
rect 33036 30982 33066 31034
rect 33066 30982 33078 31034
rect 33078 30982 33092 31034
rect 33116 30982 33130 31034
rect 33130 30982 33142 31034
rect 33142 30982 33172 31034
rect 33196 30982 33206 31034
rect 33206 30982 33252 31034
rect 32956 30980 33012 30982
rect 33036 30980 33092 30982
rect 33116 30980 33172 30982
rect 33196 30980 33252 30982
rect 32956 29946 33012 29948
rect 33036 29946 33092 29948
rect 33116 29946 33172 29948
rect 33196 29946 33252 29948
rect 32956 29894 33002 29946
rect 33002 29894 33012 29946
rect 33036 29894 33066 29946
rect 33066 29894 33078 29946
rect 33078 29894 33092 29946
rect 33116 29894 33130 29946
rect 33130 29894 33142 29946
rect 33142 29894 33172 29946
rect 33196 29894 33206 29946
rect 33206 29894 33252 29946
rect 32956 29892 33012 29894
rect 33036 29892 33092 29894
rect 33116 29892 33172 29894
rect 33196 29892 33252 29894
rect 32956 28858 33012 28860
rect 33036 28858 33092 28860
rect 33116 28858 33172 28860
rect 33196 28858 33252 28860
rect 32956 28806 33002 28858
rect 33002 28806 33012 28858
rect 33036 28806 33066 28858
rect 33066 28806 33078 28858
rect 33078 28806 33092 28858
rect 33116 28806 33130 28858
rect 33130 28806 33142 28858
rect 33142 28806 33172 28858
rect 33196 28806 33206 28858
rect 33206 28806 33252 28858
rect 32956 28804 33012 28806
rect 33036 28804 33092 28806
rect 33116 28804 33172 28806
rect 33196 28804 33252 28806
rect 33966 40452 34022 40488
rect 33966 40432 33968 40452
rect 33968 40432 34020 40452
rect 34020 40432 34022 40452
rect 32956 27770 33012 27772
rect 33036 27770 33092 27772
rect 33116 27770 33172 27772
rect 33196 27770 33252 27772
rect 32956 27718 33002 27770
rect 33002 27718 33012 27770
rect 33036 27718 33066 27770
rect 33066 27718 33078 27770
rect 33078 27718 33092 27770
rect 33116 27718 33130 27770
rect 33130 27718 33142 27770
rect 33142 27718 33172 27770
rect 33196 27718 33206 27770
rect 33206 27718 33252 27770
rect 32956 27716 33012 27718
rect 33036 27716 33092 27718
rect 33116 27716 33172 27718
rect 33196 27716 33252 27718
rect 32956 26682 33012 26684
rect 33036 26682 33092 26684
rect 33116 26682 33172 26684
rect 33196 26682 33252 26684
rect 32956 26630 33002 26682
rect 33002 26630 33012 26682
rect 33036 26630 33066 26682
rect 33066 26630 33078 26682
rect 33078 26630 33092 26682
rect 33116 26630 33130 26682
rect 33130 26630 33142 26682
rect 33142 26630 33172 26682
rect 33196 26630 33206 26682
rect 33206 26630 33252 26682
rect 32956 26628 33012 26630
rect 33036 26628 33092 26630
rect 33116 26628 33172 26630
rect 33196 26628 33252 26630
rect 32678 25336 32734 25392
rect 32956 25594 33012 25596
rect 33036 25594 33092 25596
rect 33116 25594 33172 25596
rect 33196 25594 33252 25596
rect 32956 25542 33002 25594
rect 33002 25542 33012 25594
rect 33036 25542 33066 25594
rect 33066 25542 33078 25594
rect 33078 25542 33092 25594
rect 33116 25542 33130 25594
rect 33130 25542 33142 25594
rect 33142 25542 33172 25594
rect 33196 25542 33206 25594
rect 33206 25542 33252 25594
rect 32956 25540 33012 25542
rect 33036 25540 33092 25542
rect 33116 25540 33172 25542
rect 33196 25540 33252 25542
rect 32956 24506 33012 24508
rect 33036 24506 33092 24508
rect 33116 24506 33172 24508
rect 33196 24506 33252 24508
rect 32956 24454 33002 24506
rect 33002 24454 33012 24506
rect 33036 24454 33066 24506
rect 33066 24454 33078 24506
rect 33078 24454 33092 24506
rect 33116 24454 33130 24506
rect 33130 24454 33142 24506
rect 33142 24454 33172 24506
rect 33196 24454 33206 24506
rect 33206 24454 33252 24506
rect 32956 24452 33012 24454
rect 33036 24452 33092 24454
rect 33116 24452 33172 24454
rect 33196 24452 33252 24454
rect 32956 23418 33012 23420
rect 33036 23418 33092 23420
rect 33116 23418 33172 23420
rect 33196 23418 33252 23420
rect 32956 23366 33002 23418
rect 33002 23366 33012 23418
rect 33036 23366 33066 23418
rect 33066 23366 33078 23418
rect 33078 23366 33092 23418
rect 33116 23366 33130 23418
rect 33130 23366 33142 23418
rect 33142 23366 33172 23418
rect 33196 23366 33206 23418
rect 33206 23366 33252 23418
rect 32956 23364 33012 23366
rect 33036 23364 33092 23366
rect 33116 23364 33172 23366
rect 33196 23364 33252 23366
rect 32956 22330 33012 22332
rect 33036 22330 33092 22332
rect 33116 22330 33172 22332
rect 33196 22330 33252 22332
rect 32956 22278 33002 22330
rect 33002 22278 33012 22330
rect 33036 22278 33066 22330
rect 33066 22278 33078 22330
rect 33078 22278 33092 22330
rect 33116 22278 33130 22330
rect 33130 22278 33142 22330
rect 33142 22278 33172 22330
rect 33196 22278 33206 22330
rect 33206 22278 33252 22330
rect 32956 22276 33012 22278
rect 33036 22276 33092 22278
rect 33116 22276 33172 22278
rect 33196 22276 33252 22278
rect 33690 36352 33746 36408
rect 33598 31340 33654 31376
rect 33598 31320 33600 31340
rect 33600 31320 33652 31340
rect 33652 31320 33654 31340
rect 33690 29028 33746 29064
rect 33690 29008 33692 29028
rect 33692 29008 33744 29028
rect 33744 29008 33746 29028
rect 34518 30232 34574 30288
rect 32956 21242 33012 21244
rect 33036 21242 33092 21244
rect 33116 21242 33172 21244
rect 33196 21242 33252 21244
rect 32956 21190 33002 21242
rect 33002 21190 33012 21242
rect 33036 21190 33066 21242
rect 33066 21190 33078 21242
rect 33078 21190 33092 21242
rect 33116 21190 33130 21242
rect 33130 21190 33142 21242
rect 33142 21190 33172 21242
rect 33196 21190 33206 21242
rect 33206 21190 33252 21242
rect 32956 21188 33012 21190
rect 33036 21188 33092 21190
rect 33116 21188 33172 21190
rect 33196 21188 33252 21190
rect 32956 20154 33012 20156
rect 33036 20154 33092 20156
rect 33116 20154 33172 20156
rect 33196 20154 33252 20156
rect 32956 20102 33002 20154
rect 33002 20102 33012 20154
rect 33036 20102 33066 20154
rect 33066 20102 33078 20154
rect 33078 20102 33092 20154
rect 33116 20102 33130 20154
rect 33130 20102 33142 20154
rect 33142 20102 33172 20154
rect 33196 20102 33206 20154
rect 33206 20102 33252 20154
rect 32956 20100 33012 20102
rect 33036 20100 33092 20102
rect 33116 20100 33172 20102
rect 33196 20100 33252 20102
rect 34610 26968 34666 27024
rect 35990 39516 35992 39536
rect 35992 39516 36044 39536
rect 36044 39516 36046 39536
rect 35990 39480 36046 39516
rect 35898 38664 35954 38720
rect 36174 35672 36230 35728
rect 36082 35148 36138 35184
rect 36082 35128 36084 35148
rect 36084 35128 36136 35148
rect 36136 35128 36138 35148
rect 35346 28364 35348 28384
rect 35348 28364 35400 28384
rect 35400 28364 35402 28384
rect 35346 28328 35402 28364
rect 34978 27376 35034 27432
rect 32956 19066 33012 19068
rect 33036 19066 33092 19068
rect 33116 19066 33172 19068
rect 33196 19066 33252 19068
rect 32956 19014 33002 19066
rect 33002 19014 33012 19066
rect 33036 19014 33066 19066
rect 33066 19014 33078 19066
rect 33078 19014 33092 19066
rect 33116 19014 33130 19066
rect 33130 19014 33142 19066
rect 33142 19014 33172 19066
rect 33196 19014 33206 19066
rect 33206 19014 33252 19066
rect 32956 19012 33012 19014
rect 33036 19012 33092 19014
rect 33116 19012 33172 19014
rect 33196 19012 33252 19014
rect 32956 17978 33012 17980
rect 33036 17978 33092 17980
rect 33116 17978 33172 17980
rect 33196 17978 33252 17980
rect 32956 17926 33002 17978
rect 33002 17926 33012 17978
rect 33036 17926 33066 17978
rect 33066 17926 33078 17978
rect 33078 17926 33092 17978
rect 33116 17926 33130 17978
rect 33130 17926 33142 17978
rect 33142 17926 33172 17978
rect 33196 17926 33206 17978
rect 33206 17926 33252 17978
rect 32956 17924 33012 17926
rect 33036 17924 33092 17926
rect 33116 17924 33172 17926
rect 33196 17924 33252 17926
rect 32956 16890 33012 16892
rect 33036 16890 33092 16892
rect 33116 16890 33172 16892
rect 33196 16890 33252 16892
rect 32956 16838 33002 16890
rect 33002 16838 33012 16890
rect 33036 16838 33066 16890
rect 33066 16838 33078 16890
rect 33078 16838 33092 16890
rect 33116 16838 33130 16890
rect 33130 16838 33142 16890
rect 33142 16838 33172 16890
rect 33196 16838 33206 16890
rect 33206 16838 33252 16890
rect 32956 16836 33012 16838
rect 33036 16836 33092 16838
rect 33116 16836 33172 16838
rect 33196 16836 33252 16838
rect 32956 15802 33012 15804
rect 33036 15802 33092 15804
rect 33116 15802 33172 15804
rect 33196 15802 33252 15804
rect 32956 15750 33002 15802
rect 33002 15750 33012 15802
rect 33036 15750 33066 15802
rect 33066 15750 33078 15802
rect 33078 15750 33092 15802
rect 33116 15750 33130 15802
rect 33130 15750 33142 15802
rect 33142 15750 33172 15802
rect 33196 15750 33206 15802
rect 33206 15750 33252 15802
rect 32956 15748 33012 15750
rect 33036 15748 33092 15750
rect 33116 15748 33172 15750
rect 33196 15748 33252 15750
rect 32956 14714 33012 14716
rect 33036 14714 33092 14716
rect 33116 14714 33172 14716
rect 33196 14714 33252 14716
rect 32956 14662 33002 14714
rect 33002 14662 33012 14714
rect 33036 14662 33066 14714
rect 33066 14662 33078 14714
rect 33078 14662 33092 14714
rect 33116 14662 33130 14714
rect 33130 14662 33142 14714
rect 33142 14662 33172 14714
rect 33196 14662 33206 14714
rect 33206 14662 33252 14714
rect 32956 14660 33012 14662
rect 33036 14660 33092 14662
rect 33116 14660 33172 14662
rect 33196 14660 33252 14662
rect 32956 13626 33012 13628
rect 33036 13626 33092 13628
rect 33116 13626 33172 13628
rect 33196 13626 33252 13628
rect 32956 13574 33002 13626
rect 33002 13574 33012 13626
rect 33036 13574 33066 13626
rect 33066 13574 33078 13626
rect 33078 13574 33092 13626
rect 33116 13574 33130 13626
rect 33130 13574 33142 13626
rect 33142 13574 33172 13626
rect 33196 13574 33206 13626
rect 33206 13574 33252 13626
rect 32956 13572 33012 13574
rect 33036 13572 33092 13574
rect 33116 13572 33172 13574
rect 33196 13572 33252 13574
rect 34058 16652 34114 16688
rect 34058 16632 34060 16652
rect 34060 16632 34112 16652
rect 34112 16632 34114 16652
rect 32956 12538 33012 12540
rect 33036 12538 33092 12540
rect 33116 12538 33172 12540
rect 33196 12538 33252 12540
rect 32956 12486 33002 12538
rect 33002 12486 33012 12538
rect 33036 12486 33066 12538
rect 33066 12486 33078 12538
rect 33078 12486 33092 12538
rect 33116 12486 33130 12538
rect 33130 12486 33142 12538
rect 33142 12486 33172 12538
rect 33196 12486 33206 12538
rect 33206 12486 33252 12538
rect 32956 12484 33012 12486
rect 33036 12484 33092 12486
rect 33116 12484 33172 12486
rect 33196 12484 33252 12486
rect 32956 11450 33012 11452
rect 33036 11450 33092 11452
rect 33116 11450 33172 11452
rect 33196 11450 33252 11452
rect 32956 11398 33002 11450
rect 33002 11398 33012 11450
rect 33036 11398 33066 11450
rect 33066 11398 33078 11450
rect 33078 11398 33092 11450
rect 33116 11398 33130 11450
rect 33130 11398 33142 11450
rect 33142 11398 33172 11450
rect 33196 11398 33206 11450
rect 33206 11398 33252 11450
rect 32956 11396 33012 11398
rect 33036 11396 33092 11398
rect 33116 11396 33172 11398
rect 33196 11396 33252 11398
rect 32956 10362 33012 10364
rect 33036 10362 33092 10364
rect 33116 10362 33172 10364
rect 33196 10362 33252 10364
rect 32956 10310 33002 10362
rect 33002 10310 33012 10362
rect 33036 10310 33066 10362
rect 33066 10310 33078 10362
rect 33078 10310 33092 10362
rect 33116 10310 33130 10362
rect 33130 10310 33142 10362
rect 33142 10310 33172 10362
rect 33196 10310 33206 10362
rect 33206 10310 33252 10362
rect 32956 10308 33012 10310
rect 33036 10308 33092 10310
rect 33116 10308 33172 10310
rect 33196 10308 33252 10310
rect 32956 9274 33012 9276
rect 33036 9274 33092 9276
rect 33116 9274 33172 9276
rect 33196 9274 33252 9276
rect 32956 9222 33002 9274
rect 33002 9222 33012 9274
rect 33036 9222 33066 9274
rect 33066 9222 33078 9274
rect 33078 9222 33092 9274
rect 33116 9222 33130 9274
rect 33130 9222 33142 9274
rect 33142 9222 33172 9274
rect 33196 9222 33206 9274
rect 33206 9222 33252 9274
rect 32956 9220 33012 9222
rect 33036 9220 33092 9222
rect 33116 9220 33172 9222
rect 33196 9220 33252 9222
rect 32956 8186 33012 8188
rect 33036 8186 33092 8188
rect 33116 8186 33172 8188
rect 33196 8186 33252 8188
rect 32956 8134 33002 8186
rect 33002 8134 33012 8186
rect 33036 8134 33066 8186
rect 33066 8134 33078 8186
rect 33078 8134 33092 8186
rect 33116 8134 33130 8186
rect 33130 8134 33142 8186
rect 33142 8134 33172 8186
rect 33196 8134 33206 8186
rect 33206 8134 33252 8186
rect 32956 8132 33012 8134
rect 33036 8132 33092 8134
rect 33116 8132 33172 8134
rect 33196 8132 33252 8134
rect 32956 7098 33012 7100
rect 33036 7098 33092 7100
rect 33116 7098 33172 7100
rect 33196 7098 33252 7100
rect 32956 7046 33002 7098
rect 33002 7046 33012 7098
rect 33036 7046 33066 7098
rect 33066 7046 33078 7098
rect 33078 7046 33092 7098
rect 33116 7046 33130 7098
rect 33130 7046 33142 7098
rect 33142 7046 33172 7098
rect 33196 7046 33206 7098
rect 33206 7046 33252 7098
rect 32956 7044 33012 7046
rect 33036 7044 33092 7046
rect 33116 7044 33172 7046
rect 33196 7044 33252 7046
rect 32956 6010 33012 6012
rect 33036 6010 33092 6012
rect 33116 6010 33172 6012
rect 33196 6010 33252 6012
rect 32956 5958 33002 6010
rect 33002 5958 33012 6010
rect 33036 5958 33066 6010
rect 33066 5958 33078 6010
rect 33078 5958 33092 6010
rect 33116 5958 33130 6010
rect 33130 5958 33142 6010
rect 33142 5958 33172 6010
rect 33196 5958 33206 6010
rect 33206 5958 33252 6010
rect 32956 5956 33012 5958
rect 33036 5956 33092 5958
rect 33116 5956 33172 5958
rect 33196 5956 33252 5958
rect 32956 4922 33012 4924
rect 33036 4922 33092 4924
rect 33116 4922 33172 4924
rect 33196 4922 33252 4924
rect 32956 4870 33002 4922
rect 33002 4870 33012 4922
rect 33036 4870 33066 4922
rect 33066 4870 33078 4922
rect 33078 4870 33092 4922
rect 33116 4870 33130 4922
rect 33130 4870 33142 4922
rect 33142 4870 33172 4922
rect 33196 4870 33206 4922
rect 33206 4870 33252 4922
rect 32956 4868 33012 4870
rect 33036 4868 33092 4870
rect 33116 4868 33172 4870
rect 33196 4868 33252 4870
rect 32956 3834 33012 3836
rect 33036 3834 33092 3836
rect 33116 3834 33172 3836
rect 33196 3834 33252 3836
rect 32956 3782 33002 3834
rect 33002 3782 33012 3834
rect 33036 3782 33066 3834
rect 33066 3782 33078 3834
rect 33078 3782 33092 3834
rect 33116 3782 33130 3834
rect 33130 3782 33142 3834
rect 33142 3782 33172 3834
rect 33196 3782 33206 3834
rect 33206 3782 33252 3834
rect 32956 3780 33012 3782
rect 33036 3780 33092 3782
rect 33116 3780 33172 3782
rect 33196 3780 33252 3782
rect 32956 2746 33012 2748
rect 33036 2746 33092 2748
rect 33116 2746 33172 2748
rect 33196 2746 33252 2748
rect 32956 2694 33002 2746
rect 33002 2694 33012 2746
rect 33036 2694 33066 2746
rect 33066 2694 33078 2746
rect 33078 2694 33092 2746
rect 33116 2694 33130 2746
rect 33130 2694 33142 2746
rect 33142 2694 33172 2746
rect 33196 2694 33206 2746
rect 33206 2694 33252 2746
rect 32956 2692 33012 2694
rect 33036 2692 33092 2694
rect 33116 2692 33172 2694
rect 33196 2692 33252 2694
rect 37956 54426 38012 54428
rect 38036 54426 38092 54428
rect 38116 54426 38172 54428
rect 38196 54426 38252 54428
rect 37956 54374 38002 54426
rect 38002 54374 38012 54426
rect 38036 54374 38066 54426
rect 38066 54374 38078 54426
rect 38078 54374 38092 54426
rect 38116 54374 38130 54426
rect 38130 54374 38142 54426
rect 38142 54374 38172 54426
rect 38196 54374 38206 54426
rect 38206 54374 38252 54426
rect 37956 54372 38012 54374
rect 38036 54372 38092 54374
rect 38116 54372 38172 54374
rect 38196 54372 38252 54374
rect 37956 53338 38012 53340
rect 38036 53338 38092 53340
rect 38116 53338 38172 53340
rect 38196 53338 38252 53340
rect 37956 53286 38002 53338
rect 38002 53286 38012 53338
rect 38036 53286 38066 53338
rect 38066 53286 38078 53338
rect 38078 53286 38092 53338
rect 38116 53286 38130 53338
rect 38130 53286 38142 53338
rect 38142 53286 38172 53338
rect 38196 53286 38206 53338
rect 38206 53286 38252 53338
rect 37956 53284 38012 53286
rect 38036 53284 38092 53286
rect 38116 53284 38172 53286
rect 38196 53284 38252 53286
rect 37956 52250 38012 52252
rect 38036 52250 38092 52252
rect 38116 52250 38172 52252
rect 38196 52250 38252 52252
rect 37956 52198 38002 52250
rect 38002 52198 38012 52250
rect 38036 52198 38066 52250
rect 38066 52198 38078 52250
rect 38078 52198 38092 52250
rect 38116 52198 38130 52250
rect 38130 52198 38142 52250
rect 38142 52198 38172 52250
rect 38196 52198 38206 52250
rect 38206 52198 38252 52250
rect 37956 52196 38012 52198
rect 38036 52196 38092 52198
rect 38116 52196 38172 52198
rect 38196 52196 38252 52198
rect 37956 51162 38012 51164
rect 38036 51162 38092 51164
rect 38116 51162 38172 51164
rect 38196 51162 38252 51164
rect 37956 51110 38002 51162
rect 38002 51110 38012 51162
rect 38036 51110 38066 51162
rect 38066 51110 38078 51162
rect 38078 51110 38092 51162
rect 38116 51110 38130 51162
rect 38130 51110 38142 51162
rect 38142 51110 38172 51162
rect 38196 51110 38206 51162
rect 38206 51110 38252 51162
rect 37956 51108 38012 51110
rect 38036 51108 38092 51110
rect 38116 51108 38172 51110
rect 38196 51108 38252 51110
rect 37956 50074 38012 50076
rect 38036 50074 38092 50076
rect 38116 50074 38172 50076
rect 38196 50074 38252 50076
rect 37956 50022 38002 50074
rect 38002 50022 38012 50074
rect 38036 50022 38066 50074
rect 38066 50022 38078 50074
rect 38078 50022 38092 50074
rect 38116 50022 38130 50074
rect 38130 50022 38142 50074
rect 38142 50022 38172 50074
rect 38196 50022 38206 50074
rect 38206 50022 38252 50074
rect 37956 50020 38012 50022
rect 38036 50020 38092 50022
rect 38116 50020 38172 50022
rect 38196 50020 38252 50022
rect 37956 48986 38012 48988
rect 38036 48986 38092 48988
rect 38116 48986 38172 48988
rect 38196 48986 38252 48988
rect 37956 48934 38002 48986
rect 38002 48934 38012 48986
rect 38036 48934 38066 48986
rect 38066 48934 38078 48986
rect 38078 48934 38092 48986
rect 38116 48934 38130 48986
rect 38130 48934 38142 48986
rect 38142 48934 38172 48986
rect 38196 48934 38206 48986
rect 38206 48934 38252 48986
rect 37956 48932 38012 48934
rect 38036 48932 38092 48934
rect 38116 48932 38172 48934
rect 38196 48932 38252 48934
rect 37956 47898 38012 47900
rect 38036 47898 38092 47900
rect 38116 47898 38172 47900
rect 38196 47898 38252 47900
rect 37956 47846 38002 47898
rect 38002 47846 38012 47898
rect 38036 47846 38066 47898
rect 38066 47846 38078 47898
rect 38078 47846 38092 47898
rect 38116 47846 38130 47898
rect 38130 47846 38142 47898
rect 38142 47846 38172 47898
rect 38196 47846 38206 47898
rect 38206 47846 38252 47898
rect 37956 47844 38012 47846
rect 38036 47844 38092 47846
rect 38116 47844 38172 47846
rect 38196 47844 38252 47846
rect 37956 46810 38012 46812
rect 38036 46810 38092 46812
rect 38116 46810 38172 46812
rect 38196 46810 38252 46812
rect 37956 46758 38002 46810
rect 38002 46758 38012 46810
rect 38036 46758 38066 46810
rect 38066 46758 38078 46810
rect 38078 46758 38092 46810
rect 38116 46758 38130 46810
rect 38130 46758 38142 46810
rect 38142 46758 38172 46810
rect 38196 46758 38206 46810
rect 38206 46758 38252 46810
rect 37956 46756 38012 46758
rect 38036 46756 38092 46758
rect 38116 46756 38172 46758
rect 38196 46756 38252 46758
rect 37956 45722 38012 45724
rect 38036 45722 38092 45724
rect 38116 45722 38172 45724
rect 38196 45722 38252 45724
rect 37956 45670 38002 45722
rect 38002 45670 38012 45722
rect 38036 45670 38066 45722
rect 38066 45670 38078 45722
rect 38078 45670 38092 45722
rect 38116 45670 38130 45722
rect 38130 45670 38142 45722
rect 38142 45670 38172 45722
rect 38196 45670 38206 45722
rect 38206 45670 38252 45722
rect 37956 45668 38012 45670
rect 38036 45668 38092 45670
rect 38116 45668 38172 45670
rect 38196 45668 38252 45670
rect 37956 44634 38012 44636
rect 38036 44634 38092 44636
rect 38116 44634 38172 44636
rect 38196 44634 38252 44636
rect 37956 44582 38002 44634
rect 38002 44582 38012 44634
rect 38036 44582 38066 44634
rect 38066 44582 38078 44634
rect 38078 44582 38092 44634
rect 38116 44582 38130 44634
rect 38130 44582 38142 44634
rect 38142 44582 38172 44634
rect 38196 44582 38206 44634
rect 38206 44582 38252 44634
rect 37956 44580 38012 44582
rect 38036 44580 38092 44582
rect 38116 44580 38172 44582
rect 38196 44580 38252 44582
rect 36726 39480 36782 39536
rect 36542 34040 36598 34096
rect 35990 31456 36046 31512
rect 37956 43546 38012 43548
rect 38036 43546 38092 43548
rect 38116 43546 38172 43548
rect 38196 43546 38252 43548
rect 37956 43494 38002 43546
rect 38002 43494 38012 43546
rect 38036 43494 38066 43546
rect 38066 43494 38078 43546
rect 38078 43494 38092 43546
rect 38116 43494 38130 43546
rect 38130 43494 38142 43546
rect 38142 43494 38172 43546
rect 38196 43494 38206 43546
rect 38206 43494 38252 43546
rect 37956 43492 38012 43494
rect 38036 43492 38092 43494
rect 38116 43492 38172 43494
rect 38196 43492 38252 43494
rect 37956 42458 38012 42460
rect 38036 42458 38092 42460
rect 38116 42458 38172 42460
rect 38196 42458 38252 42460
rect 37956 42406 38002 42458
rect 38002 42406 38012 42458
rect 38036 42406 38066 42458
rect 38066 42406 38078 42458
rect 38078 42406 38092 42458
rect 38116 42406 38130 42458
rect 38130 42406 38142 42458
rect 38142 42406 38172 42458
rect 38196 42406 38206 42458
rect 38206 42406 38252 42458
rect 37956 42404 38012 42406
rect 38036 42404 38092 42406
rect 38116 42404 38172 42406
rect 38196 42404 38252 42406
rect 37956 41370 38012 41372
rect 38036 41370 38092 41372
rect 38116 41370 38172 41372
rect 38196 41370 38252 41372
rect 37956 41318 38002 41370
rect 38002 41318 38012 41370
rect 38036 41318 38066 41370
rect 38066 41318 38078 41370
rect 38078 41318 38092 41370
rect 38116 41318 38130 41370
rect 38130 41318 38142 41370
rect 38142 41318 38172 41370
rect 38196 41318 38206 41370
rect 38206 41318 38252 41370
rect 37956 41316 38012 41318
rect 38036 41316 38092 41318
rect 38116 41316 38172 41318
rect 38196 41316 38252 41318
rect 37094 33904 37150 33960
rect 37956 40282 38012 40284
rect 38036 40282 38092 40284
rect 38116 40282 38172 40284
rect 38196 40282 38252 40284
rect 37956 40230 38002 40282
rect 38002 40230 38012 40282
rect 38036 40230 38066 40282
rect 38066 40230 38078 40282
rect 38078 40230 38092 40282
rect 38116 40230 38130 40282
rect 38130 40230 38142 40282
rect 38142 40230 38172 40282
rect 38196 40230 38206 40282
rect 38206 40230 38252 40282
rect 37956 40228 38012 40230
rect 38036 40228 38092 40230
rect 38116 40228 38172 40230
rect 38196 40228 38252 40230
rect 37956 39194 38012 39196
rect 38036 39194 38092 39196
rect 38116 39194 38172 39196
rect 38196 39194 38252 39196
rect 37956 39142 38002 39194
rect 38002 39142 38012 39194
rect 38036 39142 38066 39194
rect 38066 39142 38078 39194
rect 38078 39142 38092 39194
rect 38116 39142 38130 39194
rect 38130 39142 38142 39194
rect 38142 39142 38172 39194
rect 38196 39142 38206 39194
rect 38206 39142 38252 39194
rect 37956 39140 38012 39142
rect 38036 39140 38092 39142
rect 38116 39140 38172 39142
rect 38196 39140 38252 39142
rect 37956 38106 38012 38108
rect 38036 38106 38092 38108
rect 38116 38106 38172 38108
rect 38196 38106 38252 38108
rect 37956 38054 38002 38106
rect 38002 38054 38012 38106
rect 38036 38054 38066 38106
rect 38066 38054 38078 38106
rect 38078 38054 38092 38106
rect 38116 38054 38130 38106
rect 38130 38054 38142 38106
rect 38142 38054 38172 38106
rect 38196 38054 38206 38106
rect 38206 38054 38252 38106
rect 37956 38052 38012 38054
rect 38036 38052 38092 38054
rect 38116 38052 38172 38054
rect 38196 38052 38252 38054
rect 37922 37748 37924 37768
rect 37924 37748 37976 37768
rect 37976 37748 37978 37768
rect 37922 37712 37978 37748
rect 37956 37018 38012 37020
rect 38036 37018 38092 37020
rect 38116 37018 38172 37020
rect 38196 37018 38252 37020
rect 37956 36966 38002 37018
rect 38002 36966 38012 37018
rect 38036 36966 38066 37018
rect 38066 36966 38078 37018
rect 38078 36966 38092 37018
rect 38116 36966 38130 37018
rect 38130 36966 38142 37018
rect 38142 36966 38172 37018
rect 38196 36966 38206 37018
rect 38206 36966 38252 37018
rect 37956 36964 38012 36966
rect 38036 36964 38092 36966
rect 38116 36964 38172 36966
rect 38196 36964 38252 36966
rect 38014 36624 38070 36680
rect 37956 35930 38012 35932
rect 38036 35930 38092 35932
rect 38116 35930 38172 35932
rect 38196 35930 38252 35932
rect 37956 35878 38002 35930
rect 38002 35878 38012 35930
rect 38036 35878 38066 35930
rect 38066 35878 38078 35930
rect 38078 35878 38092 35930
rect 38116 35878 38130 35930
rect 38130 35878 38142 35930
rect 38142 35878 38172 35930
rect 38196 35878 38206 35930
rect 38206 35878 38252 35930
rect 37956 35876 38012 35878
rect 38036 35876 38092 35878
rect 38116 35876 38172 35878
rect 38196 35876 38252 35878
rect 38658 40432 38714 40488
rect 38658 38664 38714 38720
rect 38842 37712 38898 37768
rect 38566 36760 38622 36816
rect 37922 35148 37978 35184
rect 37922 35128 37924 35148
rect 37924 35128 37976 35148
rect 37976 35128 37978 35148
rect 37956 34842 38012 34844
rect 38036 34842 38092 34844
rect 38116 34842 38172 34844
rect 38196 34842 38252 34844
rect 37956 34790 38002 34842
rect 38002 34790 38012 34842
rect 38036 34790 38066 34842
rect 38066 34790 38078 34842
rect 38078 34790 38092 34842
rect 38116 34790 38130 34842
rect 38130 34790 38142 34842
rect 38142 34790 38172 34842
rect 38196 34790 38206 34842
rect 38206 34790 38252 34842
rect 37956 34788 38012 34790
rect 38036 34788 38092 34790
rect 38116 34788 38172 34790
rect 38196 34788 38252 34790
rect 37094 31728 37150 31784
rect 37002 31320 37058 31376
rect 36450 28464 36506 28520
rect 35162 20576 35218 20632
rect 34978 19352 35034 19408
rect 37094 26288 37150 26344
rect 38658 35012 38714 35048
rect 38658 34992 38660 35012
rect 38660 34992 38712 35012
rect 38712 34992 38714 35012
rect 39118 37712 39174 37768
rect 38934 34856 38990 34912
rect 38934 34740 38990 34776
rect 38934 34720 38936 34740
rect 38936 34720 38988 34740
rect 38988 34720 38990 34740
rect 38750 34176 38806 34232
rect 37956 33754 38012 33756
rect 38036 33754 38092 33756
rect 38116 33754 38172 33756
rect 38196 33754 38252 33756
rect 37956 33702 38002 33754
rect 38002 33702 38012 33754
rect 38036 33702 38066 33754
rect 38066 33702 38078 33754
rect 38078 33702 38092 33754
rect 38116 33702 38130 33754
rect 38130 33702 38142 33754
rect 38142 33702 38172 33754
rect 38196 33702 38206 33754
rect 38206 33702 38252 33754
rect 37956 33700 38012 33702
rect 38036 33700 38092 33702
rect 38116 33700 38172 33702
rect 38196 33700 38252 33702
rect 38658 34060 38714 34096
rect 38658 34040 38660 34060
rect 38660 34040 38712 34060
rect 38712 34040 38714 34060
rect 37830 33516 37886 33552
rect 37830 33496 37832 33516
rect 37832 33496 37884 33516
rect 37884 33496 37886 33516
rect 37956 32666 38012 32668
rect 38036 32666 38092 32668
rect 38116 32666 38172 32668
rect 38196 32666 38252 32668
rect 37956 32614 38002 32666
rect 38002 32614 38012 32666
rect 38036 32614 38066 32666
rect 38066 32614 38078 32666
rect 38078 32614 38092 32666
rect 38116 32614 38130 32666
rect 38130 32614 38142 32666
rect 38142 32614 38172 32666
rect 38196 32614 38206 32666
rect 38206 32614 38252 32666
rect 37956 32612 38012 32614
rect 38036 32612 38092 32614
rect 38116 32612 38172 32614
rect 38196 32612 38252 32614
rect 38750 33632 38806 33688
rect 38842 33496 38898 33552
rect 37278 28056 37334 28112
rect 37956 31578 38012 31580
rect 38036 31578 38092 31580
rect 38116 31578 38172 31580
rect 38196 31578 38252 31580
rect 37956 31526 38002 31578
rect 38002 31526 38012 31578
rect 38036 31526 38066 31578
rect 38066 31526 38078 31578
rect 38078 31526 38092 31578
rect 38116 31526 38130 31578
rect 38130 31526 38142 31578
rect 38142 31526 38172 31578
rect 38196 31526 38206 31578
rect 38206 31526 38252 31578
rect 37956 31524 38012 31526
rect 38036 31524 38092 31526
rect 38116 31524 38172 31526
rect 38196 31524 38252 31526
rect 38566 31884 38622 31920
rect 38566 31864 38568 31884
rect 38568 31864 38620 31884
rect 38620 31864 38622 31884
rect 38566 31728 38622 31784
rect 38474 31320 38530 31376
rect 37956 30490 38012 30492
rect 38036 30490 38092 30492
rect 38116 30490 38172 30492
rect 38196 30490 38252 30492
rect 37956 30438 38002 30490
rect 38002 30438 38012 30490
rect 38036 30438 38066 30490
rect 38066 30438 38078 30490
rect 38078 30438 38092 30490
rect 38116 30438 38130 30490
rect 38130 30438 38142 30490
rect 38142 30438 38172 30490
rect 38196 30438 38206 30490
rect 38206 30438 38252 30490
rect 37956 30436 38012 30438
rect 38036 30436 38092 30438
rect 38116 30436 38172 30438
rect 38196 30436 38252 30438
rect 37922 30268 37924 30288
rect 37924 30268 37976 30288
rect 37976 30268 37978 30288
rect 37922 30232 37978 30268
rect 37956 29402 38012 29404
rect 38036 29402 38092 29404
rect 38116 29402 38172 29404
rect 38196 29402 38252 29404
rect 37956 29350 38002 29402
rect 38002 29350 38012 29402
rect 38036 29350 38066 29402
rect 38066 29350 38078 29402
rect 38078 29350 38092 29402
rect 38116 29350 38130 29402
rect 38130 29350 38142 29402
rect 38142 29350 38172 29402
rect 38196 29350 38206 29402
rect 38206 29350 38252 29402
rect 37956 29348 38012 29350
rect 38036 29348 38092 29350
rect 38116 29348 38172 29350
rect 38196 29348 38252 29350
rect 37956 28314 38012 28316
rect 38036 28314 38092 28316
rect 38116 28314 38172 28316
rect 38196 28314 38252 28316
rect 37956 28262 38002 28314
rect 38002 28262 38012 28314
rect 38036 28262 38066 28314
rect 38066 28262 38078 28314
rect 38078 28262 38092 28314
rect 38116 28262 38130 28314
rect 38130 28262 38142 28314
rect 38142 28262 38172 28314
rect 38196 28262 38206 28314
rect 38206 28262 38252 28314
rect 37956 28260 38012 28262
rect 38036 28260 38092 28262
rect 38116 28260 38172 28262
rect 38196 28260 38252 28262
rect 37956 27226 38012 27228
rect 38036 27226 38092 27228
rect 38116 27226 38172 27228
rect 38196 27226 38252 27228
rect 37956 27174 38002 27226
rect 38002 27174 38012 27226
rect 38036 27174 38066 27226
rect 38066 27174 38078 27226
rect 38078 27174 38092 27226
rect 38116 27174 38130 27226
rect 38130 27174 38142 27226
rect 38142 27174 38172 27226
rect 38196 27174 38206 27226
rect 38206 27174 38252 27226
rect 37956 27172 38012 27174
rect 38036 27172 38092 27174
rect 38116 27172 38172 27174
rect 38196 27172 38252 27174
rect 37956 26138 38012 26140
rect 38036 26138 38092 26140
rect 38116 26138 38172 26140
rect 38196 26138 38252 26140
rect 37956 26086 38002 26138
rect 38002 26086 38012 26138
rect 38036 26086 38066 26138
rect 38066 26086 38078 26138
rect 38078 26086 38092 26138
rect 38116 26086 38130 26138
rect 38130 26086 38142 26138
rect 38142 26086 38172 26138
rect 38196 26086 38206 26138
rect 38206 26086 38252 26138
rect 37956 26084 38012 26086
rect 38036 26084 38092 26086
rect 38116 26084 38172 26086
rect 38196 26084 38252 26086
rect 37956 25050 38012 25052
rect 38036 25050 38092 25052
rect 38116 25050 38172 25052
rect 38196 25050 38252 25052
rect 37956 24998 38002 25050
rect 38002 24998 38012 25050
rect 38036 24998 38066 25050
rect 38066 24998 38078 25050
rect 38078 24998 38092 25050
rect 38116 24998 38130 25050
rect 38130 24998 38142 25050
rect 38142 24998 38172 25050
rect 38196 24998 38206 25050
rect 38206 24998 38252 25050
rect 37956 24996 38012 24998
rect 38036 24996 38092 24998
rect 38116 24996 38172 24998
rect 38196 24996 38252 24998
rect 37956 23962 38012 23964
rect 38036 23962 38092 23964
rect 38116 23962 38172 23964
rect 38196 23962 38252 23964
rect 37956 23910 38002 23962
rect 38002 23910 38012 23962
rect 38036 23910 38066 23962
rect 38066 23910 38078 23962
rect 38078 23910 38092 23962
rect 38116 23910 38130 23962
rect 38130 23910 38142 23962
rect 38142 23910 38172 23962
rect 38196 23910 38206 23962
rect 38206 23910 38252 23962
rect 37956 23908 38012 23910
rect 38036 23908 38092 23910
rect 38116 23908 38172 23910
rect 38196 23908 38252 23910
rect 38658 26288 38714 26344
rect 37956 22874 38012 22876
rect 38036 22874 38092 22876
rect 38116 22874 38172 22876
rect 38196 22874 38252 22876
rect 37956 22822 38002 22874
rect 38002 22822 38012 22874
rect 38036 22822 38066 22874
rect 38066 22822 38078 22874
rect 38078 22822 38092 22874
rect 38116 22822 38130 22874
rect 38130 22822 38142 22874
rect 38142 22822 38172 22874
rect 38196 22822 38206 22874
rect 38206 22822 38252 22874
rect 37956 22820 38012 22822
rect 38036 22820 38092 22822
rect 38116 22820 38172 22822
rect 38196 22820 38252 22822
rect 37956 21786 38012 21788
rect 38036 21786 38092 21788
rect 38116 21786 38172 21788
rect 38196 21786 38252 21788
rect 37956 21734 38002 21786
rect 38002 21734 38012 21786
rect 38036 21734 38066 21786
rect 38066 21734 38078 21786
rect 38078 21734 38092 21786
rect 38116 21734 38130 21786
rect 38130 21734 38142 21786
rect 38142 21734 38172 21786
rect 38196 21734 38206 21786
rect 38206 21734 38252 21786
rect 37956 21732 38012 21734
rect 38036 21732 38092 21734
rect 38116 21732 38172 21734
rect 38196 21732 38252 21734
rect 37956 20698 38012 20700
rect 38036 20698 38092 20700
rect 38116 20698 38172 20700
rect 38196 20698 38252 20700
rect 37956 20646 38002 20698
rect 38002 20646 38012 20698
rect 38036 20646 38066 20698
rect 38066 20646 38078 20698
rect 38078 20646 38092 20698
rect 38116 20646 38130 20698
rect 38130 20646 38142 20698
rect 38142 20646 38172 20698
rect 38196 20646 38206 20698
rect 38206 20646 38252 20698
rect 37956 20644 38012 20646
rect 38036 20644 38092 20646
rect 38116 20644 38172 20646
rect 38196 20644 38252 20646
rect 37956 19610 38012 19612
rect 38036 19610 38092 19612
rect 38116 19610 38172 19612
rect 38196 19610 38252 19612
rect 37956 19558 38002 19610
rect 38002 19558 38012 19610
rect 38036 19558 38066 19610
rect 38066 19558 38078 19610
rect 38078 19558 38092 19610
rect 38116 19558 38130 19610
rect 38130 19558 38142 19610
rect 38142 19558 38172 19610
rect 38196 19558 38206 19610
rect 38206 19558 38252 19610
rect 37956 19556 38012 19558
rect 38036 19556 38092 19558
rect 38116 19556 38172 19558
rect 38196 19556 38252 19558
rect 37956 18522 38012 18524
rect 38036 18522 38092 18524
rect 38116 18522 38172 18524
rect 38196 18522 38252 18524
rect 37956 18470 38002 18522
rect 38002 18470 38012 18522
rect 38036 18470 38066 18522
rect 38066 18470 38078 18522
rect 38078 18470 38092 18522
rect 38116 18470 38130 18522
rect 38130 18470 38142 18522
rect 38142 18470 38172 18522
rect 38196 18470 38206 18522
rect 38206 18470 38252 18522
rect 37956 18468 38012 18470
rect 38036 18468 38092 18470
rect 38116 18468 38172 18470
rect 38196 18468 38252 18470
rect 37956 17434 38012 17436
rect 38036 17434 38092 17436
rect 38116 17434 38172 17436
rect 38196 17434 38252 17436
rect 37956 17382 38002 17434
rect 38002 17382 38012 17434
rect 38036 17382 38066 17434
rect 38066 17382 38078 17434
rect 38078 17382 38092 17434
rect 38116 17382 38130 17434
rect 38130 17382 38142 17434
rect 38142 17382 38172 17434
rect 38196 17382 38206 17434
rect 38206 17382 38252 17434
rect 37956 17380 38012 17382
rect 38036 17380 38092 17382
rect 38116 17380 38172 17382
rect 38196 17380 38252 17382
rect 37956 16346 38012 16348
rect 38036 16346 38092 16348
rect 38116 16346 38172 16348
rect 38196 16346 38252 16348
rect 37956 16294 38002 16346
rect 38002 16294 38012 16346
rect 38036 16294 38066 16346
rect 38066 16294 38078 16346
rect 38078 16294 38092 16346
rect 38116 16294 38130 16346
rect 38130 16294 38142 16346
rect 38142 16294 38172 16346
rect 38196 16294 38206 16346
rect 38206 16294 38252 16346
rect 37956 16292 38012 16294
rect 38036 16292 38092 16294
rect 38116 16292 38172 16294
rect 38196 16292 38252 16294
rect 37956 15258 38012 15260
rect 38036 15258 38092 15260
rect 38116 15258 38172 15260
rect 38196 15258 38252 15260
rect 37956 15206 38002 15258
rect 38002 15206 38012 15258
rect 38036 15206 38066 15258
rect 38066 15206 38078 15258
rect 38078 15206 38092 15258
rect 38116 15206 38130 15258
rect 38130 15206 38142 15258
rect 38142 15206 38172 15258
rect 38196 15206 38206 15258
rect 38206 15206 38252 15258
rect 37956 15204 38012 15206
rect 38036 15204 38092 15206
rect 38116 15204 38172 15206
rect 38196 15204 38252 15206
rect 37956 14170 38012 14172
rect 38036 14170 38092 14172
rect 38116 14170 38172 14172
rect 38196 14170 38252 14172
rect 37956 14118 38002 14170
rect 38002 14118 38012 14170
rect 38036 14118 38066 14170
rect 38066 14118 38078 14170
rect 38078 14118 38092 14170
rect 38116 14118 38130 14170
rect 38130 14118 38142 14170
rect 38142 14118 38172 14170
rect 38196 14118 38206 14170
rect 38206 14118 38252 14170
rect 37956 14116 38012 14118
rect 38036 14116 38092 14118
rect 38116 14116 38172 14118
rect 38196 14116 38252 14118
rect 39302 36624 39358 36680
rect 39394 34992 39450 35048
rect 39670 36216 39726 36272
rect 39302 33632 39358 33688
rect 39578 34076 39580 34096
rect 39580 34076 39632 34096
rect 39632 34076 39634 34096
rect 39578 34040 39634 34076
rect 40406 41656 40462 41712
rect 40038 36760 40094 36816
rect 40038 34176 40094 34232
rect 40774 35808 40830 35864
rect 40590 32952 40646 33008
rect 42956 53882 43012 53884
rect 43036 53882 43092 53884
rect 43116 53882 43172 53884
rect 43196 53882 43252 53884
rect 42956 53830 43002 53882
rect 43002 53830 43012 53882
rect 43036 53830 43066 53882
rect 43066 53830 43078 53882
rect 43078 53830 43092 53882
rect 43116 53830 43130 53882
rect 43130 53830 43142 53882
rect 43142 53830 43172 53882
rect 43196 53830 43206 53882
rect 43206 53830 43252 53882
rect 42956 53828 43012 53830
rect 43036 53828 43092 53830
rect 43116 53828 43172 53830
rect 43196 53828 43252 53830
rect 42956 52794 43012 52796
rect 43036 52794 43092 52796
rect 43116 52794 43172 52796
rect 43196 52794 43252 52796
rect 42956 52742 43002 52794
rect 43002 52742 43012 52794
rect 43036 52742 43066 52794
rect 43066 52742 43078 52794
rect 43078 52742 43092 52794
rect 43116 52742 43130 52794
rect 43130 52742 43142 52794
rect 43142 52742 43172 52794
rect 43196 52742 43206 52794
rect 43206 52742 43252 52794
rect 42956 52740 43012 52742
rect 43036 52740 43092 52742
rect 43116 52740 43172 52742
rect 43196 52740 43252 52742
rect 42956 51706 43012 51708
rect 43036 51706 43092 51708
rect 43116 51706 43172 51708
rect 43196 51706 43252 51708
rect 42956 51654 43002 51706
rect 43002 51654 43012 51706
rect 43036 51654 43066 51706
rect 43066 51654 43078 51706
rect 43078 51654 43092 51706
rect 43116 51654 43130 51706
rect 43130 51654 43142 51706
rect 43142 51654 43172 51706
rect 43196 51654 43206 51706
rect 43206 51654 43252 51706
rect 42956 51652 43012 51654
rect 43036 51652 43092 51654
rect 43116 51652 43172 51654
rect 43196 51652 43252 51654
rect 42956 50618 43012 50620
rect 43036 50618 43092 50620
rect 43116 50618 43172 50620
rect 43196 50618 43252 50620
rect 42956 50566 43002 50618
rect 43002 50566 43012 50618
rect 43036 50566 43066 50618
rect 43066 50566 43078 50618
rect 43078 50566 43092 50618
rect 43116 50566 43130 50618
rect 43130 50566 43142 50618
rect 43142 50566 43172 50618
rect 43196 50566 43206 50618
rect 43206 50566 43252 50618
rect 42956 50564 43012 50566
rect 43036 50564 43092 50566
rect 43116 50564 43172 50566
rect 43196 50564 43252 50566
rect 42956 49530 43012 49532
rect 43036 49530 43092 49532
rect 43116 49530 43172 49532
rect 43196 49530 43252 49532
rect 42956 49478 43002 49530
rect 43002 49478 43012 49530
rect 43036 49478 43066 49530
rect 43066 49478 43078 49530
rect 43078 49478 43092 49530
rect 43116 49478 43130 49530
rect 43130 49478 43142 49530
rect 43142 49478 43172 49530
rect 43196 49478 43206 49530
rect 43206 49478 43252 49530
rect 42956 49476 43012 49478
rect 43036 49476 43092 49478
rect 43116 49476 43172 49478
rect 43196 49476 43252 49478
rect 42956 48442 43012 48444
rect 43036 48442 43092 48444
rect 43116 48442 43172 48444
rect 43196 48442 43252 48444
rect 42956 48390 43002 48442
rect 43002 48390 43012 48442
rect 43036 48390 43066 48442
rect 43066 48390 43078 48442
rect 43078 48390 43092 48442
rect 43116 48390 43130 48442
rect 43130 48390 43142 48442
rect 43142 48390 43172 48442
rect 43196 48390 43206 48442
rect 43206 48390 43252 48442
rect 42956 48388 43012 48390
rect 43036 48388 43092 48390
rect 43116 48388 43172 48390
rect 43196 48388 43252 48390
rect 42956 47354 43012 47356
rect 43036 47354 43092 47356
rect 43116 47354 43172 47356
rect 43196 47354 43252 47356
rect 42956 47302 43002 47354
rect 43002 47302 43012 47354
rect 43036 47302 43066 47354
rect 43066 47302 43078 47354
rect 43078 47302 43092 47354
rect 43116 47302 43130 47354
rect 43130 47302 43142 47354
rect 43142 47302 43172 47354
rect 43196 47302 43206 47354
rect 43206 47302 43252 47354
rect 42956 47300 43012 47302
rect 43036 47300 43092 47302
rect 43116 47300 43172 47302
rect 43196 47300 43252 47302
rect 42956 46266 43012 46268
rect 43036 46266 43092 46268
rect 43116 46266 43172 46268
rect 43196 46266 43252 46268
rect 42956 46214 43002 46266
rect 43002 46214 43012 46266
rect 43036 46214 43066 46266
rect 43066 46214 43078 46266
rect 43078 46214 43092 46266
rect 43116 46214 43130 46266
rect 43130 46214 43142 46266
rect 43142 46214 43172 46266
rect 43196 46214 43206 46266
rect 43206 46214 43252 46266
rect 42956 46212 43012 46214
rect 43036 46212 43092 46214
rect 43116 46212 43172 46214
rect 43196 46212 43252 46214
rect 42956 45178 43012 45180
rect 43036 45178 43092 45180
rect 43116 45178 43172 45180
rect 43196 45178 43252 45180
rect 42956 45126 43002 45178
rect 43002 45126 43012 45178
rect 43036 45126 43066 45178
rect 43066 45126 43078 45178
rect 43078 45126 43092 45178
rect 43116 45126 43130 45178
rect 43130 45126 43142 45178
rect 43142 45126 43172 45178
rect 43196 45126 43206 45178
rect 43206 45126 43252 45178
rect 42956 45124 43012 45126
rect 43036 45124 43092 45126
rect 43116 45124 43172 45126
rect 43196 45124 43252 45126
rect 42956 44090 43012 44092
rect 43036 44090 43092 44092
rect 43116 44090 43172 44092
rect 43196 44090 43252 44092
rect 42956 44038 43002 44090
rect 43002 44038 43012 44090
rect 43036 44038 43066 44090
rect 43066 44038 43078 44090
rect 43078 44038 43092 44090
rect 43116 44038 43130 44090
rect 43130 44038 43142 44090
rect 43142 44038 43172 44090
rect 43196 44038 43206 44090
rect 43206 44038 43252 44090
rect 42956 44036 43012 44038
rect 43036 44036 43092 44038
rect 43116 44036 43172 44038
rect 43196 44036 43252 44038
rect 41326 42064 41382 42120
rect 42956 43002 43012 43004
rect 43036 43002 43092 43004
rect 43116 43002 43172 43004
rect 43196 43002 43252 43004
rect 42956 42950 43002 43002
rect 43002 42950 43012 43002
rect 43036 42950 43066 43002
rect 43066 42950 43078 43002
rect 43078 42950 43092 43002
rect 43116 42950 43130 43002
rect 43130 42950 43142 43002
rect 43142 42950 43172 43002
rect 43196 42950 43206 43002
rect 43206 42950 43252 43002
rect 42956 42948 43012 42950
rect 43036 42948 43092 42950
rect 43116 42948 43172 42950
rect 43196 42948 43252 42950
rect 42956 41914 43012 41916
rect 43036 41914 43092 41916
rect 43116 41914 43172 41916
rect 43196 41914 43252 41916
rect 42956 41862 43002 41914
rect 43002 41862 43012 41914
rect 43036 41862 43066 41914
rect 43066 41862 43078 41914
rect 43078 41862 43092 41914
rect 43116 41862 43130 41914
rect 43130 41862 43142 41914
rect 43142 41862 43172 41914
rect 43196 41862 43206 41914
rect 43206 41862 43252 41914
rect 42956 41860 43012 41862
rect 43036 41860 43092 41862
rect 43116 41860 43172 41862
rect 43196 41860 43252 41862
rect 42956 40826 43012 40828
rect 43036 40826 43092 40828
rect 43116 40826 43172 40828
rect 43196 40826 43252 40828
rect 42956 40774 43002 40826
rect 43002 40774 43012 40826
rect 43036 40774 43066 40826
rect 43066 40774 43078 40826
rect 43078 40774 43092 40826
rect 43116 40774 43130 40826
rect 43130 40774 43142 40826
rect 43142 40774 43172 40826
rect 43196 40774 43206 40826
rect 43206 40774 43252 40826
rect 42956 40772 43012 40774
rect 43036 40772 43092 40774
rect 43116 40772 43172 40774
rect 43196 40772 43252 40774
rect 41142 35808 41198 35864
rect 41142 34720 41198 34776
rect 40866 32952 40922 33008
rect 41786 36236 41842 36272
rect 41786 36216 41788 36236
rect 41788 36216 41840 36236
rect 41840 36216 41842 36236
rect 42956 39738 43012 39740
rect 43036 39738 43092 39740
rect 43116 39738 43172 39740
rect 43196 39738 43252 39740
rect 42956 39686 43002 39738
rect 43002 39686 43012 39738
rect 43036 39686 43066 39738
rect 43066 39686 43078 39738
rect 43078 39686 43092 39738
rect 43116 39686 43130 39738
rect 43130 39686 43142 39738
rect 43142 39686 43172 39738
rect 43196 39686 43206 39738
rect 43206 39686 43252 39738
rect 42956 39684 43012 39686
rect 43036 39684 43092 39686
rect 43116 39684 43172 39686
rect 43196 39684 43252 39686
rect 42956 38650 43012 38652
rect 43036 38650 43092 38652
rect 43116 38650 43172 38652
rect 43196 38650 43252 38652
rect 42956 38598 43002 38650
rect 43002 38598 43012 38650
rect 43036 38598 43066 38650
rect 43066 38598 43078 38650
rect 43078 38598 43092 38650
rect 43116 38598 43130 38650
rect 43130 38598 43142 38650
rect 43142 38598 43172 38650
rect 43196 38598 43206 38650
rect 43206 38598 43252 38650
rect 42956 38596 43012 38598
rect 43036 38596 43092 38598
rect 43116 38596 43172 38598
rect 43196 38596 43252 38598
rect 42338 36796 42340 36816
rect 42340 36796 42392 36816
rect 42392 36796 42394 36816
rect 42338 36760 42394 36796
rect 42956 37562 43012 37564
rect 43036 37562 43092 37564
rect 43116 37562 43172 37564
rect 43196 37562 43252 37564
rect 42956 37510 43002 37562
rect 43002 37510 43012 37562
rect 43036 37510 43066 37562
rect 43066 37510 43078 37562
rect 43078 37510 43092 37562
rect 43116 37510 43130 37562
rect 43130 37510 43142 37562
rect 43142 37510 43172 37562
rect 43196 37510 43206 37562
rect 43206 37510 43252 37562
rect 42956 37508 43012 37510
rect 43036 37508 43092 37510
rect 43116 37508 43172 37510
rect 43196 37508 43252 37510
rect 42956 36474 43012 36476
rect 43036 36474 43092 36476
rect 43116 36474 43172 36476
rect 43196 36474 43252 36476
rect 42956 36422 43002 36474
rect 43002 36422 43012 36474
rect 43036 36422 43066 36474
rect 43066 36422 43078 36474
rect 43078 36422 43092 36474
rect 43116 36422 43130 36474
rect 43130 36422 43142 36474
rect 43142 36422 43172 36474
rect 43196 36422 43206 36474
rect 43206 36422 43252 36474
rect 42956 36420 43012 36422
rect 43036 36420 43092 36422
rect 43116 36420 43172 36422
rect 43196 36420 43252 36422
rect 42956 35386 43012 35388
rect 43036 35386 43092 35388
rect 43116 35386 43172 35388
rect 43196 35386 43252 35388
rect 42956 35334 43002 35386
rect 43002 35334 43012 35386
rect 43036 35334 43066 35386
rect 43066 35334 43078 35386
rect 43078 35334 43092 35386
rect 43116 35334 43130 35386
rect 43130 35334 43142 35386
rect 43142 35334 43172 35386
rect 43196 35334 43206 35386
rect 43206 35334 43252 35386
rect 42956 35332 43012 35334
rect 43036 35332 43092 35334
rect 43116 35332 43172 35334
rect 43196 35332 43252 35334
rect 42956 34298 43012 34300
rect 43036 34298 43092 34300
rect 43116 34298 43172 34300
rect 43196 34298 43252 34300
rect 42956 34246 43002 34298
rect 43002 34246 43012 34298
rect 43036 34246 43066 34298
rect 43066 34246 43078 34298
rect 43078 34246 43092 34298
rect 43116 34246 43130 34298
rect 43130 34246 43142 34298
rect 43142 34246 43172 34298
rect 43196 34246 43206 34298
rect 43206 34246 43252 34298
rect 42956 34244 43012 34246
rect 43036 34244 43092 34246
rect 43116 34244 43172 34246
rect 43196 34244 43252 34246
rect 42956 33210 43012 33212
rect 43036 33210 43092 33212
rect 43116 33210 43172 33212
rect 43196 33210 43252 33212
rect 42956 33158 43002 33210
rect 43002 33158 43012 33210
rect 43036 33158 43066 33210
rect 43066 33158 43078 33210
rect 43078 33158 43092 33210
rect 43116 33158 43130 33210
rect 43130 33158 43142 33210
rect 43142 33158 43172 33210
rect 43196 33158 43206 33210
rect 43206 33158 43252 33210
rect 42956 33156 43012 33158
rect 43036 33156 43092 33158
rect 43116 33156 43172 33158
rect 43196 33156 43252 33158
rect 42956 32122 43012 32124
rect 43036 32122 43092 32124
rect 43116 32122 43172 32124
rect 43196 32122 43252 32124
rect 42956 32070 43002 32122
rect 43002 32070 43012 32122
rect 43036 32070 43066 32122
rect 43066 32070 43078 32122
rect 43078 32070 43092 32122
rect 43116 32070 43130 32122
rect 43130 32070 43142 32122
rect 43142 32070 43172 32122
rect 43196 32070 43206 32122
rect 43206 32070 43252 32122
rect 42956 32068 43012 32070
rect 43036 32068 43092 32070
rect 43116 32068 43172 32070
rect 43196 32068 43252 32070
rect 42956 31034 43012 31036
rect 43036 31034 43092 31036
rect 43116 31034 43172 31036
rect 43196 31034 43252 31036
rect 42956 30982 43002 31034
rect 43002 30982 43012 31034
rect 43036 30982 43066 31034
rect 43066 30982 43078 31034
rect 43078 30982 43092 31034
rect 43116 30982 43130 31034
rect 43130 30982 43142 31034
rect 43142 30982 43172 31034
rect 43196 30982 43206 31034
rect 43206 30982 43252 31034
rect 42956 30980 43012 30982
rect 43036 30980 43092 30982
rect 43116 30980 43172 30982
rect 43196 30980 43252 30982
rect 47956 54426 48012 54428
rect 48036 54426 48092 54428
rect 48116 54426 48172 54428
rect 48196 54426 48252 54428
rect 47956 54374 48002 54426
rect 48002 54374 48012 54426
rect 48036 54374 48066 54426
rect 48066 54374 48078 54426
rect 48078 54374 48092 54426
rect 48116 54374 48130 54426
rect 48130 54374 48142 54426
rect 48142 54374 48172 54426
rect 48196 54374 48206 54426
rect 48206 54374 48252 54426
rect 47956 54372 48012 54374
rect 48036 54372 48092 54374
rect 48116 54372 48172 54374
rect 48196 54372 48252 54374
rect 47956 53338 48012 53340
rect 48036 53338 48092 53340
rect 48116 53338 48172 53340
rect 48196 53338 48252 53340
rect 47956 53286 48002 53338
rect 48002 53286 48012 53338
rect 48036 53286 48066 53338
rect 48066 53286 48078 53338
rect 48078 53286 48092 53338
rect 48116 53286 48130 53338
rect 48130 53286 48142 53338
rect 48142 53286 48172 53338
rect 48196 53286 48206 53338
rect 48206 53286 48252 53338
rect 47956 53284 48012 53286
rect 48036 53284 48092 53286
rect 48116 53284 48172 53286
rect 48196 53284 48252 53286
rect 47956 52250 48012 52252
rect 48036 52250 48092 52252
rect 48116 52250 48172 52252
rect 48196 52250 48252 52252
rect 47956 52198 48002 52250
rect 48002 52198 48012 52250
rect 48036 52198 48066 52250
rect 48066 52198 48078 52250
rect 48078 52198 48092 52250
rect 48116 52198 48130 52250
rect 48130 52198 48142 52250
rect 48142 52198 48172 52250
rect 48196 52198 48206 52250
rect 48206 52198 48252 52250
rect 47956 52196 48012 52198
rect 48036 52196 48092 52198
rect 48116 52196 48172 52198
rect 48196 52196 48252 52198
rect 47956 51162 48012 51164
rect 48036 51162 48092 51164
rect 48116 51162 48172 51164
rect 48196 51162 48252 51164
rect 47956 51110 48002 51162
rect 48002 51110 48012 51162
rect 48036 51110 48066 51162
rect 48066 51110 48078 51162
rect 48078 51110 48092 51162
rect 48116 51110 48130 51162
rect 48130 51110 48142 51162
rect 48142 51110 48172 51162
rect 48196 51110 48206 51162
rect 48206 51110 48252 51162
rect 47956 51108 48012 51110
rect 48036 51108 48092 51110
rect 48116 51108 48172 51110
rect 48196 51108 48252 51110
rect 47956 50074 48012 50076
rect 48036 50074 48092 50076
rect 48116 50074 48172 50076
rect 48196 50074 48252 50076
rect 47956 50022 48002 50074
rect 48002 50022 48012 50074
rect 48036 50022 48066 50074
rect 48066 50022 48078 50074
rect 48078 50022 48092 50074
rect 48116 50022 48130 50074
rect 48130 50022 48142 50074
rect 48142 50022 48172 50074
rect 48196 50022 48206 50074
rect 48206 50022 48252 50074
rect 47956 50020 48012 50022
rect 48036 50020 48092 50022
rect 48116 50020 48172 50022
rect 48196 50020 48252 50022
rect 47956 48986 48012 48988
rect 48036 48986 48092 48988
rect 48116 48986 48172 48988
rect 48196 48986 48252 48988
rect 47956 48934 48002 48986
rect 48002 48934 48012 48986
rect 48036 48934 48066 48986
rect 48066 48934 48078 48986
rect 48078 48934 48092 48986
rect 48116 48934 48130 48986
rect 48130 48934 48142 48986
rect 48142 48934 48172 48986
rect 48196 48934 48206 48986
rect 48206 48934 48252 48986
rect 47956 48932 48012 48934
rect 48036 48932 48092 48934
rect 48116 48932 48172 48934
rect 48196 48932 48252 48934
rect 47956 47898 48012 47900
rect 48036 47898 48092 47900
rect 48116 47898 48172 47900
rect 48196 47898 48252 47900
rect 47956 47846 48002 47898
rect 48002 47846 48012 47898
rect 48036 47846 48066 47898
rect 48066 47846 48078 47898
rect 48078 47846 48092 47898
rect 48116 47846 48130 47898
rect 48130 47846 48142 47898
rect 48142 47846 48172 47898
rect 48196 47846 48206 47898
rect 48206 47846 48252 47898
rect 47956 47844 48012 47846
rect 48036 47844 48092 47846
rect 48116 47844 48172 47846
rect 48196 47844 48252 47846
rect 49330 52536 49386 52592
rect 49054 51856 49110 51912
rect 49054 51176 49110 51232
rect 48962 50496 49018 50552
rect 47956 46810 48012 46812
rect 48036 46810 48092 46812
rect 48116 46810 48172 46812
rect 48196 46810 48252 46812
rect 47956 46758 48002 46810
rect 48002 46758 48012 46810
rect 48036 46758 48066 46810
rect 48066 46758 48078 46810
rect 48078 46758 48092 46810
rect 48116 46758 48130 46810
rect 48130 46758 48142 46810
rect 48142 46758 48172 46810
rect 48196 46758 48206 46810
rect 48206 46758 48252 46810
rect 47956 46756 48012 46758
rect 48036 46756 48092 46758
rect 48116 46756 48172 46758
rect 48196 46756 48252 46758
rect 47956 45722 48012 45724
rect 48036 45722 48092 45724
rect 48116 45722 48172 45724
rect 48196 45722 48252 45724
rect 47956 45670 48002 45722
rect 48002 45670 48012 45722
rect 48036 45670 48066 45722
rect 48066 45670 48078 45722
rect 48078 45670 48092 45722
rect 48116 45670 48130 45722
rect 48130 45670 48142 45722
rect 48142 45670 48172 45722
rect 48196 45670 48206 45722
rect 48206 45670 48252 45722
rect 47956 45668 48012 45670
rect 48036 45668 48092 45670
rect 48116 45668 48172 45670
rect 48196 45668 48252 45670
rect 42956 29946 43012 29948
rect 43036 29946 43092 29948
rect 43116 29946 43172 29948
rect 43196 29946 43252 29948
rect 42956 29894 43002 29946
rect 43002 29894 43012 29946
rect 43036 29894 43066 29946
rect 43066 29894 43078 29946
rect 43078 29894 43092 29946
rect 43116 29894 43130 29946
rect 43130 29894 43142 29946
rect 43142 29894 43172 29946
rect 43196 29894 43206 29946
rect 43206 29894 43252 29946
rect 42956 29892 43012 29894
rect 43036 29892 43092 29894
rect 43116 29892 43172 29894
rect 43196 29892 43252 29894
rect 42956 28858 43012 28860
rect 43036 28858 43092 28860
rect 43116 28858 43172 28860
rect 43196 28858 43252 28860
rect 42956 28806 43002 28858
rect 43002 28806 43012 28858
rect 43036 28806 43066 28858
rect 43066 28806 43078 28858
rect 43078 28806 43092 28858
rect 43116 28806 43130 28858
rect 43130 28806 43142 28858
rect 43142 28806 43172 28858
rect 43196 28806 43206 28858
rect 43206 28806 43252 28858
rect 42956 28804 43012 28806
rect 43036 28804 43092 28806
rect 43116 28804 43172 28806
rect 43196 28804 43252 28806
rect 42956 27770 43012 27772
rect 43036 27770 43092 27772
rect 43116 27770 43172 27772
rect 43196 27770 43252 27772
rect 42956 27718 43002 27770
rect 43002 27718 43012 27770
rect 43036 27718 43066 27770
rect 43066 27718 43078 27770
rect 43078 27718 43092 27770
rect 43116 27718 43130 27770
rect 43130 27718 43142 27770
rect 43142 27718 43172 27770
rect 43196 27718 43206 27770
rect 43206 27718 43252 27770
rect 42956 27716 43012 27718
rect 43036 27716 43092 27718
rect 43116 27716 43172 27718
rect 43196 27716 43252 27718
rect 42956 26682 43012 26684
rect 43036 26682 43092 26684
rect 43116 26682 43172 26684
rect 43196 26682 43252 26684
rect 42956 26630 43002 26682
rect 43002 26630 43012 26682
rect 43036 26630 43066 26682
rect 43066 26630 43078 26682
rect 43078 26630 43092 26682
rect 43116 26630 43130 26682
rect 43130 26630 43142 26682
rect 43142 26630 43172 26682
rect 43196 26630 43206 26682
rect 43206 26630 43252 26682
rect 42956 26628 43012 26630
rect 43036 26628 43092 26630
rect 43116 26628 43172 26630
rect 43196 26628 43252 26630
rect 42956 25594 43012 25596
rect 43036 25594 43092 25596
rect 43116 25594 43172 25596
rect 43196 25594 43252 25596
rect 42956 25542 43002 25594
rect 43002 25542 43012 25594
rect 43036 25542 43066 25594
rect 43066 25542 43078 25594
rect 43078 25542 43092 25594
rect 43116 25542 43130 25594
rect 43130 25542 43142 25594
rect 43142 25542 43172 25594
rect 43196 25542 43206 25594
rect 43206 25542 43252 25594
rect 42956 25540 43012 25542
rect 43036 25540 43092 25542
rect 43116 25540 43172 25542
rect 43196 25540 43252 25542
rect 46294 36624 46350 36680
rect 47956 44634 48012 44636
rect 48036 44634 48092 44636
rect 48116 44634 48172 44636
rect 48196 44634 48252 44636
rect 47956 44582 48002 44634
rect 48002 44582 48012 44634
rect 48036 44582 48066 44634
rect 48066 44582 48078 44634
rect 48078 44582 48092 44634
rect 48116 44582 48130 44634
rect 48130 44582 48142 44634
rect 48142 44582 48172 44634
rect 48196 44582 48206 44634
rect 48206 44582 48252 44634
rect 47956 44580 48012 44582
rect 48036 44580 48092 44582
rect 48116 44580 48172 44582
rect 48196 44580 48252 44582
rect 47956 43546 48012 43548
rect 48036 43546 48092 43548
rect 48116 43546 48172 43548
rect 48196 43546 48252 43548
rect 47956 43494 48002 43546
rect 48002 43494 48012 43546
rect 48036 43494 48066 43546
rect 48066 43494 48078 43546
rect 48078 43494 48092 43546
rect 48116 43494 48130 43546
rect 48130 43494 48142 43546
rect 48142 43494 48172 43546
rect 48196 43494 48206 43546
rect 48206 43494 48252 43546
rect 47956 43492 48012 43494
rect 48036 43492 48092 43494
rect 48116 43492 48172 43494
rect 48196 43492 48252 43494
rect 47956 42458 48012 42460
rect 48036 42458 48092 42460
rect 48116 42458 48172 42460
rect 48196 42458 48252 42460
rect 47956 42406 48002 42458
rect 48002 42406 48012 42458
rect 48036 42406 48066 42458
rect 48066 42406 48078 42458
rect 48078 42406 48092 42458
rect 48116 42406 48130 42458
rect 48130 42406 48142 42458
rect 48142 42406 48172 42458
rect 48196 42406 48206 42458
rect 48206 42406 48252 42458
rect 47956 42404 48012 42406
rect 48036 42404 48092 42406
rect 48116 42404 48172 42406
rect 48196 42404 48252 42406
rect 48502 44376 48558 44432
rect 48502 43732 48504 43752
rect 48504 43732 48556 43752
rect 48556 43732 48558 43752
rect 48502 43696 48558 43732
rect 48502 43016 48558 43072
rect 48502 42336 48558 42392
rect 49054 49816 49110 49872
rect 49146 49136 49202 49192
rect 49238 48456 49294 48512
rect 49054 47776 49110 47832
rect 49054 47096 49110 47152
rect 48502 41656 48558 41712
rect 47956 41370 48012 41372
rect 48036 41370 48092 41372
rect 48116 41370 48172 41372
rect 48196 41370 48252 41372
rect 47956 41318 48002 41370
rect 48002 41318 48012 41370
rect 48036 41318 48066 41370
rect 48066 41318 48078 41370
rect 48078 41318 48092 41370
rect 48116 41318 48130 41370
rect 48130 41318 48142 41370
rect 48142 41318 48172 41370
rect 48196 41318 48206 41370
rect 48206 41318 48252 41370
rect 47956 41316 48012 41318
rect 48036 41316 48092 41318
rect 48116 41316 48172 41318
rect 48196 41316 48252 41318
rect 47956 40282 48012 40284
rect 48036 40282 48092 40284
rect 48116 40282 48172 40284
rect 48196 40282 48252 40284
rect 47956 40230 48002 40282
rect 48002 40230 48012 40282
rect 48036 40230 48066 40282
rect 48066 40230 48078 40282
rect 48078 40230 48092 40282
rect 48116 40230 48130 40282
rect 48130 40230 48142 40282
rect 48142 40230 48172 40282
rect 48196 40230 48206 40282
rect 48206 40230 48252 40282
rect 47956 40228 48012 40230
rect 48036 40228 48092 40230
rect 48116 40228 48172 40230
rect 48196 40228 48252 40230
rect 47956 39194 48012 39196
rect 48036 39194 48092 39196
rect 48116 39194 48172 39196
rect 48196 39194 48252 39196
rect 47956 39142 48002 39194
rect 48002 39142 48012 39194
rect 48036 39142 48066 39194
rect 48066 39142 48078 39194
rect 48078 39142 48092 39194
rect 48116 39142 48130 39194
rect 48130 39142 48142 39194
rect 48142 39142 48172 39194
rect 48196 39142 48206 39194
rect 48206 39142 48252 39194
rect 47956 39140 48012 39142
rect 48036 39140 48092 39142
rect 48116 39140 48172 39142
rect 48196 39140 48252 39142
rect 47956 38106 48012 38108
rect 48036 38106 48092 38108
rect 48116 38106 48172 38108
rect 48196 38106 48252 38108
rect 47956 38054 48002 38106
rect 48002 38054 48012 38106
rect 48036 38054 48066 38106
rect 48066 38054 48078 38106
rect 48078 38054 48092 38106
rect 48116 38054 48130 38106
rect 48130 38054 48142 38106
rect 48142 38054 48172 38106
rect 48196 38054 48206 38106
rect 48206 38054 48252 38106
rect 47956 38052 48012 38054
rect 48036 38052 48092 38054
rect 48116 38052 48172 38054
rect 48196 38052 48252 38054
rect 47956 37018 48012 37020
rect 48036 37018 48092 37020
rect 48116 37018 48172 37020
rect 48196 37018 48252 37020
rect 47956 36966 48002 37018
rect 48002 36966 48012 37018
rect 48036 36966 48066 37018
rect 48066 36966 48078 37018
rect 48078 36966 48092 37018
rect 48116 36966 48130 37018
rect 48130 36966 48142 37018
rect 48142 36966 48172 37018
rect 48196 36966 48206 37018
rect 48206 36966 48252 37018
rect 47956 36964 48012 36966
rect 48036 36964 48092 36966
rect 48116 36964 48172 36966
rect 48196 36964 48252 36966
rect 47956 35930 48012 35932
rect 48036 35930 48092 35932
rect 48116 35930 48172 35932
rect 48196 35930 48252 35932
rect 47956 35878 48002 35930
rect 48002 35878 48012 35930
rect 48036 35878 48066 35930
rect 48066 35878 48078 35930
rect 48078 35878 48092 35930
rect 48116 35878 48130 35930
rect 48130 35878 48142 35930
rect 48142 35878 48172 35930
rect 48196 35878 48206 35930
rect 48206 35878 48252 35930
rect 47956 35876 48012 35878
rect 48036 35876 48092 35878
rect 48116 35876 48172 35878
rect 48196 35876 48252 35878
rect 47956 34842 48012 34844
rect 48036 34842 48092 34844
rect 48116 34842 48172 34844
rect 48196 34842 48252 34844
rect 47956 34790 48002 34842
rect 48002 34790 48012 34842
rect 48036 34790 48066 34842
rect 48066 34790 48078 34842
rect 48078 34790 48092 34842
rect 48116 34790 48130 34842
rect 48130 34790 48142 34842
rect 48142 34790 48172 34842
rect 48196 34790 48206 34842
rect 48206 34790 48252 34842
rect 47956 34788 48012 34790
rect 48036 34788 48092 34790
rect 48116 34788 48172 34790
rect 48196 34788 48252 34790
rect 47956 33754 48012 33756
rect 48036 33754 48092 33756
rect 48116 33754 48172 33756
rect 48196 33754 48252 33756
rect 47956 33702 48002 33754
rect 48002 33702 48012 33754
rect 48036 33702 48066 33754
rect 48066 33702 48078 33754
rect 48078 33702 48092 33754
rect 48116 33702 48130 33754
rect 48130 33702 48142 33754
rect 48142 33702 48172 33754
rect 48196 33702 48206 33754
rect 48206 33702 48252 33754
rect 47956 33700 48012 33702
rect 48036 33700 48092 33702
rect 48116 33700 48172 33702
rect 48196 33700 48252 33702
rect 47956 32666 48012 32668
rect 48036 32666 48092 32668
rect 48116 32666 48172 32668
rect 48196 32666 48252 32668
rect 47956 32614 48002 32666
rect 48002 32614 48012 32666
rect 48036 32614 48066 32666
rect 48066 32614 48078 32666
rect 48078 32614 48092 32666
rect 48116 32614 48130 32666
rect 48130 32614 48142 32666
rect 48142 32614 48172 32666
rect 48196 32614 48206 32666
rect 48206 32614 48252 32666
rect 47956 32612 48012 32614
rect 48036 32612 48092 32614
rect 48116 32612 48172 32614
rect 48196 32612 48252 32614
rect 42956 24506 43012 24508
rect 43036 24506 43092 24508
rect 43116 24506 43172 24508
rect 43196 24506 43252 24508
rect 42956 24454 43002 24506
rect 43002 24454 43012 24506
rect 43036 24454 43066 24506
rect 43066 24454 43078 24506
rect 43078 24454 43092 24506
rect 43116 24454 43130 24506
rect 43130 24454 43142 24506
rect 43142 24454 43172 24506
rect 43196 24454 43206 24506
rect 43206 24454 43252 24506
rect 42956 24452 43012 24454
rect 43036 24452 43092 24454
rect 43116 24452 43172 24454
rect 43196 24452 43252 24454
rect 42956 23418 43012 23420
rect 43036 23418 43092 23420
rect 43116 23418 43172 23420
rect 43196 23418 43252 23420
rect 42956 23366 43002 23418
rect 43002 23366 43012 23418
rect 43036 23366 43066 23418
rect 43066 23366 43078 23418
rect 43078 23366 43092 23418
rect 43116 23366 43130 23418
rect 43130 23366 43142 23418
rect 43142 23366 43172 23418
rect 43196 23366 43206 23418
rect 43206 23366 43252 23418
rect 42956 23364 43012 23366
rect 43036 23364 43092 23366
rect 43116 23364 43172 23366
rect 43196 23364 43252 23366
rect 42956 22330 43012 22332
rect 43036 22330 43092 22332
rect 43116 22330 43172 22332
rect 43196 22330 43252 22332
rect 42956 22278 43002 22330
rect 43002 22278 43012 22330
rect 43036 22278 43066 22330
rect 43066 22278 43078 22330
rect 43078 22278 43092 22330
rect 43116 22278 43130 22330
rect 43130 22278 43142 22330
rect 43142 22278 43172 22330
rect 43196 22278 43206 22330
rect 43206 22278 43252 22330
rect 42956 22276 43012 22278
rect 43036 22276 43092 22278
rect 43116 22276 43172 22278
rect 43196 22276 43252 22278
rect 42956 21242 43012 21244
rect 43036 21242 43092 21244
rect 43116 21242 43172 21244
rect 43196 21242 43252 21244
rect 42956 21190 43002 21242
rect 43002 21190 43012 21242
rect 43036 21190 43066 21242
rect 43066 21190 43078 21242
rect 43078 21190 43092 21242
rect 43116 21190 43130 21242
rect 43130 21190 43142 21242
rect 43142 21190 43172 21242
rect 43196 21190 43206 21242
rect 43206 21190 43252 21242
rect 42956 21188 43012 21190
rect 43036 21188 43092 21190
rect 43116 21188 43172 21190
rect 43196 21188 43252 21190
rect 42956 20154 43012 20156
rect 43036 20154 43092 20156
rect 43116 20154 43172 20156
rect 43196 20154 43252 20156
rect 42956 20102 43002 20154
rect 43002 20102 43012 20154
rect 43036 20102 43066 20154
rect 43066 20102 43078 20154
rect 43078 20102 43092 20154
rect 43116 20102 43130 20154
rect 43130 20102 43142 20154
rect 43142 20102 43172 20154
rect 43196 20102 43206 20154
rect 43206 20102 43252 20154
rect 42956 20100 43012 20102
rect 43036 20100 43092 20102
rect 43116 20100 43172 20102
rect 43196 20100 43252 20102
rect 42956 19066 43012 19068
rect 43036 19066 43092 19068
rect 43116 19066 43172 19068
rect 43196 19066 43252 19068
rect 42956 19014 43002 19066
rect 43002 19014 43012 19066
rect 43036 19014 43066 19066
rect 43066 19014 43078 19066
rect 43078 19014 43092 19066
rect 43116 19014 43130 19066
rect 43130 19014 43142 19066
rect 43142 19014 43172 19066
rect 43196 19014 43206 19066
rect 43206 19014 43252 19066
rect 42956 19012 43012 19014
rect 43036 19012 43092 19014
rect 43116 19012 43172 19014
rect 43196 19012 43252 19014
rect 37956 13082 38012 13084
rect 38036 13082 38092 13084
rect 38116 13082 38172 13084
rect 38196 13082 38252 13084
rect 37956 13030 38002 13082
rect 38002 13030 38012 13082
rect 38036 13030 38066 13082
rect 38066 13030 38078 13082
rect 38078 13030 38092 13082
rect 38116 13030 38130 13082
rect 38130 13030 38142 13082
rect 38142 13030 38172 13082
rect 38196 13030 38206 13082
rect 38206 13030 38252 13082
rect 37956 13028 38012 13030
rect 38036 13028 38092 13030
rect 38116 13028 38172 13030
rect 38196 13028 38252 13030
rect 37956 11994 38012 11996
rect 38036 11994 38092 11996
rect 38116 11994 38172 11996
rect 38196 11994 38252 11996
rect 37956 11942 38002 11994
rect 38002 11942 38012 11994
rect 38036 11942 38066 11994
rect 38066 11942 38078 11994
rect 38078 11942 38092 11994
rect 38116 11942 38130 11994
rect 38130 11942 38142 11994
rect 38142 11942 38172 11994
rect 38196 11942 38206 11994
rect 38206 11942 38252 11994
rect 37956 11940 38012 11942
rect 38036 11940 38092 11942
rect 38116 11940 38172 11942
rect 38196 11940 38252 11942
rect 37956 10906 38012 10908
rect 38036 10906 38092 10908
rect 38116 10906 38172 10908
rect 38196 10906 38252 10908
rect 37956 10854 38002 10906
rect 38002 10854 38012 10906
rect 38036 10854 38066 10906
rect 38066 10854 38078 10906
rect 38078 10854 38092 10906
rect 38116 10854 38130 10906
rect 38130 10854 38142 10906
rect 38142 10854 38172 10906
rect 38196 10854 38206 10906
rect 38206 10854 38252 10906
rect 37956 10852 38012 10854
rect 38036 10852 38092 10854
rect 38116 10852 38172 10854
rect 38196 10852 38252 10854
rect 37956 9818 38012 9820
rect 38036 9818 38092 9820
rect 38116 9818 38172 9820
rect 38196 9818 38252 9820
rect 37956 9766 38002 9818
rect 38002 9766 38012 9818
rect 38036 9766 38066 9818
rect 38066 9766 38078 9818
rect 38078 9766 38092 9818
rect 38116 9766 38130 9818
rect 38130 9766 38142 9818
rect 38142 9766 38172 9818
rect 38196 9766 38206 9818
rect 38206 9766 38252 9818
rect 37956 9764 38012 9766
rect 38036 9764 38092 9766
rect 38116 9764 38172 9766
rect 38196 9764 38252 9766
rect 37956 8730 38012 8732
rect 38036 8730 38092 8732
rect 38116 8730 38172 8732
rect 38196 8730 38252 8732
rect 37956 8678 38002 8730
rect 38002 8678 38012 8730
rect 38036 8678 38066 8730
rect 38066 8678 38078 8730
rect 38078 8678 38092 8730
rect 38116 8678 38130 8730
rect 38130 8678 38142 8730
rect 38142 8678 38172 8730
rect 38196 8678 38206 8730
rect 38206 8678 38252 8730
rect 37956 8676 38012 8678
rect 38036 8676 38092 8678
rect 38116 8676 38172 8678
rect 38196 8676 38252 8678
rect 37956 7642 38012 7644
rect 38036 7642 38092 7644
rect 38116 7642 38172 7644
rect 38196 7642 38252 7644
rect 37956 7590 38002 7642
rect 38002 7590 38012 7642
rect 38036 7590 38066 7642
rect 38066 7590 38078 7642
rect 38078 7590 38092 7642
rect 38116 7590 38130 7642
rect 38130 7590 38142 7642
rect 38142 7590 38172 7642
rect 38196 7590 38206 7642
rect 38206 7590 38252 7642
rect 37956 7588 38012 7590
rect 38036 7588 38092 7590
rect 38116 7588 38172 7590
rect 38196 7588 38252 7590
rect 37956 6554 38012 6556
rect 38036 6554 38092 6556
rect 38116 6554 38172 6556
rect 38196 6554 38252 6556
rect 37956 6502 38002 6554
rect 38002 6502 38012 6554
rect 38036 6502 38066 6554
rect 38066 6502 38078 6554
rect 38078 6502 38092 6554
rect 38116 6502 38130 6554
rect 38130 6502 38142 6554
rect 38142 6502 38172 6554
rect 38196 6502 38206 6554
rect 38206 6502 38252 6554
rect 37956 6500 38012 6502
rect 38036 6500 38092 6502
rect 38116 6500 38172 6502
rect 38196 6500 38252 6502
rect 37956 5466 38012 5468
rect 38036 5466 38092 5468
rect 38116 5466 38172 5468
rect 38196 5466 38252 5468
rect 37956 5414 38002 5466
rect 38002 5414 38012 5466
rect 38036 5414 38066 5466
rect 38066 5414 38078 5466
rect 38078 5414 38092 5466
rect 38116 5414 38130 5466
rect 38130 5414 38142 5466
rect 38142 5414 38172 5466
rect 38196 5414 38206 5466
rect 38206 5414 38252 5466
rect 37956 5412 38012 5414
rect 38036 5412 38092 5414
rect 38116 5412 38172 5414
rect 38196 5412 38252 5414
rect 37956 4378 38012 4380
rect 38036 4378 38092 4380
rect 38116 4378 38172 4380
rect 38196 4378 38252 4380
rect 37956 4326 38002 4378
rect 38002 4326 38012 4378
rect 38036 4326 38066 4378
rect 38066 4326 38078 4378
rect 38078 4326 38092 4378
rect 38116 4326 38130 4378
rect 38130 4326 38142 4378
rect 38142 4326 38172 4378
rect 38196 4326 38206 4378
rect 38206 4326 38252 4378
rect 37956 4324 38012 4326
rect 38036 4324 38092 4326
rect 38116 4324 38172 4326
rect 38196 4324 38252 4326
rect 38934 12280 38990 12336
rect 37956 3290 38012 3292
rect 38036 3290 38092 3292
rect 38116 3290 38172 3292
rect 38196 3290 38252 3292
rect 37956 3238 38002 3290
rect 38002 3238 38012 3290
rect 38036 3238 38066 3290
rect 38066 3238 38078 3290
rect 38078 3238 38092 3290
rect 38116 3238 38130 3290
rect 38130 3238 38142 3290
rect 38142 3238 38172 3290
rect 38196 3238 38206 3290
rect 38206 3238 38252 3290
rect 37956 3236 38012 3238
rect 38036 3236 38092 3238
rect 38116 3236 38172 3238
rect 38196 3236 38252 3238
rect 37956 2202 38012 2204
rect 38036 2202 38092 2204
rect 38116 2202 38172 2204
rect 38196 2202 38252 2204
rect 37956 2150 38002 2202
rect 38002 2150 38012 2202
rect 38036 2150 38066 2202
rect 38066 2150 38078 2202
rect 38078 2150 38092 2202
rect 38116 2150 38130 2202
rect 38130 2150 38142 2202
rect 38142 2150 38172 2202
rect 38196 2150 38206 2202
rect 38206 2150 38252 2202
rect 37956 2148 38012 2150
rect 38036 2148 38092 2150
rect 38116 2148 38172 2150
rect 38196 2148 38252 2150
rect 42956 17978 43012 17980
rect 43036 17978 43092 17980
rect 43116 17978 43172 17980
rect 43196 17978 43252 17980
rect 42956 17926 43002 17978
rect 43002 17926 43012 17978
rect 43036 17926 43066 17978
rect 43066 17926 43078 17978
rect 43078 17926 43092 17978
rect 43116 17926 43130 17978
rect 43130 17926 43142 17978
rect 43142 17926 43172 17978
rect 43196 17926 43206 17978
rect 43206 17926 43252 17978
rect 42956 17924 43012 17926
rect 43036 17924 43092 17926
rect 43116 17924 43172 17926
rect 43196 17924 43252 17926
rect 42956 16890 43012 16892
rect 43036 16890 43092 16892
rect 43116 16890 43172 16892
rect 43196 16890 43252 16892
rect 42956 16838 43002 16890
rect 43002 16838 43012 16890
rect 43036 16838 43066 16890
rect 43066 16838 43078 16890
rect 43078 16838 43092 16890
rect 43116 16838 43130 16890
rect 43130 16838 43142 16890
rect 43142 16838 43172 16890
rect 43196 16838 43206 16890
rect 43206 16838 43252 16890
rect 42956 16836 43012 16838
rect 43036 16836 43092 16838
rect 43116 16836 43172 16838
rect 43196 16836 43252 16838
rect 42956 15802 43012 15804
rect 43036 15802 43092 15804
rect 43116 15802 43172 15804
rect 43196 15802 43252 15804
rect 42956 15750 43002 15802
rect 43002 15750 43012 15802
rect 43036 15750 43066 15802
rect 43066 15750 43078 15802
rect 43078 15750 43092 15802
rect 43116 15750 43130 15802
rect 43130 15750 43142 15802
rect 43142 15750 43172 15802
rect 43196 15750 43206 15802
rect 43206 15750 43252 15802
rect 42956 15748 43012 15750
rect 43036 15748 43092 15750
rect 43116 15748 43172 15750
rect 43196 15748 43252 15750
rect 42956 14714 43012 14716
rect 43036 14714 43092 14716
rect 43116 14714 43172 14716
rect 43196 14714 43252 14716
rect 42956 14662 43002 14714
rect 43002 14662 43012 14714
rect 43036 14662 43066 14714
rect 43066 14662 43078 14714
rect 43078 14662 43092 14714
rect 43116 14662 43130 14714
rect 43130 14662 43142 14714
rect 43142 14662 43172 14714
rect 43196 14662 43206 14714
rect 43206 14662 43252 14714
rect 42956 14660 43012 14662
rect 43036 14660 43092 14662
rect 43116 14660 43172 14662
rect 43196 14660 43252 14662
rect 42956 13626 43012 13628
rect 43036 13626 43092 13628
rect 43116 13626 43172 13628
rect 43196 13626 43252 13628
rect 42956 13574 43002 13626
rect 43002 13574 43012 13626
rect 43036 13574 43066 13626
rect 43066 13574 43078 13626
rect 43078 13574 43092 13626
rect 43116 13574 43130 13626
rect 43130 13574 43142 13626
rect 43142 13574 43172 13626
rect 43196 13574 43206 13626
rect 43206 13574 43252 13626
rect 42956 13572 43012 13574
rect 43036 13572 43092 13574
rect 43116 13572 43172 13574
rect 43196 13572 43252 13574
rect 42956 12538 43012 12540
rect 43036 12538 43092 12540
rect 43116 12538 43172 12540
rect 43196 12538 43252 12540
rect 42956 12486 43002 12538
rect 43002 12486 43012 12538
rect 43036 12486 43066 12538
rect 43066 12486 43078 12538
rect 43078 12486 43092 12538
rect 43116 12486 43130 12538
rect 43130 12486 43142 12538
rect 43142 12486 43172 12538
rect 43196 12486 43206 12538
rect 43206 12486 43252 12538
rect 42956 12484 43012 12486
rect 43036 12484 43092 12486
rect 43116 12484 43172 12486
rect 43196 12484 43252 12486
rect 42956 11450 43012 11452
rect 43036 11450 43092 11452
rect 43116 11450 43172 11452
rect 43196 11450 43252 11452
rect 42956 11398 43002 11450
rect 43002 11398 43012 11450
rect 43036 11398 43066 11450
rect 43066 11398 43078 11450
rect 43078 11398 43092 11450
rect 43116 11398 43130 11450
rect 43130 11398 43142 11450
rect 43142 11398 43172 11450
rect 43196 11398 43206 11450
rect 43206 11398 43252 11450
rect 42956 11396 43012 11398
rect 43036 11396 43092 11398
rect 43116 11396 43172 11398
rect 43196 11396 43252 11398
rect 42956 10362 43012 10364
rect 43036 10362 43092 10364
rect 43116 10362 43172 10364
rect 43196 10362 43252 10364
rect 42956 10310 43002 10362
rect 43002 10310 43012 10362
rect 43036 10310 43066 10362
rect 43066 10310 43078 10362
rect 43078 10310 43092 10362
rect 43116 10310 43130 10362
rect 43130 10310 43142 10362
rect 43142 10310 43172 10362
rect 43196 10310 43206 10362
rect 43206 10310 43252 10362
rect 42956 10308 43012 10310
rect 43036 10308 43092 10310
rect 43116 10308 43172 10310
rect 43196 10308 43252 10310
rect 42956 9274 43012 9276
rect 43036 9274 43092 9276
rect 43116 9274 43172 9276
rect 43196 9274 43252 9276
rect 42956 9222 43002 9274
rect 43002 9222 43012 9274
rect 43036 9222 43066 9274
rect 43066 9222 43078 9274
rect 43078 9222 43092 9274
rect 43116 9222 43130 9274
rect 43130 9222 43142 9274
rect 43142 9222 43172 9274
rect 43196 9222 43206 9274
rect 43206 9222 43252 9274
rect 42956 9220 43012 9222
rect 43036 9220 43092 9222
rect 43116 9220 43172 9222
rect 43196 9220 43252 9222
rect 42956 8186 43012 8188
rect 43036 8186 43092 8188
rect 43116 8186 43172 8188
rect 43196 8186 43252 8188
rect 42956 8134 43002 8186
rect 43002 8134 43012 8186
rect 43036 8134 43066 8186
rect 43066 8134 43078 8186
rect 43078 8134 43092 8186
rect 43116 8134 43130 8186
rect 43130 8134 43142 8186
rect 43142 8134 43172 8186
rect 43196 8134 43206 8186
rect 43206 8134 43252 8186
rect 42956 8132 43012 8134
rect 43036 8132 43092 8134
rect 43116 8132 43172 8134
rect 43196 8132 43252 8134
rect 42956 7098 43012 7100
rect 43036 7098 43092 7100
rect 43116 7098 43172 7100
rect 43196 7098 43252 7100
rect 42956 7046 43002 7098
rect 43002 7046 43012 7098
rect 43036 7046 43066 7098
rect 43066 7046 43078 7098
rect 43078 7046 43092 7098
rect 43116 7046 43130 7098
rect 43130 7046 43142 7098
rect 43142 7046 43172 7098
rect 43196 7046 43206 7098
rect 43206 7046 43252 7098
rect 42956 7044 43012 7046
rect 43036 7044 43092 7046
rect 43116 7044 43172 7046
rect 43196 7044 43252 7046
rect 42956 6010 43012 6012
rect 43036 6010 43092 6012
rect 43116 6010 43172 6012
rect 43196 6010 43252 6012
rect 42956 5958 43002 6010
rect 43002 5958 43012 6010
rect 43036 5958 43066 6010
rect 43066 5958 43078 6010
rect 43078 5958 43092 6010
rect 43116 5958 43130 6010
rect 43130 5958 43142 6010
rect 43142 5958 43172 6010
rect 43196 5958 43206 6010
rect 43206 5958 43252 6010
rect 42956 5956 43012 5958
rect 43036 5956 43092 5958
rect 43116 5956 43172 5958
rect 43196 5956 43252 5958
rect 42956 4922 43012 4924
rect 43036 4922 43092 4924
rect 43116 4922 43172 4924
rect 43196 4922 43252 4924
rect 42956 4870 43002 4922
rect 43002 4870 43012 4922
rect 43036 4870 43066 4922
rect 43066 4870 43078 4922
rect 43078 4870 43092 4922
rect 43116 4870 43130 4922
rect 43130 4870 43142 4922
rect 43142 4870 43172 4922
rect 43196 4870 43206 4922
rect 43206 4870 43252 4922
rect 42956 4868 43012 4870
rect 43036 4868 43092 4870
rect 43116 4868 43172 4870
rect 43196 4868 43252 4870
rect 42956 3834 43012 3836
rect 43036 3834 43092 3836
rect 43116 3834 43172 3836
rect 43196 3834 43252 3836
rect 42956 3782 43002 3834
rect 43002 3782 43012 3834
rect 43036 3782 43066 3834
rect 43066 3782 43078 3834
rect 43078 3782 43092 3834
rect 43116 3782 43130 3834
rect 43130 3782 43142 3834
rect 43142 3782 43172 3834
rect 43196 3782 43206 3834
rect 43206 3782 43252 3834
rect 42956 3780 43012 3782
rect 43036 3780 43092 3782
rect 43116 3780 43172 3782
rect 43196 3780 43252 3782
rect 42956 2746 43012 2748
rect 43036 2746 43092 2748
rect 43116 2746 43172 2748
rect 43196 2746 43252 2748
rect 42956 2694 43002 2746
rect 43002 2694 43012 2746
rect 43036 2694 43066 2746
rect 43066 2694 43078 2746
rect 43078 2694 43092 2746
rect 43116 2694 43130 2746
rect 43130 2694 43142 2746
rect 43142 2694 43172 2746
rect 43196 2694 43206 2746
rect 43206 2694 43252 2746
rect 42956 2692 43012 2694
rect 43036 2692 43092 2694
rect 43116 2692 43172 2694
rect 43196 2692 43252 2694
rect 44914 3440 44970 3496
rect 47956 31578 48012 31580
rect 48036 31578 48092 31580
rect 48116 31578 48172 31580
rect 48196 31578 48252 31580
rect 47956 31526 48002 31578
rect 48002 31526 48012 31578
rect 48036 31526 48066 31578
rect 48066 31526 48078 31578
rect 48078 31526 48092 31578
rect 48116 31526 48130 31578
rect 48130 31526 48142 31578
rect 48142 31526 48172 31578
rect 48196 31526 48206 31578
rect 48206 31526 48252 31578
rect 47956 31524 48012 31526
rect 48036 31524 48092 31526
rect 48116 31524 48172 31526
rect 48196 31524 48252 31526
rect 47956 30490 48012 30492
rect 48036 30490 48092 30492
rect 48116 30490 48172 30492
rect 48196 30490 48252 30492
rect 47956 30438 48002 30490
rect 48002 30438 48012 30490
rect 48036 30438 48066 30490
rect 48066 30438 48078 30490
rect 48078 30438 48092 30490
rect 48116 30438 48130 30490
rect 48130 30438 48142 30490
rect 48142 30438 48172 30490
rect 48196 30438 48206 30490
rect 48206 30438 48252 30490
rect 47956 30436 48012 30438
rect 48036 30436 48092 30438
rect 48116 30436 48172 30438
rect 48196 30436 48252 30438
rect 47956 29402 48012 29404
rect 48036 29402 48092 29404
rect 48116 29402 48172 29404
rect 48196 29402 48252 29404
rect 47956 29350 48002 29402
rect 48002 29350 48012 29402
rect 48036 29350 48066 29402
rect 48066 29350 48078 29402
rect 48078 29350 48092 29402
rect 48116 29350 48130 29402
rect 48130 29350 48142 29402
rect 48142 29350 48172 29402
rect 48196 29350 48206 29402
rect 48206 29350 48252 29402
rect 47956 29348 48012 29350
rect 48036 29348 48092 29350
rect 48116 29348 48172 29350
rect 48196 29348 48252 29350
rect 47956 28314 48012 28316
rect 48036 28314 48092 28316
rect 48116 28314 48172 28316
rect 48196 28314 48252 28316
rect 47956 28262 48002 28314
rect 48002 28262 48012 28314
rect 48036 28262 48066 28314
rect 48066 28262 48078 28314
rect 48078 28262 48092 28314
rect 48116 28262 48130 28314
rect 48130 28262 48142 28314
rect 48142 28262 48172 28314
rect 48196 28262 48206 28314
rect 48206 28262 48252 28314
rect 47956 28260 48012 28262
rect 48036 28260 48092 28262
rect 48116 28260 48172 28262
rect 48196 28260 48252 28262
rect 47956 27226 48012 27228
rect 48036 27226 48092 27228
rect 48116 27226 48172 27228
rect 48196 27226 48252 27228
rect 47956 27174 48002 27226
rect 48002 27174 48012 27226
rect 48036 27174 48066 27226
rect 48066 27174 48078 27226
rect 48078 27174 48092 27226
rect 48116 27174 48130 27226
rect 48130 27174 48142 27226
rect 48142 27174 48172 27226
rect 48196 27174 48206 27226
rect 48206 27174 48252 27226
rect 47956 27172 48012 27174
rect 48036 27172 48092 27174
rect 48116 27172 48172 27174
rect 48196 27172 48252 27174
rect 47956 26138 48012 26140
rect 48036 26138 48092 26140
rect 48116 26138 48172 26140
rect 48196 26138 48252 26140
rect 47956 26086 48002 26138
rect 48002 26086 48012 26138
rect 48036 26086 48066 26138
rect 48066 26086 48078 26138
rect 48078 26086 48092 26138
rect 48116 26086 48130 26138
rect 48130 26086 48142 26138
rect 48142 26086 48172 26138
rect 48196 26086 48206 26138
rect 48206 26086 48252 26138
rect 47956 26084 48012 26086
rect 48036 26084 48092 26086
rect 48116 26084 48172 26086
rect 48196 26084 48252 26086
rect 47956 25050 48012 25052
rect 48036 25050 48092 25052
rect 48116 25050 48172 25052
rect 48196 25050 48252 25052
rect 47956 24998 48002 25050
rect 48002 24998 48012 25050
rect 48036 24998 48066 25050
rect 48066 24998 48078 25050
rect 48078 24998 48092 25050
rect 48116 24998 48130 25050
rect 48130 24998 48142 25050
rect 48142 24998 48172 25050
rect 48196 24998 48206 25050
rect 48206 24998 48252 25050
rect 47956 24996 48012 24998
rect 48036 24996 48092 24998
rect 48116 24996 48172 24998
rect 48196 24996 48252 24998
rect 47956 23962 48012 23964
rect 48036 23962 48092 23964
rect 48116 23962 48172 23964
rect 48196 23962 48252 23964
rect 47956 23910 48002 23962
rect 48002 23910 48012 23962
rect 48036 23910 48066 23962
rect 48066 23910 48078 23962
rect 48078 23910 48092 23962
rect 48116 23910 48130 23962
rect 48130 23910 48142 23962
rect 48142 23910 48172 23962
rect 48196 23910 48206 23962
rect 48206 23910 48252 23962
rect 47956 23908 48012 23910
rect 48036 23908 48092 23910
rect 48116 23908 48172 23910
rect 48196 23908 48252 23910
rect 47956 22874 48012 22876
rect 48036 22874 48092 22876
rect 48116 22874 48172 22876
rect 48196 22874 48252 22876
rect 47956 22822 48002 22874
rect 48002 22822 48012 22874
rect 48036 22822 48066 22874
rect 48066 22822 48078 22874
rect 48078 22822 48092 22874
rect 48116 22822 48130 22874
rect 48130 22822 48142 22874
rect 48142 22822 48172 22874
rect 48196 22822 48206 22874
rect 48206 22822 48252 22874
rect 47956 22820 48012 22822
rect 48036 22820 48092 22822
rect 48116 22820 48172 22822
rect 48196 22820 48252 22822
rect 47956 21786 48012 21788
rect 48036 21786 48092 21788
rect 48116 21786 48172 21788
rect 48196 21786 48252 21788
rect 47956 21734 48002 21786
rect 48002 21734 48012 21786
rect 48036 21734 48066 21786
rect 48066 21734 48078 21786
rect 48078 21734 48092 21786
rect 48116 21734 48130 21786
rect 48130 21734 48142 21786
rect 48142 21734 48172 21786
rect 48196 21734 48206 21786
rect 48206 21734 48252 21786
rect 47956 21732 48012 21734
rect 48036 21732 48092 21734
rect 48116 21732 48172 21734
rect 48196 21732 48252 21734
rect 47956 20698 48012 20700
rect 48036 20698 48092 20700
rect 48116 20698 48172 20700
rect 48196 20698 48252 20700
rect 47956 20646 48002 20698
rect 48002 20646 48012 20698
rect 48036 20646 48066 20698
rect 48066 20646 48078 20698
rect 48078 20646 48092 20698
rect 48116 20646 48130 20698
rect 48130 20646 48142 20698
rect 48142 20646 48172 20698
rect 48196 20646 48206 20698
rect 48206 20646 48252 20698
rect 47956 20644 48012 20646
rect 48036 20644 48092 20646
rect 48116 20644 48172 20646
rect 48196 20644 48252 20646
rect 47956 19610 48012 19612
rect 48036 19610 48092 19612
rect 48116 19610 48172 19612
rect 48196 19610 48252 19612
rect 47956 19558 48002 19610
rect 48002 19558 48012 19610
rect 48036 19558 48066 19610
rect 48066 19558 48078 19610
rect 48078 19558 48092 19610
rect 48116 19558 48130 19610
rect 48130 19558 48142 19610
rect 48142 19558 48172 19610
rect 48196 19558 48206 19610
rect 48206 19558 48252 19610
rect 47956 19556 48012 19558
rect 48036 19556 48092 19558
rect 48116 19556 48172 19558
rect 48196 19556 48252 19558
rect 47956 18522 48012 18524
rect 48036 18522 48092 18524
rect 48116 18522 48172 18524
rect 48196 18522 48252 18524
rect 47956 18470 48002 18522
rect 48002 18470 48012 18522
rect 48036 18470 48066 18522
rect 48066 18470 48078 18522
rect 48078 18470 48092 18522
rect 48116 18470 48130 18522
rect 48130 18470 48142 18522
rect 48142 18470 48172 18522
rect 48196 18470 48206 18522
rect 48206 18470 48252 18522
rect 47956 18468 48012 18470
rect 48036 18468 48092 18470
rect 48116 18468 48172 18470
rect 48196 18468 48252 18470
rect 47956 17434 48012 17436
rect 48036 17434 48092 17436
rect 48116 17434 48172 17436
rect 48196 17434 48252 17436
rect 47956 17382 48002 17434
rect 48002 17382 48012 17434
rect 48036 17382 48066 17434
rect 48066 17382 48078 17434
rect 48078 17382 48092 17434
rect 48116 17382 48130 17434
rect 48130 17382 48142 17434
rect 48142 17382 48172 17434
rect 48196 17382 48206 17434
rect 48206 17382 48252 17434
rect 47956 17380 48012 17382
rect 48036 17380 48092 17382
rect 48116 17380 48172 17382
rect 48196 17380 48252 17382
rect 47956 16346 48012 16348
rect 48036 16346 48092 16348
rect 48116 16346 48172 16348
rect 48196 16346 48252 16348
rect 47956 16294 48002 16346
rect 48002 16294 48012 16346
rect 48036 16294 48066 16346
rect 48066 16294 48078 16346
rect 48078 16294 48092 16346
rect 48116 16294 48130 16346
rect 48130 16294 48142 16346
rect 48142 16294 48172 16346
rect 48196 16294 48206 16346
rect 48206 16294 48252 16346
rect 47956 16292 48012 16294
rect 48036 16292 48092 16294
rect 48116 16292 48172 16294
rect 48196 16292 48252 16294
rect 47956 15258 48012 15260
rect 48036 15258 48092 15260
rect 48116 15258 48172 15260
rect 48196 15258 48252 15260
rect 47956 15206 48002 15258
rect 48002 15206 48012 15258
rect 48036 15206 48066 15258
rect 48066 15206 48078 15258
rect 48078 15206 48092 15258
rect 48116 15206 48130 15258
rect 48130 15206 48142 15258
rect 48142 15206 48172 15258
rect 48196 15206 48206 15258
rect 48206 15206 48252 15258
rect 47956 15204 48012 15206
rect 48036 15204 48092 15206
rect 48116 15204 48172 15206
rect 48196 15204 48252 15206
rect 47956 14170 48012 14172
rect 48036 14170 48092 14172
rect 48116 14170 48172 14172
rect 48196 14170 48252 14172
rect 47956 14118 48002 14170
rect 48002 14118 48012 14170
rect 48036 14118 48066 14170
rect 48066 14118 48078 14170
rect 48078 14118 48092 14170
rect 48116 14118 48130 14170
rect 48130 14118 48142 14170
rect 48142 14118 48172 14170
rect 48196 14118 48206 14170
rect 48206 14118 48252 14170
rect 47956 14116 48012 14118
rect 48036 14116 48092 14118
rect 48116 14116 48172 14118
rect 48196 14116 48252 14118
rect 47956 13082 48012 13084
rect 48036 13082 48092 13084
rect 48116 13082 48172 13084
rect 48196 13082 48252 13084
rect 47956 13030 48002 13082
rect 48002 13030 48012 13082
rect 48036 13030 48066 13082
rect 48066 13030 48078 13082
rect 48078 13030 48092 13082
rect 48116 13030 48130 13082
rect 48130 13030 48142 13082
rect 48142 13030 48172 13082
rect 48196 13030 48206 13082
rect 48206 13030 48252 13082
rect 47956 13028 48012 13030
rect 48036 13028 48092 13030
rect 48116 13028 48172 13030
rect 48196 13028 48252 13030
rect 47956 11994 48012 11996
rect 48036 11994 48092 11996
rect 48116 11994 48172 11996
rect 48196 11994 48252 11996
rect 47956 11942 48002 11994
rect 48002 11942 48012 11994
rect 48036 11942 48066 11994
rect 48066 11942 48078 11994
rect 48078 11942 48092 11994
rect 48116 11942 48130 11994
rect 48130 11942 48142 11994
rect 48142 11942 48172 11994
rect 48196 11942 48206 11994
rect 48206 11942 48252 11994
rect 47956 11940 48012 11942
rect 48036 11940 48092 11942
rect 48116 11940 48172 11942
rect 48196 11940 48252 11942
rect 47956 10906 48012 10908
rect 48036 10906 48092 10908
rect 48116 10906 48172 10908
rect 48196 10906 48252 10908
rect 47956 10854 48002 10906
rect 48002 10854 48012 10906
rect 48036 10854 48066 10906
rect 48066 10854 48078 10906
rect 48078 10854 48092 10906
rect 48116 10854 48130 10906
rect 48130 10854 48142 10906
rect 48142 10854 48172 10906
rect 48196 10854 48206 10906
rect 48206 10854 48252 10906
rect 47956 10852 48012 10854
rect 48036 10852 48092 10854
rect 48116 10852 48172 10854
rect 48196 10852 48252 10854
rect 47956 9818 48012 9820
rect 48036 9818 48092 9820
rect 48116 9818 48172 9820
rect 48196 9818 48252 9820
rect 47956 9766 48002 9818
rect 48002 9766 48012 9818
rect 48036 9766 48066 9818
rect 48066 9766 48078 9818
rect 48078 9766 48092 9818
rect 48116 9766 48130 9818
rect 48130 9766 48142 9818
rect 48142 9766 48172 9818
rect 48196 9766 48206 9818
rect 48206 9766 48252 9818
rect 47956 9764 48012 9766
rect 48036 9764 48092 9766
rect 48116 9764 48172 9766
rect 48196 9764 48252 9766
rect 48502 41012 48504 41032
rect 48504 41012 48556 41032
rect 48556 41012 48558 41032
rect 48502 40976 48558 41012
rect 48778 40588 48834 40624
rect 48778 40568 48780 40588
rect 48780 40568 48832 40588
rect 48832 40568 48834 40588
rect 48502 40296 48558 40352
rect 48502 39616 48558 39672
rect 48502 38936 48558 38992
rect 49146 45736 49202 45792
rect 48778 39500 48834 39536
rect 48778 39480 48780 39500
rect 48780 39480 48832 39500
rect 48832 39480 48834 39500
rect 48502 36896 48558 36952
rect 49330 46416 49386 46472
rect 49330 45056 49386 45112
rect 49330 38292 49332 38312
rect 49332 38292 49384 38312
rect 49384 38292 49386 38312
rect 49330 38256 49386 38292
rect 49330 37576 49386 37632
rect 49330 36216 49386 36272
rect 49330 35536 49386 35592
rect 49330 34856 49386 34912
rect 49330 34176 49386 34232
rect 49238 33904 49294 33960
rect 48502 32136 48558 32192
rect 48502 31456 48558 31512
rect 48502 30776 48558 30832
rect 49330 33496 49386 33552
rect 49330 32852 49332 32872
rect 49332 32852 49384 32872
rect 49384 32852 49386 32872
rect 49330 32816 49386 32852
rect 49330 30096 49386 30152
rect 48502 29416 48558 29472
rect 49330 28736 49386 28792
rect 49330 28056 49386 28112
rect 48502 27412 48504 27432
rect 48504 27412 48556 27432
rect 48556 27412 48558 27432
rect 48502 27376 48558 27412
rect 48502 26696 48558 26752
rect 48502 26016 48558 26072
rect 49330 25336 49386 25392
rect 49146 24692 49148 24712
rect 49148 24692 49200 24712
rect 49200 24692 49202 24712
rect 49146 24656 49202 24692
rect 49146 23976 49202 24032
rect 49146 23296 49202 23352
rect 49146 22616 49202 22672
rect 49146 21972 49148 21992
rect 49148 21972 49200 21992
rect 49200 21972 49202 21992
rect 49146 21936 49202 21972
rect 49146 21256 49202 21312
rect 49146 20576 49202 20632
rect 49146 19896 49202 19952
rect 49146 19216 49202 19272
rect 49146 18536 49202 18592
rect 49146 17856 49202 17912
rect 49146 17176 49202 17232
rect 49146 16516 49202 16552
rect 49146 16496 49148 16516
rect 49148 16496 49200 16516
rect 49200 16496 49202 16516
rect 49146 15816 49202 15872
rect 49146 15136 49202 15192
rect 49146 14456 49202 14512
rect 49146 13812 49148 13832
rect 49148 13812 49200 13832
rect 49200 13812 49202 13832
rect 49146 13776 49202 13812
rect 49146 13096 49202 13152
rect 49146 12416 49202 12472
rect 49146 11736 49202 11792
rect 49146 11092 49148 11112
rect 49148 11092 49200 11112
rect 49200 11092 49202 11112
rect 49146 11056 49202 11092
rect 49146 10376 49202 10432
rect 49146 9696 49202 9752
rect 49146 9016 49202 9072
rect 47956 8730 48012 8732
rect 48036 8730 48092 8732
rect 48116 8730 48172 8732
rect 48196 8730 48252 8732
rect 47956 8678 48002 8730
rect 48002 8678 48012 8730
rect 48036 8678 48066 8730
rect 48066 8678 48078 8730
rect 48078 8678 48092 8730
rect 48116 8678 48130 8730
rect 48130 8678 48142 8730
rect 48142 8678 48172 8730
rect 48196 8678 48206 8730
rect 48206 8678 48252 8730
rect 47956 8676 48012 8678
rect 48036 8676 48092 8678
rect 48116 8676 48172 8678
rect 48196 8676 48252 8678
rect 47956 7642 48012 7644
rect 48036 7642 48092 7644
rect 48116 7642 48172 7644
rect 48196 7642 48252 7644
rect 47956 7590 48002 7642
rect 48002 7590 48012 7642
rect 48036 7590 48066 7642
rect 48066 7590 48078 7642
rect 48078 7590 48092 7642
rect 48116 7590 48130 7642
rect 48130 7590 48142 7642
rect 48142 7590 48172 7642
rect 48196 7590 48206 7642
rect 48206 7590 48252 7642
rect 47956 7588 48012 7590
rect 48036 7588 48092 7590
rect 48116 7588 48172 7590
rect 48196 7588 48252 7590
rect 49146 8372 49148 8392
rect 49148 8372 49200 8392
rect 49200 8372 49202 8392
rect 49146 8336 49202 8372
rect 49146 7656 49202 7712
rect 49146 6976 49202 7032
rect 47956 6554 48012 6556
rect 48036 6554 48092 6556
rect 48116 6554 48172 6556
rect 48196 6554 48252 6556
rect 47956 6502 48002 6554
rect 48002 6502 48012 6554
rect 48036 6502 48066 6554
rect 48066 6502 48078 6554
rect 48078 6502 48092 6554
rect 48116 6502 48130 6554
rect 48130 6502 48142 6554
rect 48142 6502 48172 6554
rect 48196 6502 48206 6554
rect 48206 6502 48252 6554
rect 47956 6500 48012 6502
rect 48036 6500 48092 6502
rect 48116 6500 48172 6502
rect 48196 6500 48252 6502
rect 47956 5466 48012 5468
rect 48036 5466 48092 5468
rect 48116 5466 48172 5468
rect 48196 5466 48252 5468
rect 47956 5414 48002 5466
rect 48002 5414 48012 5466
rect 48036 5414 48066 5466
rect 48066 5414 48078 5466
rect 48078 5414 48092 5466
rect 48116 5414 48130 5466
rect 48130 5414 48142 5466
rect 48142 5414 48172 5466
rect 48196 5414 48206 5466
rect 48206 5414 48252 5466
rect 47956 5412 48012 5414
rect 48036 5412 48092 5414
rect 48116 5412 48172 5414
rect 48196 5412 48252 5414
rect 47956 4378 48012 4380
rect 48036 4378 48092 4380
rect 48116 4378 48172 4380
rect 48196 4378 48252 4380
rect 47956 4326 48002 4378
rect 48002 4326 48012 4378
rect 48036 4326 48066 4378
rect 48066 4326 48078 4378
rect 48078 4326 48092 4378
rect 48116 4326 48130 4378
rect 48130 4326 48142 4378
rect 48142 4326 48172 4378
rect 48196 4326 48206 4378
rect 48206 4326 48252 4378
rect 47956 4324 48012 4326
rect 48036 4324 48092 4326
rect 48116 4324 48172 4326
rect 48196 4324 48252 4326
rect 47956 3290 48012 3292
rect 48036 3290 48092 3292
rect 48116 3290 48172 3292
rect 48196 3290 48252 3292
rect 47956 3238 48002 3290
rect 48002 3238 48012 3290
rect 48036 3238 48066 3290
rect 48066 3238 48078 3290
rect 48078 3238 48092 3290
rect 48116 3238 48130 3290
rect 48130 3238 48142 3290
rect 48142 3238 48172 3290
rect 48196 3238 48206 3290
rect 48206 3238 48252 3290
rect 47956 3236 48012 3238
rect 48036 3236 48092 3238
rect 48116 3236 48172 3238
rect 48196 3236 48252 3238
rect 47956 2202 48012 2204
rect 48036 2202 48092 2204
rect 48116 2202 48172 2204
rect 48196 2202 48252 2204
rect 47956 2150 48002 2202
rect 48002 2150 48012 2202
rect 48036 2150 48066 2202
rect 48066 2150 48078 2202
rect 48078 2150 48092 2202
rect 48116 2150 48130 2202
rect 48130 2150 48142 2202
rect 48142 2150 48172 2202
rect 48196 2150 48206 2202
rect 48206 2150 48252 2202
rect 47956 2148 48012 2150
rect 48036 2148 48092 2150
rect 48116 2148 48172 2150
rect 48196 2148 48252 2150
rect 49146 6296 49202 6352
rect 49146 5652 49148 5672
rect 49148 5652 49200 5672
rect 49200 5652 49202 5672
rect 49146 5616 49202 5652
rect 49330 4972 49332 4992
rect 49332 4972 49384 4992
rect 49384 4972 49386 4992
rect 49330 4936 49386 4972
rect 49146 4256 49202 4312
<< metal3 >>
rect 0 55042 800 55072
rect 2773 55042 2839 55045
rect 0 55040 2839 55042
rect 0 54984 2778 55040
rect 2834 54984 2839 55040
rect 0 54982 2839 54984
rect 0 54952 800 54982
rect 2773 54979 2839 54982
rect 7946 54432 8262 54433
rect 7946 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8262 54432
rect 7946 54367 8262 54368
rect 17946 54432 18262 54433
rect 17946 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18262 54432
rect 17946 54367 18262 54368
rect 27946 54432 28262 54433
rect 27946 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28262 54432
rect 27946 54367 28262 54368
rect 37946 54432 38262 54433
rect 37946 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38262 54432
rect 37946 54367 38262 54368
rect 47946 54432 48262 54433
rect 47946 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48262 54432
rect 47946 54367 48262 54368
rect 24945 53954 25011 53957
rect 25078 53954 25084 53956
rect 24945 53952 25084 53954
rect 24945 53896 24950 53952
rect 25006 53896 25084 53952
rect 24945 53894 25084 53896
rect 24945 53891 25011 53894
rect 25078 53892 25084 53894
rect 25148 53892 25154 53956
rect 2946 53888 3262 53889
rect 2946 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3262 53888
rect 2946 53823 3262 53824
rect 12946 53888 13262 53889
rect 12946 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13262 53888
rect 12946 53823 13262 53824
rect 22946 53888 23262 53889
rect 22946 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23262 53888
rect 22946 53823 23262 53824
rect 32946 53888 33262 53889
rect 32946 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33262 53888
rect 32946 53823 33262 53824
rect 42946 53888 43262 53889
rect 42946 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43262 53888
rect 42946 53823 43262 53824
rect 7946 53344 8262 53345
rect 7946 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8262 53344
rect 7946 53279 8262 53280
rect 17946 53344 18262 53345
rect 17946 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18262 53344
rect 17946 53279 18262 53280
rect 27946 53344 28262 53345
rect 27946 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28262 53344
rect 27946 53279 28262 53280
rect 37946 53344 38262 53345
rect 37946 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38262 53344
rect 37946 53279 38262 53280
rect 47946 53344 48262 53345
rect 47946 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48262 53344
rect 47946 53279 48262 53280
rect 2946 52800 3262 52801
rect 0 52730 800 52760
rect 2946 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3262 52800
rect 2946 52735 3262 52736
rect 12946 52800 13262 52801
rect 12946 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13262 52800
rect 12946 52735 13262 52736
rect 22946 52800 23262 52801
rect 22946 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23262 52800
rect 22946 52735 23262 52736
rect 32946 52800 33262 52801
rect 32946 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33262 52800
rect 32946 52735 33262 52736
rect 42946 52800 43262 52801
rect 42946 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43262 52800
rect 42946 52735 43262 52736
rect 933 52730 999 52733
rect 0 52728 999 52730
rect 0 52672 938 52728
rect 994 52672 999 52728
rect 0 52670 999 52672
rect 0 52640 800 52670
rect 933 52667 999 52670
rect 49325 52594 49391 52597
rect 50200 52594 51000 52624
rect 49325 52592 51000 52594
rect 49325 52536 49330 52592
rect 49386 52536 51000 52592
rect 49325 52534 51000 52536
rect 49325 52531 49391 52534
rect 50200 52504 51000 52534
rect 7946 52256 8262 52257
rect 7946 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8262 52256
rect 7946 52191 8262 52192
rect 17946 52256 18262 52257
rect 17946 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18262 52256
rect 17946 52191 18262 52192
rect 27946 52256 28262 52257
rect 27946 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28262 52256
rect 27946 52191 28262 52192
rect 37946 52256 38262 52257
rect 37946 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38262 52256
rect 37946 52191 38262 52192
rect 47946 52256 48262 52257
rect 47946 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48262 52256
rect 47946 52191 48262 52192
rect 49049 51914 49115 51917
rect 50200 51914 51000 51944
rect 49049 51912 51000 51914
rect 49049 51856 49054 51912
rect 49110 51856 51000 51912
rect 49049 51854 51000 51856
rect 49049 51851 49115 51854
rect 50200 51824 51000 51854
rect 2946 51712 3262 51713
rect 2946 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3262 51712
rect 2946 51647 3262 51648
rect 12946 51712 13262 51713
rect 12946 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13262 51712
rect 12946 51647 13262 51648
rect 22946 51712 23262 51713
rect 22946 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23262 51712
rect 22946 51647 23262 51648
rect 32946 51712 33262 51713
rect 32946 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33262 51712
rect 32946 51647 33262 51648
rect 42946 51712 43262 51713
rect 42946 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43262 51712
rect 42946 51647 43262 51648
rect 49049 51234 49115 51237
rect 50200 51234 51000 51264
rect 49049 51232 51000 51234
rect 49049 51176 49054 51232
rect 49110 51176 51000 51232
rect 49049 51174 51000 51176
rect 49049 51171 49115 51174
rect 7946 51168 8262 51169
rect 7946 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8262 51168
rect 7946 51103 8262 51104
rect 17946 51168 18262 51169
rect 17946 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18262 51168
rect 17946 51103 18262 51104
rect 27946 51168 28262 51169
rect 27946 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28262 51168
rect 27946 51103 28262 51104
rect 37946 51168 38262 51169
rect 37946 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38262 51168
rect 37946 51103 38262 51104
rect 47946 51168 48262 51169
rect 47946 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48262 51168
rect 50200 51144 51000 51174
rect 47946 51103 48262 51104
rect 2946 50624 3262 50625
rect 2946 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3262 50624
rect 2946 50559 3262 50560
rect 12946 50624 13262 50625
rect 12946 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13262 50624
rect 12946 50559 13262 50560
rect 22946 50624 23262 50625
rect 22946 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23262 50624
rect 22946 50559 23262 50560
rect 32946 50624 33262 50625
rect 32946 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33262 50624
rect 32946 50559 33262 50560
rect 42946 50624 43262 50625
rect 42946 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43262 50624
rect 42946 50559 43262 50560
rect 48957 50554 49023 50557
rect 50200 50554 51000 50584
rect 48957 50552 51000 50554
rect 48957 50496 48962 50552
rect 49018 50496 51000 50552
rect 48957 50494 51000 50496
rect 48957 50491 49023 50494
rect 50200 50464 51000 50494
rect 0 50418 800 50448
rect 933 50418 999 50421
rect 0 50416 999 50418
rect 0 50360 938 50416
rect 994 50360 999 50416
rect 0 50358 999 50360
rect 0 50328 800 50358
rect 933 50355 999 50358
rect 7946 50080 8262 50081
rect 7946 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8262 50080
rect 7946 50015 8262 50016
rect 17946 50080 18262 50081
rect 17946 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18262 50080
rect 17946 50015 18262 50016
rect 27946 50080 28262 50081
rect 27946 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28262 50080
rect 27946 50015 28262 50016
rect 37946 50080 38262 50081
rect 37946 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38262 50080
rect 37946 50015 38262 50016
rect 47946 50080 48262 50081
rect 47946 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48262 50080
rect 47946 50015 48262 50016
rect 49049 49874 49115 49877
rect 50200 49874 51000 49904
rect 49049 49872 51000 49874
rect 49049 49816 49054 49872
rect 49110 49816 51000 49872
rect 49049 49814 51000 49816
rect 49049 49811 49115 49814
rect 50200 49784 51000 49814
rect 2946 49536 3262 49537
rect 2946 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3262 49536
rect 2946 49471 3262 49472
rect 12946 49536 13262 49537
rect 12946 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13262 49536
rect 12946 49471 13262 49472
rect 22946 49536 23262 49537
rect 22946 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23262 49536
rect 22946 49471 23262 49472
rect 32946 49536 33262 49537
rect 32946 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33262 49536
rect 32946 49471 33262 49472
rect 42946 49536 43262 49537
rect 42946 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43262 49536
rect 42946 49471 43262 49472
rect 49141 49194 49207 49197
rect 50200 49194 51000 49224
rect 49141 49192 51000 49194
rect 49141 49136 49146 49192
rect 49202 49136 51000 49192
rect 49141 49134 51000 49136
rect 49141 49131 49207 49134
rect 50200 49104 51000 49134
rect 7946 48992 8262 48993
rect 7946 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8262 48992
rect 7946 48927 8262 48928
rect 17946 48992 18262 48993
rect 17946 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18262 48992
rect 17946 48927 18262 48928
rect 27946 48992 28262 48993
rect 27946 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28262 48992
rect 27946 48927 28262 48928
rect 37946 48992 38262 48993
rect 37946 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38262 48992
rect 37946 48927 38262 48928
rect 47946 48992 48262 48993
rect 47946 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48262 48992
rect 47946 48927 48262 48928
rect 49233 48514 49299 48517
rect 50200 48514 51000 48544
rect 49233 48512 51000 48514
rect 49233 48456 49238 48512
rect 49294 48456 51000 48512
rect 49233 48454 51000 48456
rect 49233 48451 49299 48454
rect 2946 48448 3262 48449
rect 2946 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3262 48448
rect 2946 48383 3262 48384
rect 12946 48448 13262 48449
rect 12946 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13262 48448
rect 12946 48383 13262 48384
rect 22946 48448 23262 48449
rect 22946 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23262 48448
rect 22946 48383 23262 48384
rect 32946 48448 33262 48449
rect 32946 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33262 48448
rect 32946 48383 33262 48384
rect 42946 48448 43262 48449
rect 42946 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43262 48448
rect 50200 48424 51000 48454
rect 42946 48383 43262 48384
rect 0 48106 800 48136
rect 933 48106 999 48109
rect 0 48104 999 48106
rect 0 48048 938 48104
rect 994 48048 999 48104
rect 0 48046 999 48048
rect 0 48016 800 48046
rect 933 48043 999 48046
rect 7946 47904 8262 47905
rect 7946 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8262 47904
rect 7946 47839 8262 47840
rect 17946 47904 18262 47905
rect 17946 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18262 47904
rect 17946 47839 18262 47840
rect 27946 47904 28262 47905
rect 27946 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28262 47904
rect 27946 47839 28262 47840
rect 37946 47904 38262 47905
rect 37946 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38262 47904
rect 37946 47839 38262 47840
rect 47946 47904 48262 47905
rect 47946 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48262 47904
rect 47946 47839 48262 47840
rect 49049 47834 49115 47837
rect 50200 47834 51000 47864
rect 49049 47832 51000 47834
rect 49049 47776 49054 47832
rect 49110 47776 51000 47832
rect 49049 47774 51000 47776
rect 49049 47771 49115 47774
rect 50200 47744 51000 47774
rect 2946 47360 3262 47361
rect 2946 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3262 47360
rect 2946 47295 3262 47296
rect 12946 47360 13262 47361
rect 12946 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13262 47360
rect 12946 47295 13262 47296
rect 22946 47360 23262 47361
rect 22946 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23262 47360
rect 22946 47295 23262 47296
rect 32946 47360 33262 47361
rect 32946 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33262 47360
rect 32946 47295 33262 47296
rect 42946 47360 43262 47361
rect 42946 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43262 47360
rect 42946 47295 43262 47296
rect 49049 47154 49115 47157
rect 50200 47154 51000 47184
rect 49049 47152 51000 47154
rect 49049 47096 49054 47152
rect 49110 47096 51000 47152
rect 49049 47094 51000 47096
rect 49049 47091 49115 47094
rect 50200 47064 51000 47094
rect 7946 46816 8262 46817
rect 7946 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8262 46816
rect 7946 46751 8262 46752
rect 17946 46816 18262 46817
rect 17946 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18262 46816
rect 17946 46751 18262 46752
rect 27946 46816 28262 46817
rect 27946 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28262 46816
rect 27946 46751 28262 46752
rect 37946 46816 38262 46817
rect 37946 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38262 46816
rect 37946 46751 38262 46752
rect 47946 46816 48262 46817
rect 47946 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48262 46816
rect 47946 46751 48262 46752
rect 49325 46474 49391 46477
rect 50200 46474 51000 46504
rect 49325 46472 51000 46474
rect 49325 46416 49330 46472
rect 49386 46416 51000 46472
rect 49325 46414 51000 46416
rect 49325 46411 49391 46414
rect 50200 46384 51000 46414
rect 2946 46272 3262 46273
rect 2946 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3262 46272
rect 2946 46207 3262 46208
rect 12946 46272 13262 46273
rect 12946 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13262 46272
rect 12946 46207 13262 46208
rect 22946 46272 23262 46273
rect 22946 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23262 46272
rect 22946 46207 23262 46208
rect 32946 46272 33262 46273
rect 32946 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33262 46272
rect 32946 46207 33262 46208
rect 42946 46272 43262 46273
rect 42946 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43262 46272
rect 42946 46207 43262 46208
rect 0 45794 800 45824
rect 933 45794 999 45797
rect 0 45792 999 45794
rect 0 45736 938 45792
rect 994 45736 999 45792
rect 0 45734 999 45736
rect 0 45704 800 45734
rect 933 45731 999 45734
rect 49141 45794 49207 45797
rect 50200 45794 51000 45824
rect 49141 45792 51000 45794
rect 49141 45736 49146 45792
rect 49202 45736 51000 45792
rect 49141 45734 51000 45736
rect 49141 45731 49207 45734
rect 7946 45728 8262 45729
rect 7946 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8262 45728
rect 7946 45663 8262 45664
rect 17946 45728 18262 45729
rect 17946 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18262 45728
rect 17946 45663 18262 45664
rect 27946 45728 28262 45729
rect 27946 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28262 45728
rect 27946 45663 28262 45664
rect 37946 45728 38262 45729
rect 37946 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38262 45728
rect 37946 45663 38262 45664
rect 47946 45728 48262 45729
rect 47946 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48262 45728
rect 50200 45704 51000 45734
rect 47946 45663 48262 45664
rect 2946 45184 3262 45185
rect 2946 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3262 45184
rect 2946 45119 3262 45120
rect 12946 45184 13262 45185
rect 12946 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13262 45184
rect 12946 45119 13262 45120
rect 22946 45184 23262 45185
rect 22946 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23262 45184
rect 22946 45119 23262 45120
rect 32946 45184 33262 45185
rect 32946 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33262 45184
rect 32946 45119 33262 45120
rect 42946 45184 43262 45185
rect 42946 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43262 45184
rect 42946 45119 43262 45120
rect 49325 45114 49391 45117
rect 50200 45114 51000 45144
rect 49325 45112 51000 45114
rect 49325 45056 49330 45112
rect 49386 45056 51000 45112
rect 49325 45054 51000 45056
rect 49325 45051 49391 45054
rect 50200 45024 51000 45054
rect 7946 44640 8262 44641
rect 7946 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8262 44640
rect 7946 44575 8262 44576
rect 17946 44640 18262 44641
rect 17946 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18262 44640
rect 17946 44575 18262 44576
rect 27946 44640 28262 44641
rect 27946 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28262 44640
rect 27946 44575 28262 44576
rect 37946 44640 38262 44641
rect 37946 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38262 44640
rect 37946 44575 38262 44576
rect 47946 44640 48262 44641
rect 47946 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48262 44640
rect 47946 44575 48262 44576
rect 48497 44434 48563 44437
rect 50200 44434 51000 44464
rect 48497 44432 51000 44434
rect 48497 44376 48502 44432
rect 48558 44376 51000 44432
rect 48497 44374 51000 44376
rect 48497 44371 48563 44374
rect 50200 44344 51000 44374
rect 2946 44096 3262 44097
rect 2946 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3262 44096
rect 2946 44031 3262 44032
rect 12946 44096 13262 44097
rect 12946 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13262 44096
rect 12946 44031 13262 44032
rect 22946 44096 23262 44097
rect 22946 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23262 44096
rect 22946 44031 23262 44032
rect 32946 44096 33262 44097
rect 32946 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33262 44096
rect 32946 44031 33262 44032
rect 42946 44096 43262 44097
rect 42946 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43262 44096
rect 42946 44031 43262 44032
rect 48497 43754 48563 43757
rect 50200 43754 51000 43784
rect 48497 43752 51000 43754
rect 48497 43696 48502 43752
rect 48558 43696 51000 43752
rect 48497 43694 51000 43696
rect 48497 43691 48563 43694
rect 50200 43664 51000 43694
rect 7946 43552 8262 43553
rect 0 43482 800 43512
rect 7946 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8262 43552
rect 7946 43487 8262 43488
rect 17946 43552 18262 43553
rect 17946 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18262 43552
rect 17946 43487 18262 43488
rect 27946 43552 28262 43553
rect 27946 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28262 43552
rect 27946 43487 28262 43488
rect 37946 43552 38262 43553
rect 37946 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38262 43552
rect 37946 43487 38262 43488
rect 47946 43552 48262 43553
rect 47946 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48262 43552
rect 47946 43487 48262 43488
rect 933 43482 999 43485
rect 0 43480 999 43482
rect 0 43424 938 43480
rect 994 43424 999 43480
rect 0 43422 999 43424
rect 0 43392 800 43422
rect 933 43419 999 43422
rect 48497 43074 48563 43077
rect 50200 43074 51000 43104
rect 48497 43072 51000 43074
rect 48497 43016 48502 43072
rect 48558 43016 51000 43072
rect 48497 43014 51000 43016
rect 48497 43011 48563 43014
rect 2946 43008 3262 43009
rect 2946 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3262 43008
rect 2946 42943 3262 42944
rect 12946 43008 13262 43009
rect 12946 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13262 43008
rect 12946 42943 13262 42944
rect 22946 43008 23262 43009
rect 22946 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23262 43008
rect 22946 42943 23262 42944
rect 32946 43008 33262 43009
rect 32946 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33262 43008
rect 32946 42943 33262 42944
rect 42946 43008 43262 43009
rect 42946 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43262 43008
rect 50200 42984 51000 43014
rect 42946 42943 43262 42944
rect 7946 42464 8262 42465
rect 7946 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8262 42464
rect 7946 42399 8262 42400
rect 17946 42464 18262 42465
rect 17946 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18262 42464
rect 17946 42399 18262 42400
rect 27946 42464 28262 42465
rect 27946 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28262 42464
rect 27946 42399 28262 42400
rect 37946 42464 38262 42465
rect 37946 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38262 42464
rect 37946 42399 38262 42400
rect 47946 42464 48262 42465
rect 47946 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48262 42464
rect 47946 42399 48262 42400
rect 48497 42394 48563 42397
rect 50200 42394 51000 42424
rect 48497 42392 51000 42394
rect 48497 42336 48502 42392
rect 48558 42336 51000 42392
rect 48497 42334 51000 42336
rect 48497 42331 48563 42334
rect 50200 42304 51000 42334
rect 39982 42060 39988 42124
rect 40052 42122 40058 42124
rect 41321 42122 41387 42125
rect 40052 42120 41387 42122
rect 40052 42064 41326 42120
rect 41382 42064 41387 42120
rect 40052 42062 41387 42064
rect 40052 42060 40058 42062
rect 41321 42059 41387 42062
rect 2946 41920 3262 41921
rect 2946 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3262 41920
rect 2946 41855 3262 41856
rect 12946 41920 13262 41921
rect 12946 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13262 41920
rect 12946 41855 13262 41856
rect 22946 41920 23262 41921
rect 22946 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23262 41920
rect 22946 41855 23262 41856
rect 32946 41920 33262 41921
rect 32946 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33262 41920
rect 32946 41855 33262 41856
rect 42946 41920 43262 41921
rect 42946 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43262 41920
rect 42946 41855 43262 41856
rect 40401 41714 40467 41717
rect 40534 41714 40540 41716
rect 40401 41712 40540 41714
rect 40401 41656 40406 41712
rect 40462 41656 40540 41712
rect 40401 41654 40540 41656
rect 40401 41651 40467 41654
rect 40534 41652 40540 41654
rect 40604 41652 40610 41716
rect 48497 41714 48563 41717
rect 50200 41714 51000 41744
rect 48497 41712 51000 41714
rect 48497 41656 48502 41712
rect 48558 41656 51000 41712
rect 48497 41654 51000 41656
rect 48497 41651 48563 41654
rect 50200 41624 51000 41654
rect 7946 41376 8262 41377
rect 7946 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8262 41376
rect 7946 41311 8262 41312
rect 17946 41376 18262 41377
rect 17946 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18262 41376
rect 17946 41311 18262 41312
rect 27946 41376 28262 41377
rect 27946 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28262 41376
rect 27946 41311 28262 41312
rect 37946 41376 38262 41377
rect 37946 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38262 41376
rect 37946 41311 38262 41312
rect 47946 41376 48262 41377
rect 47946 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48262 41376
rect 47946 41311 48262 41312
rect 0 41170 800 41200
rect 1669 41170 1735 41173
rect 0 41168 1735 41170
rect 0 41112 1674 41168
rect 1730 41112 1735 41168
rect 0 41110 1735 41112
rect 0 41080 800 41110
rect 1669 41107 1735 41110
rect 48497 41034 48563 41037
rect 50200 41034 51000 41064
rect 48497 41032 51000 41034
rect 48497 40976 48502 41032
rect 48558 40976 51000 41032
rect 48497 40974 51000 40976
rect 48497 40971 48563 40974
rect 50200 40944 51000 40974
rect 2946 40832 3262 40833
rect 2946 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3262 40832
rect 2946 40767 3262 40768
rect 12946 40832 13262 40833
rect 12946 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13262 40832
rect 12946 40767 13262 40768
rect 22946 40832 23262 40833
rect 22946 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23262 40832
rect 22946 40767 23262 40768
rect 32946 40832 33262 40833
rect 32946 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33262 40832
rect 32946 40767 33262 40768
rect 42946 40832 43262 40833
rect 42946 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43262 40832
rect 42946 40767 43262 40768
rect 41270 40564 41276 40628
rect 41340 40626 41346 40628
rect 48773 40626 48839 40629
rect 41340 40624 48839 40626
rect 41340 40568 48778 40624
rect 48834 40568 48839 40624
rect 41340 40566 48839 40568
rect 41340 40564 41346 40566
rect 48773 40563 48839 40566
rect 33961 40490 34027 40493
rect 38653 40490 38719 40493
rect 33961 40488 38719 40490
rect 33961 40432 33966 40488
rect 34022 40432 38658 40488
rect 38714 40432 38719 40488
rect 33961 40430 38719 40432
rect 33961 40427 34027 40430
rect 38653 40427 38719 40430
rect 48497 40354 48563 40357
rect 50200 40354 51000 40384
rect 48497 40352 51000 40354
rect 48497 40296 48502 40352
rect 48558 40296 51000 40352
rect 48497 40294 51000 40296
rect 48497 40291 48563 40294
rect 7946 40288 8262 40289
rect 7946 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8262 40288
rect 7946 40223 8262 40224
rect 17946 40288 18262 40289
rect 17946 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18262 40288
rect 17946 40223 18262 40224
rect 27946 40288 28262 40289
rect 27946 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28262 40288
rect 27946 40223 28262 40224
rect 37946 40288 38262 40289
rect 37946 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38262 40288
rect 37946 40223 38262 40224
rect 47946 40288 48262 40289
rect 47946 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48262 40288
rect 50200 40264 51000 40294
rect 47946 40223 48262 40224
rect 27061 40082 27127 40085
rect 30414 40082 30420 40084
rect 27061 40080 30420 40082
rect 27061 40024 27066 40080
rect 27122 40024 30420 40080
rect 27061 40022 30420 40024
rect 27061 40019 27127 40022
rect 30414 40020 30420 40022
rect 30484 40082 30490 40084
rect 30741 40082 30807 40085
rect 30484 40080 30807 40082
rect 30484 40024 30746 40080
rect 30802 40024 30807 40080
rect 30484 40022 30807 40024
rect 30484 40020 30490 40022
rect 30741 40019 30807 40022
rect 2946 39744 3262 39745
rect 2946 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3262 39744
rect 2946 39679 3262 39680
rect 12946 39744 13262 39745
rect 12946 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13262 39744
rect 12946 39679 13262 39680
rect 22946 39744 23262 39745
rect 22946 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23262 39744
rect 22946 39679 23262 39680
rect 32946 39744 33262 39745
rect 32946 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33262 39744
rect 32946 39679 33262 39680
rect 42946 39744 43262 39745
rect 42946 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43262 39744
rect 42946 39679 43262 39680
rect 48497 39674 48563 39677
rect 50200 39674 51000 39704
rect 48497 39672 51000 39674
rect 48497 39616 48502 39672
rect 48558 39616 51000 39672
rect 48497 39614 51000 39616
rect 48497 39611 48563 39614
rect 50200 39584 51000 39614
rect 35985 39538 36051 39541
rect 36721 39538 36787 39541
rect 48773 39538 48839 39541
rect 35985 39536 48839 39538
rect 35985 39480 35990 39536
rect 36046 39480 36726 39536
rect 36782 39480 48778 39536
rect 48834 39480 48839 39536
rect 35985 39478 48839 39480
rect 35985 39475 36051 39478
rect 36721 39475 36787 39478
rect 48773 39475 48839 39478
rect 7946 39200 8262 39201
rect 7946 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8262 39200
rect 7946 39135 8262 39136
rect 17946 39200 18262 39201
rect 17946 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18262 39200
rect 17946 39135 18262 39136
rect 27946 39200 28262 39201
rect 27946 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28262 39200
rect 27946 39135 28262 39136
rect 37946 39200 38262 39201
rect 37946 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38262 39200
rect 37946 39135 38262 39136
rect 47946 39200 48262 39201
rect 47946 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48262 39200
rect 47946 39135 48262 39136
rect 22369 38994 22435 38997
rect 27981 38994 28047 38997
rect 22369 38992 28047 38994
rect 22369 38936 22374 38992
rect 22430 38936 27986 38992
rect 28042 38936 28047 38992
rect 22369 38934 28047 38936
rect 22369 38931 22435 38934
rect 27981 38931 28047 38934
rect 48497 38994 48563 38997
rect 50200 38994 51000 39024
rect 48497 38992 51000 38994
rect 48497 38936 48502 38992
rect 48558 38936 51000 38992
rect 48497 38934 51000 38936
rect 48497 38931 48563 38934
rect 50200 38904 51000 38934
rect 0 38858 800 38888
rect 933 38858 999 38861
rect 0 38856 999 38858
rect 0 38800 938 38856
rect 994 38800 999 38856
rect 0 38798 999 38800
rect 0 38768 800 38798
rect 933 38795 999 38798
rect 35893 38722 35959 38725
rect 38653 38722 38719 38725
rect 35893 38720 38719 38722
rect 35893 38664 35898 38720
rect 35954 38664 38658 38720
rect 38714 38664 38719 38720
rect 35893 38662 38719 38664
rect 35893 38659 35959 38662
rect 38653 38659 38719 38662
rect 2946 38656 3262 38657
rect 2946 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3262 38656
rect 2946 38591 3262 38592
rect 12946 38656 13262 38657
rect 12946 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13262 38656
rect 12946 38591 13262 38592
rect 22946 38656 23262 38657
rect 22946 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23262 38656
rect 22946 38591 23262 38592
rect 32946 38656 33262 38657
rect 32946 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33262 38656
rect 32946 38591 33262 38592
rect 42946 38656 43262 38657
rect 42946 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43262 38656
rect 42946 38591 43262 38592
rect 49325 38314 49391 38317
rect 50200 38314 51000 38344
rect 49325 38312 51000 38314
rect 49325 38256 49330 38312
rect 49386 38256 51000 38312
rect 49325 38254 51000 38256
rect 49325 38251 49391 38254
rect 50200 38224 51000 38254
rect 7946 38112 8262 38113
rect 7946 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8262 38112
rect 7946 38047 8262 38048
rect 17946 38112 18262 38113
rect 17946 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18262 38112
rect 17946 38047 18262 38048
rect 27946 38112 28262 38113
rect 27946 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28262 38112
rect 27946 38047 28262 38048
rect 37946 38112 38262 38113
rect 37946 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38262 38112
rect 37946 38047 38262 38048
rect 47946 38112 48262 38113
rect 47946 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48262 38112
rect 47946 38047 48262 38048
rect 29637 37770 29703 37773
rect 33225 37770 33291 37773
rect 29637 37768 33291 37770
rect 29637 37712 29642 37768
rect 29698 37712 33230 37768
rect 33286 37712 33291 37768
rect 29637 37710 33291 37712
rect 29637 37707 29703 37710
rect 33225 37707 33291 37710
rect 37590 37708 37596 37772
rect 37660 37770 37666 37772
rect 37917 37770 37983 37773
rect 38837 37770 38903 37773
rect 39113 37770 39179 37773
rect 37660 37768 39179 37770
rect 37660 37712 37922 37768
rect 37978 37712 38842 37768
rect 38898 37712 39118 37768
rect 39174 37712 39179 37768
rect 37660 37710 39179 37712
rect 37660 37708 37666 37710
rect 37917 37707 37983 37710
rect 38837 37707 38903 37710
rect 39113 37707 39179 37710
rect 49325 37634 49391 37637
rect 50200 37634 51000 37664
rect 49325 37632 51000 37634
rect 49325 37576 49330 37632
rect 49386 37576 51000 37632
rect 49325 37574 51000 37576
rect 49325 37571 49391 37574
rect 2946 37568 3262 37569
rect 2946 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3262 37568
rect 2946 37503 3262 37504
rect 12946 37568 13262 37569
rect 12946 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13262 37568
rect 12946 37503 13262 37504
rect 22946 37568 23262 37569
rect 22946 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23262 37568
rect 22946 37503 23262 37504
rect 32946 37568 33262 37569
rect 32946 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33262 37568
rect 32946 37503 33262 37504
rect 42946 37568 43262 37569
rect 42946 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43262 37568
rect 50200 37544 51000 37574
rect 42946 37503 43262 37504
rect 7946 37024 8262 37025
rect 7946 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8262 37024
rect 7946 36959 8262 36960
rect 17946 37024 18262 37025
rect 17946 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18262 37024
rect 17946 36959 18262 36960
rect 27946 37024 28262 37025
rect 27946 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28262 37024
rect 27946 36959 28262 36960
rect 37946 37024 38262 37025
rect 37946 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38262 37024
rect 37946 36959 38262 36960
rect 47946 37024 48262 37025
rect 47946 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48262 37024
rect 47946 36959 48262 36960
rect 27337 36954 27403 36957
rect 27797 36954 27863 36957
rect 27337 36952 27863 36954
rect 27337 36896 27342 36952
rect 27398 36896 27802 36952
rect 27858 36896 27863 36952
rect 27337 36894 27863 36896
rect 27337 36891 27403 36894
rect 27797 36891 27863 36894
rect 48497 36954 48563 36957
rect 50200 36954 51000 36984
rect 48497 36952 51000 36954
rect 48497 36896 48502 36952
rect 48558 36896 51000 36952
rect 48497 36894 51000 36896
rect 48497 36891 48563 36894
rect 50200 36864 51000 36894
rect 37774 36756 37780 36820
rect 37844 36818 37850 36820
rect 38561 36818 38627 36821
rect 37844 36816 38627 36818
rect 37844 36760 38566 36816
rect 38622 36760 38627 36816
rect 37844 36758 38627 36760
rect 37844 36756 37850 36758
rect 38561 36755 38627 36758
rect 40033 36818 40099 36821
rect 42333 36818 42399 36821
rect 40033 36816 42399 36818
rect 40033 36760 40038 36816
rect 40094 36760 42338 36816
rect 42394 36760 42399 36816
rect 40033 36758 42399 36760
rect 40033 36755 40099 36758
rect 42333 36755 42399 36758
rect 29453 36682 29519 36685
rect 31017 36682 31083 36685
rect 38009 36682 38075 36685
rect 29453 36680 38075 36682
rect 29453 36624 29458 36680
rect 29514 36624 31022 36680
rect 31078 36624 38014 36680
rect 38070 36624 38075 36680
rect 29453 36622 38075 36624
rect 29453 36619 29519 36622
rect 31017 36619 31083 36622
rect 38009 36619 38075 36622
rect 39297 36682 39363 36685
rect 46289 36682 46355 36685
rect 39297 36680 46355 36682
rect 39297 36624 39302 36680
rect 39358 36624 46294 36680
rect 46350 36624 46355 36680
rect 39297 36622 46355 36624
rect 39297 36619 39363 36622
rect 46289 36619 46355 36622
rect 0 36546 800 36576
rect 933 36546 999 36549
rect 0 36544 999 36546
rect 0 36488 938 36544
rect 994 36488 999 36544
rect 0 36486 999 36488
rect 0 36456 800 36486
rect 933 36483 999 36486
rect 2946 36480 3262 36481
rect 2946 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3262 36480
rect 2946 36415 3262 36416
rect 12946 36480 13262 36481
rect 12946 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13262 36480
rect 12946 36415 13262 36416
rect 22946 36480 23262 36481
rect 22946 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23262 36480
rect 22946 36415 23262 36416
rect 32946 36480 33262 36481
rect 32946 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33262 36480
rect 32946 36415 33262 36416
rect 42946 36480 43262 36481
rect 42946 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43262 36480
rect 42946 36415 43262 36416
rect 33685 36410 33751 36413
rect 33685 36408 41430 36410
rect 33685 36352 33690 36408
rect 33746 36352 41430 36408
rect 33685 36350 41430 36352
rect 33685 36347 33751 36350
rect 32489 36274 32555 36277
rect 39665 36274 39731 36277
rect 41370 36274 41430 36350
rect 41781 36274 41847 36277
rect 32489 36272 40786 36274
rect 32489 36216 32494 36272
rect 32550 36216 39670 36272
rect 39726 36216 40786 36272
rect 32489 36214 40786 36216
rect 41370 36272 41847 36274
rect 41370 36216 41786 36272
rect 41842 36216 41847 36272
rect 41370 36214 41847 36216
rect 32489 36211 32555 36214
rect 39665 36211 39731 36214
rect 28165 36138 28231 36141
rect 37774 36138 37780 36140
rect 28165 36136 37780 36138
rect 28165 36080 28170 36136
rect 28226 36080 37780 36136
rect 28165 36078 37780 36080
rect 28165 36075 28231 36078
rect 37774 36076 37780 36078
rect 37844 36076 37850 36140
rect 25589 36004 25655 36005
rect 25589 36000 25636 36004
rect 25700 36002 25706 36004
rect 25589 35944 25594 36000
rect 25589 35940 25636 35944
rect 25700 35942 25746 36002
rect 25700 35940 25706 35942
rect 25589 35939 25655 35940
rect 7946 35936 8262 35937
rect 7946 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8262 35936
rect 7946 35871 8262 35872
rect 17946 35936 18262 35937
rect 17946 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18262 35936
rect 17946 35871 18262 35872
rect 27946 35936 28262 35937
rect 27946 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28262 35936
rect 27946 35871 28262 35872
rect 37946 35936 38262 35937
rect 37946 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38262 35936
rect 37946 35871 38262 35872
rect 40726 35869 40786 36214
rect 41781 36211 41847 36214
rect 49325 36274 49391 36277
rect 50200 36274 51000 36304
rect 49325 36272 51000 36274
rect 49325 36216 49330 36272
rect 49386 36216 51000 36272
rect 49325 36214 51000 36216
rect 49325 36211 49391 36214
rect 50200 36184 51000 36214
rect 47946 35936 48262 35937
rect 47946 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48262 35936
rect 47946 35871 48262 35872
rect 40726 35864 40835 35869
rect 40726 35808 40774 35864
rect 40830 35808 40835 35864
rect 40726 35806 40835 35808
rect 40769 35803 40835 35806
rect 41137 35866 41203 35869
rect 41270 35866 41276 35868
rect 41137 35864 41276 35866
rect 41137 35808 41142 35864
rect 41198 35808 41276 35864
rect 41137 35806 41276 35808
rect 41137 35803 41203 35806
rect 41270 35804 41276 35806
rect 41340 35804 41346 35868
rect 25773 35730 25839 35733
rect 28758 35730 28764 35732
rect 25773 35728 28764 35730
rect 25773 35672 25778 35728
rect 25834 35672 28764 35728
rect 25773 35670 28764 35672
rect 25773 35667 25839 35670
rect 28758 35668 28764 35670
rect 28828 35730 28834 35732
rect 36169 35730 36235 35733
rect 28828 35728 36235 35730
rect 28828 35672 36174 35728
rect 36230 35672 36235 35728
rect 28828 35670 36235 35672
rect 28828 35668 28834 35670
rect 36169 35667 36235 35670
rect 32765 35594 32831 35597
rect 31710 35592 32831 35594
rect 31710 35536 32770 35592
rect 32826 35536 32831 35592
rect 31710 35534 32831 35536
rect 2946 35392 3262 35393
rect 2946 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3262 35392
rect 2946 35327 3262 35328
rect 12946 35392 13262 35393
rect 12946 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13262 35392
rect 12946 35327 13262 35328
rect 22946 35392 23262 35393
rect 22946 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23262 35392
rect 22946 35327 23262 35328
rect 24393 35322 24459 35325
rect 27705 35322 27771 35325
rect 31710 35322 31770 35534
rect 32765 35531 32831 35534
rect 49325 35594 49391 35597
rect 50200 35594 51000 35624
rect 49325 35592 51000 35594
rect 49325 35536 49330 35592
rect 49386 35536 51000 35592
rect 49325 35534 51000 35536
rect 49325 35531 49391 35534
rect 50200 35504 51000 35534
rect 32946 35392 33262 35393
rect 32946 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33262 35392
rect 32946 35327 33262 35328
rect 42946 35392 43262 35393
rect 42946 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43262 35392
rect 42946 35327 43262 35328
rect 24393 35320 31770 35322
rect 24393 35264 24398 35320
rect 24454 35264 27710 35320
rect 27766 35264 31770 35320
rect 24393 35262 31770 35264
rect 24393 35259 24459 35262
rect 27705 35259 27771 35262
rect 36077 35186 36143 35189
rect 37917 35186 37983 35189
rect 36077 35184 37983 35186
rect 36077 35128 36082 35184
rect 36138 35128 37922 35184
rect 37978 35128 37983 35184
rect 36077 35126 37983 35128
rect 36077 35123 36143 35126
rect 37917 35123 37983 35126
rect 28574 34988 28580 35052
rect 28644 35050 28650 35052
rect 28901 35050 28967 35053
rect 28644 35048 28967 35050
rect 28644 34992 28906 35048
rect 28962 34992 28967 35048
rect 28644 34990 28967 34992
rect 28644 34988 28650 34990
rect 28901 34987 28967 34990
rect 38653 35050 38719 35053
rect 39389 35050 39455 35053
rect 38653 35048 39455 35050
rect 38653 34992 38658 35048
rect 38714 34992 39394 35048
rect 39450 34992 39455 35048
rect 38653 34990 39455 34992
rect 38653 34987 38719 34990
rect 39389 34987 39455 34990
rect 38929 34916 38995 34917
rect 38878 34914 38884 34916
rect 38838 34854 38884 34914
rect 38948 34912 38995 34916
rect 38990 34856 38995 34912
rect 38878 34852 38884 34854
rect 38948 34852 38995 34856
rect 38929 34851 38995 34852
rect 49325 34914 49391 34917
rect 50200 34914 51000 34944
rect 49325 34912 51000 34914
rect 49325 34856 49330 34912
rect 49386 34856 51000 34912
rect 49325 34854 51000 34856
rect 49325 34851 49391 34854
rect 7946 34848 8262 34849
rect 7946 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8262 34848
rect 7946 34783 8262 34784
rect 17946 34848 18262 34849
rect 17946 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18262 34848
rect 17946 34783 18262 34784
rect 27946 34848 28262 34849
rect 27946 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28262 34848
rect 27946 34783 28262 34784
rect 37946 34848 38262 34849
rect 37946 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38262 34848
rect 37946 34783 38262 34784
rect 47946 34848 48262 34849
rect 47946 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48262 34848
rect 50200 34824 51000 34854
rect 47946 34783 48262 34784
rect 38929 34778 38995 34781
rect 41137 34778 41203 34781
rect 38929 34776 41203 34778
rect 38929 34720 38934 34776
rect 38990 34720 41142 34776
rect 41198 34720 41203 34776
rect 38929 34718 41203 34720
rect 38929 34715 38995 34718
rect 41137 34715 41203 34718
rect 2946 34304 3262 34305
rect 0 34234 800 34264
rect 2946 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3262 34304
rect 2946 34239 3262 34240
rect 12946 34304 13262 34305
rect 12946 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13262 34304
rect 12946 34239 13262 34240
rect 22946 34304 23262 34305
rect 22946 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23262 34304
rect 22946 34239 23262 34240
rect 32946 34304 33262 34305
rect 32946 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33262 34304
rect 32946 34239 33262 34240
rect 42946 34304 43262 34305
rect 42946 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43262 34304
rect 42946 34239 43262 34240
rect 1761 34234 1827 34237
rect 0 34232 1827 34234
rect 0 34176 1766 34232
rect 1822 34176 1827 34232
rect 0 34174 1827 34176
rect 0 34144 800 34174
rect 1761 34171 1827 34174
rect 38745 34234 38811 34237
rect 40033 34234 40099 34237
rect 38745 34232 40099 34234
rect 38745 34176 38750 34232
rect 38806 34176 40038 34232
rect 40094 34176 40099 34232
rect 38745 34174 40099 34176
rect 38745 34171 38811 34174
rect 40033 34171 40099 34174
rect 49325 34234 49391 34237
rect 50200 34234 51000 34264
rect 49325 34232 51000 34234
rect 49325 34176 49330 34232
rect 49386 34176 51000 34232
rect 49325 34174 51000 34176
rect 49325 34171 49391 34174
rect 50200 34144 51000 34174
rect 31569 34098 31635 34101
rect 36537 34098 36603 34101
rect 31569 34096 36603 34098
rect 31569 34040 31574 34096
rect 31630 34040 36542 34096
rect 36598 34040 36603 34096
rect 31569 34038 36603 34040
rect 31569 34035 31635 34038
rect 36537 34035 36603 34038
rect 38653 34098 38719 34101
rect 39573 34098 39639 34101
rect 38653 34096 39639 34098
rect 38653 34040 38658 34096
rect 38714 34040 39578 34096
rect 39634 34040 39639 34096
rect 38653 34038 39639 34040
rect 38653 34035 38719 34038
rect 39573 34035 39639 34038
rect 27981 33962 28047 33965
rect 27340 33960 28047 33962
rect 27340 33904 27986 33960
rect 28042 33904 28047 33960
rect 27340 33902 28047 33904
rect 27340 33829 27400 33902
rect 27981 33899 28047 33902
rect 37089 33962 37155 33965
rect 49233 33962 49299 33965
rect 37089 33960 49299 33962
rect 37089 33904 37094 33960
rect 37150 33904 49238 33960
rect 49294 33904 49299 33960
rect 37089 33902 49299 33904
rect 37089 33899 37155 33902
rect 49233 33899 49299 33902
rect 27337 33824 27403 33829
rect 27337 33768 27342 33824
rect 27398 33768 27403 33824
rect 27337 33763 27403 33768
rect 7946 33760 8262 33761
rect 7946 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8262 33760
rect 7946 33695 8262 33696
rect 17946 33760 18262 33761
rect 17946 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18262 33760
rect 17946 33695 18262 33696
rect 27946 33760 28262 33761
rect 27946 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28262 33760
rect 27946 33695 28262 33696
rect 37946 33760 38262 33761
rect 37946 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38262 33760
rect 37946 33695 38262 33696
rect 47946 33760 48262 33761
rect 47946 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48262 33760
rect 47946 33695 48262 33696
rect 38745 33690 38811 33693
rect 39297 33690 39363 33693
rect 38745 33688 39363 33690
rect 38745 33632 38750 33688
rect 38806 33632 39302 33688
rect 39358 33632 39363 33688
rect 38745 33630 39363 33632
rect 38745 33627 38811 33630
rect 39297 33627 39363 33630
rect 37825 33554 37891 33557
rect 38837 33556 38903 33557
rect 38837 33554 38884 33556
rect 31710 33552 37891 33554
rect 31710 33496 37830 33552
rect 37886 33496 37891 33552
rect 31710 33494 37891 33496
rect 38792 33552 38884 33554
rect 38792 33496 38842 33552
rect 38792 33494 38884 33496
rect 26969 33282 27035 33285
rect 31710 33282 31770 33494
rect 37825 33491 37891 33494
rect 38837 33492 38884 33494
rect 38948 33492 38954 33556
rect 49325 33554 49391 33557
rect 50200 33554 51000 33584
rect 49325 33552 51000 33554
rect 49325 33496 49330 33552
rect 49386 33496 51000 33552
rect 49325 33494 51000 33496
rect 38837 33491 38903 33492
rect 49325 33491 49391 33494
rect 50200 33464 51000 33494
rect 26969 33280 31770 33282
rect 26969 33224 26974 33280
rect 27030 33224 31770 33280
rect 26969 33222 31770 33224
rect 26969 33219 27035 33222
rect 2946 33216 3262 33217
rect 2946 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3262 33216
rect 2946 33151 3262 33152
rect 12946 33216 13262 33217
rect 12946 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13262 33216
rect 12946 33151 13262 33152
rect 22946 33216 23262 33217
rect 22946 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23262 33216
rect 22946 33151 23262 33152
rect 32946 33216 33262 33217
rect 32946 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33262 33216
rect 32946 33151 33262 33152
rect 42946 33216 43262 33217
rect 42946 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43262 33216
rect 42946 33151 43262 33152
rect 28717 33010 28783 33013
rect 40585 33010 40651 33013
rect 40861 33010 40927 33013
rect 28717 33008 29010 33010
rect 28717 32952 28722 33008
rect 28778 32952 29010 33008
rect 28717 32950 29010 32952
rect 28717 32947 28783 32950
rect 28950 32877 29010 32950
rect 40585 33008 40927 33010
rect 40585 32952 40590 33008
rect 40646 32952 40866 33008
rect 40922 32952 40927 33008
rect 40585 32950 40927 32952
rect 40585 32947 40651 32950
rect 40861 32947 40927 32950
rect 24209 32874 24275 32877
rect 26693 32874 26759 32877
rect 28717 32874 28783 32877
rect 24209 32872 28783 32874
rect 24209 32816 24214 32872
rect 24270 32816 26698 32872
rect 26754 32816 28722 32872
rect 28778 32816 28783 32872
rect 24209 32814 28783 32816
rect 24209 32811 24275 32814
rect 26693 32811 26759 32814
rect 28717 32811 28783 32814
rect 28901 32872 29010 32877
rect 28901 32816 28906 32872
rect 28962 32816 29010 32872
rect 28901 32814 29010 32816
rect 49325 32874 49391 32877
rect 50200 32874 51000 32904
rect 49325 32872 51000 32874
rect 49325 32816 49330 32872
rect 49386 32816 51000 32872
rect 49325 32814 51000 32816
rect 28901 32811 28967 32814
rect 49325 32811 49391 32814
rect 50200 32784 51000 32814
rect 7946 32672 8262 32673
rect 7946 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8262 32672
rect 7946 32607 8262 32608
rect 17946 32672 18262 32673
rect 17946 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18262 32672
rect 17946 32607 18262 32608
rect 27946 32672 28262 32673
rect 27946 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28262 32672
rect 27946 32607 28262 32608
rect 37946 32672 38262 32673
rect 37946 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38262 32672
rect 37946 32607 38262 32608
rect 47946 32672 48262 32673
rect 47946 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48262 32672
rect 47946 32607 48262 32608
rect 28533 32196 28599 32197
rect 28533 32192 28580 32196
rect 28644 32194 28650 32196
rect 48497 32194 48563 32197
rect 50200 32194 51000 32224
rect 28533 32136 28538 32192
rect 28533 32132 28580 32136
rect 28644 32134 28690 32194
rect 48497 32192 51000 32194
rect 48497 32136 48502 32192
rect 48558 32136 51000 32192
rect 48497 32134 51000 32136
rect 28644 32132 28650 32134
rect 28533 32131 28599 32132
rect 48497 32131 48563 32134
rect 2946 32128 3262 32129
rect 2946 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3262 32128
rect 2946 32063 3262 32064
rect 12946 32128 13262 32129
rect 12946 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13262 32128
rect 12946 32063 13262 32064
rect 22946 32128 23262 32129
rect 22946 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23262 32128
rect 22946 32063 23262 32064
rect 32946 32128 33262 32129
rect 32946 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33262 32128
rect 32946 32063 33262 32064
rect 42946 32128 43262 32129
rect 42946 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43262 32128
rect 50200 32104 51000 32134
rect 42946 32063 43262 32064
rect 0 31922 800 31952
rect 933 31922 999 31925
rect 0 31920 999 31922
rect 0 31864 938 31920
rect 994 31864 999 31920
rect 0 31862 999 31864
rect 0 31832 800 31862
rect 933 31859 999 31862
rect 37406 31860 37412 31924
rect 37476 31922 37482 31924
rect 38561 31922 38627 31925
rect 37476 31920 38627 31922
rect 37476 31864 38566 31920
rect 38622 31864 38627 31920
rect 37476 31862 38627 31864
rect 37476 31860 37482 31862
rect 38561 31859 38627 31862
rect 37089 31786 37155 31789
rect 38561 31786 38627 31789
rect 37089 31784 38627 31786
rect 37089 31728 37094 31784
rect 37150 31728 38566 31784
rect 38622 31728 38627 31784
rect 37089 31726 38627 31728
rect 37089 31723 37155 31726
rect 38561 31723 38627 31726
rect 7946 31584 8262 31585
rect 7946 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8262 31584
rect 7946 31519 8262 31520
rect 17946 31584 18262 31585
rect 17946 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18262 31584
rect 17946 31519 18262 31520
rect 27946 31584 28262 31585
rect 27946 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28262 31584
rect 27946 31519 28262 31520
rect 37946 31584 38262 31585
rect 37946 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38262 31584
rect 37946 31519 38262 31520
rect 47946 31584 48262 31585
rect 47946 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48262 31584
rect 47946 31519 48262 31520
rect 35985 31514 36051 31517
rect 48497 31514 48563 31517
rect 50200 31514 51000 31544
rect 35985 31512 37842 31514
rect 35985 31456 35990 31512
rect 36046 31456 37842 31512
rect 35985 31454 37842 31456
rect 35985 31451 36051 31454
rect 33593 31378 33659 31381
rect 36997 31378 37063 31381
rect 33593 31376 37063 31378
rect 33593 31320 33598 31376
rect 33654 31320 37002 31376
rect 37058 31320 37063 31376
rect 33593 31318 37063 31320
rect 37782 31378 37842 31454
rect 48497 31512 51000 31514
rect 48497 31456 48502 31512
rect 48558 31456 51000 31512
rect 48497 31454 51000 31456
rect 48497 31451 48563 31454
rect 50200 31424 51000 31454
rect 38469 31378 38535 31381
rect 37782 31376 38535 31378
rect 37782 31320 38474 31376
rect 38530 31320 38535 31376
rect 37782 31318 38535 31320
rect 33593 31315 33659 31318
rect 36997 31315 37063 31318
rect 38469 31315 38535 31318
rect 9765 31242 9831 31245
rect 22461 31244 22527 31245
rect 22461 31242 22508 31244
rect 9765 31240 22508 31242
rect 9765 31184 9770 31240
rect 9826 31184 22466 31240
rect 9765 31182 22508 31184
rect 9765 31179 9831 31182
rect 22461 31180 22508 31182
rect 22572 31180 22578 31244
rect 22461 31179 22527 31180
rect 2946 31040 3262 31041
rect 2946 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3262 31040
rect 2946 30975 3262 30976
rect 12946 31040 13262 31041
rect 12946 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13262 31040
rect 12946 30975 13262 30976
rect 22946 31040 23262 31041
rect 22946 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23262 31040
rect 22946 30975 23262 30976
rect 32946 31040 33262 31041
rect 32946 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33262 31040
rect 32946 30975 33262 30976
rect 42946 31040 43262 31041
rect 42946 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43262 31040
rect 42946 30975 43262 30976
rect 48497 30834 48563 30837
rect 50200 30834 51000 30864
rect 48497 30832 51000 30834
rect 48497 30776 48502 30832
rect 48558 30776 51000 30832
rect 48497 30774 51000 30776
rect 48497 30771 48563 30774
rect 50200 30744 51000 30774
rect 30189 30698 30255 30701
rect 27662 30696 30255 30698
rect 27662 30640 30194 30696
rect 30250 30640 30255 30696
rect 27662 30638 30255 30640
rect 7946 30496 8262 30497
rect 7946 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8262 30496
rect 7946 30431 8262 30432
rect 17946 30496 18262 30497
rect 17946 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18262 30496
rect 17946 30431 18262 30432
rect 25078 30364 25084 30428
rect 25148 30426 25154 30428
rect 26049 30426 26115 30429
rect 27662 30426 27722 30638
rect 30189 30635 30255 30638
rect 27946 30496 28262 30497
rect 27946 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28262 30496
rect 27946 30431 28262 30432
rect 37946 30496 38262 30497
rect 37946 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38262 30496
rect 37946 30431 38262 30432
rect 47946 30496 48262 30497
rect 47946 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48262 30496
rect 47946 30431 48262 30432
rect 25148 30424 27722 30426
rect 25148 30368 26054 30424
rect 26110 30368 27722 30424
rect 25148 30366 27722 30368
rect 25148 30364 25154 30366
rect 26049 30363 26115 30366
rect 28257 30290 28323 30293
rect 34513 30290 34579 30293
rect 28257 30288 34579 30290
rect 28257 30232 28262 30288
rect 28318 30232 34518 30288
rect 34574 30232 34579 30288
rect 28257 30230 34579 30232
rect 28257 30227 28323 30230
rect 34513 30227 34579 30230
rect 37774 30228 37780 30292
rect 37844 30290 37850 30292
rect 37917 30290 37983 30293
rect 37844 30288 37983 30290
rect 37844 30232 37922 30288
rect 37978 30232 37983 30288
rect 37844 30230 37983 30232
rect 37844 30228 37850 30230
rect 37917 30227 37983 30230
rect 22093 30154 22159 30157
rect 28758 30154 28764 30156
rect 22093 30152 28764 30154
rect 22093 30096 22098 30152
rect 22154 30096 28764 30152
rect 22093 30094 28764 30096
rect 22093 30091 22159 30094
rect 28758 30092 28764 30094
rect 28828 30154 28834 30156
rect 28901 30154 28967 30157
rect 28828 30152 28967 30154
rect 28828 30096 28906 30152
rect 28962 30096 28967 30152
rect 28828 30094 28967 30096
rect 28828 30092 28834 30094
rect 28901 30091 28967 30094
rect 30649 30154 30715 30157
rect 30782 30154 30788 30156
rect 30649 30152 30788 30154
rect 30649 30096 30654 30152
rect 30710 30096 30788 30152
rect 30649 30094 30788 30096
rect 30649 30091 30715 30094
rect 30782 30092 30788 30094
rect 30852 30092 30858 30156
rect 49325 30154 49391 30157
rect 50200 30154 51000 30184
rect 49325 30152 51000 30154
rect 49325 30096 49330 30152
rect 49386 30096 51000 30152
rect 49325 30094 51000 30096
rect 49325 30091 49391 30094
rect 50200 30064 51000 30094
rect 2946 29952 3262 29953
rect 2946 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3262 29952
rect 2946 29887 3262 29888
rect 12946 29952 13262 29953
rect 12946 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13262 29952
rect 12946 29887 13262 29888
rect 22946 29952 23262 29953
rect 22946 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23262 29952
rect 22946 29887 23262 29888
rect 32946 29952 33262 29953
rect 32946 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33262 29952
rect 32946 29887 33262 29888
rect 42946 29952 43262 29953
rect 42946 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43262 29952
rect 42946 29887 43262 29888
rect 0 29610 800 29640
rect 1301 29610 1367 29613
rect 0 29608 1367 29610
rect 0 29552 1306 29608
rect 1362 29552 1367 29608
rect 0 29550 1367 29552
rect 0 29520 800 29550
rect 1301 29547 1367 29550
rect 48497 29474 48563 29477
rect 50200 29474 51000 29504
rect 48497 29472 51000 29474
rect 48497 29416 48502 29472
rect 48558 29416 51000 29472
rect 48497 29414 51000 29416
rect 48497 29411 48563 29414
rect 7946 29408 8262 29409
rect 7946 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8262 29408
rect 7946 29343 8262 29344
rect 17946 29408 18262 29409
rect 17946 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18262 29408
rect 17946 29343 18262 29344
rect 27946 29408 28262 29409
rect 27946 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28262 29408
rect 27946 29343 28262 29344
rect 37946 29408 38262 29409
rect 37946 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38262 29408
rect 37946 29343 38262 29344
rect 47946 29408 48262 29409
rect 47946 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48262 29408
rect 50200 29384 51000 29414
rect 47946 29343 48262 29344
rect 33685 29066 33751 29069
rect 37590 29066 37596 29068
rect 33685 29064 37596 29066
rect 33685 29008 33690 29064
rect 33746 29008 37596 29064
rect 33685 29006 37596 29008
rect 33685 29003 33751 29006
rect 37590 29004 37596 29006
rect 37660 29004 37666 29068
rect 2946 28864 3262 28865
rect 2946 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3262 28864
rect 2946 28799 3262 28800
rect 12946 28864 13262 28865
rect 12946 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13262 28864
rect 12946 28799 13262 28800
rect 22946 28864 23262 28865
rect 22946 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23262 28864
rect 22946 28799 23262 28800
rect 32946 28864 33262 28865
rect 32946 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33262 28864
rect 32946 28799 33262 28800
rect 42946 28864 43262 28865
rect 42946 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43262 28864
rect 42946 28799 43262 28800
rect 49325 28794 49391 28797
rect 50200 28794 51000 28824
rect 49325 28792 51000 28794
rect 49325 28736 49330 28792
rect 49386 28736 51000 28792
rect 49325 28734 51000 28736
rect 49325 28731 49391 28734
rect 50200 28704 51000 28734
rect 36445 28522 36511 28525
rect 40534 28522 40540 28524
rect 36445 28520 40540 28522
rect 36445 28464 36450 28520
rect 36506 28464 40540 28520
rect 36445 28462 40540 28464
rect 36445 28459 36511 28462
rect 40534 28460 40540 28462
rect 40604 28460 40610 28524
rect 35198 28324 35204 28388
rect 35268 28386 35274 28388
rect 35341 28386 35407 28389
rect 35268 28384 35407 28386
rect 35268 28328 35346 28384
rect 35402 28328 35407 28384
rect 35268 28326 35407 28328
rect 35268 28324 35274 28326
rect 35341 28323 35407 28326
rect 7946 28320 8262 28321
rect 7946 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8262 28320
rect 7946 28255 8262 28256
rect 17946 28320 18262 28321
rect 17946 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18262 28320
rect 17946 28255 18262 28256
rect 27946 28320 28262 28321
rect 27946 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28262 28320
rect 27946 28255 28262 28256
rect 37946 28320 38262 28321
rect 37946 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38262 28320
rect 37946 28255 38262 28256
rect 47946 28320 48262 28321
rect 47946 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48262 28320
rect 47946 28255 48262 28256
rect 27705 28252 27771 28253
rect 27654 28250 27660 28252
rect 27614 28190 27660 28250
rect 27724 28248 27771 28252
rect 27766 28192 27771 28248
rect 27654 28188 27660 28190
rect 27724 28188 27771 28192
rect 27705 28187 27771 28188
rect 31201 28114 31267 28117
rect 37273 28114 37339 28117
rect 31201 28112 37339 28114
rect 31201 28056 31206 28112
rect 31262 28056 37278 28112
rect 37334 28056 37339 28112
rect 31201 28054 37339 28056
rect 31201 28051 31267 28054
rect 37273 28051 37339 28054
rect 49325 28114 49391 28117
rect 50200 28114 51000 28144
rect 49325 28112 51000 28114
rect 49325 28056 49330 28112
rect 49386 28056 51000 28112
rect 49325 28054 51000 28056
rect 49325 28051 49391 28054
rect 50200 28024 51000 28054
rect 2946 27776 3262 27777
rect 2946 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3262 27776
rect 2946 27711 3262 27712
rect 12946 27776 13262 27777
rect 12946 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13262 27776
rect 12946 27711 13262 27712
rect 22946 27776 23262 27777
rect 22946 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23262 27776
rect 22946 27711 23262 27712
rect 32946 27776 33262 27777
rect 32946 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33262 27776
rect 32946 27711 33262 27712
rect 42946 27776 43262 27777
rect 42946 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43262 27776
rect 42946 27711 43262 27712
rect 27061 27708 27127 27709
rect 27061 27704 27108 27708
rect 27172 27706 27178 27708
rect 27061 27648 27066 27704
rect 27061 27644 27108 27648
rect 27172 27646 27218 27706
rect 27172 27644 27178 27646
rect 27061 27643 27127 27644
rect 31569 27434 31635 27437
rect 34973 27434 35039 27437
rect 31569 27432 35039 27434
rect 31569 27376 31574 27432
rect 31630 27376 34978 27432
rect 35034 27376 35039 27432
rect 31569 27374 35039 27376
rect 31569 27371 31635 27374
rect 34973 27371 35039 27374
rect 48497 27434 48563 27437
rect 50200 27434 51000 27464
rect 48497 27432 51000 27434
rect 48497 27376 48502 27432
rect 48558 27376 51000 27432
rect 48497 27374 51000 27376
rect 48497 27371 48563 27374
rect 50200 27344 51000 27374
rect 0 27298 800 27328
rect 1301 27298 1367 27301
rect 0 27296 1367 27298
rect 0 27240 1306 27296
rect 1362 27240 1367 27296
rect 0 27238 1367 27240
rect 0 27208 800 27238
rect 1301 27235 1367 27238
rect 29453 27298 29519 27301
rect 30414 27298 30420 27300
rect 29453 27296 30420 27298
rect 29453 27240 29458 27296
rect 29514 27240 30420 27296
rect 29453 27238 30420 27240
rect 29453 27235 29519 27238
rect 30414 27236 30420 27238
rect 30484 27298 30490 27300
rect 30925 27298 30991 27301
rect 30484 27296 30991 27298
rect 30484 27240 30930 27296
rect 30986 27240 30991 27296
rect 30484 27238 30991 27240
rect 30484 27236 30490 27238
rect 30925 27235 30991 27238
rect 7946 27232 8262 27233
rect 7946 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8262 27232
rect 7946 27167 8262 27168
rect 17946 27232 18262 27233
rect 17946 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18262 27232
rect 17946 27167 18262 27168
rect 27946 27232 28262 27233
rect 27946 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28262 27232
rect 27946 27167 28262 27168
rect 37946 27232 38262 27233
rect 37946 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38262 27232
rect 37946 27167 38262 27168
rect 47946 27232 48262 27233
rect 47946 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48262 27232
rect 47946 27167 48262 27168
rect 30966 26964 30972 27028
rect 31036 27026 31042 27028
rect 31293 27026 31359 27029
rect 31036 27024 31359 27026
rect 31036 26968 31298 27024
rect 31354 26968 31359 27024
rect 31036 26966 31359 26968
rect 31036 26964 31042 26966
rect 31293 26963 31359 26966
rect 34605 27026 34671 27029
rect 37406 27026 37412 27028
rect 34605 27024 37412 27026
rect 34605 26968 34610 27024
rect 34666 26968 37412 27024
rect 34605 26966 37412 26968
rect 34605 26963 34671 26966
rect 37406 26964 37412 26966
rect 37476 27026 37482 27028
rect 38510 27026 38516 27028
rect 37476 26966 38516 27026
rect 37476 26964 37482 26966
rect 38510 26964 38516 26966
rect 38580 26964 38586 27028
rect 48497 26754 48563 26757
rect 50200 26754 51000 26784
rect 48497 26752 51000 26754
rect 48497 26696 48502 26752
rect 48558 26696 51000 26752
rect 48497 26694 51000 26696
rect 48497 26691 48563 26694
rect 2946 26688 3262 26689
rect 2946 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3262 26688
rect 2946 26623 3262 26624
rect 12946 26688 13262 26689
rect 12946 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13262 26688
rect 12946 26623 13262 26624
rect 22946 26688 23262 26689
rect 22946 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23262 26688
rect 22946 26623 23262 26624
rect 32946 26688 33262 26689
rect 32946 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33262 26688
rect 32946 26623 33262 26624
rect 42946 26688 43262 26689
rect 42946 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43262 26688
rect 50200 26664 51000 26694
rect 42946 26623 43262 26624
rect 31017 26346 31083 26349
rect 32121 26346 32187 26349
rect 32622 26346 32628 26348
rect 31017 26344 32628 26346
rect 31017 26288 31022 26344
rect 31078 26288 32126 26344
rect 32182 26288 32628 26344
rect 31017 26286 32628 26288
rect 31017 26283 31083 26286
rect 32121 26283 32187 26286
rect 32622 26284 32628 26286
rect 32692 26284 32698 26348
rect 37089 26346 37155 26349
rect 38653 26346 38719 26349
rect 39982 26346 39988 26348
rect 37089 26344 39988 26346
rect 37089 26288 37094 26344
rect 37150 26288 38658 26344
rect 38714 26288 39988 26344
rect 37089 26286 39988 26288
rect 37089 26283 37155 26286
rect 38653 26283 38719 26286
rect 39982 26284 39988 26286
rect 40052 26284 40058 26348
rect 7946 26144 8262 26145
rect 7946 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8262 26144
rect 7946 26079 8262 26080
rect 17946 26144 18262 26145
rect 17946 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18262 26144
rect 17946 26079 18262 26080
rect 27946 26144 28262 26145
rect 27946 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28262 26144
rect 27946 26079 28262 26080
rect 37946 26144 38262 26145
rect 37946 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38262 26144
rect 37946 26079 38262 26080
rect 47946 26144 48262 26145
rect 47946 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48262 26144
rect 47946 26079 48262 26080
rect 48497 26074 48563 26077
rect 50200 26074 51000 26104
rect 48497 26072 51000 26074
rect 48497 26016 48502 26072
rect 48558 26016 51000 26072
rect 48497 26014 51000 26016
rect 48497 26011 48563 26014
rect 50200 25984 51000 26014
rect 2946 25600 3262 25601
rect 2946 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3262 25600
rect 2946 25535 3262 25536
rect 12946 25600 13262 25601
rect 12946 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13262 25600
rect 12946 25535 13262 25536
rect 22946 25600 23262 25601
rect 22946 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23262 25600
rect 22946 25535 23262 25536
rect 32946 25600 33262 25601
rect 32946 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33262 25600
rect 32946 25535 33262 25536
rect 42946 25600 43262 25601
rect 42946 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43262 25600
rect 42946 25535 43262 25536
rect 32673 25394 32739 25397
rect 31710 25392 32739 25394
rect 31710 25336 32678 25392
rect 32734 25336 32739 25392
rect 31710 25334 32739 25336
rect 9581 25258 9647 25261
rect 30414 25258 30420 25260
rect 9581 25256 30420 25258
rect 9581 25200 9586 25256
rect 9642 25200 30420 25256
rect 9581 25198 30420 25200
rect 9581 25195 9647 25198
rect 30414 25196 30420 25198
rect 30484 25258 30490 25260
rect 31710 25258 31770 25334
rect 32673 25331 32739 25334
rect 49325 25394 49391 25397
rect 50200 25394 51000 25424
rect 49325 25392 51000 25394
rect 49325 25336 49330 25392
rect 49386 25336 51000 25392
rect 49325 25334 51000 25336
rect 49325 25331 49391 25334
rect 50200 25304 51000 25334
rect 30484 25198 31770 25258
rect 30484 25196 30490 25198
rect 28901 25122 28967 25125
rect 28901 25120 29010 25122
rect 28901 25064 28906 25120
rect 28962 25064 29010 25120
rect 28901 25059 29010 25064
rect 7946 25056 8262 25057
rect 0 24986 800 25016
rect 7946 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8262 25056
rect 7946 24991 8262 24992
rect 17946 25056 18262 25057
rect 17946 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18262 25056
rect 17946 24991 18262 24992
rect 27946 25056 28262 25057
rect 27946 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28262 25056
rect 27946 24991 28262 24992
rect 1301 24986 1367 24989
rect 0 24984 1367 24986
rect 0 24928 1306 24984
rect 1362 24928 1367 24984
rect 0 24926 1367 24928
rect 0 24896 800 24926
rect 1301 24923 1367 24926
rect 8845 24986 8911 24989
rect 9581 24986 9647 24989
rect 8845 24984 9647 24986
rect 8845 24928 8850 24984
rect 8906 24928 9586 24984
rect 9642 24928 9647 24984
rect 8845 24926 9647 24928
rect 8845 24923 8911 24926
rect 9581 24923 9647 24926
rect 26693 24986 26759 24989
rect 27705 24986 27771 24989
rect 28809 24986 28875 24989
rect 26693 24984 27771 24986
rect 26693 24928 26698 24984
rect 26754 24928 27710 24984
rect 27766 24928 27771 24984
rect 26693 24926 27771 24928
rect 26693 24923 26759 24926
rect 27705 24923 27771 24926
rect 28766 24984 28875 24986
rect 28766 24928 28814 24984
rect 28870 24928 28875 24984
rect 28766 24923 28875 24928
rect 26141 24850 26207 24853
rect 27613 24850 27679 24853
rect 28766 24850 28826 24923
rect 26141 24848 28826 24850
rect 26141 24792 26146 24848
rect 26202 24792 27618 24848
rect 27674 24792 28826 24848
rect 26141 24790 28826 24792
rect 26141 24787 26207 24790
rect 27613 24787 27679 24790
rect 28809 24714 28875 24717
rect 28950 24714 29010 25059
rect 37946 25056 38262 25057
rect 37946 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38262 25056
rect 37946 24991 38262 24992
rect 47946 25056 48262 25057
rect 47946 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48262 25056
rect 47946 24991 48262 24992
rect 28809 24712 29010 24714
rect 28809 24656 28814 24712
rect 28870 24656 29010 24712
rect 28809 24654 29010 24656
rect 49141 24714 49207 24717
rect 50200 24714 51000 24744
rect 49141 24712 51000 24714
rect 49141 24656 49146 24712
rect 49202 24656 51000 24712
rect 49141 24654 51000 24656
rect 28809 24651 28875 24654
rect 49141 24651 49207 24654
rect 50200 24624 51000 24654
rect 2946 24512 3262 24513
rect 2946 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3262 24512
rect 2946 24447 3262 24448
rect 12946 24512 13262 24513
rect 12946 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13262 24512
rect 12946 24447 13262 24448
rect 22946 24512 23262 24513
rect 22946 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23262 24512
rect 22946 24447 23262 24448
rect 32946 24512 33262 24513
rect 32946 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33262 24512
rect 32946 24447 33262 24448
rect 42946 24512 43262 24513
rect 42946 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43262 24512
rect 42946 24447 43262 24448
rect 25497 24306 25563 24309
rect 25630 24306 25636 24308
rect 25497 24304 25636 24306
rect 25497 24248 25502 24304
rect 25558 24248 25636 24304
rect 25497 24246 25636 24248
rect 25497 24243 25563 24246
rect 25630 24244 25636 24246
rect 25700 24244 25706 24308
rect 27705 24172 27771 24173
rect 27654 24108 27660 24172
rect 27724 24170 27771 24172
rect 27724 24168 27816 24170
rect 27766 24112 27816 24168
rect 27724 24110 27816 24112
rect 27724 24108 27771 24110
rect 27705 24107 27771 24108
rect 49141 24034 49207 24037
rect 50200 24034 51000 24064
rect 49141 24032 51000 24034
rect 49141 23976 49146 24032
rect 49202 23976 51000 24032
rect 49141 23974 51000 23976
rect 49141 23971 49207 23974
rect 7946 23968 8262 23969
rect 7946 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8262 23968
rect 7946 23903 8262 23904
rect 17946 23968 18262 23969
rect 17946 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18262 23968
rect 17946 23903 18262 23904
rect 27946 23968 28262 23969
rect 27946 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28262 23968
rect 27946 23903 28262 23904
rect 37946 23968 38262 23969
rect 37946 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38262 23968
rect 37946 23903 38262 23904
rect 47946 23968 48262 23969
rect 47946 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48262 23968
rect 50200 23944 51000 23974
rect 47946 23903 48262 23904
rect 22134 23564 22140 23628
rect 22204 23626 22210 23628
rect 22461 23626 22527 23629
rect 23381 23626 23447 23629
rect 22204 23624 23447 23626
rect 22204 23568 22466 23624
rect 22522 23568 23386 23624
rect 23442 23568 23447 23624
rect 22204 23566 23447 23568
rect 22204 23564 22210 23566
rect 22461 23563 22527 23566
rect 23381 23563 23447 23566
rect 26233 23626 26299 23629
rect 28901 23626 28967 23629
rect 26233 23624 28967 23626
rect 26233 23568 26238 23624
rect 26294 23568 28906 23624
rect 28962 23568 28967 23624
rect 26233 23566 28967 23568
rect 26233 23563 26299 23566
rect 28901 23563 28967 23566
rect 23381 23490 23447 23493
rect 28533 23490 28599 23493
rect 29913 23490 29979 23493
rect 23381 23488 29979 23490
rect 23381 23432 23386 23488
rect 23442 23432 28538 23488
rect 28594 23432 29918 23488
rect 29974 23432 29979 23488
rect 23381 23430 29979 23432
rect 23381 23427 23447 23430
rect 28533 23427 28599 23430
rect 29913 23427 29979 23430
rect 2946 23424 3262 23425
rect 2946 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3262 23424
rect 2946 23359 3262 23360
rect 12946 23424 13262 23425
rect 12946 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13262 23424
rect 12946 23359 13262 23360
rect 22946 23424 23262 23425
rect 22946 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23262 23424
rect 22946 23359 23262 23360
rect 32946 23424 33262 23425
rect 32946 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33262 23424
rect 32946 23359 33262 23360
rect 42946 23424 43262 23425
rect 42946 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43262 23424
rect 42946 23359 43262 23360
rect 49141 23354 49207 23357
rect 50200 23354 51000 23384
rect 49141 23352 51000 23354
rect 49141 23296 49146 23352
rect 49202 23296 51000 23352
rect 49141 23294 51000 23296
rect 49141 23291 49207 23294
rect 50200 23264 51000 23294
rect 22502 22884 22508 22948
rect 22572 22946 22578 22948
rect 25037 22946 25103 22949
rect 22572 22944 25103 22946
rect 22572 22888 25042 22944
rect 25098 22888 25103 22944
rect 22572 22886 25103 22888
rect 22572 22884 22578 22886
rect 25037 22883 25103 22886
rect 7946 22880 8262 22881
rect 7946 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8262 22880
rect 7946 22815 8262 22816
rect 17946 22880 18262 22881
rect 17946 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18262 22880
rect 17946 22815 18262 22816
rect 27946 22880 28262 22881
rect 27946 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28262 22880
rect 27946 22815 28262 22816
rect 37946 22880 38262 22881
rect 37946 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38262 22880
rect 37946 22815 38262 22816
rect 47946 22880 48262 22881
rect 47946 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48262 22880
rect 47946 22815 48262 22816
rect 0 22674 800 22704
rect 1301 22674 1367 22677
rect 0 22672 1367 22674
rect 0 22616 1306 22672
rect 1362 22616 1367 22672
rect 0 22614 1367 22616
rect 0 22584 800 22614
rect 1301 22611 1367 22614
rect 8937 22674 9003 22677
rect 30373 22674 30439 22677
rect 8937 22672 30439 22674
rect 8937 22616 8942 22672
rect 8998 22616 30378 22672
rect 30434 22616 30439 22672
rect 8937 22614 30439 22616
rect 8937 22611 9003 22614
rect 30373 22611 30439 22614
rect 49141 22674 49207 22677
rect 50200 22674 51000 22704
rect 49141 22672 51000 22674
rect 49141 22616 49146 22672
rect 49202 22616 51000 22672
rect 49141 22614 51000 22616
rect 49141 22611 49207 22614
rect 50200 22584 51000 22614
rect 25957 22538 26023 22541
rect 27797 22538 27863 22541
rect 25957 22536 27863 22538
rect 25957 22480 25962 22536
rect 26018 22480 27802 22536
rect 27858 22480 27863 22536
rect 25957 22478 27863 22480
rect 25957 22475 26023 22478
rect 27797 22475 27863 22478
rect 2946 22336 3262 22337
rect 2946 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3262 22336
rect 2946 22271 3262 22272
rect 12946 22336 13262 22337
rect 12946 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13262 22336
rect 12946 22271 13262 22272
rect 22946 22336 23262 22337
rect 22946 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23262 22336
rect 22946 22271 23262 22272
rect 32946 22336 33262 22337
rect 32946 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33262 22336
rect 32946 22271 33262 22272
rect 42946 22336 43262 22337
rect 42946 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43262 22336
rect 42946 22271 43262 22272
rect 8937 22130 9003 22133
rect 9397 22130 9463 22133
rect 8937 22128 9463 22130
rect 8937 22072 8942 22128
rect 8998 22072 9402 22128
rect 9458 22072 9463 22128
rect 8937 22070 9463 22072
rect 8937 22067 9003 22070
rect 9397 22067 9463 22070
rect 28533 21994 28599 21997
rect 30782 21994 30788 21996
rect 28533 21992 30788 21994
rect 28533 21936 28538 21992
rect 28594 21936 30788 21992
rect 28533 21934 30788 21936
rect 28533 21931 28599 21934
rect 30782 21932 30788 21934
rect 30852 21932 30858 21996
rect 49141 21994 49207 21997
rect 50200 21994 51000 22024
rect 49141 21992 51000 21994
rect 49141 21936 49146 21992
rect 49202 21936 51000 21992
rect 49141 21934 51000 21936
rect 49141 21931 49207 21934
rect 50200 21904 51000 21934
rect 7946 21792 8262 21793
rect 7946 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8262 21792
rect 7946 21727 8262 21728
rect 17946 21792 18262 21793
rect 17946 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18262 21792
rect 17946 21727 18262 21728
rect 27946 21792 28262 21793
rect 27946 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28262 21792
rect 27946 21727 28262 21728
rect 37946 21792 38262 21793
rect 37946 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38262 21792
rect 37946 21727 38262 21728
rect 47946 21792 48262 21793
rect 47946 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48262 21792
rect 47946 21727 48262 21728
rect 49141 21314 49207 21317
rect 50200 21314 51000 21344
rect 49141 21312 51000 21314
rect 49141 21256 49146 21312
rect 49202 21256 51000 21312
rect 49141 21254 51000 21256
rect 49141 21251 49207 21254
rect 2946 21248 3262 21249
rect 2946 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3262 21248
rect 2946 21183 3262 21184
rect 12946 21248 13262 21249
rect 12946 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13262 21248
rect 12946 21183 13262 21184
rect 22946 21248 23262 21249
rect 22946 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23262 21248
rect 22946 21183 23262 21184
rect 32946 21248 33262 21249
rect 32946 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33262 21248
rect 32946 21183 33262 21184
rect 42946 21248 43262 21249
rect 42946 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43262 21248
rect 50200 21224 51000 21254
rect 42946 21183 43262 21184
rect 7946 20704 8262 20705
rect 7946 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8262 20704
rect 7946 20639 8262 20640
rect 17946 20704 18262 20705
rect 17946 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18262 20704
rect 17946 20639 18262 20640
rect 27946 20704 28262 20705
rect 27946 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28262 20704
rect 27946 20639 28262 20640
rect 37946 20704 38262 20705
rect 37946 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38262 20704
rect 37946 20639 38262 20640
rect 47946 20704 48262 20705
rect 47946 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48262 20704
rect 47946 20639 48262 20640
rect 30465 20636 30531 20637
rect 30414 20572 30420 20636
rect 30484 20634 30531 20636
rect 35157 20636 35223 20637
rect 30484 20632 30576 20634
rect 30526 20576 30576 20632
rect 30484 20574 30576 20576
rect 35157 20632 35204 20636
rect 35268 20634 35274 20636
rect 49141 20634 49207 20637
rect 50200 20634 51000 20664
rect 35157 20576 35162 20632
rect 30484 20572 30531 20574
rect 30465 20571 30531 20572
rect 35157 20572 35204 20576
rect 35268 20574 35314 20634
rect 49141 20632 51000 20634
rect 49141 20576 49146 20632
rect 49202 20576 51000 20632
rect 49141 20574 51000 20576
rect 35268 20572 35274 20574
rect 35157 20571 35223 20572
rect 49141 20571 49207 20574
rect 50200 20544 51000 20574
rect 22553 20498 22619 20501
rect 23289 20498 23355 20501
rect 22553 20496 23355 20498
rect 22553 20440 22558 20496
rect 22614 20440 23294 20496
rect 23350 20440 23355 20496
rect 22553 20438 23355 20440
rect 22553 20435 22619 20438
rect 23289 20435 23355 20438
rect 0 20362 800 20392
rect 1301 20362 1367 20365
rect 0 20360 1367 20362
rect 0 20304 1306 20360
rect 1362 20304 1367 20360
rect 0 20302 1367 20304
rect 0 20272 800 20302
rect 1301 20299 1367 20302
rect 2946 20160 3262 20161
rect 2946 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3262 20160
rect 2946 20095 3262 20096
rect 12946 20160 13262 20161
rect 12946 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13262 20160
rect 12946 20095 13262 20096
rect 22946 20160 23262 20161
rect 22946 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23262 20160
rect 22946 20095 23262 20096
rect 32946 20160 33262 20161
rect 32946 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33262 20160
rect 32946 20095 33262 20096
rect 42946 20160 43262 20161
rect 42946 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43262 20160
rect 42946 20095 43262 20096
rect 49141 19954 49207 19957
rect 50200 19954 51000 19984
rect 49141 19952 51000 19954
rect 49141 19896 49146 19952
rect 49202 19896 51000 19952
rect 49141 19894 51000 19896
rect 49141 19891 49207 19894
rect 50200 19864 51000 19894
rect 7946 19616 8262 19617
rect 7946 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8262 19616
rect 7946 19551 8262 19552
rect 17946 19616 18262 19617
rect 17946 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18262 19616
rect 17946 19551 18262 19552
rect 27946 19616 28262 19617
rect 27946 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28262 19616
rect 27946 19551 28262 19552
rect 37946 19616 38262 19617
rect 37946 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38262 19616
rect 37946 19551 38262 19552
rect 47946 19616 48262 19617
rect 47946 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48262 19616
rect 47946 19551 48262 19552
rect 29085 19410 29151 19413
rect 34973 19410 35039 19413
rect 29085 19408 35039 19410
rect 29085 19352 29090 19408
rect 29146 19352 34978 19408
rect 35034 19352 35039 19408
rect 29085 19350 35039 19352
rect 29085 19347 29151 19350
rect 34973 19347 35039 19350
rect 27061 19274 27127 19277
rect 28533 19274 28599 19277
rect 27061 19272 28599 19274
rect 27061 19216 27066 19272
rect 27122 19216 28538 19272
rect 28594 19216 28599 19272
rect 27061 19214 28599 19216
rect 27061 19211 27127 19214
rect 28533 19211 28599 19214
rect 32806 19212 32812 19276
rect 32876 19274 32882 19276
rect 38510 19274 38516 19276
rect 32876 19214 38516 19274
rect 32876 19212 32882 19214
rect 38510 19212 38516 19214
rect 38580 19212 38586 19276
rect 49141 19274 49207 19277
rect 50200 19274 51000 19304
rect 49141 19272 51000 19274
rect 49141 19216 49146 19272
rect 49202 19216 51000 19272
rect 49141 19214 51000 19216
rect 49141 19211 49207 19214
rect 50200 19184 51000 19214
rect 2946 19072 3262 19073
rect 2946 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3262 19072
rect 2946 19007 3262 19008
rect 12946 19072 13262 19073
rect 12946 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13262 19072
rect 12946 19007 13262 19008
rect 22946 19072 23262 19073
rect 22946 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23262 19072
rect 22946 19007 23262 19008
rect 32946 19072 33262 19073
rect 32946 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33262 19072
rect 32946 19007 33262 19008
rect 42946 19072 43262 19073
rect 42946 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43262 19072
rect 42946 19007 43262 19008
rect 22686 18804 22692 18868
rect 22756 18866 22762 18868
rect 22829 18866 22895 18869
rect 22756 18864 22895 18866
rect 22756 18808 22834 18864
rect 22890 18808 22895 18864
rect 22756 18806 22895 18808
rect 22756 18804 22762 18806
rect 22829 18803 22895 18806
rect 49141 18594 49207 18597
rect 50200 18594 51000 18624
rect 49141 18592 51000 18594
rect 49141 18536 49146 18592
rect 49202 18536 51000 18592
rect 49141 18534 51000 18536
rect 49141 18531 49207 18534
rect 7946 18528 8262 18529
rect 7946 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8262 18528
rect 7946 18463 8262 18464
rect 17946 18528 18262 18529
rect 17946 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18262 18528
rect 17946 18463 18262 18464
rect 27946 18528 28262 18529
rect 27946 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28262 18528
rect 27946 18463 28262 18464
rect 37946 18528 38262 18529
rect 37946 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38262 18528
rect 37946 18463 38262 18464
rect 47946 18528 48262 18529
rect 47946 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48262 18528
rect 50200 18504 51000 18534
rect 47946 18463 48262 18464
rect 0 18050 800 18080
rect 1301 18050 1367 18053
rect 0 18048 1367 18050
rect 0 17992 1306 18048
rect 1362 17992 1367 18048
rect 0 17990 1367 17992
rect 0 17960 800 17990
rect 1301 17987 1367 17990
rect 29085 18050 29151 18053
rect 30966 18050 30972 18052
rect 29085 18048 30972 18050
rect 29085 17992 29090 18048
rect 29146 17992 30972 18048
rect 29085 17990 30972 17992
rect 29085 17987 29151 17990
rect 30966 17988 30972 17990
rect 31036 17988 31042 18052
rect 2946 17984 3262 17985
rect 2946 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3262 17984
rect 2946 17919 3262 17920
rect 12946 17984 13262 17985
rect 12946 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13262 17984
rect 12946 17919 13262 17920
rect 22946 17984 23262 17985
rect 22946 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23262 17984
rect 22946 17919 23262 17920
rect 32946 17984 33262 17985
rect 32946 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33262 17984
rect 32946 17919 33262 17920
rect 42946 17984 43262 17985
rect 42946 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43262 17984
rect 42946 17919 43262 17920
rect 49141 17914 49207 17917
rect 50200 17914 51000 17944
rect 49141 17912 51000 17914
rect 49141 17856 49146 17912
rect 49202 17856 51000 17912
rect 49141 17854 51000 17856
rect 49141 17851 49207 17854
rect 50200 17824 51000 17854
rect 7946 17440 8262 17441
rect 7946 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8262 17440
rect 7946 17375 8262 17376
rect 17946 17440 18262 17441
rect 17946 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18262 17440
rect 17946 17375 18262 17376
rect 27946 17440 28262 17441
rect 27946 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28262 17440
rect 27946 17375 28262 17376
rect 37946 17440 38262 17441
rect 37946 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38262 17440
rect 37946 17375 38262 17376
rect 47946 17440 48262 17441
rect 47946 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48262 17440
rect 47946 17375 48262 17376
rect 28809 17370 28875 17373
rect 32806 17370 32812 17372
rect 28809 17368 32812 17370
rect 28809 17312 28814 17368
rect 28870 17312 32812 17368
rect 28809 17310 32812 17312
rect 28809 17307 28875 17310
rect 32806 17308 32812 17310
rect 32876 17308 32882 17372
rect 49141 17234 49207 17237
rect 50200 17234 51000 17264
rect 49141 17232 51000 17234
rect 49141 17176 49146 17232
rect 49202 17176 51000 17232
rect 49141 17174 51000 17176
rect 49141 17171 49207 17174
rect 50200 17144 51000 17174
rect 2946 16896 3262 16897
rect 2946 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3262 16896
rect 2946 16831 3262 16832
rect 12946 16896 13262 16897
rect 12946 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13262 16896
rect 12946 16831 13262 16832
rect 22946 16896 23262 16897
rect 22946 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23262 16896
rect 22946 16831 23262 16832
rect 32946 16896 33262 16897
rect 32946 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33262 16896
rect 32946 16831 33262 16832
rect 42946 16896 43262 16897
rect 42946 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43262 16896
rect 42946 16831 43262 16832
rect 32622 16628 32628 16692
rect 32692 16690 32698 16692
rect 34053 16690 34119 16693
rect 32692 16688 34119 16690
rect 32692 16632 34058 16688
rect 34114 16632 34119 16688
rect 32692 16630 34119 16632
rect 32692 16628 32698 16630
rect 34053 16627 34119 16630
rect 49141 16554 49207 16557
rect 50200 16554 51000 16584
rect 49141 16552 51000 16554
rect 49141 16496 49146 16552
rect 49202 16496 51000 16552
rect 49141 16494 51000 16496
rect 49141 16491 49207 16494
rect 50200 16464 51000 16494
rect 7946 16352 8262 16353
rect 7946 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8262 16352
rect 7946 16287 8262 16288
rect 17946 16352 18262 16353
rect 17946 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18262 16352
rect 17946 16287 18262 16288
rect 27946 16352 28262 16353
rect 27946 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28262 16352
rect 27946 16287 28262 16288
rect 37946 16352 38262 16353
rect 37946 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38262 16352
rect 37946 16287 38262 16288
rect 47946 16352 48262 16353
rect 47946 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48262 16352
rect 47946 16287 48262 16288
rect 49141 15874 49207 15877
rect 50200 15874 51000 15904
rect 49141 15872 51000 15874
rect 49141 15816 49146 15872
rect 49202 15816 51000 15872
rect 49141 15814 51000 15816
rect 49141 15811 49207 15814
rect 2946 15808 3262 15809
rect 0 15738 800 15768
rect 2946 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3262 15808
rect 2946 15743 3262 15744
rect 12946 15808 13262 15809
rect 12946 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13262 15808
rect 12946 15743 13262 15744
rect 22946 15808 23262 15809
rect 22946 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23262 15808
rect 22946 15743 23262 15744
rect 32946 15808 33262 15809
rect 32946 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33262 15808
rect 32946 15743 33262 15744
rect 42946 15808 43262 15809
rect 42946 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43262 15808
rect 50200 15784 51000 15814
rect 42946 15743 43262 15744
rect 1301 15738 1367 15741
rect 0 15736 1367 15738
rect 0 15680 1306 15736
rect 1362 15680 1367 15736
rect 0 15678 1367 15680
rect 0 15648 800 15678
rect 1301 15675 1367 15678
rect 7946 15264 8262 15265
rect 7946 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8262 15264
rect 7946 15199 8262 15200
rect 17946 15264 18262 15265
rect 17946 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18262 15264
rect 17946 15199 18262 15200
rect 27946 15264 28262 15265
rect 27946 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28262 15264
rect 27946 15199 28262 15200
rect 37946 15264 38262 15265
rect 37946 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38262 15264
rect 37946 15199 38262 15200
rect 47946 15264 48262 15265
rect 47946 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48262 15264
rect 47946 15199 48262 15200
rect 49141 15194 49207 15197
rect 50200 15194 51000 15224
rect 49141 15192 51000 15194
rect 49141 15136 49146 15192
rect 49202 15136 51000 15192
rect 49141 15134 51000 15136
rect 49141 15131 49207 15134
rect 50200 15104 51000 15134
rect 2946 14720 3262 14721
rect 2946 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3262 14720
rect 2946 14655 3262 14656
rect 12946 14720 13262 14721
rect 12946 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13262 14720
rect 12946 14655 13262 14656
rect 22946 14720 23262 14721
rect 22946 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23262 14720
rect 22946 14655 23262 14656
rect 32946 14720 33262 14721
rect 32946 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33262 14720
rect 32946 14655 33262 14656
rect 42946 14720 43262 14721
rect 42946 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43262 14720
rect 42946 14655 43262 14656
rect 49141 14514 49207 14517
rect 50200 14514 51000 14544
rect 49141 14512 51000 14514
rect 49141 14456 49146 14512
rect 49202 14456 51000 14512
rect 49141 14454 51000 14456
rect 49141 14451 49207 14454
rect 50200 14424 51000 14454
rect 7946 14176 8262 14177
rect 7946 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8262 14176
rect 7946 14111 8262 14112
rect 17946 14176 18262 14177
rect 17946 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18262 14176
rect 17946 14111 18262 14112
rect 27946 14176 28262 14177
rect 27946 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28262 14176
rect 27946 14111 28262 14112
rect 37946 14176 38262 14177
rect 37946 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38262 14176
rect 37946 14111 38262 14112
rect 47946 14176 48262 14177
rect 47946 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48262 14176
rect 47946 14111 48262 14112
rect 49141 13834 49207 13837
rect 50200 13834 51000 13864
rect 49141 13832 51000 13834
rect 49141 13776 49146 13832
rect 49202 13776 51000 13832
rect 49141 13774 51000 13776
rect 49141 13771 49207 13774
rect 50200 13744 51000 13774
rect 2946 13632 3262 13633
rect 2946 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3262 13632
rect 2946 13567 3262 13568
rect 12946 13632 13262 13633
rect 12946 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13262 13632
rect 12946 13567 13262 13568
rect 22946 13632 23262 13633
rect 22946 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23262 13632
rect 22946 13567 23262 13568
rect 32946 13632 33262 13633
rect 32946 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33262 13632
rect 32946 13567 33262 13568
rect 42946 13632 43262 13633
rect 42946 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43262 13632
rect 42946 13567 43262 13568
rect 0 13426 800 13456
rect 2773 13426 2839 13429
rect 0 13424 2839 13426
rect 0 13368 2778 13424
rect 2834 13368 2839 13424
rect 0 13366 2839 13368
rect 0 13336 800 13366
rect 2773 13363 2839 13366
rect 49141 13154 49207 13157
rect 50200 13154 51000 13184
rect 49141 13152 51000 13154
rect 49141 13096 49146 13152
rect 49202 13096 51000 13152
rect 49141 13094 51000 13096
rect 49141 13091 49207 13094
rect 7946 13088 8262 13089
rect 7946 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8262 13088
rect 7946 13023 8262 13024
rect 17946 13088 18262 13089
rect 17946 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18262 13088
rect 17946 13023 18262 13024
rect 27946 13088 28262 13089
rect 27946 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28262 13088
rect 27946 13023 28262 13024
rect 37946 13088 38262 13089
rect 37946 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38262 13088
rect 37946 13023 38262 13024
rect 47946 13088 48262 13089
rect 47946 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48262 13088
rect 50200 13064 51000 13094
rect 47946 13023 48262 13024
rect 28809 12610 28875 12613
rect 28766 12608 28875 12610
rect 28766 12552 28814 12608
rect 28870 12552 28875 12608
rect 28766 12547 28875 12552
rect 2946 12544 3262 12545
rect 2946 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3262 12544
rect 2946 12479 3262 12480
rect 12946 12544 13262 12545
rect 12946 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13262 12544
rect 12946 12479 13262 12480
rect 22946 12544 23262 12545
rect 22946 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23262 12544
rect 22946 12479 23262 12480
rect 28533 12474 28599 12477
rect 28766 12474 28826 12547
rect 32946 12544 33262 12545
rect 32946 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33262 12544
rect 32946 12479 33262 12480
rect 42946 12544 43262 12545
rect 42946 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43262 12544
rect 42946 12479 43262 12480
rect 28533 12472 28826 12474
rect 28533 12416 28538 12472
rect 28594 12416 28826 12472
rect 28533 12414 28826 12416
rect 49141 12474 49207 12477
rect 50200 12474 51000 12504
rect 49141 12472 51000 12474
rect 49141 12416 49146 12472
rect 49202 12416 51000 12472
rect 49141 12414 51000 12416
rect 28533 12411 28599 12414
rect 49141 12411 49207 12414
rect 50200 12384 51000 12414
rect 38510 12276 38516 12340
rect 38580 12338 38586 12340
rect 38929 12338 38995 12341
rect 38580 12336 38995 12338
rect 38580 12280 38934 12336
rect 38990 12280 38995 12336
rect 38580 12278 38995 12280
rect 38580 12276 38586 12278
rect 38929 12275 38995 12278
rect 7946 12000 8262 12001
rect 7946 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8262 12000
rect 7946 11935 8262 11936
rect 17946 12000 18262 12001
rect 17946 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18262 12000
rect 17946 11935 18262 11936
rect 27946 12000 28262 12001
rect 27946 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28262 12000
rect 27946 11935 28262 11936
rect 37946 12000 38262 12001
rect 37946 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38262 12000
rect 37946 11935 38262 11936
rect 47946 12000 48262 12001
rect 47946 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48262 12000
rect 47946 11935 48262 11936
rect 49141 11794 49207 11797
rect 50200 11794 51000 11824
rect 49141 11792 51000 11794
rect 49141 11736 49146 11792
rect 49202 11736 51000 11792
rect 49141 11734 51000 11736
rect 49141 11731 49207 11734
rect 50200 11704 51000 11734
rect 2946 11456 3262 11457
rect 2946 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3262 11456
rect 2946 11391 3262 11392
rect 12946 11456 13262 11457
rect 12946 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13262 11456
rect 12946 11391 13262 11392
rect 22946 11456 23262 11457
rect 22946 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23262 11456
rect 22946 11391 23262 11392
rect 32946 11456 33262 11457
rect 32946 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33262 11456
rect 32946 11391 33262 11392
rect 42946 11456 43262 11457
rect 42946 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43262 11456
rect 42946 11391 43262 11392
rect 0 11114 800 11144
rect 3325 11114 3391 11117
rect 0 11112 3391 11114
rect 0 11056 3330 11112
rect 3386 11056 3391 11112
rect 0 11054 3391 11056
rect 0 11024 800 11054
rect 3325 11051 3391 11054
rect 49141 11114 49207 11117
rect 50200 11114 51000 11144
rect 49141 11112 51000 11114
rect 49141 11056 49146 11112
rect 49202 11056 51000 11112
rect 49141 11054 51000 11056
rect 49141 11051 49207 11054
rect 50200 11024 51000 11054
rect 7946 10912 8262 10913
rect 7946 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8262 10912
rect 7946 10847 8262 10848
rect 17946 10912 18262 10913
rect 17946 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18262 10912
rect 17946 10847 18262 10848
rect 27946 10912 28262 10913
rect 27946 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28262 10912
rect 27946 10847 28262 10848
rect 37946 10912 38262 10913
rect 37946 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38262 10912
rect 37946 10847 38262 10848
rect 47946 10912 48262 10913
rect 47946 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48262 10912
rect 47946 10847 48262 10848
rect 49141 10434 49207 10437
rect 50200 10434 51000 10464
rect 49141 10432 51000 10434
rect 49141 10376 49146 10432
rect 49202 10376 51000 10432
rect 49141 10374 51000 10376
rect 49141 10371 49207 10374
rect 2946 10368 3262 10369
rect 2946 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3262 10368
rect 2946 10303 3262 10304
rect 12946 10368 13262 10369
rect 12946 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13262 10368
rect 12946 10303 13262 10304
rect 22946 10368 23262 10369
rect 22946 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23262 10368
rect 22946 10303 23262 10304
rect 32946 10368 33262 10369
rect 32946 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33262 10368
rect 32946 10303 33262 10304
rect 42946 10368 43262 10369
rect 42946 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43262 10368
rect 50200 10344 51000 10374
rect 42946 10303 43262 10304
rect 7946 9824 8262 9825
rect 7946 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8262 9824
rect 7946 9759 8262 9760
rect 17946 9824 18262 9825
rect 17946 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18262 9824
rect 17946 9759 18262 9760
rect 27946 9824 28262 9825
rect 27946 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28262 9824
rect 27946 9759 28262 9760
rect 37946 9824 38262 9825
rect 37946 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38262 9824
rect 37946 9759 38262 9760
rect 47946 9824 48262 9825
rect 47946 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48262 9824
rect 47946 9759 48262 9760
rect 49141 9754 49207 9757
rect 50200 9754 51000 9784
rect 49141 9752 51000 9754
rect 49141 9696 49146 9752
rect 49202 9696 51000 9752
rect 49141 9694 51000 9696
rect 49141 9691 49207 9694
rect 50200 9664 51000 9694
rect 2946 9280 3262 9281
rect 2946 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3262 9280
rect 2946 9215 3262 9216
rect 12946 9280 13262 9281
rect 12946 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13262 9280
rect 12946 9215 13262 9216
rect 22946 9280 23262 9281
rect 22946 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23262 9280
rect 22946 9215 23262 9216
rect 32946 9280 33262 9281
rect 32946 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33262 9280
rect 32946 9215 33262 9216
rect 42946 9280 43262 9281
rect 42946 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43262 9280
rect 42946 9215 43262 9216
rect 49141 9074 49207 9077
rect 50200 9074 51000 9104
rect 49141 9072 51000 9074
rect 49141 9016 49146 9072
rect 49202 9016 51000 9072
rect 49141 9014 51000 9016
rect 49141 9011 49207 9014
rect 50200 8984 51000 9014
rect 0 8802 800 8832
rect 3325 8802 3391 8805
rect 0 8800 3391 8802
rect 0 8744 3330 8800
rect 3386 8744 3391 8800
rect 0 8742 3391 8744
rect 0 8712 800 8742
rect 3325 8739 3391 8742
rect 7946 8736 8262 8737
rect 7946 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8262 8736
rect 7946 8671 8262 8672
rect 17946 8736 18262 8737
rect 17946 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18262 8736
rect 17946 8671 18262 8672
rect 27946 8736 28262 8737
rect 27946 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28262 8736
rect 27946 8671 28262 8672
rect 37946 8736 38262 8737
rect 37946 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38262 8736
rect 37946 8671 38262 8672
rect 47946 8736 48262 8737
rect 47946 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48262 8736
rect 47946 8671 48262 8672
rect 49141 8394 49207 8397
rect 50200 8394 51000 8424
rect 49141 8392 51000 8394
rect 49141 8336 49146 8392
rect 49202 8336 51000 8392
rect 49141 8334 51000 8336
rect 49141 8331 49207 8334
rect 50200 8304 51000 8334
rect 2946 8192 3262 8193
rect 2946 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3262 8192
rect 2946 8127 3262 8128
rect 12946 8192 13262 8193
rect 12946 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13262 8192
rect 12946 8127 13262 8128
rect 22946 8192 23262 8193
rect 22946 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23262 8192
rect 22946 8127 23262 8128
rect 32946 8192 33262 8193
rect 32946 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33262 8192
rect 32946 8127 33262 8128
rect 42946 8192 43262 8193
rect 42946 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43262 8192
rect 42946 8127 43262 8128
rect 49141 7714 49207 7717
rect 50200 7714 51000 7744
rect 49141 7712 51000 7714
rect 49141 7656 49146 7712
rect 49202 7656 51000 7712
rect 49141 7654 51000 7656
rect 49141 7651 49207 7654
rect 7946 7648 8262 7649
rect 7946 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8262 7648
rect 7946 7583 8262 7584
rect 17946 7648 18262 7649
rect 17946 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18262 7648
rect 17946 7583 18262 7584
rect 27946 7648 28262 7649
rect 27946 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28262 7648
rect 27946 7583 28262 7584
rect 37946 7648 38262 7649
rect 37946 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38262 7648
rect 37946 7583 38262 7584
rect 47946 7648 48262 7649
rect 47946 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48262 7648
rect 50200 7624 51000 7654
rect 47946 7583 48262 7584
rect 2946 7104 3262 7105
rect 2946 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3262 7104
rect 2946 7039 3262 7040
rect 12946 7104 13262 7105
rect 12946 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13262 7104
rect 12946 7039 13262 7040
rect 22946 7104 23262 7105
rect 22946 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23262 7104
rect 22946 7039 23262 7040
rect 32946 7104 33262 7105
rect 32946 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33262 7104
rect 32946 7039 33262 7040
rect 42946 7104 43262 7105
rect 42946 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43262 7104
rect 42946 7039 43262 7040
rect 49141 7034 49207 7037
rect 50200 7034 51000 7064
rect 49141 7032 51000 7034
rect 49141 6976 49146 7032
rect 49202 6976 51000 7032
rect 49141 6974 51000 6976
rect 49141 6971 49207 6974
rect 50200 6944 51000 6974
rect 7946 6560 8262 6561
rect 0 6490 800 6520
rect 7946 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8262 6560
rect 7946 6495 8262 6496
rect 17946 6560 18262 6561
rect 17946 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18262 6560
rect 17946 6495 18262 6496
rect 27946 6560 28262 6561
rect 27946 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28262 6560
rect 27946 6495 28262 6496
rect 37946 6560 38262 6561
rect 37946 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38262 6560
rect 37946 6495 38262 6496
rect 47946 6560 48262 6561
rect 47946 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48262 6560
rect 47946 6495 48262 6496
rect 3417 6490 3483 6493
rect 0 6488 3483 6490
rect 0 6432 3422 6488
rect 3478 6432 3483 6488
rect 0 6430 3483 6432
rect 0 6400 800 6430
rect 3417 6427 3483 6430
rect 49141 6354 49207 6357
rect 50200 6354 51000 6384
rect 49141 6352 51000 6354
rect 49141 6296 49146 6352
rect 49202 6296 51000 6352
rect 49141 6294 51000 6296
rect 49141 6291 49207 6294
rect 50200 6264 51000 6294
rect 2946 6016 3262 6017
rect 2946 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3262 6016
rect 2946 5951 3262 5952
rect 12946 6016 13262 6017
rect 12946 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13262 6016
rect 12946 5951 13262 5952
rect 22946 6016 23262 6017
rect 22946 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23262 6016
rect 22946 5951 23262 5952
rect 32946 6016 33262 6017
rect 32946 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33262 6016
rect 32946 5951 33262 5952
rect 42946 6016 43262 6017
rect 42946 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43262 6016
rect 42946 5951 43262 5952
rect 49141 5674 49207 5677
rect 50200 5674 51000 5704
rect 49141 5672 51000 5674
rect 49141 5616 49146 5672
rect 49202 5616 51000 5672
rect 49141 5614 51000 5616
rect 49141 5611 49207 5614
rect 50200 5584 51000 5614
rect 7946 5472 8262 5473
rect 7946 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8262 5472
rect 7946 5407 8262 5408
rect 17946 5472 18262 5473
rect 17946 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18262 5472
rect 17946 5407 18262 5408
rect 27946 5472 28262 5473
rect 27946 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28262 5472
rect 27946 5407 28262 5408
rect 37946 5472 38262 5473
rect 37946 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38262 5472
rect 37946 5407 38262 5408
rect 47946 5472 48262 5473
rect 47946 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48262 5472
rect 47946 5407 48262 5408
rect 49325 4994 49391 4997
rect 50200 4994 51000 5024
rect 49325 4992 51000 4994
rect 49325 4936 49330 4992
rect 49386 4936 51000 4992
rect 49325 4934 51000 4936
rect 49325 4931 49391 4934
rect 2946 4928 3262 4929
rect 2946 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3262 4928
rect 2946 4863 3262 4864
rect 12946 4928 13262 4929
rect 12946 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13262 4928
rect 12946 4863 13262 4864
rect 22946 4928 23262 4929
rect 22946 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23262 4928
rect 22946 4863 23262 4864
rect 32946 4928 33262 4929
rect 32946 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33262 4928
rect 32946 4863 33262 4864
rect 42946 4928 43262 4929
rect 42946 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43262 4928
rect 50200 4904 51000 4934
rect 42946 4863 43262 4864
rect 7946 4384 8262 4385
rect 7946 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8262 4384
rect 7946 4319 8262 4320
rect 17946 4384 18262 4385
rect 17946 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18262 4384
rect 17946 4319 18262 4320
rect 27946 4384 28262 4385
rect 27946 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28262 4384
rect 27946 4319 28262 4320
rect 37946 4384 38262 4385
rect 37946 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38262 4384
rect 37946 4319 38262 4320
rect 47946 4384 48262 4385
rect 47946 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48262 4384
rect 47946 4319 48262 4320
rect 49141 4314 49207 4317
rect 50200 4314 51000 4344
rect 49141 4312 51000 4314
rect 49141 4256 49146 4312
rect 49202 4256 51000 4312
rect 49141 4254 51000 4256
rect 49141 4251 49207 4254
rect 50200 4224 51000 4254
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 2946 3840 3262 3841
rect 2946 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3262 3840
rect 2946 3775 3262 3776
rect 12946 3840 13262 3841
rect 12946 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13262 3840
rect 12946 3775 13262 3776
rect 22946 3840 23262 3841
rect 22946 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23262 3840
rect 22946 3775 23262 3776
rect 32946 3840 33262 3841
rect 32946 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33262 3840
rect 32946 3775 33262 3776
rect 42946 3840 43262 3841
rect 42946 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43262 3840
rect 42946 3775 43262 3776
rect 27102 3436 27108 3500
rect 27172 3498 27178 3500
rect 44909 3498 44975 3501
rect 27172 3496 44975 3498
rect 27172 3440 44914 3496
rect 44970 3440 44975 3496
rect 27172 3438 44975 3440
rect 27172 3436 27178 3438
rect 44909 3435 44975 3438
rect 7946 3296 8262 3297
rect 7946 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8262 3296
rect 7946 3231 8262 3232
rect 17946 3296 18262 3297
rect 17946 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18262 3296
rect 17946 3231 18262 3232
rect 27946 3296 28262 3297
rect 27946 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28262 3296
rect 27946 3231 28262 3232
rect 37946 3296 38262 3297
rect 37946 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38262 3296
rect 37946 3231 38262 3232
rect 47946 3296 48262 3297
rect 47946 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48262 3296
rect 47946 3231 48262 3232
rect 5717 2954 5783 2957
rect 22502 2954 22508 2956
rect 5717 2952 22508 2954
rect 5717 2896 5722 2952
rect 5778 2896 22508 2952
rect 5717 2894 22508 2896
rect 5717 2891 5783 2894
rect 22502 2892 22508 2894
rect 22572 2892 22578 2956
rect 2946 2752 3262 2753
rect 2946 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3262 2752
rect 2946 2687 3262 2688
rect 12946 2752 13262 2753
rect 12946 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13262 2752
rect 12946 2687 13262 2688
rect 22946 2752 23262 2753
rect 22946 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23262 2752
rect 22946 2687 23262 2688
rect 32946 2752 33262 2753
rect 32946 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33262 2752
rect 32946 2687 33262 2688
rect 42946 2752 43262 2753
rect 42946 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43262 2752
rect 42946 2687 43262 2688
rect 13629 2682 13695 2685
rect 22134 2682 22140 2684
rect 13629 2680 22140 2682
rect 13629 2624 13634 2680
rect 13690 2624 22140 2680
rect 13629 2622 22140 2624
rect 13629 2619 13695 2622
rect 22134 2620 22140 2622
rect 22204 2620 22210 2684
rect 9489 2546 9555 2549
rect 22686 2546 22692 2548
rect 9489 2544 22692 2546
rect 9489 2488 9494 2544
rect 9550 2488 22692 2544
rect 9489 2486 22692 2488
rect 9489 2483 9555 2486
rect 22686 2484 22692 2486
rect 22756 2484 22762 2548
rect 4981 2410 5047 2413
rect 21081 2410 21147 2413
rect 4981 2408 21147 2410
rect 4981 2352 4986 2408
rect 5042 2352 21086 2408
rect 21142 2352 21147 2408
rect 4981 2350 21147 2352
rect 4981 2347 5047 2350
rect 21081 2347 21147 2350
rect 7946 2208 8262 2209
rect 7946 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8262 2208
rect 7946 2143 8262 2144
rect 17946 2208 18262 2209
rect 17946 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18262 2208
rect 17946 2143 18262 2144
rect 27946 2208 28262 2209
rect 27946 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28262 2208
rect 27946 2143 28262 2144
rect 37946 2208 38262 2209
rect 37946 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38262 2208
rect 37946 2143 38262 2144
rect 47946 2208 48262 2209
rect 47946 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48262 2208
rect 47946 2143 48262 2144
rect 0 1866 800 1896
rect 2773 1866 2839 1869
rect 0 1864 2839 1866
rect 0 1808 2778 1864
rect 2834 1808 2839 1864
rect 0 1806 2839 1808
rect 0 1776 800 1806
rect 2773 1803 2839 1806
<< via3 >>
rect 7952 54428 8016 54432
rect 7952 54372 7956 54428
rect 7956 54372 8012 54428
rect 8012 54372 8016 54428
rect 7952 54368 8016 54372
rect 8032 54428 8096 54432
rect 8032 54372 8036 54428
rect 8036 54372 8092 54428
rect 8092 54372 8096 54428
rect 8032 54368 8096 54372
rect 8112 54428 8176 54432
rect 8112 54372 8116 54428
rect 8116 54372 8172 54428
rect 8172 54372 8176 54428
rect 8112 54368 8176 54372
rect 8192 54428 8256 54432
rect 8192 54372 8196 54428
rect 8196 54372 8252 54428
rect 8252 54372 8256 54428
rect 8192 54368 8256 54372
rect 17952 54428 18016 54432
rect 17952 54372 17956 54428
rect 17956 54372 18012 54428
rect 18012 54372 18016 54428
rect 17952 54368 18016 54372
rect 18032 54428 18096 54432
rect 18032 54372 18036 54428
rect 18036 54372 18092 54428
rect 18092 54372 18096 54428
rect 18032 54368 18096 54372
rect 18112 54428 18176 54432
rect 18112 54372 18116 54428
rect 18116 54372 18172 54428
rect 18172 54372 18176 54428
rect 18112 54368 18176 54372
rect 18192 54428 18256 54432
rect 18192 54372 18196 54428
rect 18196 54372 18252 54428
rect 18252 54372 18256 54428
rect 18192 54368 18256 54372
rect 27952 54428 28016 54432
rect 27952 54372 27956 54428
rect 27956 54372 28012 54428
rect 28012 54372 28016 54428
rect 27952 54368 28016 54372
rect 28032 54428 28096 54432
rect 28032 54372 28036 54428
rect 28036 54372 28092 54428
rect 28092 54372 28096 54428
rect 28032 54368 28096 54372
rect 28112 54428 28176 54432
rect 28112 54372 28116 54428
rect 28116 54372 28172 54428
rect 28172 54372 28176 54428
rect 28112 54368 28176 54372
rect 28192 54428 28256 54432
rect 28192 54372 28196 54428
rect 28196 54372 28252 54428
rect 28252 54372 28256 54428
rect 28192 54368 28256 54372
rect 37952 54428 38016 54432
rect 37952 54372 37956 54428
rect 37956 54372 38012 54428
rect 38012 54372 38016 54428
rect 37952 54368 38016 54372
rect 38032 54428 38096 54432
rect 38032 54372 38036 54428
rect 38036 54372 38092 54428
rect 38092 54372 38096 54428
rect 38032 54368 38096 54372
rect 38112 54428 38176 54432
rect 38112 54372 38116 54428
rect 38116 54372 38172 54428
rect 38172 54372 38176 54428
rect 38112 54368 38176 54372
rect 38192 54428 38256 54432
rect 38192 54372 38196 54428
rect 38196 54372 38252 54428
rect 38252 54372 38256 54428
rect 38192 54368 38256 54372
rect 47952 54428 48016 54432
rect 47952 54372 47956 54428
rect 47956 54372 48012 54428
rect 48012 54372 48016 54428
rect 47952 54368 48016 54372
rect 48032 54428 48096 54432
rect 48032 54372 48036 54428
rect 48036 54372 48092 54428
rect 48092 54372 48096 54428
rect 48032 54368 48096 54372
rect 48112 54428 48176 54432
rect 48112 54372 48116 54428
rect 48116 54372 48172 54428
rect 48172 54372 48176 54428
rect 48112 54368 48176 54372
rect 48192 54428 48256 54432
rect 48192 54372 48196 54428
rect 48196 54372 48252 54428
rect 48252 54372 48256 54428
rect 48192 54368 48256 54372
rect 25084 53892 25148 53956
rect 2952 53884 3016 53888
rect 2952 53828 2956 53884
rect 2956 53828 3012 53884
rect 3012 53828 3016 53884
rect 2952 53824 3016 53828
rect 3032 53884 3096 53888
rect 3032 53828 3036 53884
rect 3036 53828 3092 53884
rect 3092 53828 3096 53884
rect 3032 53824 3096 53828
rect 3112 53884 3176 53888
rect 3112 53828 3116 53884
rect 3116 53828 3172 53884
rect 3172 53828 3176 53884
rect 3112 53824 3176 53828
rect 3192 53884 3256 53888
rect 3192 53828 3196 53884
rect 3196 53828 3252 53884
rect 3252 53828 3256 53884
rect 3192 53824 3256 53828
rect 12952 53884 13016 53888
rect 12952 53828 12956 53884
rect 12956 53828 13012 53884
rect 13012 53828 13016 53884
rect 12952 53824 13016 53828
rect 13032 53884 13096 53888
rect 13032 53828 13036 53884
rect 13036 53828 13092 53884
rect 13092 53828 13096 53884
rect 13032 53824 13096 53828
rect 13112 53884 13176 53888
rect 13112 53828 13116 53884
rect 13116 53828 13172 53884
rect 13172 53828 13176 53884
rect 13112 53824 13176 53828
rect 13192 53884 13256 53888
rect 13192 53828 13196 53884
rect 13196 53828 13252 53884
rect 13252 53828 13256 53884
rect 13192 53824 13256 53828
rect 22952 53884 23016 53888
rect 22952 53828 22956 53884
rect 22956 53828 23012 53884
rect 23012 53828 23016 53884
rect 22952 53824 23016 53828
rect 23032 53884 23096 53888
rect 23032 53828 23036 53884
rect 23036 53828 23092 53884
rect 23092 53828 23096 53884
rect 23032 53824 23096 53828
rect 23112 53884 23176 53888
rect 23112 53828 23116 53884
rect 23116 53828 23172 53884
rect 23172 53828 23176 53884
rect 23112 53824 23176 53828
rect 23192 53884 23256 53888
rect 23192 53828 23196 53884
rect 23196 53828 23252 53884
rect 23252 53828 23256 53884
rect 23192 53824 23256 53828
rect 32952 53884 33016 53888
rect 32952 53828 32956 53884
rect 32956 53828 33012 53884
rect 33012 53828 33016 53884
rect 32952 53824 33016 53828
rect 33032 53884 33096 53888
rect 33032 53828 33036 53884
rect 33036 53828 33092 53884
rect 33092 53828 33096 53884
rect 33032 53824 33096 53828
rect 33112 53884 33176 53888
rect 33112 53828 33116 53884
rect 33116 53828 33172 53884
rect 33172 53828 33176 53884
rect 33112 53824 33176 53828
rect 33192 53884 33256 53888
rect 33192 53828 33196 53884
rect 33196 53828 33252 53884
rect 33252 53828 33256 53884
rect 33192 53824 33256 53828
rect 42952 53884 43016 53888
rect 42952 53828 42956 53884
rect 42956 53828 43012 53884
rect 43012 53828 43016 53884
rect 42952 53824 43016 53828
rect 43032 53884 43096 53888
rect 43032 53828 43036 53884
rect 43036 53828 43092 53884
rect 43092 53828 43096 53884
rect 43032 53824 43096 53828
rect 43112 53884 43176 53888
rect 43112 53828 43116 53884
rect 43116 53828 43172 53884
rect 43172 53828 43176 53884
rect 43112 53824 43176 53828
rect 43192 53884 43256 53888
rect 43192 53828 43196 53884
rect 43196 53828 43252 53884
rect 43252 53828 43256 53884
rect 43192 53824 43256 53828
rect 7952 53340 8016 53344
rect 7952 53284 7956 53340
rect 7956 53284 8012 53340
rect 8012 53284 8016 53340
rect 7952 53280 8016 53284
rect 8032 53340 8096 53344
rect 8032 53284 8036 53340
rect 8036 53284 8092 53340
rect 8092 53284 8096 53340
rect 8032 53280 8096 53284
rect 8112 53340 8176 53344
rect 8112 53284 8116 53340
rect 8116 53284 8172 53340
rect 8172 53284 8176 53340
rect 8112 53280 8176 53284
rect 8192 53340 8256 53344
rect 8192 53284 8196 53340
rect 8196 53284 8252 53340
rect 8252 53284 8256 53340
rect 8192 53280 8256 53284
rect 17952 53340 18016 53344
rect 17952 53284 17956 53340
rect 17956 53284 18012 53340
rect 18012 53284 18016 53340
rect 17952 53280 18016 53284
rect 18032 53340 18096 53344
rect 18032 53284 18036 53340
rect 18036 53284 18092 53340
rect 18092 53284 18096 53340
rect 18032 53280 18096 53284
rect 18112 53340 18176 53344
rect 18112 53284 18116 53340
rect 18116 53284 18172 53340
rect 18172 53284 18176 53340
rect 18112 53280 18176 53284
rect 18192 53340 18256 53344
rect 18192 53284 18196 53340
rect 18196 53284 18252 53340
rect 18252 53284 18256 53340
rect 18192 53280 18256 53284
rect 27952 53340 28016 53344
rect 27952 53284 27956 53340
rect 27956 53284 28012 53340
rect 28012 53284 28016 53340
rect 27952 53280 28016 53284
rect 28032 53340 28096 53344
rect 28032 53284 28036 53340
rect 28036 53284 28092 53340
rect 28092 53284 28096 53340
rect 28032 53280 28096 53284
rect 28112 53340 28176 53344
rect 28112 53284 28116 53340
rect 28116 53284 28172 53340
rect 28172 53284 28176 53340
rect 28112 53280 28176 53284
rect 28192 53340 28256 53344
rect 28192 53284 28196 53340
rect 28196 53284 28252 53340
rect 28252 53284 28256 53340
rect 28192 53280 28256 53284
rect 37952 53340 38016 53344
rect 37952 53284 37956 53340
rect 37956 53284 38012 53340
rect 38012 53284 38016 53340
rect 37952 53280 38016 53284
rect 38032 53340 38096 53344
rect 38032 53284 38036 53340
rect 38036 53284 38092 53340
rect 38092 53284 38096 53340
rect 38032 53280 38096 53284
rect 38112 53340 38176 53344
rect 38112 53284 38116 53340
rect 38116 53284 38172 53340
rect 38172 53284 38176 53340
rect 38112 53280 38176 53284
rect 38192 53340 38256 53344
rect 38192 53284 38196 53340
rect 38196 53284 38252 53340
rect 38252 53284 38256 53340
rect 38192 53280 38256 53284
rect 47952 53340 48016 53344
rect 47952 53284 47956 53340
rect 47956 53284 48012 53340
rect 48012 53284 48016 53340
rect 47952 53280 48016 53284
rect 48032 53340 48096 53344
rect 48032 53284 48036 53340
rect 48036 53284 48092 53340
rect 48092 53284 48096 53340
rect 48032 53280 48096 53284
rect 48112 53340 48176 53344
rect 48112 53284 48116 53340
rect 48116 53284 48172 53340
rect 48172 53284 48176 53340
rect 48112 53280 48176 53284
rect 48192 53340 48256 53344
rect 48192 53284 48196 53340
rect 48196 53284 48252 53340
rect 48252 53284 48256 53340
rect 48192 53280 48256 53284
rect 2952 52796 3016 52800
rect 2952 52740 2956 52796
rect 2956 52740 3012 52796
rect 3012 52740 3016 52796
rect 2952 52736 3016 52740
rect 3032 52796 3096 52800
rect 3032 52740 3036 52796
rect 3036 52740 3092 52796
rect 3092 52740 3096 52796
rect 3032 52736 3096 52740
rect 3112 52796 3176 52800
rect 3112 52740 3116 52796
rect 3116 52740 3172 52796
rect 3172 52740 3176 52796
rect 3112 52736 3176 52740
rect 3192 52796 3256 52800
rect 3192 52740 3196 52796
rect 3196 52740 3252 52796
rect 3252 52740 3256 52796
rect 3192 52736 3256 52740
rect 12952 52796 13016 52800
rect 12952 52740 12956 52796
rect 12956 52740 13012 52796
rect 13012 52740 13016 52796
rect 12952 52736 13016 52740
rect 13032 52796 13096 52800
rect 13032 52740 13036 52796
rect 13036 52740 13092 52796
rect 13092 52740 13096 52796
rect 13032 52736 13096 52740
rect 13112 52796 13176 52800
rect 13112 52740 13116 52796
rect 13116 52740 13172 52796
rect 13172 52740 13176 52796
rect 13112 52736 13176 52740
rect 13192 52796 13256 52800
rect 13192 52740 13196 52796
rect 13196 52740 13252 52796
rect 13252 52740 13256 52796
rect 13192 52736 13256 52740
rect 22952 52796 23016 52800
rect 22952 52740 22956 52796
rect 22956 52740 23012 52796
rect 23012 52740 23016 52796
rect 22952 52736 23016 52740
rect 23032 52796 23096 52800
rect 23032 52740 23036 52796
rect 23036 52740 23092 52796
rect 23092 52740 23096 52796
rect 23032 52736 23096 52740
rect 23112 52796 23176 52800
rect 23112 52740 23116 52796
rect 23116 52740 23172 52796
rect 23172 52740 23176 52796
rect 23112 52736 23176 52740
rect 23192 52796 23256 52800
rect 23192 52740 23196 52796
rect 23196 52740 23252 52796
rect 23252 52740 23256 52796
rect 23192 52736 23256 52740
rect 32952 52796 33016 52800
rect 32952 52740 32956 52796
rect 32956 52740 33012 52796
rect 33012 52740 33016 52796
rect 32952 52736 33016 52740
rect 33032 52796 33096 52800
rect 33032 52740 33036 52796
rect 33036 52740 33092 52796
rect 33092 52740 33096 52796
rect 33032 52736 33096 52740
rect 33112 52796 33176 52800
rect 33112 52740 33116 52796
rect 33116 52740 33172 52796
rect 33172 52740 33176 52796
rect 33112 52736 33176 52740
rect 33192 52796 33256 52800
rect 33192 52740 33196 52796
rect 33196 52740 33252 52796
rect 33252 52740 33256 52796
rect 33192 52736 33256 52740
rect 42952 52796 43016 52800
rect 42952 52740 42956 52796
rect 42956 52740 43012 52796
rect 43012 52740 43016 52796
rect 42952 52736 43016 52740
rect 43032 52796 43096 52800
rect 43032 52740 43036 52796
rect 43036 52740 43092 52796
rect 43092 52740 43096 52796
rect 43032 52736 43096 52740
rect 43112 52796 43176 52800
rect 43112 52740 43116 52796
rect 43116 52740 43172 52796
rect 43172 52740 43176 52796
rect 43112 52736 43176 52740
rect 43192 52796 43256 52800
rect 43192 52740 43196 52796
rect 43196 52740 43252 52796
rect 43252 52740 43256 52796
rect 43192 52736 43256 52740
rect 7952 52252 8016 52256
rect 7952 52196 7956 52252
rect 7956 52196 8012 52252
rect 8012 52196 8016 52252
rect 7952 52192 8016 52196
rect 8032 52252 8096 52256
rect 8032 52196 8036 52252
rect 8036 52196 8092 52252
rect 8092 52196 8096 52252
rect 8032 52192 8096 52196
rect 8112 52252 8176 52256
rect 8112 52196 8116 52252
rect 8116 52196 8172 52252
rect 8172 52196 8176 52252
rect 8112 52192 8176 52196
rect 8192 52252 8256 52256
rect 8192 52196 8196 52252
rect 8196 52196 8252 52252
rect 8252 52196 8256 52252
rect 8192 52192 8256 52196
rect 17952 52252 18016 52256
rect 17952 52196 17956 52252
rect 17956 52196 18012 52252
rect 18012 52196 18016 52252
rect 17952 52192 18016 52196
rect 18032 52252 18096 52256
rect 18032 52196 18036 52252
rect 18036 52196 18092 52252
rect 18092 52196 18096 52252
rect 18032 52192 18096 52196
rect 18112 52252 18176 52256
rect 18112 52196 18116 52252
rect 18116 52196 18172 52252
rect 18172 52196 18176 52252
rect 18112 52192 18176 52196
rect 18192 52252 18256 52256
rect 18192 52196 18196 52252
rect 18196 52196 18252 52252
rect 18252 52196 18256 52252
rect 18192 52192 18256 52196
rect 27952 52252 28016 52256
rect 27952 52196 27956 52252
rect 27956 52196 28012 52252
rect 28012 52196 28016 52252
rect 27952 52192 28016 52196
rect 28032 52252 28096 52256
rect 28032 52196 28036 52252
rect 28036 52196 28092 52252
rect 28092 52196 28096 52252
rect 28032 52192 28096 52196
rect 28112 52252 28176 52256
rect 28112 52196 28116 52252
rect 28116 52196 28172 52252
rect 28172 52196 28176 52252
rect 28112 52192 28176 52196
rect 28192 52252 28256 52256
rect 28192 52196 28196 52252
rect 28196 52196 28252 52252
rect 28252 52196 28256 52252
rect 28192 52192 28256 52196
rect 37952 52252 38016 52256
rect 37952 52196 37956 52252
rect 37956 52196 38012 52252
rect 38012 52196 38016 52252
rect 37952 52192 38016 52196
rect 38032 52252 38096 52256
rect 38032 52196 38036 52252
rect 38036 52196 38092 52252
rect 38092 52196 38096 52252
rect 38032 52192 38096 52196
rect 38112 52252 38176 52256
rect 38112 52196 38116 52252
rect 38116 52196 38172 52252
rect 38172 52196 38176 52252
rect 38112 52192 38176 52196
rect 38192 52252 38256 52256
rect 38192 52196 38196 52252
rect 38196 52196 38252 52252
rect 38252 52196 38256 52252
rect 38192 52192 38256 52196
rect 47952 52252 48016 52256
rect 47952 52196 47956 52252
rect 47956 52196 48012 52252
rect 48012 52196 48016 52252
rect 47952 52192 48016 52196
rect 48032 52252 48096 52256
rect 48032 52196 48036 52252
rect 48036 52196 48092 52252
rect 48092 52196 48096 52252
rect 48032 52192 48096 52196
rect 48112 52252 48176 52256
rect 48112 52196 48116 52252
rect 48116 52196 48172 52252
rect 48172 52196 48176 52252
rect 48112 52192 48176 52196
rect 48192 52252 48256 52256
rect 48192 52196 48196 52252
rect 48196 52196 48252 52252
rect 48252 52196 48256 52252
rect 48192 52192 48256 52196
rect 2952 51708 3016 51712
rect 2952 51652 2956 51708
rect 2956 51652 3012 51708
rect 3012 51652 3016 51708
rect 2952 51648 3016 51652
rect 3032 51708 3096 51712
rect 3032 51652 3036 51708
rect 3036 51652 3092 51708
rect 3092 51652 3096 51708
rect 3032 51648 3096 51652
rect 3112 51708 3176 51712
rect 3112 51652 3116 51708
rect 3116 51652 3172 51708
rect 3172 51652 3176 51708
rect 3112 51648 3176 51652
rect 3192 51708 3256 51712
rect 3192 51652 3196 51708
rect 3196 51652 3252 51708
rect 3252 51652 3256 51708
rect 3192 51648 3256 51652
rect 12952 51708 13016 51712
rect 12952 51652 12956 51708
rect 12956 51652 13012 51708
rect 13012 51652 13016 51708
rect 12952 51648 13016 51652
rect 13032 51708 13096 51712
rect 13032 51652 13036 51708
rect 13036 51652 13092 51708
rect 13092 51652 13096 51708
rect 13032 51648 13096 51652
rect 13112 51708 13176 51712
rect 13112 51652 13116 51708
rect 13116 51652 13172 51708
rect 13172 51652 13176 51708
rect 13112 51648 13176 51652
rect 13192 51708 13256 51712
rect 13192 51652 13196 51708
rect 13196 51652 13252 51708
rect 13252 51652 13256 51708
rect 13192 51648 13256 51652
rect 22952 51708 23016 51712
rect 22952 51652 22956 51708
rect 22956 51652 23012 51708
rect 23012 51652 23016 51708
rect 22952 51648 23016 51652
rect 23032 51708 23096 51712
rect 23032 51652 23036 51708
rect 23036 51652 23092 51708
rect 23092 51652 23096 51708
rect 23032 51648 23096 51652
rect 23112 51708 23176 51712
rect 23112 51652 23116 51708
rect 23116 51652 23172 51708
rect 23172 51652 23176 51708
rect 23112 51648 23176 51652
rect 23192 51708 23256 51712
rect 23192 51652 23196 51708
rect 23196 51652 23252 51708
rect 23252 51652 23256 51708
rect 23192 51648 23256 51652
rect 32952 51708 33016 51712
rect 32952 51652 32956 51708
rect 32956 51652 33012 51708
rect 33012 51652 33016 51708
rect 32952 51648 33016 51652
rect 33032 51708 33096 51712
rect 33032 51652 33036 51708
rect 33036 51652 33092 51708
rect 33092 51652 33096 51708
rect 33032 51648 33096 51652
rect 33112 51708 33176 51712
rect 33112 51652 33116 51708
rect 33116 51652 33172 51708
rect 33172 51652 33176 51708
rect 33112 51648 33176 51652
rect 33192 51708 33256 51712
rect 33192 51652 33196 51708
rect 33196 51652 33252 51708
rect 33252 51652 33256 51708
rect 33192 51648 33256 51652
rect 42952 51708 43016 51712
rect 42952 51652 42956 51708
rect 42956 51652 43012 51708
rect 43012 51652 43016 51708
rect 42952 51648 43016 51652
rect 43032 51708 43096 51712
rect 43032 51652 43036 51708
rect 43036 51652 43092 51708
rect 43092 51652 43096 51708
rect 43032 51648 43096 51652
rect 43112 51708 43176 51712
rect 43112 51652 43116 51708
rect 43116 51652 43172 51708
rect 43172 51652 43176 51708
rect 43112 51648 43176 51652
rect 43192 51708 43256 51712
rect 43192 51652 43196 51708
rect 43196 51652 43252 51708
rect 43252 51652 43256 51708
rect 43192 51648 43256 51652
rect 7952 51164 8016 51168
rect 7952 51108 7956 51164
rect 7956 51108 8012 51164
rect 8012 51108 8016 51164
rect 7952 51104 8016 51108
rect 8032 51164 8096 51168
rect 8032 51108 8036 51164
rect 8036 51108 8092 51164
rect 8092 51108 8096 51164
rect 8032 51104 8096 51108
rect 8112 51164 8176 51168
rect 8112 51108 8116 51164
rect 8116 51108 8172 51164
rect 8172 51108 8176 51164
rect 8112 51104 8176 51108
rect 8192 51164 8256 51168
rect 8192 51108 8196 51164
rect 8196 51108 8252 51164
rect 8252 51108 8256 51164
rect 8192 51104 8256 51108
rect 17952 51164 18016 51168
rect 17952 51108 17956 51164
rect 17956 51108 18012 51164
rect 18012 51108 18016 51164
rect 17952 51104 18016 51108
rect 18032 51164 18096 51168
rect 18032 51108 18036 51164
rect 18036 51108 18092 51164
rect 18092 51108 18096 51164
rect 18032 51104 18096 51108
rect 18112 51164 18176 51168
rect 18112 51108 18116 51164
rect 18116 51108 18172 51164
rect 18172 51108 18176 51164
rect 18112 51104 18176 51108
rect 18192 51164 18256 51168
rect 18192 51108 18196 51164
rect 18196 51108 18252 51164
rect 18252 51108 18256 51164
rect 18192 51104 18256 51108
rect 27952 51164 28016 51168
rect 27952 51108 27956 51164
rect 27956 51108 28012 51164
rect 28012 51108 28016 51164
rect 27952 51104 28016 51108
rect 28032 51164 28096 51168
rect 28032 51108 28036 51164
rect 28036 51108 28092 51164
rect 28092 51108 28096 51164
rect 28032 51104 28096 51108
rect 28112 51164 28176 51168
rect 28112 51108 28116 51164
rect 28116 51108 28172 51164
rect 28172 51108 28176 51164
rect 28112 51104 28176 51108
rect 28192 51164 28256 51168
rect 28192 51108 28196 51164
rect 28196 51108 28252 51164
rect 28252 51108 28256 51164
rect 28192 51104 28256 51108
rect 37952 51164 38016 51168
rect 37952 51108 37956 51164
rect 37956 51108 38012 51164
rect 38012 51108 38016 51164
rect 37952 51104 38016 51108
rect 38032 51164 38096 51168
rect 38032 51108 38036 51164
rect 38036 51108 38092 51164
rect 38092 51108 38096 51164
rect 38032 51104 38096 51108
rect 38112 51164 38176 51168
rect 38112 51108 38116 51164
rect 38116 51108 38172 51164
rect 38172 51108 38176 51164
rect 38112 51104 38176 51108
rect 38192 51164 38256 51168
rect 38192 51108 38196 51164
rect 38196 51108 38252 51164
rect 38252 51108 38256 51164
rect 38192 51104 38256 51108
rect 47952 51164 48016 51168
rect 47952 51108 47956 51164
rect 47956 51108 48012 51164
rect 48012 51108 48016 51164
rect 47952 51104 48016 51108
rect 48032 51164 48096 51168
rect 48032 51108 48036 51164
rect 48036 51108 48092 51164
rect 48092 51108 48096 51164
rect 48032 51104 48096 51108
rect 48112 51164 48176 51168
rect 48112 51108 48116 51164
rect 48116 51108 48172 51164
rect 48172 51108 48176 51164
rect 48112 51104 48176 51108
rect 48192 51164 48256 51168
rect 48192 51108 48196 51164
rect 48196 51108 48252 51164
rect 48252 51108 48256 51164
rect 48192 51104 48256 51108
rect 2952 50620 3016 50624
rect 2952 50564 2956 50620
rect 2956 50564 3012 50620
rect 3012 50564 3016 50620
rect 2952 50560 3016 50564
rect 3032 50620 3096 50624
rect 3032 50564 3036 50620
rect 3036 50564 3092 50620
rect 3092 50564 3096 50620
rect 3032 50560 3096 50564
rect 3112 50620 3176 50624
rect 3112 50564 3116 50620
rect 3116 50564 3172 50620
rect 3172 50564 3176 50620
rect 3112 50560 3176 50564
rect 3192 50620 3256 50624
rect 3192 50564 3196 50620
rect 3196 50564 3252 50620
rect 3252 50564 3256 50620
rect 3192 50560 3256 50564
rect 12952 50620 13016 50624
rect 12952 50564 12956 50620
rect 12956 50564 13012 50620
rect 13012 50564 13016 50620
rect 12952 50560 13016 50564
rect 13032 50620 13096 50624
rect 13032 50564 13036 50620
rect 13036 50564 13092 50620
rect 13092 50564 13096 50620
rect 13032 50560 13096 50564
rect 13112 50620 13176 50624
rect 13112 50564 13116 50620
rect 13116 50564 13172 50620
rect 13172 50564 13176 50620
rect 13112 50560 13176 50564
rect 13192 50620 13256 50624
rect 13192 50564 13196 50620
rect 13196 50564 13252 50620
rect 13252 50564 13256 50620
rect 13192 50560 13256 50564
rect 22952 50620 23016 50624
rect 22952 50564 22956 50620
rect 22956 50564 23012 50620
rect 23012 50564 23016 50620
rect 22952 50560 23016 50564
rect 23032 50620 23096 50624
rect 23032 50564 23036 50620
rect 23036 50564 23092 50620
rect 23092 50564 23096 50620
rect 23032 50560 23096 50564
rect 23112 50620 23176 50624
rect 23112 50564 23116 50620
rect 23116 50564 23172 50620
rect 23172 50564 23176 50620
rect 23112 50560 23176 50564
rect 23192 50620 23256 50624
rect 23192 50564 23196 50620
rect 23196 50564 23252 50620
rect 23252 50564 23256 50620
rect 23192 50560 23256 50564
rect 32952 50620 33016 50624
rect 32952 50564 32956 50620
rect 32956 50564 33012 50620
rect 33012 50564 33016 50620
rect 32952 50560 33016 50564
rect 33032 50620 33096 50624
rect 33032 50564 33036 50620
rect 33036 50564 33092 50620
rect 33092 50564 33096 50620
rect 33032 50560 33096 50564
rect 33112 50620 33176 50624
rect 33112 50564 33116 50620
rect 33116 50564 33172 50620
rect 33172 50564 33176 50620
rect 33112 50560 33176 50564
rect 33192 50620 33256 50624
rect 33192 50564 33196 50620
rect 33196 50564 33252 50620
rect 33252 50564 33256 50620
rect 33192 50560 33256 50564
rect 42952 50620 43016 50624
rect 42952 50564 42956 50620
rect 42956 50564 43012 50620
rect 43012 50564 43016 50620
rect 42952 50560 43016 50564
rect 43032 50620 43096 50624
rect 43032 50564 43036 50620
rect 43036 50564 43092 50620
rect 43092 50564 43096 50620
rect 43032 50560 43096 50564
rect 43112 50620 43176 50624
rect 43112 50564 43116 50620
rect 43116 50564 43172 50620
rect 43172 50564 43176 50620
rect 43112 50560 43176 50564
rect 43192 50620 43256 50624
rect 43192 50564 43196 50620
rect 43196 50564 43252 50620
rect 43252 50564 43256 50620
rect 43192 50560 43256 50564
rect 7952 50076 8016 50080
rect 7952 50020 7956 50076
rect 7956 50020 8012 50076
rect 8012 50020 8016 50076
rect 7952 50016 8016 50020
rect 8032 50076 8096 50080
rect 8032 50020 8036 50076
rect 8036 50020 8092 50076
rect 8092 50020 8096 50076
rect 8032 50016 8096 50020
rect 8112 50076 8176 50080
rect 8112 50020 8116 50076
rect 8116 50020 8172 50076
rect 8172 50020 8176 50076
rect 8112 50016 8176 50020
rect 8192 50076 8256 50080
rect 8192 50020 8196 50076
rect 8196 50020 8252 50076
rect 8252 50020 8256 50076
rect 8192 50016 8256 50020
rect 17952 50076 18016 50080
rect 17952 50020 17956 50076
rect 17956 50020 18012 50076
rect 18012 50020 18016 50076
rect 17952 50016 18016 50020
rect 18032 50076 18096 50080
rect 18032 50020 18036 50076
rect 18036 50020 18092 50076
rect 18092 50020 18096 50076
rect 18032 50016 18096 50020
rect 18112 50076 18176 50080
rect 18112 50020 18116 50076
rect 18116 50020 18172 50076
rect 18172 50020 18176 50076
rect 18112 50016 18176 50020
rect 18192 50076 18256 50080
rect 18192 50020 18196 50076
rect 18196 50020 18252 50076
rect 18252 50020 18256 50076
rect 18192 50016 18256 50020
rect 27952 50076 28016 50080
rect 27952 50020 27956 50076
rect 27956 50020 28012 50076
rect 28012 50020 28016 50076
rect 27952 50016 28016 50020
rect 28032 50076 28096 50080
rect 28032 50020 28036 50076
rect 28036 50020 28092 50076
rect 28092 50020 28096 50076
rect 28032 50016 28096 50020
rect 28112 50076 28176 50080
rect 28112 50020 28116 50076
rect 28116 50020 28172 50076
rect 28172 50020 28176 50076
rect 28112 50016 28176 50020
rect 28192 50076 28256 50080
rect 28192 50020 28196 50076
rect 28196 50020 28252 50076
rect 28252 50020 28256 50076
rect 28192 50016 28256 50020
rect 37952 50076 38016 50080
rect 37952 50020 37956 50076
rect 37956 50020 38012 50076
rect 38012 50020 38016 50076
rect 37952 50016 38016 50020
rect 38032 50076 38096 50080
rect 38032 50020 38036 50076
rect 38036 50020 38092 50076
rect 38092 50020 38096 50076
rect 38032 50016 38096 50020
rect 38112 50076 38176 50080
rect 38112 50020 38116 50076
rect 38116 50020 38172 50076
rect 38172 50020 38176 50076
rect 38112 50016 38176 50020
rect 38192 50076 38256 50080
rect 38192 50020 38196 50076
rect 38196 50020 38252 50076
rect 38252 50020 38256 50076
rect 38192 50016 38256 50020
rect 47952 50076 48016 50080
rect 47952 50020 47956 50076
rect 47956 50020 48012 50076
rect 48012 50020 48016 50076
rect 47952 50016 48016 50020
rect 48032 50076 48096 50080
rect 48032 50020 48036 50076
rect 48036 50020 48092 50076
rect 48092 50020 48096 50076
rect 48032 50016 48096 50020
rect 48112 50076 48176 50080
rect 48112 50020 48116 50076
rect 48116 50020 48172 50076
rect 48172 50020 48176 50076
rect 48112 50016 48176 50020
rect 48192 50076 48256 50080
rect 48192 50020 48196 50076
rect 48196 50020 48252 50076
rect 48252 50020 48256 50076
rect 48192 50016 48256 50020
rect 2952 49532 3016 49536
rect 2952 49476 2956 49532
rect 2956 49476 3012 49532
rect 3012 49476 3016 49532
rect 2952 49472 3016 49476
rect 3032 49532 3096 49536
rect 3032 49476 3036 49532
rect 3036 49476 3092 49532
rect 3092 49476 3096 49532
rect 3032 49472 3096 49476
rect 3112 49532 3176 49536
rect 3112 49476 3116 49532
rect 3116 49476 3172 49532
rect 3172 49476 3176 49532
rect 3112 49472 3176 49476
rect 3192 49532 3256 49536
rect 3192 49476 3196 49532
rect 3196 49476 3252 49532
rect 3252 49476 3256 49532
rect 3192 49472 3256 49476
rect 12952 49532 13016 49536
rect 12952 49476 12956 49532
rect 12956 49476 13012 49532
rect 13012 49476 13016 49532
rect 12952 49472 13016 49476
rect 13032 49532 13096 49536
rect 13032 49476 13036 49532
rect 13036 49476 13092 49532
rect 13092 49476 13096 49532
rect 13032 49472 13096 49476
rect 13112 49532 13176 49536
rect 13112 49476 13116 49532
rect 13116 49476 13172 49532
rect 13172 49476 13176 49532
rect 13112 49472 13176 49476
rect 13192 49532 13256 49536
rect 13192 49476 13196 49532
rect 13196 49476 13252 49532
rect 13252 49476 13256 49532
rect 13192 49472 13256 49476
rect 22952 49532 23016 49536
rect 22952 49476 22956 49532
rect 22956 49476 23012 49532
rect 23012 49476 23016 49532
rect 22952 49472 23016 49476
rect 23032 49532 23096 49536
rect 23032 49476 23036 49532
rect 23036 49476 23092 49532
rect 23092 49476 23096 49532
rect 23032 49472 23096 49476
rect 23112 49532 23176 49536
rect 23112 49476 23116 49532
rect 23116 49476 23172 49532
rect 23172 49476 23176 49532
rect 23112 49472 23176 49476
rect 23192 49532 23256 49536
rect 23192 49476 23196 49532
rect 23196 49476 23252 49532
rect 23252 49476 23256 49532
rect 23192 49472 23256 49476
rect 32952 49532 33016 49536
rect 32952 49476 32956 49532
rect 32956 49476 33012 49532
rect 33012 49476 33016 49532
rect 32952 49472 33016 49476
rect 33032 49532 33096 49536
rect 33032 49476 33036 49532
rect 33036 49476 33092 49532
rect 33092 49476 33096 49532
rect 33032 49472 33096 49476
rect 33112 49532 33176 49536
rect 33112 49476 33116 49532
rect 33116 49476 33172 49532
rect 33172 49476 33176 49532
rect 33112 49472 33176 49476
rect 33192 49532 33256 49536
rect 33192 49476 33196 49532
rect 33196 49476 33252 49532
rect 33252 49476 33256 49532
rect 33192 49472 33256 49476
rect 42952 49532 43016 49536
rect 42952 49476 42956 49532
rect 42956 49476 43012 49532
rect 43012 49476 43016 49532
rect 42952 49472 43016 49476
rect 43032 49532 43096 49536
rect 43032 49476 43036 49532
rect 43036 49476 43092 49532
rect 43092 49476 43096 49532
rect 43032 49472 43096 49476
rect 43112 49532 43176 49536
rect 43112 49476 43116 49532
rect 43116 49476 43172 49532
rect 43172 49476 43176 49532
rect 43112 49472 43176 49476
rect 43192 49532 43256 49536
rect 43192 49476 43196 49532
rect 43196 49476 43252 49532
rect 43252 49476 43256 49532
rect 43192 49472 43256 49476
rect 7952 48988 8016 48992
rect 7952 48932 7956 48988
rect 7956 48932 8012 48988
rect 8012 48932 8016 48988
rect 7952 48928 8016 48932
rect 8032 48988 8096 48992
rect 8032 48932 8036 48988
rect 8036 48932 8092 48988
rect 8092 48932 8096 48988
rect 8032 48928 8096 48932
rect 8112 48988 8176 48992
rect 8112 48932 8116 48988
rect 8116 48932 8172 48988
rect 8172 48932 8176 48988
rect 8112 48928 8176 48932
rect 8192 48988 8256 48992
rect 8192 48932 8196 48988
rect 8196 48932 8252 48988
rect 8252 48932 8256 48988
rect 8192 48928 8256 48932
rect 17952 48988 18016 48992
rect 17952 48932 17956 48988
rect 17956 48932 18012 48988
rect 18012 48932 18016 48988
rect 17952 48928 18016 48932
rect 18032 48988 18096 48992
rect 18032 48932 18036 48988
rect 18036 48932 18092 48988
rect 18092 48932 18096 48988
rect 18032 48928 18096 48932
rect 18112 48988 18176 48992
rect 18112 48932 18116 48988
rect 18116 48932 18172 48988
rect 18172 48932 18176 48988
rect 18112 48928 18176 48932
rect 18192 48988 18256 48992
rect 18192 48932 18196 48988
rect 18196 48932 18252 48988
rect 18252 48932 18256 48988
rect 18192 48928 18256 48932
rect 27952 48988 28016 48992
rect 27952 48932 27956 48988
rect 27956 48932 28012 48988
rect 28012 48932 28016 48988
rect 27952 48928 28016 48932
rect 28032 48988 28096 48992
rect 28032 48932 28036 48988
rect 28036 48932 28092 48988
rect 28092 48932 28096 48988
rect 28032 48928 28096 48932
rect 28112 48988 28176 48992
rect 28112 48932 28116 48988
rect 28116 48932 28172 48988
rect 28172 48932 28176 48988
rect 28112 48928 28176 48932
rect 28192 48988 28256 48992
rect 28192 48932 28196 48988
rect 28196 48932 28252 48988
rect 28252 48932 28256 48988
rect 28192 48928 28256 48932
rect 37952 48988 38016 48992
rect 37952 48932 37956 48988
rect 37956 48932 38012 48988
rect 38012 48932 38016 48988
rect 37952 48928 38016 48932
rect 38032 48988 38096 48992
rect 38032 48932 38036 48988
rect 38036 48932 38092 48988
rect 38092 48932 38096 48988
rect 38032 48928 38096 48932
rect 38112 48988 38176 48992
rect 38112 48932 38116 48988
rect 38116 48932 38172 48988
rect 38172 48932 38176 48988
rect 38112 48928 38176 48932
rect 38192 48988 38256 48992
rect 38192 48932 38196 48988
rect 38196 48932 38252 48988
rect 38252 48932 38256 48988
rect 38192 48928 38256 48932
rect 47952 48988 48016 48992
rect 47952 48932 47956 48988
rect 47956 48932 48012 48988
rect 48012 48932 48016 48988
rect 47952 48928 48016 48932
rect 48032 48988 48096 48992
rect 48032 48932 48036 48988
rect 48036 48932 48092 48988
rect 48092 48932 48096 48988
rect 48032 48928 48096 48932
rect 48112 48988 48176 48992
rect 48112 48932 48116 48988
rect 48116 48932 48172 48988
rect 48172 48932 48176 48988
rect 48112 48928 48176 48932
rect 48192 48988 48256 48992
rect 48192 48932 48196 48988
rect 48196 48932 48252 48988
rect 48252 48932 48256 48988
rect 48192 48928 48256 48932
rect 2952 48444 3016 48448
rect 2952 48388 2956 48444
rect 2956 48388 3012 48444
rect 3012 48388 3016 48444
rect 2952 48384 3016 48388
rect 3032 48444 3096 48448
rect 3032 48388 3036 48444
rect 3036 48388 3092 48444
rect 3092 48388 3096 48444
rect 3032 48384 3096 48388
rect 3112 48444 3176 48448
rect 3112 48388 3116 48444
rect 3116 48388 3172 48444
rect 3172 48388 3176 48444
rect 3112 48384 3176 48388
rect 3192 48444 3256 48448
rect 3192 48388 3196 48444
rect 3196 48388 3252 48444
rect 3252 48388 3256 48444
rect 3192 48384 3256 48388
rect 12952 48444 13016 48448
rect 12952 48388 12956 48444
rect 12956 48388 13012 48444
rect 13012 48388 13016 48444
rect 12952 48384 13016 48388
rect 13032 48444 13096 48448
rect 13032 48388 13036 48444
rect 13036 48388 13092 48444
rect 13092 48388 13096 48444
rect 13032 48384 13096 48388
rect 13112 48444 13176 48448
rect 13112 48388 13116 48444
rect 13116 48388 13172 48444
rect 13172 48388 13176 48444
rect 13112 48384 13176 48388
rect 13192 48444 13256 48448
rect 13192 48388 13196 48444
rect 13196 48388 13252 48444
rect 13252 48388 13256 48444
rect 13192 48384 13256 48388
rect 22952 48444 23016 48448
rect 22952 48388 22956 48444
rect 22956 48388 23012 48444
rect 23012 48388 23016 48444
rect 22952 48384 23016 48388
rect 23032 48444 23096 48448
rect 23032 48388 23036 48444
rect 23036 48388 23092 48444
rect 23092 48388 23096 48444
rect 23032 48384 23096 48388
rect 23112 48444 23176 48448
rect 23112 48388 23116 48444
rect 23116 48388 23172 48444
rect 23172 48388 23176 48444
rect 23112 48384 23176 48388
rect 23192 48444 23256 48448
rect 23192 48388 23196 48444
rect 23196 48388 23252 48444
rect 23252 48388 23256 48444
rect 23192 48384 23256 48388
rect 32952 48444 33016 48448
rect 32952 48388 32956 48444
rect 32956 48388 33012 48444
rect 33012 48388 33016 48444
rect 32952 48384 33016 48388
rect 33032 48444 33096 48448
rect 33032 48388 33036 48444
rect 33036 48388 33092 48444
rect 33092 48388 33096 48444
rect 33032 48384 33096 48388
rect 33112 48444 33176 48448
rect 33112 48388 33116 48444
rect 33116 48388 33172 48444
rect 33172 48388 33176 48444
rect 33112 48384 33176 48388
rect 33192 48444 33256 48448
rect 33192 48388 33196 48444
rect 33196 48388 33252 48444
rect 33252 48388 33256 48444
rect 33192 48384 33256 48388
rect 42952 48444 43016 48448
rect 42952 48388 42956 48444
rect 42956 48388 43012 48444
rect 43012 48388 43016 48444
rect 42952 48384 43016 48388
rect 43032 48444 43096 48448
rect 43032 48388 43036 48444
rect 43036 48388 43092 48444
rect 43092 48388 43096 48444
rect 43032 48384 43096 48388
rect 43112 48444 43176 48448
rect 43112 48388 43116 48444
rect 43116 48388 43172 48444
rect 43172 48388 43176 48444
rect 43112 48384 43176 48388
rect 43192 48444 43256 48448
rect 43192 48388 43196 48444
rect 43196 48388 43252 48444
rect 43252 48388 43256 48444
rect 43192 48384 43256 48388
rect 7952 47900 8016 47904
rect 7952 47844 7956 47900
rect 7956 47844 8012 47900
rect 8012 47844 8016 47900
rect 7952 47840 8016 47844
rect 8032 47900 8096 47904
rect 8032 47844 8036 47900
rect 8036 47844 8092 47900
rect 8092 47844 8096 47900
rect 8032 47840 8096 47844
rect 8112 47900 8176 47904
rect 8112 47844 8116 47900
rect 8116 47844 8172 47900
rect 8172 47844 8176 47900
rect 8112 47840 8176 47844
rect 8192 47900 8256 47904
rect 8192 47844 8196 47900
rect 8196 47844 8252 47900
rect 8252 47844 8256 47900
rect 8192 47840 8256 47844
rect 17952 47900 18016 47904
rect 17952 47844 17956 47900
rect 17956 47844 18012 47900
rect 18012 47844 18016 47900
rect 17952 47840 18016 47844
rect 18032 47900 18096 47904
rect 18032 47844 18036 47900
rect 18036 47844 18092 47900
rect 18092 47844 18096 47900
rect 18032 47840 18096 47844
rect 18112 47900 18176 47904
rect 18112 47844 18116 47900
rect 18116 47844 18172 47900
rect 18172 47844 18176 47900
rect 18112 47840 18176 47844
rect 18192 47900 18256 47904
rect 18192 47844 18196 47900
rect 18196 47844 18252 47900
rect 18252 47844 18256 47900
rect 18192 47840 18256 47844
rect 27952 47900 28016 47904
rect 27952 47844 27956 47900
rect 27956 47844 28012 47900
rect 28012 47844 28016 47900
rect 27952 47840 28016 47844
rect 28032 47900 28096 47904
rect 28032 47844 28036 47900
rect 28036 47844 28092 47900
rect 28092 47844 28096 47900
rect 28032 47840 28096 47844
rect 28112 47900 28176 47904
rect 28112 47844 28116 47900
rect 28116 47844 28172 47900
rect 28172 47844 28176 47900
rect 28112 47840 28176 47844
rect 28192 47900 28256 47904
rect 28192 47844 28196 47900
rect 28196 47844 28252 47900
rect 28252 47844 28256 47900
rect 28192 47840 28256 47844
rect 37952 47900 38016 47904
rect 37952 47844 37956 47900
rect 37956 47844 38012 47900
rect 38012 47844 38016 47900
rect 37952 47840 38016 47844
rect 38032 47900 38096 47904
rect 38032 47844 38036 47900
rect 38036 47844 38092 47900
rect 38092 47844 38096 47900
rect 38032 47840 38096 47844
rect 38112 47900 38176 47904
rect 38112 47844 38116 47900
rect 38116 47844 38172 47900
rect 38172 47844 38176 47900
rect 38112 47840 38176 47844
rect 38192 47900 38256 47904
rect 38192 47844 38196 47900
rect 38196 47844 38252 47900
rect 38252 47844 38256 47900
rect 38192 47840 38256 47844
rect 47952 47900 48016 47904
rect 47952 47844 47956 47900
rect 47956 47844 48012 47900
rect 48012 47844 48016 47900
rect 47952 47840 48016 47844
rect 48032 47900 48096 47904
rect 48032 47844 48036 47900
rect 48036 47844 48092 47900
rect 48092 47844 48096 47900
rect 48032 47840 48096 47844
rect 48112 47900 48176 47904
rect 48112 47844 48116 47900
rect 48116 47844 48172 47900
rect 48172 47844 48176 47900
rect 48112 47840 48176 47844
rect 48192 47900 48256 47904
rect 48192 47844 48196 47900
rect 48196 47844 48252 47900
rect 48252 47844 48256 47900
rect 48192 47840 48256 47844
rect 2952 47356 3016 47360
rect 2952 47300 2956 47356
rect 2956 47300 3012 47356
rect 3012 47300 3016 47356
rect 2952 47296 3016 47300
rect 3032 47356 3096 47360
rect 3032 47300 3036 47356
rect 3036 47300 3092 47356
rect 3092 47300 3096 47356
rect 3032 47296 3096 47300
rect 3112 47356 3176 47360
rect 3112 47300 3116 47356
rect 3116 47300 3172 47356
rect 3172 47300 3176 47356
rect 3112 47296 3176 47300
rect 3192 47356 3256 47360
rect 3192 47300 3196 47356
rect 3196 47300 3252 47356
rect 3252 47300 3256 47356
rect 3192 47296 3256 47300
rect 12952 47356 13016 47360
rect 12952 47300 12956 47356
rect 12956 47300 13012 47356
rect 13012 47300 13016 47356
rect 12952 47296 13016 47300
rect 13032 47356 13096 47360
rect 13032 47300 13036 47356
rect 13036 47300 13092 47356
rect 13092 47300 13096 47356
rect 13032 47296 13096 47300
rect 13112 47356 13176 47360
rect 13112 47300 13116 47356
rect 13116 47300 13172 47356
rect 13172 47300 13176 47356
rect 13112 47296 13176 47300
rect 13192 47356 13256 47360
rect 13192 47300 13196 47356
rect 13196 47300 13252 47356
rect 13252 47300 13256 47356
rect 13192 47296 13256 47300
rect 22952 47356 23016 47360
rect 22952 47300 22956 47356
rect 22956 47300 23012 47356
rect 23012 47300 23016 47356
rect 22952 47296 23016 47300
rect 23032 47356 23096 47360
rect 23032 47300 23036 47356
rect 23036 47300 23092 47356
rect 23092 47300 23096 47356
rect 23032 47296 23096 47300
rect 23112 47356 23176 47360
rect 23112 47300 23116 47356
rect 23116 47300 23172 47356
rect 23172 47300 23176 47356
rect 23112 47296 23176 47300
rect 23192 47356 23256 47360
rect 23192 47300 23196 47356
rect 23196 47300 23252 47356
rect 23252 47300 23256 47356
rect 23192 47296 23256 47300
rect 32952 47356 33016 47360
rect 32952 47300 32956 47356
rect 32956 47300 33012 47356
rect 33012 47300 33016 47356
rect 32952 47296 33016 47300
rect 33032 47356 33096 47360
rect 33032 47300 33036 47356
rect 33036 47300 33092 47356
rect 33092 47300 33096 47356
rect 33032 47296 33096 47300
rect 33112 47356 33176 47360
rect 33112 47300 33116 47356
rect 33116 47300 33172 47356
rect 33172 47300 33176 47356
rect 33112 47296 33176 47300
rect 33192 47356 33256 47360
rect 33192 47300 33196 47356
rect 33196 47300 33252 47356
rect 33252 47300 33256 47356
rect 33192 47296 33256 47300
rect 42952 47356 43016 47360
rect 42952 47300 42956 47356
rect 42956 47300 43012 47356
rect 43012 47300 43016 47356
rect 42952 47296 43016 47300
rect 43032 47356 43096 47360
rect 43032 47300 43036 47356
rect 43036 47300 43092 47356
rect 43092 47300 43096 47356
rect 43032 47296 43096 47300
rect 43112 47356 43176 47360
rect 43112 47300 43116 47356
rect 43116 47300 43172 47356
rect 43172 47300 43176 47356
rect 43112 47296 43176 47300
rect 43192 47356 43256 47360
rect 43192 47300 43196 47356
rect 43196 47300 43252 47356
rect 43252 47300 43256 47356
rect 43192 47296 43256 47300
rect 7952 46812 8016 46816
rect 7952 46756 7956 46812
rect 7956 46756 8012 46812
rect 8012 46756 8016 46812
rect 7952 46752 8016 46756
rect 8032 46812 8096 46816
rect 8032 46756 8036 46812
rect 8036 46756 8092 46812
rect 8092 46756 8096 46812
rect 8032 46752 8096 46756
rect 8112 46812 8176 46816
rect 8112 46756 8116 46812
rect 8116 46756 8172 46812
rect 8172 46756 8176 46812
rect 8112 46752 8176 46756
rect 8192 46812 8256 46816
rect 8192 46756 8196 46812
rect 8196 46756 8252 46812
rect 8252 46756 8256 46812
rect 8192 46752 8256 46756
rect 17952 46812 18016 46816
rect 17952 46756 17956 46812
rect 17956 46756 18012 46812
rect 18012 46756 18016 46812
rect 17952 46752 18016 46756
rect 18032 46812 18096 46816
rect 18032 46756 18036 46812
rect 18036 46756 18092 46812
rect 18092 46756 18096 46812
rect 18032 46752 18096 46756
rect 18112 46812 18176 46816
rect 18112 46756 18116 46812
rect 18116 46756 18172 46812
rect 18172 46756 18176 46812
rect 18112 46752 18176 46756
rect 18192 46812 18256 46816
rect 18192 46756 18196 46812
rect 18196 46756 18252 46812
rect 18252 46756 18256 46812
rect 18192 46752 18256 46756
rect 27952 46812 28016 46816
rect 27952 46756 27956 46812
rect 27956 46756 28012 46812
rect 28012 46756 28016 46812
rect 27952 46752 28016 46756
rect 28032 46812 28096 46816
rect 28032 46756 28036 46812
rect 28036 46756 28092 46812
rect 28092 46756 28096 46812
rect 28032 46752 28096 46756
rect 28112 46812 28176 46816
rect 28112 46756 28116 46812
rect 28116 46756 28172 46812
rect 28172 46756 28176 46812
rect 28112 46752 28176 46756
rect 28192 46812 28256 46816
rect 28192 46756 28196 46812
rect 28196 46756 28252 46812
rect 28252 46756 28256 46812
rect 28192 46752 28256 46756
rect 37952 46812 38016 46816
rect 37952 46756 37956 46812
rect 37956 46756 38012 46812
rect 38012 46756 38016 46812
rect 37952 46752 38016 46756
rect 38032 46812 38096 46816
rect 38032 46756 38036 46812
rect 38036 46756 38092 46812
rect 38092 46756 38096 46812
rect 38032 46752 38096 46756
rect 38112 46812 38176 46816
rect 38112 46756 38116 46812
rect 38116 46756 38172 46812
rect 38172 46756 38176 46812
rect 38112 46752 38176 46756
rect 38192 46812 38256 46816
rect 38192 46756 38196 46812
rect 38196 46756 38252 46812
rect 38252 46756 38256 46812
rect 38192 46752 38256 46756
rect 47952 46812 48016 46816
rect 47952 46756 47956 46812
rect 47956 46756 48012 46812
rect 48012 46756 48016 46812
rect 47952 46752 48016 46756
rect 48032 46812 48096 46816
rect 48032 46756 48036 46812
rect 48036 46756 48092 46812
rect 48092 46756 48096 46812
rect 48032 46752 48096 46756
rect 48112 46812 48176 46816
rect 48112 46756 48116 46812
rect 48116 46756 48172 46812
rect 48172 46756 48176 46812
rect 48112 46752 48176 46756
rect 48192 46812 48256 46816
rect 48192 46756 48196 46812
rect 48196 46756 48252 46812
rect 48252 46756 48256 46812
rect 48192 46752 48256 46756
rect 2952 46268 3016 46272
rect 2952 46212 2956 46268
rect 2956 46212 3012 46268
rect 3012 46212 3016 46268
rect 2952 46208 3016 46212
rect 3032 46268 3096 46272
rect 3032 46212 3036 46268
rect 3036 46212 3092 46268
rect 3092 46212 3096 46268
rect 3032 46208 3096 46212
rect 3112 46268 3176 46272
rect 3112 46212 3116 46268
rect 3116 46212 3172 46268
rect 3172 46212 3176 46268
rect 3112 46208 3176 46212
rect 3192 46268 3256 46272
rect 3192 46212 3196 46268
rect 3196 46212 3252 46268
rect 3252 46212 3256 46268
rect 3192 46208 3256 46212
rect 12952 46268 13016 46272
rect 12952 46212 12956 46268
rect 12956 46212 13012 46268
rect 13012 46212 13016 46268
rect 12952 46208 13016 46212
rect 13032 46268 13096 46272
rect 13032 46212 13036 46268
rect 13036 46212 13092 46268
rect 13092 46212 13096 46268
rect 13032 46208 13096 46212
rect 13112 46268 13176 46272
rect 13112 46212 13116 46268
rect 13116 46212 13172 46268
rect 13172 46212 13176 46268
rect 13112 46208 13176 46212
rect 13192 46268 13256 46272
rect 13192 46212 13196 46268
rect 13196 46212 13252 46268
rect 13252 46212 13256 46268
rect 13192 46208 13256 46212
rect 22952 46268 23016 46272
rect 22952 46212 22956 46268
rect 22956 46212 23012 46268
rect 23012 46212 23016 46268
rect 22952 46208 23016 46212
rect 23032 46268 23096 46272
rect 23032 46212 23036 46268
rect 23036 46212 23092 46268
rect 23092 46212 23096 46268
rect 23032 46208 23096 46212
rect 23112 46268 23176 46272
rect 23112 46212 23116 46268
rect 23116 46212 23172 46268
rect 23172 46212 23176 46268
rect 23112 46208 23176 46212
rect 23192 46268 23256 46272
rect 23192 46212 23196 46268
rect 23196 46212 23252 46268
rect 23252 46212 23256 46268
rect 23192 46208 23256 46212
rect 32952 46268 33016 46272
rect 32952 46212 32956 46268
rect 32956 46212 33012 46268
rect 33012 46212 33016 46268
rect 32952 46208 33016 46212
rect 33032 46268 33096 46272
rect 33032 46212 33036 46268
rect 33036 46212 33092 46268
rect 33092 46212 33096 46268
rect 33032 46208 33096 46212
rect 33112 46268 33176 46272
rect 33112 46212 33116 46268
rect 33116 46212 33172 46268
rect 33172 46212 33176 46268
rect 33112 46208 33176 46212
rect 33192 46268 33256 46272
rect 33192 46212 33196 46268
rect 33196 46212 33252 46268
rect 33252 46212 33256 46268
rect 33192 46208 33256 46212
rect 42952 46268 43016 46272
rect 42952 46212 42956 46268
rect 42956 46212 43012 46268
rect 43012 46212 43016 46268
rect 42952 46208 43016 46212
rect 43032 46268 43096 46272
rect 43032 46212 43036 46268
rect 43036 46212 43092 46268
rect 43092 46212 43096 46268
rect 43032 46208 43096 46212
rect 43112 46268 43176 46272
rect 43112 46212 43116 46268
rect 43116 46212 43172 46268
rect 43172 46212 43176 46268
rect 43112 46208 43176 46212
rect 43192 46268 43256 46272
rect 43192 46212 43196 46268
rect 43196 46212 43252 46268
rect 43252 46212 43256 46268
rect 43192 46208 43256 46212
rect 7952 45724 8016 45728
rect 7952 45668 7956 45724
rect 7956 45668 8012 45724
rect 8012 45668 8016 45724
rect 7952 45664 8016 45668
rect 8032 45724 8096 45728
rect 8032 45668 8036 45724
rect 8036 45668 8092 45724
rect 8092 45668 8096 45724
rect 8032 45664 8096 45668
rect 8112 45724 8176 45728
rect 8112 45668 8116 45724
rect 8116 45668 8172 45724
rect 8172 45668 8176 45724
rect 8112 45664 8176 45668
rect 8192 45724 8256 45728
rect 8192 45668 8196 45724
rect 8196 45668 8252 45724
rect 8252 45668 8256 45724
rect 8192 45664 8256 45668
rect 17952 45724 18016 45728
rect 17952 45668 17956 45724
rect 17956 45668 18012 45724
rect 18012 45668 18016 45724
rect 17952 45664 18016 45668
rect 18032 45724 18096 45728
rect 18032 45668 18036 45724
rect 18036 45668 18092 45724
rect 18092 45668 18096 45724
rect 18032 45664 18096 45668
rect 18112 45724 18176 45728
rect 18112 45668 18116 45724
rect 18116 45668 18172 45724
rect 18172 45668 18176 45724
rect 18112 45664 18176 45668
rect 18192 45724 18256 45728
rect 18192 45668 18196 45724
rect 18196 45668 18252 45724
rect 18252 45668 18256 45724
rect 18192 45664 18256 45668
rect 27952 45724 28016 45728
rect 27952 45668 27956 45724
rect 27956 45668 28012 45724
rect 28012 45668 28016 45724
rect 27952 45664 28016 45668
rect 28032 45724 28096 45728
rect 28032 45668 28036 45724
rect 28036 45668 28092 45724
rect 28092 45668 28096 45724
rect 28032 45664 28096 45668
rect 28112 45724 28176 45728
rect 28112 45668 28116 45724
rect 28116 45668 28172 45724
rect 28172 45668 28176 45724
rect 28112 45664 28176 45668
rect 28192 45724 28256 45728
rect 28192 45668 28196 45724
rect 28196 45668 28252 45724
rect 28252 45668 28256 45724
rect 28192 45664 28256 45668
rect 37952 45724 38016 45728
rect 37952 45668 37956 45724
rect 37956 45668 38012 45724
rect 38012 45668 38016 45724
rect 37952 45664 38016 45668
rect 38032 45724 38096 45728
rect 38032 45668 38036 45724
rect 38036 45668 38092 45724
rect 38092 45668 38096 45724
rect 38032 45664 38096 45668
rect 38112 45724 38176 45728
rect 38112 45668 38116 45724
rect 38116 45668 38172 45724
rect 38172 45668 38176 45724
rect 38112 45664 38176 45668
rect 38192 45724 38256 45728
rect 38192 45668 38196 45724
rect 38196 45668 38252 45724
rect 38252 45668 38256 45724
rect 38192 45664 38256 45668
rect 47952 45724 48016 45728
rect 47952 45668 47956 45724
rect 47956 45668 48012 45724
rect 48012 45668 48016 45724
rect 47952 45664 48016 45668
rect 48032 45724 48096 45728
rect 48032 45668 48036 45724
rect 48036 45668 48092 45724
rect 48092 45668 48096 45724
rect 48032 45664 48096 45668
rect 48112 45724 48176 45728
rect 48112 45668 48116 45724
rect 48116 45668 48172 45724
rect 48172 45668 48176 45724
rect 48112 45664 48176 45668
rect 48192 45724 48256 45728
rect 48192 45668 48196 45724
rect 48196 45668 48252 45724
rect 48252 45668 48256 45724
rect 48192 45664 48256 45668
rect 2952 45180 3016 45184
rect 2952 45124 2956 45180
rect 2956 45124 3012 45180
rect 3012 45124 3016 45180
rect 2952 45120 3016 45124
rect 3032 45180 3096 45184
rect 3032 45124 3036 45180
rect 3036 45124 3092 45180
rect 3092 45124 3096 45180
rect 3032 45120 3096 45124
rect 3112 45180 3176 45184
rect 3112 45124 3116 45180
rect 3116 45124 3172 45180
rect 3172 45124 3176 45180
rect 3112 45120 3176 45124
rect 3192 45180 3256 45184
rect 3192 45124 3196 45180
rect 3196 45124 3252 45180
rect 3252 45124 3256 45180
rect 3192 45120 3256 45124
rect 12952 45180 13016 45184
rect 12952 45124 12956 45180
rect 12956 45124 13012 45180
rect 13012 45124 13016 45180
rect 12952 45120 13016 45124
rect 13032 45180 13096 45184
rect 13032 45124 13036 45180
rect 13036 45124 13092 45180
rect 13092 45124 13096 45180
rect 13032 45120 13096 45124
rect 13112 45180 13176 45184
rect 13112 45124 13116 45180
rect 13116 45124 13172 45180
rect 13172 45124 13176 45180
rect 13112 45120 13176 45124
rect 13192 45180 13256 45184
rect 13192 45124 13196 45180
rect 13196 45124 13252 45180
rect 13252 45124 13256 45180
rect 13192 45120 13256 45124
rect 22952 45180 23016 45184
rect 22952 45124 22956 45180
rect 22956 45124 23012 45180
rect 23012 45124 23016 45180
rect 22952 45120 23016 45124
rect 23032 45180 23096 45184
rect 23032 45124 23036 45180
rect 23036 45124 23092 45180
rect 23092 45124 23096 45180
rect 23032 45120 23096 45124
rect 23112 45180 23176 45184
rect 23112 45124 23116 45180
rect 23116 45124 23172 45180
rect 23172 45124 23176 45180
rect 23112 45120 23176 45124
rect 23192 45180 23256 45184
rect 23192 45124 23196 45180
rect 23196 45124 23252 45180
rect 23252 45124 23256 45180
rect 23192 45120 23256 45124
rect 32952 45180 33016 45184
rect 32952 45124 32956 45180
rect 32956 45124 33012 45180
rect 33012 45124 33016 45180
rect 32952 45120 33016 45124
rect 33032 45180 33096 45184
rect 33032 45124 33036 45180
rect 33036 45124 33092 45180
rect 33092 45124 33096 45180
rect 33032 45120 33096 45124
rect 33112 45180 33176 45184
rect 33112 45124 33116 45180
rect 33116 45124 33172 45180
rect 33172 45124 33176 45180
rect 33112 45120 33176 45124
rect 33192 45180 33256 45184
rect 33192 45124 33196 45180
rect 33196 45124 33252 45180
rect 33252 45124 33256 45180
rect 33192 45120 33256 45124
rect 42952 45180 43016 45184
rect 42952 45124 42956 45180
rect 42956 45124 43012 45180
rect 43012 45124 43016 45180
rect 42952 45120 43016 45124
rect 43032 45180 43096 45184
rect 43032 45124 43036 45180
rect 43036 45124 43092 45180
rect 43092 45124 43096 45180
rect 43032 45120 43096 45124
rect 43112 45180 43176 45184
rect 43112 45124 43116 45180
rect 43116 45124 43172 45180
rect 43172 45124 43176 45180
rect 43112 45120 43176 45124
rect 43192 45180 43256 45184
rect 43192 45124 43196 45180
rect 43196 45124 43252 45180
rect 43252 45124 43256 45180
rect 43192 45120 43256 45124
rect 7952 44636 8016 44640
rect 7952 44580 7956 44636
rect 7956 44580 8012 44636
rect 8012 44580 8016 44636
rect 7952 44576 8016 44580
rect 8032 44636 8096 44640
rect 8032 44580 8036 44636
rect 8036 44580 8092 44636
rect 8092 44580 8096 44636
rect 8032 44576 8096 44580
rect 8112 44636 8176 44640
rect 8112 44580 8116 44636
rect 8116 44580 8172 44636
rect 8172 44580 8176 44636
rect 8112 44576 8176 44580
rect 8192 44636 8256 44640
rect 8192 44580 8196 44636
rect 8196 44580 8252 44636
rect 8252 44580 8256 44636
rect 8192 44576 8256 44580
rect 17952 44636 18016 44640
rect 17952 44580 17956 44636
rect 17956 44580 18012 44636
rect 18012 44580 18016 44636
rect 17952 44576 18016 44580
rect 18032 44636 18096 44640
rect 18032 44580 18036 44636
rect 18036 44580 18092 44636
rect 18092 44580 18096 44636
rect 18032 44576 18096 44580
rect 18112 44636 18176 44640
rect 18112 44580 18116 44636
rect 18116 44580 18172 44636
rect 18172 44580 18176 44636
rect 18112 44576 18176 44580
rect 18192 44636 18256 44640
rect 18192 44580 18196 44636
rect 18196 44580 18252 44636
rect 18252 44580 18256 44636
rect 18192 44576 18256 44580
rect 27952 44636 28016 44640
rect 27952 44580 27956 44636
rect 27956 44580 28012 44636
rect 28012 44580 28016 44636
rect 27952 44576 28016 44580
rect 28032 44636 28096 44640
rect 28032 44580 28036 44636
rect 28036 44580 28092 44636
rect 28092 44580 28096 44636
rect 28032 44576 28096 44580
rect 28112 44636 28176 44640
rect 28112 44580 28116 44636
rect 28116 44580 28172 44636
rect 28172 44580 28176 44636
rect 28112 44576 28176 44580
rect 28192 44636 28256 44640
rect 28192 44580 28196 44636
rect 28196 44580 28252 44636
rect 28252 44580 28256 44636
rect 28192 44576 28256 44580
rect 37952 44636 38016 44640
rect 37952 44580 37956 44636
rect 37956 44580 38012 44636
rect 38012 44580 38016 44636
rect 37952 44576 38016 44580
rect 38032 44636 38096 44640
rect 38032 44580 38036 44636
rect 38036 44580 38092 44636
rect 38092 44580 38096 44636
rect 38032 44576 38096 44580
rect 38112 44636 38176 44640
rect 38112 44580 38116 44636
rect 38116 44580 38172 44636
rect 38172 44580 38176 44636
rect 38112 44576 38176 44580
rect 38192 44636 38256 44640
rect 38192 44580 38196 44636
rect 38196 44580 38252 44636
rect 38252 44580 38256 44636
rect 38192 44576 38256 44580
rect 47952 44636 48016 44640
rect 47952 44580 47956 44636
rect 47956 44580 48012 44636
rect 48012 44580 48016 44636
rect 47952 44576 48016 44580
rect 48032 44636 48096 44640
rect 48032 44580 48036 44636
rect 48036 44580 48092 44636
rect 48092 44580 48096 44636
rect 48032 44576 48096 44580
rect 48112 44636 48176 44640
rect 48112 44580 48116 44636
rect 48116 44580 48172 44636
rect 48172 44580 48176 44636
rect 48112 44576 48176 44580
rect 48192 44636 48256 44640
rect 48192 44580 48196 44636
rect 48196 44580 48252 44636
rect 48252 44580 48256 44636
rect 48192 44576 48256 44580
rect 2952 44092 3016 44096
rect 2952 44036 2956 44092
rect 2956 44036 3012 44092
rect 3012 44036 3016 44092
rect 2952 44032 3016 44036
rect 3032 44092 3096 44096
rect 3032 44036 3036 44092
rect 3036 44036 3092 44092
rect 3092 44036 3096 44092
rect 3032 44032 3096 44036
rect 3112 44092 3176 44096
rect 3112 44036 3116 44092
rect 3116 44036 3172 44092
rect 3172 44036 3176 44092
rect 3112 44032 3176 44036
rect 3192 44092 3256 44096
rect 3192 44036 3196 44092
rect 3196 44036 3252 44092
rect 3252 44036 3256 44092
rect 3192 44032 3256 44036
rect 12952 44092 13016 44096
rect 12952 44036 12956 44092
rect 12956 44036 13012 44092
rect 13012 44036 13016 44092
rect 12952 44032 13016 44036
rect 13032 44092 13096 44096
rect 13032 44036 13036 44092
rect 13036 44036 13092 44092
rect 13092 44036 13096 44092
rect 13032 44032 13096 44036
rect 13112 44092 13176 44096
rect 13112 44036 13116 44092
rect 13116 44036 13172 44092
rect 13172 44036 13176 44092
rect 13112 44032 13176 44036
rect 13192 44092 13256 44096
rect 13192 44036 13196 44092
rect 13196 44036 13252 44092
rect 13252 44036 13256 44092
rect 13192 44032 13256 44036
rect 22952 44092 23016 44096
rect 22952 44036 22956 44092
rect 22956 44036 23012 44092
rect 23012 44036 23016 44092
rect 22952 44032 23016 44036
rect 23032 44092 23096 44096
rect 23032 44036 23036 44092
rect 23036 44036 23092 44092
rect 23092 44036 23096 44092
rect 23032 44032 23096 44036
rect 23112 44092 23176 44096
rect 23112 44036 23116 44092
rect 23116 44036 23172 44092
rect 23172 44036 23176 44092
rect 23112 44032 23176 44036
rect 23192 44092 23256 44096
rect 23192 44036 23196 44092
rect 23196 44036 23252 44092
rect 23252 44036 23256 44092
rect 23192 44032 23256 44036
rect 32952 44092 33016 44096
rect 32952 44036 32956 44092
rect 32956 44036 33012 44092
rect 33012 44036 33016 44092
rect 32952 44032 33016 44036
rect 33032 44092 33096 44096
rect 33032 44036 33036 44092
rect 33036 44036 33092 44092
rect 33092 44036 33096 44092
rect 33032 44032 33096 44036
rect 33112 44092 33176 44096
rect 33112 44036 33116 44092
rect 33116 44036 33172 44092
rect 33172 44036 33176 44092
rect 33112 44032 33176 44036
rect 33192 44092 33256 44096
rect 33192 44036 33196 44092
rect 33196 44036 33252 44092
rect 33252 44036 33256 44092
rect 33192 44032 33256 44036
rect 42952 44092 43016 44096
rect 42952 44036 42956 44092
rect 42956 44036 43012 44092
rect 43012 44036 43016 44092
rect 42952 44032 43016 44036
rect 43032 44092 43096 44096
rect 43032 44036 43036 44092
rect 43036 44036 43092 44092
rect 43092 44036 43096 44092
rect 43032 44032 43096 44036
rect 43112 44092 43176 44096
rect 43112 44036 43116 44092
rect 43116 44036 43172 44092
rect 43172 44036 43176 44092
rect 43112 44032 43176 44036
rect 43192 44092 43256 44096
rect 43192 44036 43196 44092
rect 43196 44036 43252 44092
rect 43252 44036 43256 44092
rect 43192 44032 43256 44036
rect 7952 43548 8016 43552
rect 7952 43492 7956 43548
rect 7956 43492 8012 43548
rect 8012 43492 8016 43548
rect 7952 43488 8016 43492
rect 8032 43548 8096 43552
rect 8032 43492 8036 43548
rect 8036 43492 8092 43548
rect 8092 43492 8096 43548
rect 8032 43488 8096 43492
rect 8112 43548 8176 43552
rect 8112 43492 8116 43548
rect 8116 43492 8172 43548
rect 8172 43492 8176 43548
rect 8112 43488 8176 43492
rect 8192 43548 8256 43552
rect 8192 43492 8196 43548
rect 8196 43492 8252 43548
rect 8252 43492 8256 43548
rect 8192 43488 8256 43492
rect 17952 43548 18016 43552
rect 17952 43492 17956 43548
rect 17956 43492 18012 43548
rect 18012 43492 18016 43548
rect 17952 43488 18016 43492
rect 18032 43548 18096 43552
rect 18032 43492 18036 43548
rect 18036 43492 18092 43548
rect 18092 43492 18096 43548
rect 18032 43488 18096 43492
rect 18112 43548 18176 43552
rect 18112 43492 18116 43548
rect 18116 43492 18172 43548
rect 18172 43492 18176 43548
rect 18112 43488 18176 43492
rect 18192 43548 18256 43552
rect 18192 43492 18196 43548
rect 18196 43492 18252 43548
rect 18252 43492 18256 43548
rect 18192 43488 18256 43492
rect 27952 43548 28016 43552
rect 27952 43492 27956 43548
rect 27956 43492 28012 43548
rect 28012 43492 28016 43548
rect 27952 43488 28016 43492
rect 28032 43548 28096 43552
rect 28032 43492 28036 43548
rect 28036 43492 28092 43548
rect 28092 43492 28096 43548
rect 28032 43488 28096 43492
rect 28112 43548 28176 43552
rect 28112 43492 28116 43548
rect 28116 43492 28172 43548
rect 28172 43492 28176 43548
rect 28112 43488 28176 43492
rect 28192 43548 28256 43552
rect 28192 43492 28196 43548
rect 28196 43492 28252 43548
rect 28252 43492 28256 43548
rect 28192 43488 28256 43492
rect 37952 43548 38016 43552
rect 37952 43492 37956 43548
rect 37956 43492 38012 43548
rect 38012 43492 38016 43548
rect 37952 43488 38016 43492
rect 38032 43548 38096 43552
rect 38032 43492 38036 43548
rect 38036 43492 38092 43548
rect 38092 43492 38096 43548
rect 38032 43488 38096 43492
rect 38112 43548 38176 43552
rect 38112 43492 38116 43548
rect 38116 43492 38172 43548
rect 38172 43492 38176 43548
rect 38112 43488 38176 43492
rect 38192 43548 38256 43552
rect 38192 43492 38196 43548
rect 38196 43492 38252 43548
rect 38252 43492 38256 43548
rect 38192 43488 38256 43492
rect 47952 43548 48016 43552
rect 47952 43492 47956 43548
rect 47956 43492 48012 43548
rect 48012 43492 48016 43548
rect 47952 43488 48016 43492
rect 48032 43548 48096 43552
rect 48032 43492 48036 43548
rect 48036 43492 48092 43548
rect 48092 43492 48096 43548
rect 48032 43488 48096 43492
rect 48112 43548 48176 43552
rect 48112 43492 48116 43548
rect 48116 43492 48172 43548
rect 48172 43492 48176 43548
rect 48112 43488 48176 43492
rect 48192 43548 48256 43552
rect 48192 43492 48196 43548
rect 48196 43492 48252 43548
rect 48252 43492 48256 43548
rect 48192 43488 48256 43492
rect 2952 43004 3016 43008
rect 2952 42948 2956 43004
rect 2956 42948 3012 43004
rect 3012 42948 3016 43004
rect 2952 42944 3016 42948
rect 3032 43004 3096 43008
rect 3032 42948 3036 43004
rect 3036 42948 3092 43004
rect 3092 42948 3096 43004
rect 3032 42944 3096 42948
rect 3112 43004 3176 43008
rect 3112 42948 3116 43004
rect 3116 42948 3172 43004
rect 3172 42948 3176 43004
rect 3112 42944 3176 42948
rect 3192 43004 3256 43008
rect 3192 42948 3196 43004
rect 3196 42948 3252 43004
rect 3252 42948 3256 43004
rect 3192 42944 3256 42948
rect 12952 43004 13016 43008
rect 12952 42948 12956 43004
rect 12956 42948 13012 43004
rect 13012 42948 13016 43004
rect 12952 42944 13016 42948
rect 13032 43004 13096 43008
rect 13032 42948 13036 43004
rect 13036 42948 13092 43004
rect 13092 42948 13096 43004
rect 13032 42944 13096 42948
rect 13112 43004 13176 43008
rect 13112 42948 13116 43004
rect 13116 42948 13172 43004
rect 13172 42948 13176 43004
rect 13112 42944 13176 42948
rect 13192 43004 13256 43008
rect 13192 42948 13196 43004
rect 13196 42948 13252 43004
rect 13252 42948 13256 43004
rect 13192 42944 13256 42948
rect 22952 43004 23016 43008
rect 22952 42948 22956 43004
rect 22956 42948 23012 43004
rect 23012 42948 23016 43004
rect 22952 42944 23016 42948
rect 23032 43004 23096 43008
rect 23032 42948 23036 43004
rect 23036 42948 23092 43004
rect 23092 42948 23096 43004
rect 23032 42944 23096 42948
rect 23112 43004 23176 43008
rect 23112 42948 23116 43004
rect 23116 42948 23172 43004
rect 23172 42948 23176 43004
rect 23112 42944 23176 42948
rect 23192 43004 23256 43008
rect 23192 42948 23196 43004
rect 23196 42948 23252 43004
rect 23252 42948 23256 43004
rect 23192 42944 23256 42948
rect 32952 43004 33016 43008
rect 32952 42948 32956 43004
rect 32956 42948 33012 43004
rect 33012 42948 33016 43004
rect 32952 42944 33016 42948
rect 33032 43004 33096 43008
rect 33032 42948 33036 43004
rect 33036 42948 33092 43004
rect 33092 42948 33096 43004
rect 33032 42944 33096 42948
rect 33112 43004 33176 43008
rect 33112 42948 33116 43004
rect 33116 42948 33172 43004
rect 33172 42948 33176 43004
rect 33112 42944 33176 42948
rect 33192 43004 33256 43008
rect 33192 42948 33196 43004
rect 33196 42948 33252 43004
rect 33252 42948 33256 43004
rect 33192 42944 33256 42948
rect 42952 43004 43016 43008
rect 42952 42948 42956 43004
rect 42956 42948 43012 43004
rect 43012 42948 43016 43004
rect 42952 42944 43016 42948
rect 43032 43004 43096 43008
rect 43032 42948 43036 43004
rect 43036 42948 43092 43004
rect 43092 42948 43096 43004
rect 43032 42944 43096 42948
rect 43112 43004 43176 43008
rect 43112 42948 43116 43004
rect 43116 42948 43172 43004
rect 43172 42948 43176 43004
rect 43112 42944 43176 42948
rect 43192 43004 43256 43008
rect 43192 42948 43196 43004
rect 43196 42948 43252 43004
rect 43252 42948 43256 43004
rect 43192 42944 43256 42948
rect 7952 42460 8016 42464
rect 7952 42404 7956 42460
rect 7956 42404 8012 42460
rect 8012 42404 8016 42460
rect 7952 42400 8016 42404
rect 8032 42460 8096 42464
rect 8032 42404 8036 42460
rect 8036 42404 8092 42460
rect 8092 42404 8096 42460
rect 8032 42400 8096 42404
rect 8112 42460 8176 42464
rect 8112 42404 8116 42460
rect 8116 42404 8172 42460
rect 8172 42404 8176 42460
rect 8112 42400 8176 42404
rect 8192 42460 8256 42464
rect 8192 42404 8196 42460
rect 8196 42404 8252 42460
rect 8252 42404 8256 42460
rect 8192 42400 8256 42404
rect 17952 42460 18016 42464
rect 17952 42404 17956 42460
rect 17956 42404 18012 42460
rect 18012 42404 18016 42460
rect 17952 42400 18016 42404
rect 18032 42460 18096 42464
rect 18032 42404 18036 42460
rect 18036 42404 18092 42460
rect 18092 42404 18096 42460
rect 18032 42400 18096 42404
rect 18112 42460 18176 42464
rect 18112 42404 18116 42460
rect 18116 42404 18172 42460
rect 18172 42404 18176 42460
rect 18112 42400 18176 42404
rect 18192 42460 18256 42464
rect 18192 42404 18196 42460
rect 18196 42404 18252 42460
rect 18252 42404 18256 42460
rect 18192 42400 18256 42404
rect 27952 42460 28016 42464
rect 27952 42404 27956 42460
rect 27956 42404 28012 42460
rect 28012 42404 28016 42460
rect 27952 42400 28016 42404
rect 28032 42460 28096 42464
rect 28032 42404 28036 42460
rect 28036 42404 28092 42460
rect 28092 42404 28096 42460
rect 28032 42400 28096 42404
rect 28112 42460 28176 42464
rect 28112 42404 28116 42460
rect 28116 42404 28172 42460
rect 28172 42404 28176 42460
rect 28112 42400 28176 42404
rect 28192 42460 28256 42464
rect 28192 42404 28196 42460
rect 28196 42404 28252 42460
rect 28252 42404 28256 42460
rect 28192 42400 28256 42404
rect 37952 42460 38016 42464
rect 37952 42404 37956 42460
rect 37956 42404 38012 42460
rect 38012 42404 38016 42460
rect 37952 42400 38016 42404
rect 38032 42460 38096 42464
rect 38032 42404 38036 42460
rect 38036 42404 38092 42460
rect 38092 42404 38096 42460
rect 38032 42400 38096 42404
rect 38112 42460 38176 42464
rect 38112 42404 38116 42460
rect 38116 42404 38172 42460
rect 38172 42404 38176 42460
rect 38112 42400 38176 42404
rect 38192 42460 38256 42464
rect 38192 42404 38196 42460
rect 38196 42404 38252 42460
rect 38252 42404 38256 42460
rect 38192 42400 38256 42404
rect 47952 42460 48016 42464
rect 47952 42404 47956 42460
rect 47956 42404 48012 42460
rect 48012 42404 48016 42460
rect 47952 42400 48016 42404
rect 48032 42460 48096 42464
rect 48032 42404 48036 42460
rect 48036 42404 48092 42460
rect 48092 42404 48096 42460
rect 48032 42400 48096 42404
rect 48112 42460 48176 42464
rect 48112 42404 48116 42460
rect 48116 42404 48172 42460
rect 48172 42404 48176 42460
rect 48112 42400 48176 42404
rect 48192 42460 48256 42464
rect 48192 42404 48196 42460
rect 48196 42404 48252 42460
rect 48252 42404 48256 42460
rect 48192 42400 48256 42404
rect 39988 42060 40052 42124
rect 2952 41916 3016 41920
rect 2952 41860 2956 41916
rect 2956 41860 3012 41916
rect 3012 41860 3016 41916
rect 2952 41856 3016 41860
rect 3032 41916 3096 41920
rect 3032 41860 3036 41916
rect 3036 41860 3092 41916
rect 3092 41860 3096 41916
rect 3032 41856 3096 41860
rect 3112 41916 3176 41920
rect 3112 41860 3116 41916
rect 3116 41860 3172 41916
rect 3172 41860 3176 41916
rect 3112 41856 3176 41860
rect 3192 41916 3256 41920
rect 3192 41860 3196 41916
rect 3196 41860 3252 41916
rect 3252 41860 3256 41916
rect 3192 41856 3256 41860
rect 12952 41916 13016 41920
rect 12952 41860 12956 41916
rect 12956 41860 13012 41916
rect 13012 41860 13016 41916
rect 12952 41856 13016 41860
rect 13032 41916 13096 41920
rect 13032 41860 13036 41916
rect 13036 41860 13092 41916
rect 13092 41860 13096 41916
rect 13032 41856 13096 41860
rect 13112 41916 13176 41920
rect 13112 41860 13116 41916
rect 13116 41860 13172 41916
rect 13172 41860 13176 41916
rect 13112 41856 13176 41860
rect 13192 41916 13256 41920
rect 13192 41860 13196 41916
rect 13196 41860 13252 41916
rect 13252 41860 13256 41916
rect 13192 41856 13256 41860
rect 22952 41916 23016 41920
rect 22952 41860 22956 41916
rect 22956 41860 23012 41916
rect 23012 41860 23016 41916
rect 22952 41856 23016 41860
rect 23032 41916 23096 41920
rect 23032 41860 23036 41916
rect 23036 41860 23092 41916
rect 23092 41860 23096 41916
rect 23032 41856 23096 41860
rect 23112 41916 23176 41920
rect 23112 41860 23116 41916
rect 23116 41860 23172 41916
rect 23172 41860 23176 41916
rect 23112 41856 23176 41860
rect 23192 41916 23256 41920
rect 23192 41860 23196 41916
rect 23196 41860 23252 41916
rect 23252 41860 23256 41916
rect 23192 41856 23256 41860
rect 32952 41916 33016 41920
rect 32952 41860 32956 41916
rect 32956 41860 33012 41916
rect 33012 41860 33016 41916
rect 32952 41856 33016 41860
rect 33032 41916 33096 41920
rect 33032 41860 33036 41916
rect 33036 41860 33092 41916
rect 33092 41860 33096 41916
rect 33032 41856 33096 41860
rect 33112 41916 33176 41920
rect 33112 41860 33116 41916
rect 33116 41860 33172 41916
rect 33172 41860 33176 41916
rect 33112 41856 33176 41860
rect 33192 41916 33256 41920
rect 33192 41860 33196 41916
rect 33196 41860 33252 41916
rect 33252 41860 33256 41916
rect 33192 41856 33256 41860
rect 42952 41916 43016 41920
rect 42952 41860 42956 41916
rect 42956 41860 43012 41916
rect 43012 41860 43016 41916
rect 42952 41856 43016 41860
rect 43032 41916 43096 41920
rect 43032 41860 43036 41916
rect 43036 41860 43092 41916
rect 43092 41860 43096 41916
rect 43032 41856 43096 41860
rect 43112 41916 43176 41920
rect 43112 41860 43116 41916
rect 43116 41860 43172 41916
rect 43172 41860 43176 41916
rect 43112 41856 43176 41860
rect 43192 41916 43256 41920
rect 43192 41860 43196 41916
rect 43196 41860 43252 41916
rect 43252 41860 43256 41916
rect 43192 41856 43256 41860
rect 40540 41652 40604 41716
rect 7952 41372 8016 41376
rect 7952 41316 7956 41372
rect 7956 41316 8012 41372
rect 8012 41316 8016 41372
rect 7952 41312 8016 41316
rect 8032 41372 8096 41376
rect 8032 41316 8036 41372
rect 8036 41316 8092 41372
rect 8092 41316 8096 41372
rect 8032 41312 8096 41316
rect 8112 41372 8176 41376
rect 8112 41316 8116 41372
rect 8116 41316 8172 41372
rect 8172 41316 8176 41372
rect 8112 41312 8176 41316
rect 8192 41372 8256 41376
rect 8192 41316 8196 41372
rect 8196 41316 8252 41372
rect 8252 41316 8256 41372
rect 8192 41312 8256 41316
rect 17952 41372 18016 41376
rect 17952 41316 17956 41372
rect 17956 41316 18012 41372
rect 18012 41316 18016 41372
rect 17952 41312 18016 41316
rect 18032 41372 18096 41376
rect 18032 41316 18036 41372
rect 18036 41316 18092 41372
rect 18092 41316 18096 41372
rect 18032 41312 18096 41316
rect 18112 41372 18176 41376
rect 18112 41316 18116 41372
rect 18116 41316 18172 41372
rect 18172 41316 18176 41372
rect 18112 41312 18176 41316
rect 18192 41372 18256 41376
rect 18192 41316 18196 41372
rect 18196 41316 18252 41372
rect 18252 41316 18256 41372
rect 18192 41312 18256 41316
rect 27952 41372 28016 41376
rect 27952 41316 27956 41372
rect 27956 41316 28012 41372
rect 28012 41316 28016 41372
rect 27952 41312 28016 41316
rect 28032 41372 28096 41376
rect 28032 41316 28036 41372
rect 28036 41316 28092 41372
rect 28092 41316 28096 41372
rect 28032 41312 28096 41316
rect 28112 41372 28176 41376
rect 28112 41316 28116 41372
rect 28116 41316 28172 41372
rect 28172 41316 28176 41372
rect 28112 41312 28176 41316
rect 28192 41372 28256 41376
rect 28192 41316 28196 41372
rect 28196 41316 28252 41372
rect 28252 41316 28256 41372
rect 28192 41312 28256 41316
rect 37952 41372 38016 41376
rect 37952 41316 37956 41372
rect 37956 41316 38012 41372
rect 38012 41316 38016 41372
rect 37952 41312 38016 41316
rect 38032 41372 38096 41376
rect 38032 41316 38036 41372
rect 38036 41316 38092 41372
rect 38092 41316 38096 41372
rect 38032 41312 38096 41316
rect 38112 41372 38176 41376
rect 38112 41316 38116 41372
rect 38116 41316 38172 41372
rect 38172 41316 38176 41372
rect 38112 41312 38176 41316
rect 38192 41372 38256 41376
rect 38192 41316 38196 41372
rect 38196 41316 38252 41372
rect 38252 41316 38256 41372
rect 38192 41312 38256 41316
rect 47952 41372 48016 41376
rect 47952 41316 47956 41372
rect 47956 41316 48012 41372
rect 48012 41316 48016 41372
rect 47952 41312 48016 41316
rect 48032 41372 48096 41376
rect 48032 41316 48036 41372
rect 48036 41316 48092 41372
rect 48092 41316 48096 41372
rect 48032 41312 48096 41316
rect 48112 41372 48176 41376
rect 48112 41316 48116 41372
rect 48116 41316 48172 41372
rect 48172 41316 48176 41372
rect 48112 41312 48176 41316
rect 48192 41372 48256 41376
rect 48192 41316 48196 41372
rect 48196 41316 48252 41372
rect 48252 41316 48256 41372
rect 48192 41312 48256 41316
rect 2952 40828 3016 40832
rect 2952 40772 2956 40828
rect 2956 40772 3012 40828
rect 3012 40772 3016 40828
rect 2952 40768 3016 40772
rect 3032 40828 3096 40832
rect 3032 40772 3036 40828
rect 3036 40772 3092 40828
rect 3092 40772 3096 40828
rect 3032 40768 3096 40772
rect 3112 40828 3176 40832
rect 3112 40772 3116 40828
rect 3116 40772 3172 40828
rect 3172 40772 3176 40828
rect 3112 40768 3176 40772
rect 3192 40828 3256 40832
rect 3192 40772 3196 40828
rect 3196 40772 3252 40828
rect 3252 40772 3256 40828
rect 3192 40768 3256 40772
rect 12952 40828 13016 40832
rect 12952 40772 12956 40828
rect 12956 40772 13012 40828
rect 13012 40772 13016 40828
rect 12952 40768 13016 40772
rect 13032 40828 13096 40832
rect 13032 40772 13036 40828
rect 13036 40772 13092 40828
rect 13092 40772 13096 40828
rect 13032 40768 13096 40772
rect 13112 40828 13176 40832
rect 13112 40772 13116 40828
rect 13116 40772 13172 40828
rect 13172 40772 13176 40828
rect 13112 40768 13176 40772
rect 13192 40828 13256 40832
rect 13192 40772 13196 40828
rect 13196 40772 13252 40828
rect 13252 40772 13256 40828
rect 13192 40768 13256 40772
rect 22952 40828 23016 40832
rect 22952 40772 22956 40828
rect 22956 40772 23012 40828
rect 23012 40772 23016 40828
rect 22952 40768 23016 40772
rect 23032 40828 23096 40832
rect 23032 40772 23036 40828
rect 23036 40772 23092 40828
rect 23092 40772 23096 40828
rect 23032 40768 23096 40772
rect 23112 40828 23176 40832
rect 23112 40772 23116 40828
rect 23116 40772 23172 40828
rect 23172 40772 23176 40828
rect 23112 40768 23176 40772
rect 23192 40828 23256 40832
rect 23192 40772 23196 40828
rect 23196 40772 23252 40828
rect 23252 40772 23256 40828
rect 23192 40768 23256 40772
rect 32952 40828 33016 40832
rect 32952 40772 32956 40828
rect 32956 40772 33012 40828
rect 33012 40772 33016 40828
rect 32952 40768 33016 40772
rect 33032 40828 33096 40832
rect 33032 40772 33036 40828
rect 33036 40772 33092 40828
rect 33092 40772 33096 40828
rect 33032 40768 33096 40772
rect 33112 40828 33176 40832
rect 33112 40772 33116 40828
rect 33116 40772 33172 40828
rect 33172 40772 33176 40828
rect 33112 40768 33176 40772
rect 33192 40828 33256 40832
rect 33192 40772 33196 40828
rect 33196 40772 33252 40828
rect 33252 40772 33256 40828
rect 33192 40768 33256 40772
rect 42952 40828 43016 40832
rect 42952 40772 42956 40828
rect 42956 40772 43012 40828
rect 43012 40772 43016 40828
rect 42952 40768 43016 40772
rect 43032 40828 43096 40832
rect 43032 40772 43036 40828
rect 43036 40772 43092 40828
rect 43092 40772 43096 40828
rect 43032 40768 43096 40772
rect 43112 40828 43176 40832
rect 43112 40772 43116 40828
rect 43116 40772 43172 40828
rect 43172 40772 43176 40828
rect 43112 40768 43176 40772
rect 43192 40828 43256 40832
rect 43192 40772 43196 40828
rect 43196 40772 43252 40828
rect 43252 40772 43256 40828
rect 43192 40768 43256 40772
rect 41276 40564 41340 40628
rect 7952 40284 8016 40288
rect 7952 40228 7956 40284
rect 7956 40228 8012 40284
rect 8012 40228 8016 40284
rect 7952 40224 8016 40228
rect 8032 40284 8096 40288
rect 8032 40228 8036 40284
rect 8036 40228 8092 40284
rect 8092 40228 8096 40284
rect 8032 40224 8096 40228
rect 8112 40284 8176 40288
rect 8112 40228 8116 40284
rect 8116 40228 8172 40284
rect 8172 40228 8176 40284
rect 8112 40224 8176 40228
rect 8192 40284 8256 40288
rect 8192 40228 8196 40284
rect 8196 40228 8252 40284
rect 8252 40228 8256 40284
rect 8192 40224 8256 40228
rect 17952 40284 18016 40288
rect 17952 40228 17956 40284
rect 17956 40228 18012 40284
rect 18012 40228 18016 40284
rect 17952 40224 18016 40228
rect 18032 40284 18096 40288
rect 18032 40228 18036 40284
rect 18036 40228 18092 40284
rect 18092 40228 18096 40284
rect 18032 40224 18096 40228
rect 18112 40284 18176 40288
rect 18112 40228 18116 40284
rect 18116 40228 18172 40284
rect 18172 40228 18176 40284
rect 18112 40224 18176 40228
rect 18192 40284 18256 40288
rect 18192 40228 18196 40284
rect 18196 40228 18252 40284
rect 18252 40228 18256 40284
rect 18192 40224 18256 40228
rect 27952 40284 28016 40288
rect 27952 40228 27956 40284
rect 27956 40228 28012 40284
rect 28012 40228 28016 40284
rect 27952 40224 28016 40228
rect 28032 40284 28096 40288
rect 28032 40228 28036 40284
rect 28036 40228 28092 40284
rect 28092 40228 28096 40284
rect 28032 40224 28096 40228
rect 28112 40284 28176 40288
rect 28112 40228 28116 40284
rect 28116 40228 28172 40284
rect 28172 40228 28176 40284
rect 28112 40224 28176 40228
rect 28192 40284 28256 40288
rect 28192 40228 28196 40284
rect 28196 40228 28252 40284
rect 28252 40228 28256 40284
rect 28192 40224 28256 40228
rect 37952 40284 38016 40288
rect 37952 40228 37956 40284
rect 37956 40228 38012 40284
rect 38012 40228 38016 40284
rect 37952 40224 38016 40228
rect 38032 40284 38096 40288
rect 38032 40228 38036 40284
rect 38036 40228 38092 40284
rect 38092 40228 38096 40284
rect 38032 40224 38096 40228
rect 38112 40284 38176 40288
rect 38112 40228 38116 40284
rect 38116 40228 38172 40284
rect 38172 40228 38176 40284
rect 38112 40224 38176 40228
rect 38192 40284 38256 40288
rect 38192 40228 38196 40284
rect 38196 40228 38252 40284
rect 38252 40228 38256 40284
rect 38192 40224 38256 40228
rect 47952 40284 48016 40288
rect 47952 40228 47956 40284
rect 47956 40228 48012 40284
rect 48012 40228 48016 40284
rect 47952 40224 48016 40228
rect 48032 40284 48096 40288
rect 48032 40228 48036 40284
rect 48036 40228 48092 40284
rect 48092 40228 48096 40284
rect 48032 40224 48096 40228
rect 48112 40284 48176 40288
rect 48112 40228 48116 40284
rect 48116 40228 48172 40284
rect 48172 40228 48176 40284
rect 48112 40224 48176 40228
rect 48192 40284 48256 40288
rect 48192 40228 48196 40284
rect 48196 40228 48252 40284
rect 48252 40228 48256 40284
rect 48192 40224 48256 40228
rect 30420 40020 30484 40084
rect 2952 39740 3016 39744
rect 2952 39684 2956 39740
rect 2956 39684 3012 39740
rect 3012 39684 3016 39740
rect 2952 39680 3016 39684
rect 3032 39740 3096 39744
rect 3032 39684 3036 39740
rect 3036 39684 3092 39740
rect 3092 39684 3096 39740
rect 3032 39680 3096 39684
rect 3112 39740 3176 39744
rect 3112 39684 3116 39740
rect 3116 39684 3172 39740
rect 3172 39684 3176 39740
rect 3112 39680 3176 39684
rect 3192 39740 3256 39744
rect 3192 39684 3196 39740
rect 3196 39684 3252 39740
rect 3252 39684 3256 39740
rect 3192 39680 3256 39684
rect 12952 39740 13016 39744
rect 12952 39684 12956 39740
rect 12956 39684 13012 39740
rect 13012 39684 13016 39740
rect 12952 39680 13016 39684
rect 13032 39740 13096 39744
rect 13032 39684 13036 39740
rect 13036 39684 13092 39740
rect 13092 39684 13096 39740
rect 13032 39680 13096 39684
rect 13112 39740 13176 39744
rect 13112 39684 13116 39740
rect 13116 39684 13172 39740
rect 13172 39684 13176 39740
rect 13112 39680 13176 39684
rect 13192 39740 13256 39744
rect 13192 39684 13196 39740
rect 13196 39684 13252 39740
rect 13252 39684 13256 39740
rect 13192 39680 13256 39684
rect 22952 39740 23016 39744
rect 22952 39684 22956 39740
rect 22956 39684 23012 39740
rect 23012 39684 23016 39740
rect 22952 39680 23016 39684
rect 23032 39740 23096 39744
rect 23032 39684 23036 39740
rect 23036 39684 23092 39740
rect 23092 39684 23096 39740
rect 23032 39680 23096 39684
rect 23112 39740 23176 39744
rect 23112 39684 23116 39740
rect 23116 39684 23172 39740
rect 23172 39684 23176 39740
rect 23112 39680 23176 39684
rect 23192 39740 23256 39744
rect 23192 39684 23196 39740
rect 23196 39684 23252 39740
rect 23252 39684 23256 39740
rect 23192 39680 23256 39684
rect 32952 39740 33016 39744
rect 32952 39684 32956 39740
rect 32956 39684 33012 39740
rect 33012 39684 33016 39740
rect 32952 39680 33016 39684
rect 33032 39740 33096 39744
rect 33032 39684 33036 39740
rect 33036 39684 33092 39740
rect 33092 39684 33096 39740
rect 33032 39680 33096 39684
rect 33112 39740 33176 39744
rect 33112 39684 33116 39740
rect 33116 39684 33172 39740
rect 33172 39684 33176 39740
rect 33112 39680 33176 39684
rect 33192 39740 33256 39744
rect 33192 39684 33196 39740
rect 33196 39684 33252 39740
rect 33252 39684 33256 39740
rect 33192 39680 33256 39684
rect 42952 39740 43016 39744
rect 42952 39684 42956 39740
rect 42956 39684 43012 39740
rect 43012 39684 43016 39740
rect 42952 39680 43016 39684
rect 43032 39740 43096 39744
rect 43032 39684 43036 39740
rect 43036 39684 43092 39740
rect 43092 39684 43096 39740
rect 43032 39680 43096 39684
rect 43112 39740 43176 39744
rect 43112 39684 43116 39740
rect 43116 39684 43172 39740
rect 43172 39684 43176 39740
rect 43112 39680 43176 39684
rect 43192 39740 43256 39744
rect 43192 39684 43196 39740
rect 43196 39684 43252 39740
rect 43252 39684 43256 39740
rect 43192 39680 43256 39684
rect 7952 39196 8016 39200
rect 7952 39140 7956 39196
rect 7956 39140 8012 39196
rect 8012 39140 8016 39196
rect 7952 39136 8016 39140
rect 8032 39196 8096 39200
rect 8032 39140 8036 39196
rect 8036 39140 8092 39196
rect 8092 39140 8096 39196
rect 8032 39136 8096 39140
rect 8112 39196 8176 39200
rect 8112 39140 8116 39196
rect 8116 39140 8172 39196
rect 8172 39140 8176 39196
rect 8112 39136 8176 39140
rect 8192 39196 8256 39200
rect 8192 39140 8196 39196
rect 8196 39140 8252 39196
rect 8252 39140 8256 39196
rect 8192 39136 8256 39140
rect 17952 39196 18016 39200
rect 17952 39140 17956 39196
rect 17956 39140 18012 39196
rect 18012 39140 18016 39196
rect 17952 39136 18016 39140
rect 18032 39196 18096 39200
rect 18032 39140 18036 39196
rect 18036 39140 18092 39196
rect 18092 39140 18096 39196
rect 18032 39136 18096 39140
rect 18112 39196 18176 39200
rect 18112 39140 18116 39196
rect 18116 39140 18172 39196
rect 18172 39140 18176 39196
rect 18112 39136 18176 39140
rect 18192 39196 18256 39200
rect 18192 39140 18196 39196
rect 18196 39140 18252 39196
rect 18252 39140 18256 39196
rect 18192 39136 18256 39140
rect 27952 39196 28016 39200
rect 27952 39140 27956 39196
rect 27956 39140 28012 39196
rect 28012 39140 28016 39196
rect 27952 39136 28016 39140
rect 28032 39196 28096 39200
rect 28032 39140 28036 39196
rect 28036 39140 28092 39196
rect 28092 39140 28096 39196
rect 28032 39136 28096 39140
rect 28112 39196 28176 39200
rect 28112 39140 28116 39196
rect 28116 39140 28172 39196
rect 28172 39140 28176 39196
rect 28112 39136 28176 39140
rect 28192 39196 28256 39200
rect 28192 39140 28196 39196
rect 28196 39140 28252 39196
rect 28252 39140 28256 39196
rect 28192 39136 28256 39140
rect 37952 39196 38016 39200
rect 37952 39140 37956 39196
rect 37956 39140 38012 39196
rect 38012 39140 38016 39196
rect 37952 39136 38016 39140
rect 38032 39196 38096 39200
rect 38032 39140 38036 39196
rect 38036 39140 38092 39196
rect 38092 39140 38096 39196
rect 38032 39136 38096 39140
rect 38112 39196 38176 39200
rect 38112 39140 38116 39196
rect 38116 39140 38172 39196
rect 38172 39140 38176 39196
rect 38112 39136 38176 39140
rect 38192 39196 38256 39200
rect 38192 39140 38196 39196
rect 38196 39140 38252 39196
rect 38252 39140 38256 39196
rect 38192 39136 38256 39140
rect 47952 39196 48016 39200
rect 47952 39140 47956 39196
rect 47956 39140 48012 39196
rect 48012 39140 48016 39196
rect 47952 39136 48016 39140
rect 48032 39196 48096 39200
rect 48032 39140 48036 39196
rect 48036 39140 48092 39196
rect 48092 39140 48096 39196
rect 48032 39136 48096 39140
rect 48112 39196 48176 39200
rect 48112 39140 48116 39196
rect 48116 39140 48172 39196
rect 48172 39140 48176 39196
rect 48112 39136 48176 39140
rect 48192 39196 48256 39200
rect 48192 39140 48196 39196
rect 48196 39140 48252 39196
rect 48252 39140 48256 39196
rect 48192 39136 48256 39140
rect 2952 38652 3016 38656
rect 2952 38596 2956 38652
rect 2956 38596 3012 38652
rect 3012 38596 3016 38652
rect 2952 38592 3016 38596
rect 3032 38652 3096 38656
rect 3032 38596 3036 38652
rect 3036 38596 3092 38652
rect 3092 38596 3096 38652
rect 3032 38592 3096 38596
rect 3112 38652 3176 38656
rect 3112 38596 3116 38652
rect 3116 38596 3172 38652
rect 3172 38596 3176 38652
rect 3112 38592 3176 38596
rect 3192 38652 3256 38656
rect 3192 38596 3196 38652
rect 3196 38596 3252 38652
rect 3252 38596 3256 38652
rect 3192 38592 3256 38596
rect 12952 38652 13016 38656
rect 12952 38596 12956 38652
rect 12956 38596 13012 38652
rect 13012 38596 13016 38652
rect 12952 38592 13016 38596
rect 13032 38652 13096 38656
rect 13032 38596 13036 38652
rect 13036 38596 13092 38652
rect 13092 38596 13096 38652
rect 13032 38592 13096 38596
rect 13112 38652 13176 38656
rect 13112 38596 13116 38652
rect 13116 38596 13172 38652
rect 13172 38596 13176 38652
rect 13112 38592 13176 38596
rect 13192 38652 13256 38656
rect 13192 38596 13196 38652
rect 13196 38596 13252 38652
rect 13252 38596 13256 38652
rect 13192 38592 13256 38596
rect 22952 38652 23016 38656
rect 22952 38596 22956 38652
rect 22956 38596 23012 38652
rect 23012 38596 23016 38652
rect 22952 38592 23016 38596
rect 23032 38652 23096 38656
rect 23032 38596 23036 38652
rect 23036 38596 23092 38652
rect 23092 38596 23096 38652
rect 23032 38592 23096 38596
rect 23112 38652 23176 38656
rect 23112 38596 23116 38652
rect 23116 38596 23172 38652
rect 23172 38596 23176 38652
rect 23112 38592 23176 38596
rect 23192 38652 23256 38656
rect 23192 38596 23196 38652
rect 23196 38596 23252 38652
rect 23252 38596 23256 38652
rect 23192 38592 23256 38596
rect 32952 38652 33016 38656
rect 32952 38596 32956 38652
rect 32956 38596 33012 38652
rect 33012 38596 33016 38652
rect 32952 38592 33016 38596
rect 33032 38652 33096 38656
rect 33032 38596 33036 38652
rect 33036 38596 33092 38652
rect 33092 38596 33096 38652
rect 33032 38592 33096 38596
rect 33112 38652 33176 38656
rect 33112 38596 33116 38652
rect 33116 38596 33172 38652
rect 33172 38596 33176 38652
rect 33112 38592 33176 38596
rect 33192 38652 33256 38656
rect 33192 38596 33196 38652
rect 33196 38596 33252 38652
rect 33252 38596 33256 38652
rect 33192 38592 33256 38596
rect 42952 38652 43016 38656
rect 42952 38596 42956 38652
rect 42956 38596 43012 38652
rect 43012 38596 43016 38652
rect 42952 38592 43016 38596
rect 43032 38652 43096 38656
rect 43032 38596 43036 38652
rect 43036 38596 43092 38652
rect 43092 38596 43096 38652
rect 43032 38592 43096 38596
rect 43112 38652 43176 38656
rect 43112 38596 43116 38652
rect 43116 38596 43172 38652
rect 43172 38596 43176 38652
rect 43112 38592 43176 38596
rect 43192 38652 43256 38656
rect 43192 38596 43196 38652
rect 43196 38596 43252 38652
rect 43252 38596 43256 38652
rect 43192 38592 43256 38596
rect 7952 38108 8016 38112
rect 7952 38052 7956 38108
rect 7956 38052 8012 38108
rect 8012 38052 8016 38108
rect 7952 38048 8016 38052
rect 8032 38108 8096 38112
rect 8032 38052 8036 38108
rect 8036 38052 8092 38108
rect 8092 38052 8096 38108
rect 8032 38048 8096 38052
rect 8112 38108 8176 38112
rect 8112 38052 8116 38108
rect 8116 38052 8172 38108
rect 8172 38052 8176 38108
rect 8112 38048 8176 38052
rect 8192 38108 8256 38112
rect 8192 38052 8196 38108
rect 8196 38052 8252 38108
rect 8252 38052 8256 38108
rect 8192 38048 8256 38052
rect 17952 38108 18016 38112
rect 17952 38052 17956 38108
rect 17956 38052 18012 38108
rect 18012 38052 18016 38108
rect 17952 38048 18016 38052
rect 18032 38108 18096 38112
rect 18032 38052 18036 38108
rect 18036 38052 18092 38108
rect 18092 38052 18096 38108
rect 18032 38048 18096 38052
rect 18112 38108 18176 38112
rect 18112 38052 18116 38108
rect 18116 38052 18172 38108
rect 18172 38052 18176 38108
rect 18112 38048 18176 38052
rect 18192 38108 18256 38112
rect 18192 38052 18196 38108
rect 18196 38052 18252 38108
rect 18252 38052 18256 38108
rect 18192 38048 18256 38052
rect 27952 38108 28016 38112
rect 27952 38052 27956 38108
rect 27956 38052 28012 38108
rect 28012 38052 28016 38108
rect 27952 38048 28016 38052
rect 28032 38108 28096 38112
rect 28032 38052 28036 38108
rect 28036 38052 28092 38108
rect 28092 38052 28096 38108
rect 28032 38048 28096 38052
rect 28112 38108 28176 38112
rect 28112 38052 28116 38108
rect 28116 38052 28172 38108
rect 28172 38052 28176 38108
rect 28112 38048 28176 38052
rect 28192 38108 28256 38112
rect 28192 38052 28196 38108
rect 28196 38052 28252 38108
rect 28252 38052 28256 38108
rect 28192 38048 28256 38052
rect 37952 38108 38016 38112
rect 37952 38052 37956 38108
rect 37956 38052 38012 38108
rect 38012 38052 38016 38108
rect 37952 38048 38016 38052
rect 38032 38108 38096 38112
rect 38032 38052 38036 38108
rect 38036 38052 38092 38108
rect 38092 38052 38096 38108
rect 38032 38048 38096 38052
rect 38112 38108 38176 38112
rect 38112 38052 38116 38108
rect 38116 38052 38172 38108
rect 38172 38052 38176 38108
rect 38112 38048 38176 38052
rect 38192 38108 38256 38112
rect 38192 38052 38196 38108
rect 38196 38052 38252 38108
rect 38252 38052 38256 38108
rect 38192 38048 38256 38052
rect 47952 38108 48016 38112
rect 47952 38052 47956 38108
rect 47956 38052 48012 38108
rect 48012 38052 48016 38108
rect 47952 38048 48016 38052
rect 48032 38108 48096 38112
rect 48032 38052 48036 38108
rect 48036 38052 48092 38108
rect 48092 38052 48096 38108
rect 48032 38048 48096 38052
rect 48112 38108 48176 38112
rect 48112 38052 48116 38108
rect 48116 38052 48172 38108
rect 48172 38052 48176 38108
rect 48112 38048 48176 38052
rect 48192 38108 48256 38112
rect 48192 38052 48196 38108
rect 48196 38052 48252 38108
rect 48252 38052 48256 38108
rect 48192 38048 48256 38052
rect 37596 37708 37660 37772
rect 2952 37564 3016 37568
rect 2952 37508 2956 37564
rect 2956 37508 3012 37564
rect 3012 37508 3016 37564
rect 2952 37504 3016 37508
rect 3032 37564 3096 37568
rect 3032 37508 3036 37564
rect 3036 37508 3092 37564
rect 3092 37508 3096 37564
rect 3032 37504 3096 37508
rect 3112 37564 3176 37568
rect 3112 37508 3116 37564
rect 3116 37508 3172 37564
rect 3172 37508 3176 37564
rect 3112 37504 3176 37508
rect 3192 37564 3256 37568
rect 3192 37508 3196 37564
rect 3196 37508 3252 37564
rect 3252 37508 3256 37564
rect 3192 37504 3256 37508
rect 12952 37564 13016 37568
rect 12952 37508 12956 37564
rect 12956 37508 13012 37564
rect 13012 37508 13016 37564
rect 12952 37504 13016 37508
rect 13032 37564 13096 37568
rect 13032 37508 13036 37564
rect 13036 37508 13092 37564
rect 13092 37508 13096 37564
rect 13032 37504 13096 37508
rect 13112 37564 13176 37568
rect 13112 37508 13116 37564
rect 13116 37508 13172 37564
rect 13172 37508 13176 37564
rect 13112 37504 13176 37508
rect 13192 37564 13256 37568
rect 13192 37508 13196 37564
rect 13196 37508 13252 37564
rect 13252 37508 13256 37564
rect 13192 37504 13256 37508
rect 22952 37564 23016 37568
rect 22952 37508 22956 37564
rect 22956 37508 23012 37564
rect 23012 37508 23016 37564
rect 22952 37504 23016 37508
rect 23032 37564 23096 37568
rect 23032 37508 23036 37564
rect 23036 37508 23092 37564
rect 23092 37508 23096 37564
rect 23032 37504 23096 37508
rect 23112 37564 23176 37568
rect 23112 37508 23116 37564
rect 23116 37508 23172 37564
rect 23172 37508 23176 37564
rect 23112 37504 23176 37508
rect 23192 37564 23256 37568
rect 23192 37508 23196 37564
rect 23196 37508 23252 37564
rect 23252 37508 23256 37564
rect 23192 37504 23256 37508
rect 32952 37564 33016 37568
rect 32952 37508 32956 37564
rect 32956 37508 33012 37564
rect 33012 37508 33016 37564
rect 32952 37504 33016 37508
rect 33032 37564 33096 37568
rect 33032 37508 33036 37564
rect 33036 37508 33092 37564
rect 33092 37508 33096 37564
rect 33032 37504 33096 37508
rect 33112 37564 33176 37568
rect 33112 37508 33116 37564
rect 33116 37508 33172 37564
rect 33172 37508 33176 37564
rect 33112 37504 33176 37508
rect 33192 37564 33256 37568
rect 33192 37508 33196 37564
rect 33196 37508 33252 37564
rect 33252 37508 33256 37564
rect 33192 37504 33256 37508
rect 42952 37564 43016 37568
rect 42952 37508 42956 37564
rect 42956 37508 43012 37564
rect 43012 37508 43016 37564
rect 42952 37504 43016 37508
rect 43032 37564 43096 37568
rect 43032 37508 43036 37564
rect 43036 37508 43092 37564
rect 43092 37508 43096 37564
rect 43032 37504 43096 37508
rect 43112 37564 43176 37568
rect 43112 37508 43116 37564
rect 43116 37508 43172 37564
rect 43172 37508 43176 37564
rect 43112 37504 43176 37508
rect 43192 37564 43256 37568
rect 43192 37508 43196 37564
rect 43196 37508 43252 37564
rect 43252 37508 43256 37564
rect 43192 37504 43256 37508
rect 7952 37020 8016 37024
rect 7952 36964 7956 37020
rect 7956 36964 8012 37020
rect 8012 36964 8016 37020
rect 7952 36960 8016 36964
rect 8032 37020 8096 37024
rect 8032 36964 8036 37020
rect 8036 36964 8092 37020
rect 8092 36964 8096 37020
rect 8032 36960 8096 36964
rect 8112 37020 8176 37024
rect 8112 36964 8116 37020
rect 8116 36964 8172 37020
rect 8172 36964 8176 37020
rect 8112 36960 8176 36964
rect 8192 37020 8256 37024
rect 8192 36964 8196 37020
rect 8196 36964 8252 37020
rect 8252 36964 8256 37020
rect 8192 36960 8256 36964
rect 17952 37020 18016 37024
rect 17952 36964 17956 37020
rect 17956 36964 18012 37020
rect 18012 36964 18016 37020
rect 17952 36960 18016 36964
rect 18032 37020 18096 37024
rect 18032 36964 18036 37020
rect 18036 36964 18092 37020
rect 18092 36964 18096 37020
rect 18032 36960 18096 36964
rect 18112 37020 18176 37024
rect 18112 36964 18116 37020
rect 18116 36964 18172 37020
rect 18172 36964 18176 37020
rect 18112 36960 18176 36964
rect 18192 37020 18256 37024
rect 18192 36964 18196 37020
rect 18196 36964 18252 37020
rect 18252 36964 18256 37020
rect 18192 36960 18256 36964
rect 27952 37020 28016 37024
rect 27952 36964 27956 37020
rect 27956 36964 28012 37020
rect 28012 36964 28016 37020
rect 27952 36960 28016 36964
rect 28032 37020 28096 37024
rect 28032 36964 28036 37020
rect 28036 36964 28092 37020
rect 28092 36964 28096 37020
rect 28032 36960 28096 36964
rect 28112 37020 28176 37024
rect 28112 36964 28116 37020
rect 28116 36964 28172 37020
rect 28172 36964 28176 37020
rect 28112 36960 28176 36964
rect 28192 37020 28256 37024
rect 28192 36964 28196 37020
rect 28196 36964 28252 37020
rect 28252 36964 28256 37020
rect 28192 36960 28256 36964
rect 37952 37020 38016 37024
rect 37952 36964 37956 37020
rect 37956 36964 38012 37020
rect 38012 36964 38016 37020
rect 37952 36960 38016 36964
rect 38032 37020 38096 37024
rect 38032 36964 38036 37020
rect 38036 36964 38092 37020
rect 38092 36964 38096 37020
rect 38032 36960 38096 36964
rect 38112 37020 38176 37024
rect 38112 36964 38116 37020
rect 38116 36964 38172 37020
rect 38172 36964 38176 37020
rect 38112 36960 38176 36964
rect 38192 37020 38256 37024
rect 38192 36964 38196 37020
rect 38196 36964 38252 37020
rect 38252 36964 38256 37020
rect 38192 36960 38256 36964
rect 47952 37020 48016 37024
rect 47952 36964 47956 37020
rect 47956 36964 48012 37020
rect 48012 36964 48016 37020
rect 47952 36960 48016 36964
rect 48032 37020 48096 37024
rect 48032 36964 48036 37020
rect 48036 36964 48092 37020
rect 48092 36964 48096 37020
rect 48032 36960 48096 36964
rect 48112 37020 48176 37024
rect 48112 36964 48116 37020
rect 48116 36964 48172 37020
rect 48172 36964 48176 37020
rect 48112 36960 48176 36964
rect 48192 37020 48256 37024
rect 48192 36964 48196 37020
rect 48196 36964 48252 37020
rect 48252 36964 48256 37020
rect 48192 36960 48256 36964
rect 37780 36756 37844 36820
rect 2952 36476 3016 36480
rect 2952 36420 2956 36476
rect 2956 36420 3012 36476
rect 3012 36420 3016 36476
rect 2952 36416 3016 36420
rect 3032 36476 3096 36480
rect 3032 36420 3036 36476
rect 3036 36420 3092 36476
rect 3092 36420 3096 36476
rect 3032 36416 3096 36420
rect 3112 36476 3176 36480
rect 3112 36420 3116 36476
rect 3116 36420 3172 36476
rect 3172 36420 3176 36476
rect 3112 36416 3176 36420
rect 3192 36476 3256 36480
rect 3192 36420 3196 36476
rect 3196 36420 3252 36476
rect 3252 36420 3256 36476
rect 3192 36416 3256 36420
rect 12952 36476 13016 36480
rect 12952 36420 12956 36476
rect 12956 36420 13012 36476
rect 13012 36420 13016 36476
rect 12952 36416 13016 36420
rect 13032 36476 13096 36480
rect 13032 36420 13036 36476
rect 13036 36420 13092 36476
rect 13092 36420 13096 36476
rect 13032 36416 13096 36420
rect 13112 36476 13176 36480
rect 13112 36420 13116 36476
rect 13116 36420 13172 36476
rect 13172 36420 13176 36476
rect 13112 36416 13176 36420
rect 13192 36476 13256 36480
rect 13192 36420 13196 36476
rect 13196 36420 13252 36476
rect 13252 36420 13256 36476
rect 13192 36416 13256 36420
rect 22952 36476 23016 36480
rect 22952 36420 22956 36476
rect 22956 36420 23012 36476
rect 23012 36420 23016 36476
rect 22952 36416 23016 36420
rect 23032 36476 23096 36480
rect 23032 36420 23036 36476
rect 23036 36420 23092 36476
rect 23092 36420 23096 36476
rect 23032 36416 23096 36420
rect 23112 36476 23176 36480
rect 23112 36420 23116 36476
rect 23116 36420 23172 36476
rect 23172 36420 23176 36476
rect 23112 36416 23176 36420
rect 23192 36476 23256 36480
rect 23192 36420 23196 36476
rect 23196 36420 23252 36476
rect 23252 36420 23256 36476
rect 23192 36416 23256 36420
rect 32952 36476 33016 36480
rect 32952 36420 32956 36476
rect 32956 36420 33012 36476
rect 33012 36420 33016 36476
rect 32952 36416 33016 36420
rect 33032 36476 33096 36480
rect 33032 36420 33036 36476
rect 33036 36420 33092 36476
rect 33092 36420 33096 36476
rect 33032 36416 33096 36420
rect 33112 36476 33176 36480
rect 33112 36420 33116 36476
rect 33116 36420 33172 36476
rect 33172 36420 33176 36476
rect 33112 36416 33176 36420
rect 33192 36476 33256 36480
rect 33192 36420 33196 36476
rect 33196 36420 33252 36476
rect 33252 36420 33256 36476
rect 33192 36416 33256 36420
rect 42952 36476 43016 36480
rect 42952 36420 42956 36476
rect 42956 36420 43012 36476
rect 43012 36420 43016 36476
rect 42952 36416 43016 36420
rect 43032 36476 43096 36480
rect 43032 36420 43036 36476
rect 43036 36420 43092 36476
rect 43092 36420 43096 36476
rect 43032 36416 43096 36420
rect 43112 36476 43176 36480
rect 43112 36420 43116 36476
rect 43116 36420 43172 36476
rect 43172 36420 43176 36476
rect 43112 36416 43176 36420
rect 43192 36476 43256 36480
rect 43192 36420 43196 36476
rect 43196 36420 43252 36476
rect 43252 36420 43256 36476
rect 43192 36416 43256 36420
rect 37780 36076 37844 36140
rect 25636 36000 25700 36004
rect 25636 35944 25650 36000
rect 25650 35944 25700 36000
rect 25636 35940 25700 35944
rect 7952 35932 8016 35936
rect 7952 35876 7956 35932
rect 7956 35876 8012 35932
rect 8012 35876 8016 35932
rect 7952 35872 8016 35876
rect 8032 35932 8096 35936
rect 8032 35876 8036 35932
rect 8036 35876 8092 35932
rect 8092 35876 8096 35932
rect 8032 35872 8096 35876
rect 8112 35932 8176 35936
rect 8112 35876 8116 35932
rect 8116 35876 8172 35932
rect 8172 35876 8176 35932
rect 8112 35872 8176 35876
rect 8192 35932 8256 35936
rect 8192 35876 8196 35932
rect 8196 35876 8252 35932
rect 8252 35876 8256 35932
rect 8192 35872 8256 35876
rect 17952 35932 18016 35936
rect 17952 35876 17956 35932
rect 17956 35876 18012 35932
rect 18012 35876 18016 35932
rect 17952 35872 18016 35876
rect 18032 35932 18096 35936
rect 18032 35876 18036 35932
rect 18036 35876 18092 35932
rect 18092 35876 18096 35932
rect 18032 35872 18096 35876
rect 18112 35932 18176 35936
rect 18112 35876 18116 35932
rect 18116 35876 18172 35932
rect 18172 35876 18176 35932
rect 18112 35872 18176 35876
rect 18192 35932 18256 35936
rect 18192 35876 18196 35932
rect 18196 35876 18252 35932
rect 18252 35876 18256 35932
rect 18192 35872 18256 35876
rect 27952 35932 28016 35936
rect 27952 35876 27956 35932
rect 27956 35876 28012 35932
rect 28012 35876 28016 35932
rect 27952 35872 28016 35876
rect 28032 35932 28096 35936
rect 28032 35876 28036 35932
rect 28036 35876 28092 35932
rect 28092 35876 28096 35932
rect 28032 35872 28096 35876
rect 28112 35932 28176 35936
rect 28112 35876 28116 35932
rect 28116 35876 28172 35932
rect 28172 35876 28176 35932
rect 28112 35872 28176 35876
rect 28192 35932 28256 35936
rect 28192 35876 28196 35932
rect 28196 35876 28252 35932
rect 28252 35876 28256 35932
rect 28192 35872 28256 35876
rect 37952 35932 38016 35936
rect 37952 35876 37956 35932
rect 37956 35876 38012 35932
rect 38012 35876 38016 35932
rect 37952 35872 38016 35876
rect 38032 35932 38096 35936
rect 38032 35876 38036 35932
rect 38036 35876 38092 35932
rect 38092 35876 38096 35932
rect 38032 35872 38096 35876
rect 38112 35932 38176 35936
rect 38112 35876 38116 35932
rect 38116 35876 38172 35932
rect 38172 35876 38176 35932
rect 38112 35872 38176 35876
rect 38192 35932 38256 35936
rect 38192 35876 38196 35932
rect 38196 35876 38252 35932
rect 38252 35876 38256 35932
rect 38192 35872 38256 35876
rect 47952 35932 48016 35936
rect 47952 35876 47956 35932
rect 47956 35876 48012 35932
rect 48012 35876 48016 35932
rect 47952 35872 48016 35876
rect 48032 35932 48096 35936
rect 48032 35876 48036 35932
rect 48036 35876 48092 35932
rect 48092 35876 48096 35932
rect 48032 35872 48096 35876
rect 48112 35932 48176 35936
rect 48112 35876 48116 35932
rect 48116 35876 48172 35932
rect 48172 35876 48176 35932
rect 48112 35872 48176 35876
rect 48192 35932 48256 35936
rect 48192 35876 48196 35932
rect 48196 35876 48252 35932
rect 48252 35876 48256 35932
rect 48192 35872 48256 35876
rect 41276 35804 41340 35868
rect 28764 35668 28828 35732
rect 2952 35388 3016 35392
rect 2952 35332 2956 35388
rect 2956 35332 3012 35388
rect 3012 35332 3016 35388
rect 2952 35328 3016 35332
rect 3032 35388 3096 35392
rect 3032 35332 3036 35388
rect 3036 35332 3092 35388
rect 3092 35332 3096 35388
rect 3032 35328 3096 35332
rect 3112 35388 3176 35392
rect 3112 35332 3116 35388
rect 3116 35332 3172 35388
rect 3172 35332 3176 35388
rect 3112 35328 3176 35332
rect 3192 35388 3256 35392
rect 3192 35332 3196 35388
rect 3196 35332 3252 35388
rect 3252 35332 3256 35388
rect 3192 35328 3256 35332
rect 12952 35388 13016 35392
rect 12952 35332 12956 35388
rect 12956 35332 13012 35388
rect 13012 35332 13016 35388
rect 12952 35328 13016 35332
rect 13032 35388 13096 35392
rect 13032 35332 13036 35388
rect 13036 35332 13092 35388
rect 13092 35332 13096 35388
rect 13032 35328 13096 35332
rect 13112 35388 13176 35392
rect 13112 35332 13116 35388
rect 13116 35332 13172 35388
rect 13172 35332 13176 35388
rect 13112 35328 13176 35332
rect 13192 35388 13256 35392
rect 13192 35332 13196 35388
rect 13196 35332 13252 35388
rect 13252 35332 13256 35388
rect 13192 35328 13256 35332
rect 22952 35388 23016 35392
rect 22952 35332 22956 35388
rect 22956 35332 23012 35388
rect 23012 35332 23016 35388
rect 22952 35328 23016 35332
rect 23032 35388 23096 35392
rect 23032 35332 23036 35388
rect 23036 35332 23092 35388
rect 23092 35332 23096 35388
rect 23032 35328 23096 35332
rect 23112 35388 23176 35392
rect 23112 35332 23116 35388
rect 23116 35332 23172 35388
rect 23172 35332 23176 35388
rect 23112 35328 23176 35332
rect 23192 35388 23256 35392
rect 23192 35332 23196 35388
rect 23196 35332 23252 35388
rect 23252 35332 23256 35388
rect 23192 35328 23256 35332
rect 32952 35388 33016 35392
rect 32952 35332 32956 35388
rect 32956 35332 33012 35388
rect 33012 35332 33016 35388
rect 32952 35328 33016 35332
rect 33032 35388 33096 35392
rect 33032 35332 33036 35388
rect 33036 35332 33092 35388
rect 33092 35332 33096 35388
rect 33032 35328 33096 35332
rect 33112 35388 33176 35392
rect 33112 35332 33116 35388
rect 33116 35332 33172 35388
rect 33172 35332 33176 35388
rect 33112 35328 33176 35332
rect 33192 35388 33256 35392
rect 33192 35332 33196 35388
rect 33196 35332 33252 35388
rect 33252 35332 33256 35388
rect 33192 35328 33256 35332
rect 42952 35388 43016 35392
rect 42952 35332 42956 35388
rect 42956 35332 43012 35388
rect 43012 35332 43016 35388
rect 42952 35328 43016 35332
rect 43032 35388 43096 35392
rect 43032 35332 43036 35388
rect 43036 35332 43092 35388
rect 43092 35332 43096 35388
rect 43032 35328 43096 35332
rect 43112 35388 43176 35392
rect 43112 35332 43116 35388
rect 43116 35332 43172 35388
rect 43172 35332 43176 35388
rect 43112 35328 43176 35332
rect 43192 35388 43256 35392
rect 43192 35332 43196 35388
rect 43196 35332 43252 35388
rect 43252 35332 43256 35388
rect 43192 35328 43256 35332
rect 28580 34988 28644 35052
rect 38884 34912 38948 34916
rect 38884 34856 38934 34912
rect 38934 34856 38948 34912
rect 38884 34852 38948 34856
rect 7952 34844 8016 34848
rect 7952 34788 7956 34844
rect 7956 34788 8012 34844
rect 8012 34788 8016 34844
rect 7952 34784 8016 34788
rect 8032 34844 8096 34848
rect 8032 34788 8036 34844
rect 8036 34788 8092 34844
rect 8092 34788 8096 34844
rect 8032 34784 8096 34788
rect 8112 34844 8176 34848
rect 8112 34788 8116 34844
rect 8116 34788 8172 34844
rect 8172 34788 8176 34844
rect 8112 34784 8176 34788
rect 8192 34844 8256 34848
rect 8192 34788 8196 34844
rect 8196 34788 8252 34844
rect 8252 34788 8256 34844
rect 8192 34784 8256 34788
rect 17952 34844 18016 34848
rect 17952 34788 17956 34844
rect 17956 34788 18012 34844
rect 18012 34788 18016 34844
rect 17952 34784 18016 34788
rect 18032 34844 18096 34848
rect 18032 34788 18036 34844
rect 18036 34788 18092 34844
rect 18092 34788 18096 34844
rect 18032 34784 18096 34788
rect 18112 34844 18176 34848
rect 18112 34788 18116 34844
rect 18116 34788 18172 34844
rect 18172 34788 18176 34844
rect 18112 34784 18176 34788
rect 18192 34844 18256 34848
rect 18192 34788 18196 34844
rect 18196 34788 18252 34844
rect 18252 34788 18256 34844
rect 18192 34784 18256 34788
rect 27952 34844 28016 34848
rect 27952 34788 27956 34844
rect 27956 34788 28012 34844
rect 28012 34788 28016 34844
rect 27952 34784 28016 34788
rect 28032 34844 28096 34848
rect 28032 34788 28036 34844
rect 28036 34788 28092 34844
rect 28092 34788 28096 34844
rect 28032 34784 28096 34788
rect 28112 34844 28176 34848
rect 28112 34788 28116 34844
rect 28116 34788 28172 34844
rect 28172 34788 28176 34844
rect 28112 34784 28176 34788
rect 28192 34844 28256 34848
rect 28192 34788 28196 34844
rect 28196 34788 28252 34844
rect 28252 34788 28256 34844
rect 28192 34784 28256 34788
rect 37952 34844 38016 34848
rect 37952 34788 37956 34844
rect 37956 34788 38012 34844
rect 38012 34788 38016 34844
rect 37952 34784 38016 34788
rect 38032 34844 38096 34848
rect 38032 34788 38036 34844
rect 38036 34788 38092 34844
rect 38092 34788 38096 34844
rect 38032 34784 38096 34788
rect 38112 34844 38176 34848
rect 38112 34788 38116 34844
rect 38116 34788 38172 34844
rect 38172 34788 38176 34844
rect 38112 34784 38176 34788
rect 38192 34844 38256 34848
rect 38192 34788 38196 34844
rect 38196 34788 38252 34844
rect 38252 34788 38256 34844
rect 38192 34784 38256 34788
rect 47952 34844 48016 34848
rect 47952 34788 47956 34844
rect 47956 34788 48012 34844
rect 48012 34788 48016 34844
rect 47952 34784 48016 34788
rect 48032 34844 48096 34848
rect 48032 34788 48036 34844
rect 48036 34788 48092 34844
rect 48092 34788 48096 34844
rect 48032 34784 48096 34788
rect 48112 34844 48176 34848
rect 48112 34788 48116 34844
rect 48116 34788 48172 34844
rect 48172 34788 48176 34844
rect 48112 34784 48176 34788
rect 48192 34844 48256 34848
rect 48192 34788 48196 34844
rect 48196 34788 48252 34844
rect 48252 34788 48256 34844
rect 48192 34784 48256 34788
rect 2952 34300 3016 34304
rect 2952 34244 2956 34300
rect 2956 34244 3012 34300
rect 3012 34244 3016 34300
rect 2952 34240 3016 34244
rect 3032 34300 3096 34304
rect 3032 34244 3036 34300
rect 3036 34244 3092 34300
rect 3092 34244 3096 34300
rect 3032 34240 3096 34244
rect 3112 34300 3176 34304
rect 3112 34244 3116 34300
rect 3116 34244 3172 34300
rect 3172 34244 3176 34300
rect 3112 34240 3176 34244
rect 3192 34300 3256 34304
rect 3192 34244 3196 34300
rect 3196 34244 3252 34300
rect 3252 34244 3256 34300
rect 3192 34240 3256 34244
rect 12952 34300 13016 34304
rect 12952 34244 12956 34300
rect 12956 34244 13012 34300
rect 13012 34244 13016 34300
rect 12952 34240 13016 34244
rect 13032 34300 13096 34304
rect 13032 34244 13036 34300
rect 13036 34244 13092 34300
rect 13092 34244 13096 34300
rect 13032 34240 13096 34244
rect 13112 34300 13176 34304
rect 13112 34244 13116 34300
rect 13116 34244 13172 34300
rect 13172 34244 13176 34300
rect 13112 34240 13176 34244
rect 13192 34300 13256 34304
rect 13192 34244 13196 34300
rect 13196 34244 13252 34300
rect 13252 34244 13256 34300
rect 13192 34240 13256 34244
rect 22952 34300 23016 34304
rect 22952 34244 22956 34300
rect 22956 34244 23012 34300
rect 23012 34244 23016 34300
rect 22952 34240 23016 34244
rect 23032 34300 23096 34304
rect 23032 34244 23036 34300
rect 23036 34244 23092 34300
rect 23092 34244 23096 34300
rect 23032 34240 23096 34244
rect 23112 34300 23176 34304
rect 23112 34244 23116 34300
rect 23116 34244 23172 34300
rect 23172 34244 23176 34300
rect 23112 34240 23176 34244
rect 23192 34300 23256 34304
rect 23192 34244 23196 34300
rect 23196 34244 23252 34300
rect 23252 34244 23256 34300
rect 23192 34240 23256 34244
rect 32952 34300 33016 34304
rect 32952 34244 32956 34300
rect 32956 34244 33012 34300
rect 33012 34244 33016 34300
rect 32952 34240 33016 34244
rect 33032 34300 33096 34304
rect 33032 34244 33036 34300
rect 33036 34244 33092 34300
rect 33092 34244 33096 34300
rect 33032 34240 33096 34244
rect 33112 34300 33176 34304
rect 33112 34244 33116 34300
rect 33116 34244 33172 34300
rect 33172 34244 33176 34300
rect 33112 34240 33176 34244
rect 33192 34300 33256 34304
rect 33192 34244 33196 34300
rect 33196 34244 33252 34300
rect 33252 34244 33256 34300
rect 33192 34240 33256 34244
rect 42952 34300 43016 34304
rect 42952 34244 42956 34300
rect 42956 34244 43012 34300
rect 43012 34244 43016 34300
rect 42952 34240 43016 34244
rect 43032 34300 43096 34304
rect 43032 34244 43036 34300
rect 43036 34244 43092 34300
rect 43092 34244 43096 34300
rect 43032 34240 43096 34244
rect 43112 34300 43176 34304
rect 43112 34244 43116 34300
rect 43116 34244 43172 34300
rect 43172 34244 43176 34300
rect 43112 34240 43176 34244
rect 43192 34300 43256 34304
rect 43192 34244 43196 34300
rect 43196 34244 43252 34300
rect 43252 34244 43256 34300
rect 43192 34240 43256 34244
rect 7952 33756 8016 33760
rect 7952 33700 7956 33756
rect 7956 33700 8012 33756
rect 8012 33700 8016 33756
rect 7952 33696 8016 33700
rect 8032 33756 8096 33760
rect 8032 33700 8036 33756
rect 8036 33700 8092 33756
rect 8092 33700 8096 33756
rect 8032 33696 8096 33700
rect 8112 33756 8176 33760
rect 8112 33700 8116 33756
rect 8116 33700 8172 33756
rect 8172 33700 8176 33756
rect 8112 33696 8176 33700
rect 8192 33756 8256 33760
rect 8192 33700 8196 33756
rect 8196 33700 8252 33756
rect 8252 33700 8256 33756
rect 8192 33696 8256 33700
rect 17952 33756 18016 33760
rect 17952 33700 17956 33756
rect 17956 33700 18012 33756
rect 18012 33700 18016 33756
rect 17952 33696 18016 33700
rect 18032 33756 18096 33760
rect 18032 33700 18036 33756
rect 18036 33700 18092 33756
rect 18092 33700 18096 33756
rect 18032 33696 18096 33700
rect 18112 33756 18176 33760
rect 18112 33700 18116 33756
rect 18116 33700 18172 33756
rect 18172 33700 18176 33756
rect 18112 33696 18176 33700
rect 18192 33756 18256 33760
rect 18192 33700 18196 33756
rect 18196 33700 18252 33756
rect 18252 33700 18256 33756
rect 18192 33696 18256 33700
rect 27952 33756 28016 33760
rect 27952 33700 27956 33756
rect 27956 33700 28012 33756
rect 28012 33700 28016 33756
rect 27952 33696 28016 33700
rect 28032 33756 28096 33760
rect 28032 33700 28036 33756
rect 28036 33700 28092 33756
rect 28092 33700 28096 33756
rect 28032 33696 28096 33700
rect 28112 33756 28176 33760
rect 28112 33700 28116 33756
rect 28116 33700 28172 33756
rect 28172 33700 28176 33756
rect 28112 33696 28176 33700
rect 28192 33756 28256 33760
rect 28192 33700 28196 33756
rect 28196 33700 28252 33756
rect 28252 33700 28256 33756
rect 28192 33696 28256 33700
rect 37952 33756 38016 33760
rect 37952 33700 37956 33756
rect 37956 33700 38012 33756
rect 38012 33700 38016 33756
rect 37952 33696 38016 33700
rect 38032 33756 38096 33760
rect 38032 33700 38036 33756
rect 38036 33700 38092 33756
rect 38092 33700 38096 33756
rect 38032 33696 38096 33700
rect 38112 33756 38176 33760
rect 38112 33700 38116 33756
rect 38116 33700 38172 33756
rect 38172 33700 38176 33756
rect 38112 33696 38176 33700
rect 38192 33756 38256 33760
rect 38192 33700 38196 33756
rect 38196 33700 38252 33756
rect 38252 33700 38256 33756
rect 38192 33696 38256 33700
rect 47952 33756 48016 33760
rect 47952 33700 47956 33756
rect 47956 33700 48012 33756
rect 48012 33700 48016 33756
rect 47952 33696 48016 33700
rect 48032 33756 48096 33760
rect 48032 33700 48036 33756
rect 48036 33700 48092 33756
rect 48092 33700 48096 33756
rect 48032 33696 48096 33700
rect 48112 33756 48176 33760
rect 48112 33700 48116 33756
rect 48116 33700 48172 33756
rect 48172 33700 48176 33756
rect 48112 33696 48176 33700
rect 48192 33756 48256 33760
rect 48192 33700 48196 33756
rect 48196 33700 48252 33756
rect 48252 33700 48256 33756
rect 48192 33696 48256 33700
rect 38884 33552 38948 33556
rect 38884 33496 38898 33552
rect 38898 33496 38948 33552
rect 38884 33492 38948 33496
rect 2952 33212 3016 33216
rect 2952 33156 2956 33212
rect 2956 33156 3012 33212
rect 3012 33156 3016 33212
rect 2952 33152 3016 33156
rect 3032 33212 3096 33216
rect 3032 33156 3036 33212
rect 3036 33156 3092 33212
rect 3092 33156 3096 33212
rect 3032 33152 3096 33156
rect 3112 33212 3176 33216
rect 3112 33156 3116 33212
rect 3116 33156 3172 33212
rect 3172 33156 3176 33212
rect 3112 33152 3176 33156
rect 3192 33212 3256 33216
rect 3192 33156 3196 33212
rect 3196 33156 3252 33212
rect 3252 33156 3256 33212
rect 3192 33152 3256 33156
rect 12952 33212 13016 33216
rect 12952 33156 12956 33212
rect 12956 33156 13012 33212
rect 13012 33156 13016 33212
rect 12952 33152 13016 33156
rect 13032 33212 13096 33216
rect 13032 33156 13036 33212
rect 13036 33156 13092 33212
rect 13092 33156 13096 33212
rect 13032 33152 13096 33156
rect 13112 33212 13176 33216
rect 13112 33156 13116 33212
rect 13116 33156 13172 33212
rect 13172 33156 13176 33212
rect 13112 33152 13176 33156
rect 13192 33212 13256 33216
rect 13192 33156 13196 33212
rect 13196 33156 13252 33212
rect 13252 33156 13256 33212
rect 13192 33152 13256 33156
rect 22952 33212 23016 33216
rect 22952 33156 22956 33212
rect 22956 33156 23012 33212
rect 23012 33156 23016 33212
rect 22952 33152 23016 33156
rect 23032 33212 23096 33216
rect 23032 33156 23036 33212
rect 23036 33156 23092 33212
rect 23092 33156 23096 33212
rect 23032 33152 23096 33156
rect 23112 33212 23176 33216
rect 23112 33156 23116 33212
rect 23116 33156 23172 33212
rect 23172 33156 23176 33212
rect 23112 33152 23176 33156
rect 23192 33212 23256 33216
rect 23192 33156 23196 33212
rect 23196 33156 23252 33212
rect 23252 33156 23256 33212
rect 23192 33152 23256 33156
rect 32952 33212 33016 33216
rect 32952 33156 32956 33212
rect 32956 33156 33012 33212
rect 33012 33156 33016 33212
rect 32952 33152 33016 33156
rect 33032 33212 33096 33216
rect 33032 33156 33036 33212
rect 33036 33156 33092 33212
rect 33092 33156 33096 33212
rect 33032 33152 33096 33156
rect 33112 33212 33176 33216
rect 33112 33156 33116 33212
rect 33116 33156 33172 33212
rect 33172 33156 33176 33212
rect 33112 33152 33176 33156
rect 33192 33212 33256 33216
rect 33192 33156 33196 33212
rect 33196 33156 33252 33212
rect 33252 33156 33256 33212
rect 33192 33152 33256 33156
rect 42952 33212 43016 33216
rect 42952 33156 42956 33212
rect 42956 33156 43012 33212
rect 43012 33156 43016 33212
rect 42952 33152 43016 33156
rect 43032 33212 43096 33216
rect 43032 33156 43036 33212
rect 43036 33156 43092 33212
rect 43092 33156 43096 33212
rect 43032 33152 43096 33156
rect 43112 33212 43176 33216
rect 43112 33156 43116 33212
rect 43116 33156 43172 33212
rect 43172 33156 43176 33212
rect 43112 33152 43176 33156
rect 43192 33212 43256 33216
rect 43192 33156 43196 33212
rect 43196 33156 43252 33212
rect 43252 33156 43256 33212
rect 43192 33152 43256 33156
rect 7952 32668 8016 32672
rect 7952 32612 7956 32668
rect 7956 32612 8012 32668
rect 8012 32612 8016 32668
rect 7952 32608 8016 32612
rect 8032 32668 8096 32672
rect 8032 32612 8036 32668
rect 8036 32612 8092 32668
rect 8092 32612 8096 32668
rect 8032 32608 8096 32612
rect 8112 32668 8176 32672
rect 8112 32612 8116 32668
rect 8116 32612 8172 32668
rect 8172 32612 8176 32668
rect 8112 32608 8176 32612
rect 8192 32668 8256 32672
rect 8192 32612 8196 32668
rect 8196 32612 8252 32668
rect 8252 32612 8256 32668
rect 8192 32608 8256 32612
rect 17952 32668 18016 32672
rect 17952 32612 17956 32668
rect 17956 32612 18012 32668
rect 18012 32612 18016 32668
rect 17952 32608 18016 32612
rect 18032 32668 18096 32672
rect 18032 32612 18036 32668
rect 18036 32612 18092 32668
rect 18092 32612 18096 32668
rect 18032 32608 18096 32612
rect 18112 32668 18176 32672
rect 18112 32612 18116 32668
rect 18116 32612 18172 32668
rect 18172 32612 18176 32668
rect 18112 32608 18176 32612
rect 18192 32668 18256 32672
rect 18192 32612 18196 32668
rect 18196 32612 18252 32668
rect 18252 32612 18256 32668
rect 18192 32608 18256 32612
rect 27952 32668 28016 32672
rect 27952 32612 27956 32668
rect 27956 32612 28012 32668
rect 28012 32612 28016 32668
rect 27952 32608 28016 32612
rect 28032 32668 28096 32672
rect 28032 32612 28036 32668
rect 28036 32612 28092 32668
rect 28092 32612 28096 32668
rect 28032 32608 28096 32612
rect 28112 32668 28176 32672
rect 28112 32612 28116 32668
rect 28116 32612 28172 32668
rect 28172 32612 28176 32668
rect 28112 32608 28176 32612
rect 28192 32668 28256 32672
rect 28192 32612 28196 32668
rect 28196 32612 28252 32668
rect 28252 32612 28256 32668
rect 28192 32608 28256 32612
rect 37952 32668 38016 32672
rect 37952 32612 37956 32668
rect 37956 32612 38012 32668
rect 38012 32612 38016 32668
rect 37952 32608 38016 32612
rect 38032 32668 38096 32672
rect 38032 32612 38036 32668
rect 38036 32612 38092 32668
rect 38092 32612 38096 32668
rect 38032 32608 38096 32612
rect 38112 32668 38176 32672
rect 38112 32612 38116 32668
rect 38116 32612 38172 32668
rect 38172 32612 38176 32668
rect 38112 32608 38176 32612
rect 38192 32668 38256 32672
rect 38192 32612 38196 32668
rect 38196 32612 38252 32668
rect 38252 32612 38256 32668
rect 38192 32608 38256 32612
rect 47952 32668 48016 32672
rect 47952 32612 47956 32668
rect 47956 32612 48012 32668
rect 48012 32612 48016 32668
rect 47952 32608 48016 32612
rect 48032 32668 48096 32672
rect 48032 32612 48036 32668
rect 48036 32612 48092 32668
rect 48092 32612 48096 32668
rect 48032 32608 48096 32612
rect 48112 32668 48176 32672
rect 48112 32612 48116 32668
rect 48116 32612 48172 32668
rect 48172 32612 48176 32668
rect 48112 32608 48176 32612
rect 48192 32668 48256 32672
rect 48192 32612 48196 32668
rect 48196 32612 48252 32668
rect 48252 32612 48256 32668
rect 48192 32608 48256 32612
rect 28580 32192 28644 32196
rect 28580 32136 28594 32192
rect 28594 32136 28644 32192
rect 28580 32132 28644 32136
rect 2952 32124 3016 32128
rect 2952 32068 2956 32124
rect 2956 32068 3012 32124
rect 3012 32068 3016 32124
rect 2952 32064 3016 32068
rect 3032 32124 3096 32128
rect 3032 32068 3036 32124
rect 3036 32068 3092 32124
rect 3092 32068 3096 32124
rect 3032 32064 3096 32068
rect 3112 32124 3176 32128
rect 3112 32068 3116 32124
rect 3116 32068 3172 32124
rect 3172 32068 3176 32124
rect 3112 32064 3176 32068
rect 3192 32124 3256 32128
rect 3192 32068 3196 32124
rect 3196 32068 3252 32124
rect 3252 32068 3256 32124
rect 3192 32064 3256 32068
rect 12952 32124 13016 32128
rect 12952 32068 12956 32124
rect 12956 32068 13012 32124
rect 13012 32068 13016 32124
rect 12952 32064 13016 32068
rect 13032 32124 13096 32128
rect 13032 32068 13036 32124
rect 13036 32068 13092 32124
rect 13092 32068 13096 32124
rect 13032 32064 13096 32068
rect 13112 32124 13176 32128
rect 13112 32068 13116 32124
rect 13116 32068 13172 32124
rect 13172 32068 13176 32124
rect 13112 32064 13176 32068
rect 13192 32124 13256 32128
rect 13192 32068 13196 32124
rect 13196 32068 13252 32124
rect 13252 32068 13256 32124
rect 13192 32064 13256 32068
rect 22952 32124 23016 32128
rect 22952 32068 22956 32124
rect 22956 32068 23012 32124
rect 23012 32068 23016 32124
rect 22952 32064 23016 32068
rect 23032 32124 23096 32128
rect 23032 32068 23036 32124
rect 23036 32068 23092 32124
rect 23092 32068 23096 32124
rect 23032 32064 23096 32068
rect 23112 32124 23176 32128
rect 23112 32068 23116 32124
rect 23116 32068 23172 32124
rect 23172 32068 23176 32124
rect 23112 32064 23176 32068
rect 23192 32124 23256 32128
rect 23192 32068 23196 32124
rect 23196 32068 23252 32124
rect 23252 32068 23256 32124
rect 23192 32064 23256 32068
rect 32952 32124 33016 32128
rect 32952 32068 32956 32124
rect 32956 32068 33012 32124
rect 33012 32068 33016 32124
rect 32952 32064 33016 32068
rect 33032 32124 33096 32128
rect 33032 32068 33036 32124
rect 33036 32068 33092 32124
rect 33092 32068 33096 32124
rect 33032 32064 33096 32068
rect 33112 32124 33176 32128
rect 33112 32068 33116 32124
rect 33116 32068 33172 32124
rect 33172 32068 33176 32124
rect 33112 32064 33176 32068
rect 33192 32124 33256 32128
rect 33192 32068 33196 32124
rect 33196 32068 33252 32124
rect 33252 32068 33256 32124
rect 33192 32064 33256 32068
rect 42952 32124 43016 32128
rect 42952 32068 42956 32124
rect 42956 32068 43012 32124
rect 43012 32068 43016 32124
rect 42952 32064 43016 32068
rect 43032 32124 43096 32128
rect 43032 32068 43036 32124
rect 43036 32068 43092 32124
rect 43092 32068 43096 32124
rect 43032 32064 43096 32068
rect 43112 32124 43176 32128
rect 43112 32068 43116 32124
rect 43116 32068 43172 32124
rect 43172 32068 43176 32124
rect 43112 32064 43176 32068
rect 43192 32124 43256 32128
rect 43192 32068 43196 32124
rect 43196 32068 43252 32124
rect 43252 32068 43256 32124
rect 43192 32064 43256 32068
rect 37412 31860 37476 31924
rect 7952 31580 8016 31584
rect 7952 31524 7956 31580
rect 7956 31524 8012 31580
rect 8012 31524 8016 31580
rect 7952 31520 8016 31524
rect 8032 31580 8096 31584
rect 8032 31524 8036 31580
rect 8036 31524 8092 31580
rect 8092 31524 8096 31580
rect 8032 31520 8096 31524
rect 8112 31580 8176 31584
rect 8112 31524 8116 31580
rect 8116 31524 8172 31580
rect 8172 31524 8176 31580
rect 8112 31520 8176 31524
rect 8192 31580 8256 31584
rect 8192 31524 8196 31580
rect 8196 31524 8252 31580
rect 8252 31524 8256 31580
rect 8192 31520 8256 31524
rect 17952 31580 18016 31584
rect 17952 31524 17956 31580
rect 17956 31524 18012 31580
rect 18012 31524 18016 31580
rect 17952 31520 18016 31524
rect 18032 31580 18096 31584
rect 18032 31524 18036 31580
rect 18036 31524 18092 31580
rect 18092 31524 18096 31580
rect 18032 31520 18096 31524
rect 18112 31580 18176 31584
rect 18112 31524 18116 31580
rect 18116 31524 18172 31580
rect 18172 31524 18176 31580
rect 18112 31520 18176 31524
rect 18192 31580 18256 31584
rect 18192 31524 18196 31580
rect 18196 31524 18252 31580
rect 18252 31524 18256 31580
rect 18192 31520 18256 31524
rect 27952 31580 28016 31584
rect 27952 31524 27956 31580
rect 27956 31524 28012 31580
rect 28012 31524 28016 31580
rect 27952 31520 28016 31524
rect 28032 31580 28096 31584
rect 28032 31524 28036 31580
rect 28036 31524 28092 31580
rect 28092 31524 28096 31580
rect 28032 31520 28096 31524
rect 28112 31580 28176 31584
rect 28112 31524 28116 31580
rect 28116 31524 28172 31580
rect 28172 31524 28176 31580
rect 28112 31520 28176 31524
rect 28192 31580 28256 31584
rect 28192 31524 28196 31580
rect 28196 31524 28252 31580
rect 28252 31524 28256 31580
rect 28192 31520 28256 31524
rect 37952 31580 38016 31584
rect 37952 31524 37956 31580
rect 37956 31524 38012 31580
rect 38012 31524 38016 31580
rect 37952 31520 38016 31524
rect 38032 31580 38096 31584
rect 38032 31524 38036 31580
rect 38036 31524 38092 31580
rect 38092 31524 38096 31580
rect 38032 31520 38096 31524
rect 38112 31580 38176 31584
rect 38112 31524 38116 31580
rect 38116 31524 38172 31580
rect 38172 31524 38176 31580
rect 38112 31520 38176 31524
rect 38192 31580 38256 31584
rect 38192 31524 38196 31580
rect 38196 31524 38252 31580
rect 38252 31524 38256 31580
rect 38192 31520 38256 31524
rect 47952 31580 48016 31584
rect 47952 31524 47956 31580
rect 47956 31524 48012 31580
rect 48012 31524 48016 31580
rect 47952 31520 48016 31524
rect 48032 31580 48096 31584
rect 48032 31524 48036 31580
rect 48036 31524 48092 31580
rect 48092 31524 48096 31580
rect 48032 31520 48096 31524
rect 48112 31580 48176 31584
rect 48112 31524 48116 31580
rect 48116 31524 48172 31580
rect 48172 31524 48176 31580
rect 48112 31520 48176 31524
rect 48192 31580 48256 31584
rect 48192 31524 48196 31580
rect 48196 31524 48252 31580
rect 48252 31524 48256 31580
rect 48192 31520 48256 31524
rect 22508 31240 22572 31244
rect 22508 31184 22522 31240
rect 22522 31184 22572 31240
rect 22508 31180 22572 31184
rect 2952 31036 3016 31040
rect 2952 30980 2956 31036
rect 2956 30980 3012 31036
rect 3012 30980 3016 31036
rect 2952 30976 3016 30980
rect 3032 31036 3096 31040
rect 3032 30980 3036 31036
rect 3036 30980 3092 31036
rect 3092 30980 3096 31036
rect 3032 30976 3096 30980
rect 3112 31036 3176 31040
rect 3112 30980 3116 31036
rect 3116 30980 3172 31036
rect 3172 30980 3176 31036
rect 3112 30976 3176 30980
rect 3192 31036 3256 31040
rect 3192 30980 3196 31036
rect 3196 30980 3252 31036
rect 3252 30980 3256 31036
rect 3192 30976 3256 30980
rect 12952 31036 13016 31040
rect 12952 30980 12956 31036
rect 12956 30980 13012 31036
rect 13012 30980 13016 31036
rect 12952 30976 13016 30980
rect 13032 31036 13096 31040
rect 13032 30980 13036 31036
rect 13036 30980 13092 31036
rect 13092 30980 13096 31036
rect 13032 30976 13096 30980
rect 13112 31036 13176 31040
rect 13112 30980 13116 31036
rect 13116 30980 13172 31036
rect 13172 30980 13176 31036
rect 13112 30976 13176 30980
rect 13192 31036 13256 31040
rect 13192 30980 13196 31036
rect 13196 30980 13252 31036
rect 13252 30980 13256 31036
rect 13192 30976 13256 30980
rect 22952 31036 23016 31040
rect 22952 30980 22956 31036
rect 22956 30980 23012 31036
rect 23012 30980 23016 31036
rect 22952 30976 23016 30980
rect 23032 31036 23096 31040
rect 23032 30980 23036 31036
rect 23036 30980 23092 31036
rect 23092 30980 23096 31036
rect 23032 30976 23096 30980
rect 23112 31036 23176 31040
rect 23112 30980 23116 31036
rect 23116 30980 23172 31036
rect 23172 30980 23176 31036
rect 23112 30976 23176 30980
rect 23192 31036 23256 31040
rect 23192 30980 23196 31036
rect 23196 30980 23252 31036
rect 23252 30980 23256 31036
rect 23192 30976 23256 30980
rect 32952 31036 33016 31040
rect 32952 30980 32956 31036
rect 32956 30980 33012 31036
rect 33012 30980 33016 31036
rect 32952 30976 33016 30980
rect 33032 31036 33096 31040
rect 33032 30980 33036 31036
rect 33036 30980 33092 31036
rect 33092 30980 33096 31036
rect 33032 30976 33096 30980
rect 33112 31036 33176 31040
rect 33112 30980 33116 31036
rect 33116 30980 33172 31036
rect 33172 30980 33176 31036
rect 33112 30976 33176 30980
rect 33192 31036 33256 31040
rect 33192 30980 33196 31036
rect 33196 30980 33252 31036
rect 33252 30980 33256 31036
rect 33192 30976 33256 30980
rect 42952 31036 43016 31040
rect 42952 30980 42956 31036
rect 42956 30980 43012 31036
rect 43012 30980 43016 31036
rect 42952 30976 43016 30980
rect 43032 31036 43096 31040
rect 43032 30980 43036 31036
rect 43036 30980 43092 31036
rect 43092 30980 43096 31036
rect 43032 30976 43096 30980
rect 43112 31036 43176 31040
rect 43112 30980 43116 31036
rect 43116 30980 43172 31036
rect 43172 30980 43176 31036
rect 43112 30976 43176 30980
rect 43192 31036 43256 31040
rect 43192 30980 43196 31036
rect 43196 30980 43252 31036
rect 43252 30980 43256 31036
rect 43192 30976 43256 30980
rect 7952 30492 8016 30496
rect 7952 30436 7956 30492
rect 7956 30436 8012 30492
rect 8012 30436 8016 30492
rect 7952 30432 8016 30436
rect 8032 30492 8096 30496
rect 8032 30436 8036 30492
rect 8036 30436 8092 30492
rect 8092 30436 8096 30492
rect 8032 30432 8096 30436
rect 8112 30492 8176 30496
rect 8112 30436 8116 30492
rect 8116 30436 8172 30492
rect 8172 30436 8176 30492
rect 8112 30432 8176 30436
rect 8192 30492 8256 30496
rect 8192 30436 8196 30492
rect 8196 30436 8252 30492
rect 8252 30436 8256 30492
rect 8192 30432 8256 30436
rect 17952 30492 18016 30496
rect 17952 30436 17956 30492
rect 17956 30436 18012 30492
rect 18012 30436 18016 30492
rect 17952 30432 18016 30436
rect 18032 30492 18096 30496
rect 18032 30436 18036 30492
rect 18036 30436 18092 30492
rect 18092 30436 18096 30492
rect 18032 30432 18096 30436
rect 18112 30492 18176 30496
rect 18112 30436 18116 30492
rect 18116 30436 18172 30492
rect 18172 30436 18176 30492
rect 18112 30432 18176 30436
rect 18192 30492 18256 30496
rect 18192 30436 18196 30492
rect 18196 30436 18252 30492
rect 18252 30436 18256 30492
rect 18192 30432 18256 30436
rect 25084 30364 25148 30428
rect 27952 30492 28016 30496
rect 27952 30436 27956 30492
rect 27956 30436 28012 30492
rect 28012 30436 28016 30492
rect 27952 30432 28016 30436
rect 28032 30492 28096 30496
rect 28032 30436 28036 30492
rect 28036 30436 28092 30492
rect 28092 30436 28096 30492
rect 28032 30432 28096 30436
rect 28112 30492 28176 30496
rect 28112 30436 28116 30492
rect 28116 30436 28172 30492
rect 28172 30436 28176 30492
rect 28112 30432 28176 30436
rect 28192 30492 28256 30496
rect 28192 30436 28196 30492
rect 28196 30436 28252 30492
rect 28252 30436 28256 30492
rect 28192 30432 28256 30436
rect 37952 30492 38016 30496
rect 37952 30436 37956 30492
rect 37956 30436 38012 30492
rect 38012 30436 38016 30492
rect 37952 30432 38016 30436
rect 38032 30492 38096 30496
rect 38032 30436 38036 30492
rect 38036 30436 38092 30492
rect 38092 30436 38096 30492
rect 38032 30432 38096 30436
rect 38112 30492 38176 30496
rect 38112 30436 38116 30492
rect 38116 30436 38172 30492
rect 38172 30436 38176 30492
rect 38112 30432 38176 30436
rect 38192 30492 38256 30496
rect 38192 30436 38196 30492
rect 38196 30436 38252 30492
rect 38252 30436 38256 30492
rect 38192 30432 38256 30436
rect 47952 30492 48016 30496
rect 47952 30436 47956 30492
rect 47956 30436 48012 30492
rect 48012 30436 48016 30492
rect 47952 30432 48016 30436
rect 48032 30492 48096 30496
rect 48032 30436 48036 30492
rect 48036 30436 48092 30492
rect 48092 30436 48096 30492
rect 48032 30432 48096 30436
rect 48112 30492 48176 30496
rect 48112 30436 48116 30492
rect 48116 30436 48172 30492
rect 48172 30436 48176 30492
rect 48112 30432 48176 30436
rect 48192 30492 48256 30496
rect 48192 30436 48196 30492
rect 48196 30436 48252 30492
rect 48252 30436 48256 30492
rect 48192 30432 48256 30436
rect 37780 30228 37844 30292
rect 28764 30092 28828 30156
rect 30788 30092 30852 30156
rect 2952 29948 3016 29952
rect 2952 29892 2956 29948
rect 2956 29892 3012 29948
rect 3012 29892 3016 29948
rect 2952 29888 3016 29892
rect 3032 29948 3096 29952
rect 3032 29892 3036 29948
rect 3036 29892 3092 29948
rect 3092 29892 3096 29948
rect 3032 29888 3096 29892
rect 3112 29948 3176 29952
rect 3112 29892 3116 29948
rect 3116 29892 3172 29948
rect 3172 29892 3176 29948
rect 3112 29888 3176 29892
rect 3192 29948 3256 29952
rect 3192 29892 3196 29948
rect 3196 29892 3252 29948
rect 3252 29892 3256 29948
rect 3192 29888 3256 29892
rect 12952 29948 13016 29952
rect 12952 29892 12956 29948
rect 12956 29892 13012 29948
rect 13012 29892 13016 29948
rect 12952 29888 13016 29892
rect 13032 29948 13096 29952
rect 13032 29892 13036 29948
rect 13036 29892 13092 29948
rect 13092 29892 13096 29948
rect 13032 29888 13096 29892
rect 13112 29948 13176 29952
rect 13112 29892 13116 29948
rect 13116 29892 13172 29948
rect 13172 29892 13176 29948
rect 13112 29888 13176 29892
rect 13192 29948 13256 29952
rect 13192 29892 13196 29948
rect 13196 29892 13252 29948
rect 13252 29892 13256 29948
rect 13192 29888 13256 29892
rect 22952 29948 23016 29952
rect 22952 29892 22956 29948
rect 22956 29892 23012 29948
rect 23012 29892 23016 29948
rect 22952 29888 23016 29892
rect 23032 29948 23096 29952
rect 23032 29892 23036 29948
rect 23036 29892 23092 29948
rect 23092 29892 23096 29948
rect 23032 29888 23096 29892
rect 23112 29948 23176 29952
rect 23112 29892 23116 29948
rect 23116 29892 23172 29948
rect 23172 29892 23176 29948
rect 23112 29888 23176 29892
rect 23192 29948 23256 29952
rect 23192 29892 23196 29948
rect 23196 29892 23252 29948
rect 23252 29892 23256 29948
rect 23192 29888 23256 29892
rect 32952 29948 33016 29952
rect 32952 29892 32956 29948
rect 32956 29892 33012 29948
rect 33012 29892 33016 29948
rect 32952 29888 33016 29892
rect 33032 29948 33096 29952
rect 33032 29892 33036 29948
rect 33036 29892 33092 29948
rect 33092 29892 33096 29948
rect 33032 29888 33096 29892
rect 33112 29948 33176 29952
rect 33112 29892 33116 29948
rect 33116 29892 33172 29948
rect 33172 29892 33176 29948
rect 33112 29888 33176 29892
rect 33192 29948 33256 29952
rect 33192 29892 33196 29948
rect 33196 29892 33252 29948
rect 33252 29892 33256 29948
rect 33192 29888 33256 29892
rect 42952 29948 43016 29952
rect 42952 29892 42956 29948
rect 42956 29892 43012 29948
rect 43012 29892 43016 29948
rect 42952 29888 43016 29892
rect 43032 29948 43096 29952
rect 43032 29892 43036 29948
rect 43036 29892 43092 29948
rect 43092 29892 43096 29948
rect 43032 29888 43096 29892
rect 43112 29948 43176 29952
rect 43112 29892 43116 29948
rect 43116 29892 43172 29948
rect 43172 29892 43176 29948
rect 43112 29888 43176 29892
rect 43192 29948 43256 29952
rect 43192 29892 43196 29948
rect 43196 29892 43252 29948
rect 43252 29892 43256 29948
rect 43192 29888 43256 29892
rect 7952 29404 8016 29408
rect 7952 29348 7956 29404
rect 7956 29348 8012 29404
rect 8012 29348 8016 29404
rect 7952 29344 8016 29348
rect 8032 29404 8096 29408
rect 8032 29348 8036 29404
rect 8036 29348 8092 29404
rect 8092 29348 8096 29404
rect 8032 29344 8096 29348
rect 8112 29404 8176 29408
rect 8112 29348 8116 29404
rect 8116 29348 8172 29404
rect 8172 29348 8176 29404
rect 8112 29344 8176 29348
rect 8192 29404 8256 29408
rect 8192 29348 8196 29404
rect 8196 29348 8252 29404
rect 8252 29348 8256 29404
rect 8192 29344 8256 29348
rect 17952 29404 18016 29408
rect 17952 29348 17956 29404
rect 17956 29348 18012 29404
rect 18012 29348 18016 29404
rect 17952 29344 18016 29348
rect 18032 29404 18096 29408
rect 18032 29348 18036 29404
rect 18036 29348 18092 29404
rect 18092 29348 18096 29404
rect 18032 29344 18096 29348
rect 18112 29404 18176 29408
rect 18112 29348 18116 29404
rect 18116 29348 18172 29404
rect 18172 29348 18176 29404
rect 18112 29344 18176 29348
rect 18192 29404 18256 29408
rect 18192 29348 18196 29404
rect 18196 29348 18252 29404
rect 18252 29348 18256 29404
rect 18192 29344 18256 29348
rect 27952 29404 28016 29408
rect 27952 29348 27956 29404
rect 27956 29348 28012 29404
rect 28012 29348 28016 29404
rect 27952 29344 28016 29348
rect 28032 29404 28096 29408
rect 28032 29348 28036 29404
rect 28036 29348 28092 29404
rect 28092 29348 28096 29404
rect 28032 29344 28096 29348
rect 28112 29404 28176 29408
rect 28112 29348 28116 29404
rect 28116 29348 28172 29404
rect 28172 29348 28176 29404
rect 28112 29344 28176 29348
rect 28192 29404 28256 29408
rect 28192 29348 28196 29404
rect 28196 29348 28252 29404
rect 28252 29348 28256 29404
rect 28192 29344 28256 29348
rect 37952 29404 38016 29408
rect 37952 29348 37956 29404
rect 37956 29348 38012 29404
rect 38012 29348 38016 29404
rect 37952 29344 38016 29348
rect 38032 29404 38096 29408
rect 38032 29348 38036 29404
rect 38036 29348 38092 29404
rect 38092 29348 38096 29404
rect 38032 29344 38096 29348
rect 38112 29404 38176 29408
rect 38112 29348 38116 29404
rect 38116 29348 38172 29404
rect 38172 29348 38176 29404
rect 38112 29344 38176 29348
rect 38192 29404 38256 29408
rect 38192 29348 38196 29404
rect 38196 29348 38252 29404
rect 38252 29348 38256 29404
rect 38192 29344 38256 29348
rect 47952 29404 48016 29408
rect 47952 29348 47956 29404
rect 47956 29348 48012 29404
rect 48012 29348 48016 29404
rect 47952 29344 48016 29348
rect 48032 29404 48096 29408
rect 48032 29348 48036 29404
rect 48036 29348 48092 29404
rect 48092 29348 48096 29404
rect 48032 29344 48096 29348
rect 48112 29404 48176 29408
rect 48112 29348 48116 29404
rect 48116 29348 48172 29404
rect 48172 29348 48176 29404
rect 48112 29344 48176 29348
rect 48192 29404 48256 29408
rect 48192 29348 48196 29404
rect 48196 29348 48252 29404
rect 48252 29348 48256 29404
rect 48192 29344 48256 29348
rect 37596 29004 37660 29068
rect 2952 28860 3016 28864
rect 2952 28804 2956 28860
rect 2956 28804 3012 28860
rect 3012 28804 3016 28860
rect 2952 28800 3016 28804
rect 3032 28860 3096 28864
rect 3032 28804 3036 28860
rect 3036 28804 3092 28860
rect 3092 28804 3096 28860
rect 3032 28800 3096 28804
rect 3112 28860 3176 28864
rect 3112 28804 3116 28860
rect 3116 28804 3172 28860
rect 3172 28804 3176 28860
rect 3112 28800 3176 28804
rect 3192 28860 3256 28864
rect 3192 28804 3196 28860
rect 3196 28804 3252 28860
rect 3252 28804 3256 28860
rect 3192 28800 3256 28804
rect 12952 28860 13016 28864
rect 12952 28804 12956 28860
rect 12956 28804 13012 28860
rect 13012 28804 13016 28860
rect 12952 28800 13016 28804
rect 13032 28860 13096 28864
rect 13032 28804 13036 28860
rect 13036 28804 13092 28860
rect 13092 28804 13096 28860
rect 13032 28800 13096 28804
rect 13112 28860 13176 28864
rect 13112 28804 13116 28860
rect 13116 28804 13172 28860
rect 13172 28804 13176 28860
rect 13112 28800 13176 28804
rect 13192 28860 13256 28864
rect 13192 28804 13196 28860
rect 13196 28804 13252 28860
rect 13252 28804 13256 28860
rect 13192 28800 13256 28804
rect 22952 28860 23016 28864
rect 22952 28804 22956 28860
rect 22956 28804 23012 28860
rect 23012 28804 23016 28860
rect 22952 28800 23016 28804
rect 23032 28860 23096 28864
rect 23032 28804 23036 28860
rect 23036 28804 23092 28860
rect 23092 28804 23096 28860
rect 23032 28800 23096 28804
rect 23112 28860 23176 28864
rect 23112 28804 23116 28860
rect 23116 28804 23172 28860
rect 23172 28804 23176 28860
rect 23112 28800 23176 28804
rect 23192 28860 23256 28864
rect 23192 28804 23196 28860
rect 23196 28804 23252 28860
rect 23252 28804 23256 28860
rect 23192 28800 23256 28804
rect 32952 28860 33016 28864
rect 32952 28804 32956 28860
rect 32956 28804 33012 28860
rect 33012 28804 33016 28860
rect 32952 28800 33016 28804
rect 33032 28860 33096 28864
rect 33032 28804 33036 28860
rect 33036 28804 33092 28860
rect 33092 28804 33096 28860
rect 33032 28800 33096 28804
rect 33112 28860 33176 28864
rect 33112 28804 33116 28860
rect 33116 28804 33172 28860
rect 33172 28804 33176 28860
rect 33112 28800 33176 28804
rect 33192 28860 33256 28864
rect 33192 28804 33196 28860
rect 33196 28804 33252 28860
rect 33252 28804 33256 28860
rect 33192 28800 33256 28804
rect 42952 28860 43016 28864
rect 42952 28804 42956 28860
rect 42956 28804 43012 28860
rect 43012 28804 43016 28860
rect 42952 28800 43016 28804
rect 43032 28860 43096 28864
rect 43032 28804 43036 28860
rect 43036 28804 43092 28860
rect 43092 28804 43096 28860
rect 43032 28800 43096 28804
rect 43112 28860 43176 28864
rect 43112 28804 43116 28860
rect 43116 28804 43172 28860
rect 43172 28804 43176 28860
rect 43112 28800 43176 28804
rect 43192 28860 43256 28864
rect 43192 28804 43196 28860
rect 43196 28804 43252 28860
rect 43252 28804 43256 28860
rect 43192 28800 43256 28804
rect 40540 28460 40604 28524
rect 35204 28324 35268 28388
rect 7952 28316 8016 28320
rect 7952 28260 7956 28316
rect 7956 28260 8012 28316
rect 8012 28260 8016 28316
rect 7952 28256 8016 28260
rect 8032 28316 8096 28320
rect 8032 28260 8036 28316
rect 8036 28260 8092 28316
rect 8092 28260 8096 28316
rect 8032 28256 8096 28260
rect 8112 28316 8176 28320
rect 8112 28260 8116 28316
rect 8116 28260 8172 28316
rect 8172 28260 8176 28316
rect 8112 28256 8176 28260
rect 8192 28316 8256 28320
rect 8192 28260 8196 28316
rect 8196 28260 8252 28316
rect 8252 28260 8256 28316
rect 8192 28256 8256 28260
rect 17952 28316 18016 28320
rect 17952 28260 17956 28316
rect 17956 28260 18012 28316
rect 18012 28260 18016 28316
rect 17952 28256 18016 28260
rect 18032 28316 18096 28320
rect 18032 28260 18036 28316
rect 18036 28260 18092 28316
rect 18092 28260 18096 28316
rect 18032 28256 18096 28260
rect 18112 28316 18176 28320
rect 18112 28260 18116 28316
rect 18116 28260 18172 28316
rect 18172 28260 18176 28316
rect 18112 28256 18176 28260
rect 18192 28316 18256 28320
rect 18192 28260 18196 28316
rect 18196 28260 18252 28316
rect 18252 28260 18256 28316
rect 18192 28256 18256 28260
rect 27952 28316 28016 28320
rect 27952 28260 27956 28316
rect 27956 28260 28012 28316
rect 28012 28260 28016 28316
rect 27952 28256 28016 28260
rect 28032 28316 28096 28320
rect 28032 28260 28036 28316
rect 28036 28260 28092 28316
rect 28092 28260 28096 28316
rect 28032 28256 28096 28260
rect 28112 28316 28176 28320
rect 28112 28260 28116 28316
rect 28116 28260 28172 28316
rect 28172 28260 28176 28316
rect 28112 28256 28176 28260
rect 28192 28316 28256 28320
rect 28192 28260 28196 28316
rect 28196 28260 28252 28316
rect 28252 28260 28256 28316
rect 28192 28256 28256 28260
rect 37952 28316 38016 28320
rect 37952 28260 37956 28316
rect 37956 28260 38012 28316
rect 38012 28260 38016 28316
rect 37952 28256 38016 28260
rect 38032 28316 38096 28320
rect 38032 28260 38036 28316
rect 38036 28260 38092 28316
rect 38092 28260 38096 28316
rect 38032 28256 38096 28260
rect 38112 28316 38176 28320
rect 38112 28260 38116 28316
rect 38116 28260 38172 28316
rect 38172 28260 38176 28316
rect 38112 28256 38176 28260
rect 38192 28316 38256 28320
rect 38192 28260 38196 28316
rect 38196 28260 38252 28316
rect 38252 28260 38256 28316
rect 38192 28256 38256 28260
rect 47952 28316 48016 28320
rect 47952 28260 47956 28316
rect 47956 28260 48012 28316
rect 48012 28260 48016 28316
rect 47952 28256 48016 28260
rect 48032 28316 48096 28320
rect 48032 28260 48036 28316
rect 48036 28260 48092 28316
rect 48092 28260 48096 28316
rect 48032 28256 48096 28260
rect 48112 28316 48176 28320
rect 48112 28260 48116 28316
rect 48116 28260 48172 28316
rect 48172 28260 48176 28316
rect 48112 28256 48176 28260
rect 48192 28316 48256 28320
rect 48192 28260 48196 28316
rect 48196 28260 48252 28316
rect 48252 28260 48256 28316
rect 48192 28256 48256 28260
rect 27660 28248 27724 28252
rect 27660 28192 27710 28248
rect 27710 28192 27724 28248
rect 27660 28188 27724 28192
rect 2952 27772 3016 27776
rect 2952 27716 2956 27772
rect 2956 27716 3012 27772
rect 3012 27716 3016 27772
rect 2952 27712 3016 27716
rect 3032 27772 3096 27776
rect 3032 27716 3036 27772
rect 3036 27716 3092 27772
rect 3092 27716 3096 27772
rect 3032 27712 3096 27716
rect 3112 27772 3176 27776
rect 3112 27716 3116 27772
rect 3116 27716 3172 27772
rect 3172 27716 3176 27772
rect 3112 27712 3176 27716
rect 3192 27772 3256 27776
rect 3192 27716 3196 27772
rect 3196 27716 3252 27772
rect 3252 27716 3256 27772
rect 3192 27712 3256 27716
rect 12952 27772 13016 27776
rect 12952 27716 12956 27772
rect 12956 27716 13012 27772
rect 13012 27716 13016 27772
rect 12952 27712 13016 27716
rect 13032 27772 13096 27776
rect 13032 27716 13036 27772
rect 13036 27716 13092 27772
rect 13092 27716 13096 27772
rect 13032 27712 13096 27716
rect 13112 27772 13176 27776
rect 13112 27716 13116 27772
rect 13116 27716 13172 27772
rect 13172 27716 13176 27772
rect 13112 27712 13176 27716
rect 13192 27772 13256 27776
rect 13192 27716 13196 27772
rect 13196 27716 13252 27772
rect 13252 27716 13256 27772
rect 13192 27712 13256 27716
rect 22952 27772 23016 27776
rect 22952 27716 22956 27772
rect 22956 27716 23012 27772
rect 23012 27716 23016 27772
rect 22952 27712 23016 27716
rect 23032 27772 23096 27776
rect 23032 27716 23036 27772
rect 23036 27716 23092 27772
rect 23092 27716 23096 27772
rect 23032 27712 23096 27716
rect 23112 27772 23176 27776
rect 23112 27716 23116 27772
rect 23116 27716 23172 27772
rect 23172 27716 23176 27772
rect 23112 27712 23176 27716
rect 23192 27772 23256 27776
rect 23192 27716 23196 27772
rect 23196 27716 23252 27772
rect 23252 27716 23256 27772
rect 23192 27712 23256 27716
rect 32952 27772 33016 27776
rect 32952 27716 32956 27772
rect 32956 27716 33012 27772
rect 33012 27716 33016 27772
rect 32952 27712 33016 27716
rect 33032 27772 33096 27776
rect 33032 27716 33036 27772
rect 33036 27716 33092 27772
rect 33092 27716 33096 27772
rect 33032 27712 33096 27716
rect 33112 27772 33176 27776
rect 33112 27716 33116 27772
rect 33116 27716 33172 27772
rect 33172 27716 33176 27772
rect 33112 27712 33176 27716
rect 33192 27772 33256 27776
rect 33192 27716 33196 27772
rect 33196 27716 33252 27772
rect 33252 27716 33256 27772
rect 33192 27712 33256 27716
rect 42952 27772 43016 27776
rect 42952 27716 42956 27772
rect 42956 27716 43012 27772
rect 43012 27716 43016 27772
rect 42952 27712 43016 27716
rect 43032 27772 43096 27776
rect 43032 27716 43036 27772
rect 43036 27716 43092 27772
rect 43092 27716 43096 27772
rect 43032 27712 43096 27716
rect 43112 27772 43176 27776
rect 43112 27716 43116 27772
rect 43116 27716 43172 27772
rect 43172 27716 43176 27772
rect 43112 27712 43176 27716
rect 43192 27772 43256 27776
rect 43192 27716 43196 27772
rect 43196 27716 43252 27772
rect 43252 27716 43256 27772
rect 43192 27712 43256 27716
rect 27108 27704 27172 27708
rect 27108 27648 27122 27704
rect 27122 27648 27172 27704
rect 27108 27644 27172 27648
rect 30420 27236 30484 27300
rect 7952 27228 8016 27232
rect 7952 27172 7956 27228
rect 7956 27172 8012 27228
rect 8012 27172 8016 27228
rect 7952 27168 8016 27172
rect 8032 27228 8096 27232
rect 8032 27172 8036 27228
rect 8036 27172 8092 27228
rect 8092 27172 8096 27228
rect 8032 27168 8096 27172
rect 8112 27228 8176 27232
rect 8112 27172 8116 27228
rect 8116 27172 8172 27228
rect 8172 27172 8176 27228
rect 8112 27168 8176 27172
rect 8192 27228 8256 27232
rect 8192 27172 8196 27228
rect 8196 27172 8252 27228
rect 8252 27172 8256 27228
rect 8192 27168 8256 27172
rect 17952 27228 18016 27232
rect 17952 27172 17956 27228
rect 17956 27172 18012 27228
rect 18012 27172 18016 27228
rect 17952 27168 18016 27172
rect 18032 27228 18096 27232
rect 18032 27172 18036 27228
rect 18036 27172 18092 27228
rect 18092 27172 18096 27228
rect 18032 27168 18096 27172
rect 18112 27228 18176 27232
rect 18112 27172 18116 27228
rect 18116 27172 18172 27228
rect 18172 27172 18176 27228
rect 18112 27168 18176 27172
rect 18192 27228 18256 27232
rect 18192 27172 18196 27228
rect 18196 27172 18252 27228
rect 18252 27172 18256 27228
rect 18192 27168 18256 27172
rect 27952 27228 28016 27232
rect 27952 27172 27956 27228
rect 27956 27172 28012 27228
rect 28012 27172 28016 27228
rect 27952 27168 28016 27172
rect 28032 27228 28096 27232
rect 28032 27172 28036 27228
rect 28036 27172 28092 27228
rect 28092 27172 28096 27228
rect 28032 27168 28096 27172
rect 28112 27228 28176 27232
rect 28112 27172 28116 27228
rect 28116 27172 28172 27228
rect 28172 27172 28176 27228
rect 28112 27168 28176 27172
rect 28192 27228 28256 27232
rect 28192 27172 28196 27228
rect 28196 27172 28252 27228
rect 28252 27172 28256 27228
rect 28192 27168 28256 27172
rect 37952 27228 38016 27232
rect 37952 27172 37956 27228
rect 37956 27172 38012 27228
rect 38012 27172 38016 27228
rect 37952 27168 38016 27172
rect 38032 27228 38096 27232
rect 38032 27172 38036 27228
rect 38036 27172 38092 27228
rect 38092 27172 38096 27228
rect 38032 27168 38096 27172
rect 38112 27228 38176 27232
rect 38112 27172 38116 27228
rect 38116 27172 38172 27228
rect 38172 27172 38176 27228
rect 38112 27168 38176 27172
rect 38192 27228 38256 27232
rect 38192 27172 38196 27228
rect 38196 27172 38252 27228
rect 38252 27172 38256 27228
rect 38192 27168 38256 27172
rect 47952 27228 48016 27232
rect 47952 27172 47956 27228
rect 47956 27172 48012 27228
rect 48012 27172 48016 27228
rect 47952 27168 48016 27172
rect 48032 27228 48096 27232
rect 48032 27172 48036 27228
rect 48036 27172 48092 27228
rect 48092 27172 48096 27228
rect 48032 27168 48096 27172
rect 48112 27228 48176 27232
rect 48112 27172 48116 27228
rect 48116 27172 48172 27228
rect 48172 27172 48176 27228
rect 48112 27168 48176 27172
rect 48192 27228 48256 27232
rect 48192 27172 48196 27228
rect 48196 27172 48252 27228
rect 48252 27172 48256 27228
rect 48192 27168 48256 27172
rect 30972 26964 31036 27028
rect 37412 26964 37476 27028
rect 38516 26964 38580 27028
rect 2952 26684 3016 26688
rect 2952 26628 2956 26684
rect 2956 26628 3012 26684
rect 3012 26628 3016 26684
rect 2952 26624 3016 26628
rect 3032 26684 3096 26688
rect 3032 26628 3036 26684
rect 3036 26628 3092 26684
rect 3092 26628 3096 26684
rect 3032 26624 3096 26628
rect 3112 26684 3176 26688
rect 3112 26628 3116 26684
rect 3116 26628 3172 26684
rect 3172 26628 3176 26684
rect 3112 26624 3176 26628
rect 3192 26684 3256 26688
rect 3192 26628 3196 26684
rect 3196 26628 3252 26684
rect 3252 26628 3256 26684
rect 3192 26624 3256 26628
rect 12952 26684 13016 26688
rect 12952 26628 12956 26684
rect 12956 26628 13012 26684
rect 13012 26628 13016 26684
rect 12952 26624 13016 26628
rect 13032 26684 13096 26688
rect 13032 26628 13036 26684
rect 13036 26628 13092 26684
rect 13092 26628 13096 26684
rect 13032 26624 13096 26628
rect 13112 26684 13176 26688
rect 13112 26628 13116 26684
rect 13116 26628 13172 26684
rect 13172 26628 13176 26684
rect 13112 26624 13176 26628
rect 13192 26684 13256 26688
rect 13192 26628 13196 26684
rect 13196 26628 13252 26684
rect 13252 26628 13256 26684
rect 13192 26624 13256 26628
rect 22952 26684 23016 26688
rect 22952 26628 22956 26684
rect 22956 26628 23012 26684
rect 23012 26628 23016 26684
rect 22952 26624 23016 26628
rect 23032 26684 23096 26688
rect 23032 26628 23036 26684
rect 23036 26628 23092 26684
rect 23092 26628 23096 26684
rect 23032 26624 23096 26628
rect 23112 26684 23176 26688
rect 23112 26628 23116 26684
rect 23116 26628 23172 26684
rect 23172 26628 23176 26684
rect 23112 26624 23176 26628
rect 23192 26684 23256 26688
rect 23192 26628 23196 26684
rect 23196 26628 23252 26684
rect 23252 26628 23256 26684
rect 23192 26624 23256 26628
rect 32952 26684 33016 26688
rect 32952 26628 32956 26684
rect 32956 26628 33012 26684
rect 33012 26628 33016 26684
rect 32952 26624 33016 26628
rect 33032 26684 33096 26688
rect 33032 26628 33036 26684
rect 33036 26628 33092 26684
rect 33092 26628 33096 26684
rect 33032 26624 33096 26628
rect 33112 26684 33176 26688
rect 33112 26628 33116 26684
rect 33116 26628 33172 26684
rect 33172 26628 33176 26684
rect 33112 26624 33176 26628
rect 33192 26684 33256 26688
rect 33192 26628 33196 26684
rect 33196 26628 33252 26684
rect 33252 26628 33256 26684
rect 33192 26624 33256 26628
rect 42952 26684 43016 26688
rect 42952 26628 42956 26684
rect 42956 26628 43012 26684
rect 43012 26628 43016 26684
rect 42952 26624 43016 26628
rect 43032 26684 43096 26688
rect 43032 26628 43036 26684
rect 43036 26628 43092 26684
rect 43092 26628 43096 26684
rect 43032 26624 43096 26628
rect 43112 26684 43176 26688
rect 43112 26628 43116 26684
rect 43116 26628 43172 26684
rect 43172 26628 43176 26684
rect 43112 26624 43176 26628
rect 43192 26684 43256 26688
rect 43192 26628 43196 26684
rect 43196 26628 43252 26684
rect 43252 26628 43256 26684
rect 43192 26624 43256 26628
rect 32628 26284 32692 26348
rect 39988 26284 40052 26348
rect 7952 26140 8016 26144
rect 7952 26084 7956 26140
rect 7956 26084 8012 26140
rect 8012 26084 8016 26140
rect 7952 26080 8016 26084
rect 8032 26140 8096 26144
rect 8032 26084 8036 26140
rect 8036 26084 8092 26140
rect 8092 26084 8096 26140
rect 8032 26080 8096 26084
rect 8112 26140 8176 26144
rect 8112 26084 8116 26140
rect 8116 26084 8172 26140
rect 8172 26084 8176 26140
rect 8112 26080 8176 26084
rect 8192 26140 8256 26144
rect 8192 26084 8196 26140
rect 8196 26084 8252 26140
rect 8252 26084 8256 26140
rect 8192 26080 8256 26084
rect 17952 26140 18016 26144
rect 17952 26084 17956 26140
rect 17956 26084 18012 26140
rect 18012 26084 18016 26140
rect 17952 26080 18016 26084
rect 18032 26140 18096 26144
rect 18032 26084 18036 26140
rect 18036 26084 18092 26140
rect 18092 26084 18096 26140
rect 18032 26080 18096 26084
rect 18112 26140 18176 26144
rect 18112 26084 18116 26140
rect 18116 26084 18172 26140
rect 18172 26084 18176 26140
rect 18112 26080 18176 26084
rect 18192 26140 18256 26144
rect 18192 26084 18196 26140
rect 18196 26084 18252 26140
rect 18252 26084 18256 26140
rect 18192 26080 18256 26084
rect 27952 26140 28016 26144
rect 27952 26084 27956 26140
rect 27956 26084 28012 26140
rect 28012 26084 28016 26140
rect 27952 26080 28016 26084
rect 28032 26140 28096 26144
rect 28032 26084 28036 26140
rect 28036 26084 28092 26140
rect 28092 26084 28096 26140
rect 28032 26080 28096 26084
rect 28112 26140 28176 26144
rect 28112 26084 28116 26140
rect 28116 26084 28172 26140
rect 28172 26084 28176 26140
rect 28112 26080 28176 26084
rect 28192 26140 28256 26144
rect 28192 26084 28196 26140
rect 28196 26084 28252 26140
rect 28252 26084 28256 26140
rect 28192 26080 28256 26084
rect 37952 26140 38016 26144
rect 37952 26084 37956 26140
rect 37956 26084 38012 26140
rect 38012 26084 38016 26140
rect 37952 26080 38016 26084
rect 38032 26140 38096 26144
rect 38032 26084 38036 26140
rect 38036 26084 38092 26140
rect 38092 26084 38096 26140
rect 38032 26080 38096 26084
rect 38112 26140 38176 26144
rect 38112 26084 38116 26140
rect 38116 26084 38172 26140
rect 38172 26084 38176 26140
rect 38112 26080 38176 26084
rect 38192 26140 38256 26144
rect 38192 26084 38196 26140
rect 38196 26084 38252 26140
rect 38252 26084 38256 26140
rect 38192 26080 38256 26084
rect 47952 26140 48016 26144
rect 47952 26084 47956 26140
rect 47956 26084 48012 26140
rect 48012 26084 48016 26140
rect 47952 26080 48016 26084
rect 48032 26140 48096 26144
rect 48032 26084 48036 26140
rect 48036 26084 48092 26140
rect 48092 26084 48096 26140
rect 48032 26080 48096 26084
rect 48112 26140 48176 26144
rect 48112 26084 48116 26140
rect 48116 26084 48172 26140
rect 48172 26084 48176 26140
rect 48112 26080 48176 26084
rect 48192 26140 48256 26144
rect 48192 26084 48196 26140
rect 48196 26084 48252 26140
rect 48252 26084 48256 26140
rect 48192 26080 48256 26084
rect 2952 25596 3016 25600
rect 2952 25540 2956 25596
rect 2956 25540 3012 25596
rect 3012 25540 3016 25596
rect 2952 25536 3016 25540
rect 3032 25596 3096 25600
rect 3032 25540 3036 25596
rect 3036 25540 3092 25596
rect 3092 25540 3096 25596
rect 3032 25536 3096 25540
rect 3112 25596 3176 25600
rect 3112 25540 3116 25596
rect 3116 25540 3172 25596
rect 3172 25540 3176 25596
rect 3112 25536 3176 25540
rect 3192 25596 3256 25600
rect 3192 25540 3196 25596
rect 3196 25540 3252 25596
rect 3252 25540 3256 25596
rect 3192 25536 3256 25540
rect 12952 25596 13016 25600
rect 12952 25540 12956 25596
rect 12956 25540 13012 25596
rect 13012 25540 13016 25596
rect 12952 25536 13016 25540
rect 13032 25596 13096 25600
rect 13032 25540 13036 25596
rect 13036 25540 13092 25596
rect 13092 25540 13096 25596
rect 13032 25536 13096 25540
rect 13112 25596 13176 25600
rect 13112 25540 13116 25596
rect 13116 25540 13172 25596
rect 13172 25540 13176 25596
rect 13112 25536 13176 25540
rect 13192 25596 13256 25600
rect 13192 25540 13196 25596
rect 13196 25540 13252 25596
rect 13252 25540 13256 25596
rect 13192 25536 13256 25540
rect 22952 25596 23016 25600
rect 22952 25540 22956 25596
rect 22956 25540 23012 25596
rect 23012 25540 23016 25596
rect 22952 25536 23016 25540
rect 23032 25596 23096 25600
rect 23032 25540 23036 25596
rect 23036 25540 23092 25596
rect 23092 25540 23096 25596
rect 23032 25536 23096 25540
rect 23112 25596 23176 25600
rect 23112 25540 23116 25596
rect 23116 25540 23172 25596
rect 23172 25540 23176 25596
rect 23112 25536 23176 25540
rect 23192 25596 23256 25600
rect 23192 25540 23196 25596
rect 23196 25540 23252 25596
rect 23252 25540 23256 25596
rect 23192 25536 23256 25540
rect 32952 25596 33016 25600
rect 32952 25540 32956 25596
rect 32956 25540 33012 25596
rect 33012 25540 33016 25596
rect 32952 25536 33016 25540
rect 33032 25596 33096 25600
rect 33032 25540 33036 25596
rect 33036 25540 33092 25596
rect 33092 25540 33096 25596
rect 33032 25536 33096 25540
rect 33112 25596 33176 25600
rect 33112 25540 33116 25596
rect 33116 25540 33172 25596
rect 33172 25540 33176 25596
rect 33112 25536 33176 25540
rect 33192 25596 33256 25600
rect 33192 25540 33196 25596
rect 33196 25540 33252 25596
rect 33252 25540 33256 25596
rect 33192 25536 33256 25540
rect 42952 25596 43016 25600
rect 42952 25540 42956 25596
rect 42956 25540 43012 25596
rect 43012 25540 43016 25596
rect 42952 25536 43016 25540
rect 43032 25596 43096 25600
rect 43032 25540 43036 25596
rect 43036 25540 43092 25596
rect 43092 25540 43096 25596
rect 43032 25536 43096 25540
rect 43112 25596 43176 25600
rect 43112 25540 43116 25596
rect 43116 25540 43172 25596
rect 43172 25540 43176 25596
rect 43112 25536 43176 25540
rect 43192 25596 43256 25600
rect 43192 25540 43196 25596
rect 43196 25540 43252 25596
rect 43252 25540 43256 25596
rect 43192 25536 43256 25540
rect 30420 25196 30484 25260
rect 7952 25052 8016 25056
rect 7952 24996 7956 25052
rect 7956 24996 8012 25052
rect 8012 24996 8016 25052
rect 7952 24992 8016 24996
rect 8032 25052 8096 25056
rect 8032 24996 8036 25052
rect 8036 24996 8092 25052
rect 8092 24996 8096 25052
rect 8032 24992 8096 24996
rect 8112 25052 8176 25056
rect 8112 24996 8116 25052
rect 8116 24996 8172 25052
rect 8172 24996 8176 25052
rect 8112 24992 8176 24996
rect 8192 25052 8256 25056
rect 8192 24996 8196 25052
rect 8196 24996 8252 25052
rect 8252 24996 8256 25052
rect 8192 24992 8256 24996
rect 17952 25052 18016 25056
rect 17952 24996 17956 25052
rect 17956 24996 18012 25052
rect 18012 24996 18016 25052
rect 17952 24992 18016 24996
rect 18032 25052 18096 25056
rect 18032 24996 18036 25052
rect 18036 24996 18092 25052
rect 18092 24996 18096 25052
rect 18032 24992 18096 24996
rect 18112 25052 18176 25056
rect 18112 24996 18116 25052
rect 18116 24996 18172 25052
rect 18172 24996 18176 25052
rect 18112 24992 18176 24996
rect 18192 25052 18256 25056
rect 18192 24996 18196 25052
rect 18196 24996 18252 25052
rect 18252 24996 18256 25052
rect 18192 24992 18256 24996
rect 27952 25052 28016 25056
rect 27952 24996 27956 25052
rect 27956 24996 28012 25052
rect 28012 24996 28016 25052
rect 27952 24992 28016 24996
rect 28032 25052 28096 25056
rect 28032 24996 28036 25052
rect 28036 24996 28092 25052
rect 28092 24996 28096 25052
rect 28032 24992 28096 24996
rect 28112 25052 28176 25056
rect 28112 24996 28116 25052
rect 28116 24996 28172 25052
rect 28172 24996 28176 25052
rect 28112 24992 28176 24996
rect 28192 25052 28256 25056
rect 28192 24996 28196 25052
rect 28196 24996 28252 25052
rect 28252 24996 28256 25052
rect 28192 24992 28256 24996
rect 37952 25052 38016 25056
rect 37952 24996 37956 25052
rect 37956 24996 38012 25052
rect 38012 24996 38016 25052
rect 37952 24992 38016 24996
rect 38032 25052 38096 25056
rect 38032 24996 38036 25052
rect 38036 24996 38092 25052
rect 38092 24996 38096 25052
rect 38032 24992 38096 24996
rect 38112 25052 38176 25056
rect 38112 24996 38116 25052
rect 38116 24996 38172 25052
rect 38172 24996 38176 25052
rect 38112 24992 38176 24996
rect 38192 25052 38256 25056
rect 38192 24996 38196 25052
rect 38196 24996 38252 25052
rect 38252 24996 38256 25052
rect 38192 24992 38256 24996
rect 47952 25052 48016 25056
rect 47952 24996 47956 25052
rect 47956 24996 48012 25052
rect 48012 24996 48016 25052
rect 47952 24992 48016 24996
rect 48032 25052 48096 25056
rect 48032 24996 48036 25052
rect 48036 24996 48092 25052
rect 48092 24996 48096 25052
rect 48032 24992 48096 24996
rect 48112 25052 48176 25056
rect 48112 24996 48116 25052
rect 48116 24996 48172 25052
rect 48172 24996 48176 25052
rect 48112 24992 48176 24996
rect 48192 25052 48256 25056
rect 48192 24996 48196 25052
rect 48196 24996 48252 25052
rect 48252 24996 48256 25052
rect 48192 24992 48256 24996
rect 2952 24508 3016 24512
rect 2952 24452 2956 24508
rect 2956 24452 3012 24508
rect 3012 24452 3016 24508
rect 2952 24448 3016 24452
rect 3032 24508 3096 24512
rect 3032 24452 3036 24508
rect 3036 24452 3092 24508
rect 3092 24452 3096 24508
rect 3032 24448 3096 24452
rect 3112 24508 3176 24512
rect 3112 24452 3116 24508
rect 3116 24452 3172 24508
rect 3172 24452 3176 24508
rect 3112 24448 3176 24452
rect 3192 24508 3256 24512
rect 3192 24452 3196 24508
rect 3196 24452 3252 24508
rect 3252 24452 3256 24508
rect 3192 24448 3256 24452
rect 12952 24508 13016 24512
rect 12952 24452 12956 24508
rect 12956 24452 13012 24508
rect 13012 24452 13016 24508
rect 12952 24448 13016 24452
rect 13032 24508 13096 24512
rect 13032 24452 13036 24508
rect 13036 24452 13092 24508
rect 13092 24452 13096 24508
rect 13032 24448 13096 24452
rect 13112 24508 13176 24512
rect 13112 24452 13116 24508
rect 13116 24452 13172 24508
rect 13172 24452 13176 24508
rect 13112 24448 13176 24452
rect 13192 24508 13256 24512
rect 13192 24452 13196 24508
rect 13196 24452 13252 24508
rect 13252 24452 13256 24508
rect 13192 24448 13256 24452
rect 22952 24508 23016 24512
rect 22952 24452 22956 24508
rect 22956 24452 23012 24508
rect 23012 24452 23016 24508
rect 22952 24448 23016 24452
rect 23032 24508 23096 24512
rect 23032 24452 23036 24508
rect 23036 24452 23092 24508
rect 23092 24452 23096 24508
rect 23032 24448 23096 24452
rect 23112 24508 23176 24512
rect 23112 24452 23116 24508
rect 23116 24452 23172 24508
rect 23172 24452 23176 24508
rect 23112 24448 23176 24452
rect 23192 24508 23256 24512
rect 23192 24452 23196 24508
rect 23196 24452 23252 24508
rect 23252 24452 23256 24508
rect 23192 24448 23256 24452
rect 32952 24508 33016 24512
rect 32952 24452 32956 24508
rect 32956 24452 33012 24508
rect 33012 24452 33016 24508
rect 32952 24448 33016 24452
rect 33032 24508 33096 24512
rect 33032 24452 33036 24508
rect 33036 24452 33092 24508
rect 33092 24452 33096 24508
rect 33032 24448 33096 24452
rect 33112 24508 33176 24512
rect 33112 24452 33116 24508
rect 33116 24452 33172 24508
rect 33172 24452 33176 24508
rect 33112 24448 33176 24452
rect 33192 24508 33256 24512
rect 33192 24452 33196 24508
rect 33196 24452 33252 24508
rect 33252 24452 33256 24508
rect 33192 24448 33256 24452
rect 42952 24508 43016 24512
rect 42952 24452 42956 24508
rect 42956 24452 43012 24508
rect 43012 24452 43016 24508
rect 42952 24448 43016 24452
rect 43032 24508 43096 24512
rect 43032 24452 43036 24508
rect 43036 24452 43092 24508
rect 43092 24452 43096 24508
rect 43032 24448 43096 24452
rect 43112 24508 43176 24512
rect 43112 24452 43116 24508
rect 43116 24452 43172 24508
rect 43172 24452 43176 24508
rect 43112 24448 43176 24452
rect 43192 24508 43256 24512
rect 43192 24452 43196 24508
rect 43196 24452 43252 24508
rect 43252 24452 43256 24508
rect 43192 24448 43256 24452
rect 25636 24244 25700 24308
rect 27660 24168 27724 24172
rect 27660 24112 27710 24168
rect 27710 24112 27724 24168
rect 27660 24108 27724 24112
rect 7952 23964 8016 23968
rect 7952 23908 7956 23964
rect 7956 23908 8012 23964
rect 8012 23908 8016 23964
rect 7952 23904 8016 23908
rect 8032 23964 8096 23968
rect 8032 23908 8036 23964
rect 8036 23908 8092 23964
rect 8092 23908 8096 23964
rect 8032 23904 8096 23908
rect 8112 23964 8176 23968
rect 8112 23908 8116 23964
rect 8116 23908 8172 23964
rect 8172 23908 8176 23964
rect 8112 23904 8176 23908
rect 8192 23964 8256 23968
rect 8192 23908 8196 23964
rect 8196 23908 8252 23964
rect 8252 23908 8256 23964
rect 8192 23904 8256 23908
rect 17952 23964 18016 23968
rect 17952 23908 17956 23964
rect 17956 23908 18012 23964
rect 18012 23908 18016 23964
rect 17952 23904 18016 23908
rect 18032 23964 18096 23968
rect 18032 23908 18036 23964
rect 18036 23908 18092 23964
rect 18092 23908 18096 23964
rect 18032 23904 18096 23908
rect 18112 23964 18176 23968
rect 18112 23908 18116 23964
rect 18116 23908 18172 23964
rect 18172 23908 18176 23964
rect 18112 23904 18176 23908
rect 18192 23964 18256 23968
rect 18192 23908 18196 23964
rect 18196 23908 18252 23964
rect 18252 23908 18256 23964
rect 18192 23904 18256 23908
rect 27952 23964 28016 23968
rect 27952 23908 27956 23964
rect 27956 23908 28012 23964
rect 28012 23908 28016 23964
rect 27952 23904 28016 23908
rect 28032 23964 28096 23968
rect 28032 23908 28036 23964
rect 28036 23908 28092 23964
rect 28092 23908 28096 23964
rect 28032 23904 28096 23908
rect 28112 23964 28176 23968
rect 28112 23908 28116 23964
rect 28116 23908 28172 23964
rect 28172 23908 28176 23964
rect 28112 23904 28176 23908
rect 28192 23964 28256 23968
rect 28192 23908 28196 23964
rect 28196 23908 28252 23964
rect 28252 23908 28256 23964
rect 28192 23904 28256 23908
rect 37952 23964 38016 23968
rect 37952 23908 37956 23964
rect 37956 23908 38012 23964
rect 38012 23908 38016 23964
rect 37952 23904 38016 23908
rect 38032 23964 38096 23968
rect 38032 23908 38036 23964
rect 38036 23908 38092 23964
rect 38092 23908 38096 23964
rect 38032 23904 38096 23908
rect 38112 23964 38176 23968
rect 38112 23908 38116 23964
rect 38116 23908 38172 23964
rect 38172 23908 38176 23964
rect 38112 23904 38176 23908
rect 38192 23964 38256 23968
rect 38192 23908 38196 23964
rect 38196 23908 38252 23964
rect 38252 23908 38256 23964
rect 38192 23904 38256 23908
rect 47952 23964 48016 23968
rect 47952 23908 47956 23964
rect 47956 23908 48012 23964
rect 48012 23908 48016 23964
rect 47952 23904 48016 23908
rect 48032 23964 48096 23968
rect 48032 23908 48036 23964
rect 48036 23908 48092 23964
rect 48092 23908 48096 23964
rect 48032 23904 48096 23908
rect 48112 23964 48176 23968
rect 48112 23908 48116 23964
rect 48116 23908 48172 23964
rect 48172 23908 48176 23964
rect 48112 23904 48176 23908
rect 48192 23964 48256 23968
rect 48192 23908 48196 23964
rect 48196 23908 48252 23964
rect 48252 23908 48256 23964
rect 48192 23904 48256 23908
rect 22140 23564 22204 23628
rect 2952 23420 3016 23424
rect 2952 23364 2956 23420
rect 2956 23364 3012 23420
rect 3012 23364 3016 23420
rect 2952 23360 3016 23364
rect 3032 23420 3096 23424
rect 3032 23364 3036 23420
rect 3036 23364 3092 23420
rect 3092 23364 3096 23420
rect 3032 23360 3096 23364
rect 3112 23420 3176 23424
rect 3112 23364 3116 23420
rect 3116 23364 3172 23420
rect 3172 23364 3176 23420
rect 3112 23360 3176 23364
rect 3192 23420 3256 23424
rect 3192 23364 3196 23420
rect 3196 23364 3252 23420
rect 3252 23364 3256 23420
rect 3192 23360 3256 23364
rect 12952 23420 13016 23424
rect 12952 23364 12956 23420
rect 12956 23364 13012 23420
rect 13012 23364 13016 23420
rect 12952 23360 13016 23364
rect 13032 23420 13096 23424
rect 13032 23364 13036 23420
rect 13036 23364 13092 23420
rect 13092 23364 13096 23420
rect 13032 23360 13096 23364
rect 13112 23420 13176 23424
rect 13112 23364 13116 23420
rect 13116 23364 13172 23420
rect 13172 23364 13176 23420
rect 13112 23360 13176 23364
rect 13192 23420 13256 23424
rect 13192 23364 13196 23420
rect 13196 23364 13252 23420
rect 13252 23364 13256 23420
rect 13192 23360 13256 23364
rect 22952 23420 23016 23424
rect 22952 23364 22956 23420
rect 22956 23364 23012 23420
rect 23012 23364 23016 23420
rect 22952 23360 23016 23364
rect 23032 23420 23096 23424
rect 23032 23364 23036 23420
rect 23036 23364 23092 23420
rect 23092 23364 23096 23420
rect 23032 23360 23096 23364
rect 23112 23420 23176 23424
rect 23112 23364 23116 23420
rect 23116 23364 23172 23420
rect 23172 23364 23176 23420
rect 23112 23360 23176 23364
rect 23192 23420 23256 23424
rect 23192 23364 23196 23420
rect 23196 23364 23252 23420
rect 23252 23364 23256 23420
rect 23192 23360 23256 23364
rect 32952 23420 33016 23424
rect 32952 23364 32956 23420
rect 32956 23364 33012 23420
rect 33012 23364 33016 23420
rect 32952 23360 33016 23364
rect 33032 23420 33096 23424
rect 33032 23364 33036 23420
rect 33036 23364 33092 23420
rect 33092 23364 33096 23420
rect 33032 23360 33096 23364
rect 33112 23420 33176 23424
rect 33112 23364 33116 23420
rect 33116 23364 33172 23420
rect 33172 23364 33176 23420
rect 33112 23360 33176 23364
rect 33192 23420 33256 23424
rect 33192 23364 33196 23420
rect 33196 23364 33252 23420
rect 33252 23364 33256 23420
rect 33192 23360 33256 23364
rect 42952 23420 43016 23424
rect 42952 23364 42956 23420
rect 42956 23364 43012 23420
rect 43012 23364 43016 23420
rect 42952 23360 43016 23364
rect 43032 23420 43096 23424
rect 43032 23364 43036 23420
rect 43036 23364 43092 23420
rect 43092 23364 43096 23420
rect 43032 23360 43096 23364
rect 43112 23420 43176 23424
rect 43112 23364 43116 23420
rect 43116 23364 43172 23420
rect 43172 23364 43176 23420
rect 43112 23360 43176 23364
rect 43192 23420 43256 23424
rect 43192 23364 43196 23420
rect 43196 23364 43252 23420
rect 43252 23364 43256 23420
rect 43192 23360 43256 23364
rect 22508 22884 22572 22948
rect 7952 22876 8016 22880
rect 7952 22820 7956 22876
rect 7956 22820 8012 22876
rect 8012 22820 8016 22876
rect 7952 22816 8016 22820
rect 8032 22876 8096 22880
rect 8032 22820 8036 22876
rect 8036 22820 8092 22876
rect 8092 22820 8096 22876
rect 8032 22816 8096 22820
rect 8112 22876 8176 22880
rect 8112 22820 8116 22876
rect 8116 22820 8172 22876
rect 8172 22820 8176 22876
rect 8112 22816 8176 22820
rect 8192 22876 8256 22880
rect 8192 22820 8196 22876
rect 8196 22820 8252 22876
rect 8252 22820 8256 22876
rect 8192 22816 8256 22820
rect 17952 22876 18016 22880
rect 17952 22820 17956 22876
rect 17956 22820 18012 22876
rect 18012 22820 18016 22876
rect 17952 22816 18016 22820
rect 18032 22876 18096 22880
rect 18032 22820 18036 22876
rect 18036 22820 18092 22876
rect 18092 22820 18096 22876
rect 18032 22816 18096 22820
rect 18112 22876 18176 22880
rect 18112 22820 18116 22876
rect 18116 22820 18172 22876
rect 18172 22820 18176 22876
rect 18112 22816 18176 22820
rect 18192 22876 18256 22880
rect 18192 22820 18196 22876
rect 18196 22820 18252 22876
rect 18252 22820 18256 22876
rect 18192 22816 18256 22820
rect 27952 22876 28016 22880
rect 27952 22820 27956 22876
rect 27956 22820 28012 22876
rect 28012 22820 28016 22876
rect 27952 22816 28016 22820
rect 28032 22876 28096 22880
rect 28032 22820 28036 22876
rect 28036 22820 28092 22876
rect 28092 22820 28096 22876
rect 28032 22816 28096 22820
rect 28112 22876 28176 22880
rect 28112 22820 28116 22876
rect 28116 22820 28172 22876
rect 28172 22820 28176 22876
rect 28112 22816 28176 22820
rect 28192 22876 28256 22880
rect 28192 22820 28196 22876
rect 28196 22820 28252 22876
rect 28252 22820 28256 22876
rect 28192 22816 28256 22820
rect 37952 22876 38016 22880
rect 37952 22820 37956 22876
rect 37956 22820 38012 22876
rect 38012 22820 38016 22876
rect 37952 22816 38016 22820
rect 38032 22876 38096 22880
rect 38032 22820 38036 22876
rect 38036 22820 38092 22876
rect 38092 22820 38096 22876
rect 38032 22816 38096 22820
rect 38112 22876 38176 22880
rect 38112 22820 38116 22876
rect 38116 22820 38172 22876
rect 38172 22820 38176 22876
rect 38112 22816 38176 22820
rect 38192 22876 38256 22880
rect 38192 22820 38196 22876
rect 38196 22820 38252 22876
rect 38252 22820 38256 22876
rect 38192 22816 38256 22820
rect 47952 22876 48016 22880
rect 47952 22820 47956 22876
rect 47956 22820 48012 22876
rect 48012 22820 48016 22876
rect 47952 22816 48016 22820
rect 48032 22876 48096 22880
rect 48032 22820 48036 22876
rect 48036 22820 48092 22876
rect 48092 22820 48096 22876
rect 48032 22816 48096 22820
rect 48112 22876 48176 22880
rect 48112 22820 48116 22876
rect 48116 22820 48172 22876
rect 48172 22820 48176 22876
rect 48112 22816 48176 22820
rect 48192 22876 48256 22880
rect 48192 22820 48196 22876
rect 48196 22820 48252 22876
rect 48252 22820 48256 22876
rect 48192 22816 48256 22820
rect 2952 22332 3016 22336
rect 2952 22276 2956 22332
rect 2956 22276 3012 22332
rect 3012 22276 3016 22332
rect 2952 22272 3016 22276
rect 3032 22332 3096 22336
rect 3032 22276 3036 22332
rect 3036 22276 3092 22332
rect 3092 22276 3096 22332
rect 3032 22272 3096 22276
rect 3112 22332 3176 22336
rect 3112 22276 3116 22332
rect 3116 22276 3172 22332
rect 3172 22276 3176 22332
rect 3112 22272 3176 22276
rect 3192 22332 3256 22336
rect 3192 22276 3196 22332
rect 3196 22276 3252 22332
rect 3252 22276 3256 22332
rect 3192 22272 3256 22276
rect 12952 22332 13016 22336
rect 12952 22276 12956 22332
rect 12956 22276 13012 22332
rect 13012 22276 13016 22332
rect 12952 22272 13016 22276
rect 13032 22332 13096 22336
rect 13032 22276 13036 22332
rect 13036 22276 13092 22332
rect 13092 22276 13096 22332
rect 13032 22272 13096 22276
rect 13112 22332 13176 22336
rect 13112 22276 13116 22332
rect 13116 22276 13172 22332
rect 13172 22276 13176 22332
rect 13112 22272 13176 22276
rect 13192 22332 13256 22336
rect 13192 22276 13196 22332
rect 13196 22276 13252 22332
rect 13252 22276 13256 22332
rect 13192 22272 13256 22276
rect 22952 22332 23016 22336
rect 22952 22276 22956 22332
rect 22956 22276 23012 22332
rect 23012 22276 23016 22332
rect 22952 22272 23016 22276
rect 23032 22332 23096 22336
rect 23032 22276 23036 22332
rect 23036 22276 23092 22332
rect 23092 22276 23096 22332
rect 23032 22272 23096 22276
rect 23112 22332 23176 22336
rect 23112 22276 23116 22332
rect 23116 22276 23172 22332
rect 23172 22276 23176 22332
rect 23112 22272 23176 22276
rect 23192 22332 23256 22336
rect 23192 22276 23196 22332
rect 23196 22276 23252 22332
rect 23252 22276 23256 22332
rect 23192 22272 23256 22276
rect 32952 22332 33016 22336
rect 32952 22276 32956 22332
rect 32956 22276 33012 22332
rect 33012 22276 33016 22332
rect 32952 22272 33016 22276
rect 33032 22332 33096 22336
rect 33032 22276 33036 22332
rect 33036 22276 33092 22332
rect 33092 22276 33096 22332
rect 33032 22272 33096 22276
rect 33112 22332 33176 22336
rect 33112 22276 33116 22332
rect 33116 22276 33172 22332
rect 33172 22276 33176 22332
rect 33112 22272 33176 22276
rect 33192 22332 33256 22336
rect 33192 22276 33196 22332
rect 33196 22276 33252 22332
rect 33252 22276 33256 22332
rect 33192 22272 33256 22276
rect 42952 22332 43016 22336
rect 42952 22276 42956 22332
rect 42956 22276 43012 22332
rect 43012 22276 43016 22332
rect 42952 22272 43016 22276
rect 43032 22332 43096 22336
rect 43032 22276 43036 22332
rect 43036 22276 43092 22332
rect 43092 22276 43096 22332
rect 43032 22272 43096 22276
rect 43112 22332 43176 22336
rect 43112 22276 43116 22332
rect 43116 22276 43172 22332
rect 43172 22276 43176 22332
rect 43112 22272 43176 22276
rect 43192 22332 43256 22336
rect 43192 22276 43196 22332
rect 43196 22276 43252 22332
rect 43252 22276 43256 22332
rect 43192 22272 43256 22276
rect 30788 21932 30852 21996
rect 7952 21788 8016 21792
rect 7952 21732 7956 21788
rect 7956 21732 8012 21788
rect 8012 21732 8016 21788
rect 7952 21728 8016 21732
rect 8032 21788 8096 21792
rect 8032 21732 8036 21788
rect 8036 21732 8092 21788
rect 8092 21732 8096 21788
rect 8032 21728 8096 21732
rect 8112 21788 8176 21792
rect 8112 21732 8116 21788
rect 8116 21732 8172 21788
rect 8172 21732 8176 21788
rect 8112 21728 8176 21732
rect 8192 21788 8256 21792
rect 8192 21732 8196 21788
rect 8196 21732 8252 21788
rect 8252 21732 8256 21788
rect 8192 21728 8256 21732
rect 17952 21788 18016 21792
rect 17952 21732 17956 21788
rect 17956 21732 18012 21788
rect 18012 21732 18016 21788
rect 17952 21728 18016 21732
rect 18032 21788 18096 21792
rect 18032 21732 18036 21788
rect 18036 21732 18092 21788
rect 18092 21732 18096 21788
rect 18032 21728 18096 21732
rect 18112 21788 18176 21792
rect 18112 21732 18116 21788
rect 18116 21732 18172 21788
rect 18172 21732 18176 21788
rect 18112 21728 18176 21732
rect 18192 21788 18256 21792
rect 18192 21732 18196 21788
rect 18196 21732 18252 21788
rect 18252 21732 18256 21788
rect 18192 21728 18256 21732
rect 27952 21788 28016 21792
rect 27952 21732 27956 21788
rect 27956 21732 28012 21788
rect 28012 21732 28016 21788
rect 27952 21728 28016 21732
rect 28032 21788 28096 21792
rect 28032 21732 28036 21788
rect 28036 21732 28092 21788
rect 28092 21732 28096 21788
rect 28032 21728 28096 21732
rect 28112 21788 28176 21792
rect 28112 21732 28116 21788
rect 28116 21732 28172 21788
rect 28172 21732 28176 21788
rect 28112 21728 28176 21732
rect 28192 21788 28256 21792
rect 28192 21732 28196 21788
rect 28196 21732 28252 21788
rect 28252 21732 28256 21788
rect 28192 21728 28256 21732
rect 37952 21788 38016 21792
rect 37952 21732 37956 21788
rect 37956 21732 38012 21788
rect 38012 21732 38016 21788
rect 37952 21728 38016 21732
rect 38032 21788 38096 21792
rect 38032 21732 38036 21788
rect 38036 21732 38092 21788
rect 38092 21732 38096 21788
rect 38032 21728 38096 21732
rect 38112 21788 38176 21792
rect 38112 21732 38116 21788
rect 38116 21732 38172 21788
rect 38172 21732 38176 21788
rect 38112 21728 38176 21732
rect 38192 21788 38256 21792
rect 38192 21732 38196 21788
rect 38196 21732 38252 21788
rect 38252 21732 38256 21788
rect 38192 21728 38256 21732
rect 47952 21788 48016 21792
rect 47952 21732 47956 21788
rect 47956 21732 48012 21788
rect 48012 21732 48016 21788
rect 47952 21728 48016 21732
rect 48032 21788 48096 21792
rect 48032 21732 48036 21788
rect 48036 21732 48092 21788
rect 48092 21732 48096 21788
rect 48032 21728 48096 21732
rect 48112 21788 48176 21792
rect 48112 21732 48116 21788
rect 48116 21732 48172 21788
rect 48172 21732 48176 21788
rect 48112 21728 48176 21732
rect 48192 21788 48256 21792
rect 48192 21732 48196 21788
rect 48196 21732 48252 21788
rect 48252 21732 48256 21788
rect 48192 21728 48256 21732
rect 2952 21244 3016 21248
rect 2952 21188 2956 21244
rect 2956 21188 3012 21244
rect 3012 21188 3016 21244
rect 2952 21184 3016 21188
rect 3032 21244 3096 21248
rect 3032 21188 3036 21244
rect 3036 21188 3092 21244
rect 3092 21188 3096 21244
rect 3032 21184 3096 21188
rect 3112 21244 3176 21248
rect 3112 21188 3116 21244
rect 3116 21188 3172 21244
rect 3172 21188 3176 21244
rect 3112 21184 3176 21188
rect 3192 21244 3256 21248
rect 3192 21188 3196 21244
rect 3196 21188 3252 21244
rect 3252 21188 3256 21244
rect 3192 21184 3256 21188
rect 12952 21244 13016 21248
rect 12952 21188 12956 21244
rect 12956 21188 13012 21244
rect 13012 21188 13016 21244
rect 12952 21184 13016 21188
rect 13032 21244 13096 21248
rect 13032 21188 13036 21244
rect 13036 21188 13092 21244
rect 13092 21188 13096 21244
rect 13032 21184 13096 21188
rect 13112 21244 13176 21248
rect 13112 21188 13116 21244
rect 13116 21188 13172 21244
rect 13172 21188 13176 21244
rect 13112 21184 13176 21188
rect 13192 21244 13256 21248
rect 13192 21188 13196 21244
rect 13196 21188 13252 21244
rect 13252 21188 13256 21244
rect 13192 21184 13256 21188
rect 22952 21244 23016 21248
rect 22952 21188 22956 21244
rect 22956 21188 23012 21244
rect 23012 21188 23016 21244
rect 22952 21184 23016 21188
rect 23032 21244 23096 21248
rect 23032 21188 23036 21244
rect 23036 21188 23092 21244
rect 23092 21188 23096 21244
rect 23032 21184 23096 21188
rect 23112 21244 23176 21248
rect 23112 21188 23116 21244
rect 23116 21188 23172 21244
rect 23172 21188 23176 21244
rect 23112 21184 23176 21188
rect 23192 21244 23256 21248
rect 23192 21188 23196 21244
rect 23196 21188 23252 21244
rect 23252 21188 23256 21244
rect 23192 21184 23256 21188
rect 32952 21244 33016 21248
rect 32952 21188 32956 21244
rect 32956 21188 33012 21244
rect 33012 21188 33016 21244
rect 32952 21184 33016 21188
rect 33032 21244 33096 21248
rect 33032 21188 33036 21244
rect 33036 21188 33092 21244
rect 33092 21188 33096 21244
rect 33032 21184 33096 21188
rect 33112 21244 33176 21248
rect 33112 21188 33116 21244
rect 33116 21188 33172 21244
rect 33172 21188 33176 21244
rect 33112 21184 33176 21188
rect 33192 21244 33256 21248
rect 33192 21188 33196 21244
rect 33196 21188 33252 21244
rect 33252 21188 33256 21244
rect 33192 21184 33256 21188
rect 42952 21244 43016 21248
rect 42952 21188 42956 21244
rect 42956 21188 43012 21244
rect 43012 21188 43016 21244
rect 42952 21184 43016 21188
rect 43032 21244 43096 21248
rect 43032 21188 43036 21244
rect 43036 21188 43092 21244
rect 43092 21188 43096 21244
rect 43032 21184 43096 21188
rect 43112 21244 43176 21248
rect 43112 21188 43116 21244
rect 43116 21188 43172 21244
rect 43172 21188 43176 21244
rect 43112 21184 43176 21188
rect 43192 21244 43256 21248
rect 43192 21188 43196 21244
rect 43196 21188 43252 21244
rect 43252 21188 43256 21244
rect 43192 21184 43256 21188
rect 7952 20700 8016 20704
rect 7952 20644 7956 20700
rect 7956 20644 8012 20700
rect 8012 20644 8016 20700
rect 7952 20640 8016 20644
rect 8032 20700 8096 20704
rect 8032 20644 8036 20700
rect 8036 20644 8092 20700
rect 8092 20644 8096 20700
rect 8032 20640 8096 20644
rect 8112 20700 8176 20704
rect 8112 20644 8116 20700
rect 8116 20644 8172 20700
rect 8172 20644 8176 20700
rect 8112 20640 8176 20644
rect 8192 20700 8256 20704
rect 8192 20644 8196 20700
rect 8196 20644 8252 20700
rect 8252 20644 8256 20700
rect 8192 20640 8256 20644
rect 17952 20700 18016 20704
rect 17952 20644 17956 20700
rect 17956 20644 18012 20700
rect 18012 20644 18016 20700
rect 17952 20640 18016 20644
rect 18032 20700 18096 20704
rect 18032 20644 18036 20700
rect 18036 20644 18092 20700
rect 18092 20644 18096 20700
rect 18032 20640 18096 20644
rect 18112 20700 18176 20704
rect 18112 20644 18116 20700
rect 18116 20644 18172 20700
rect 18172 20644 18176 20700
rect 18112 20640 18176 20644
rect 18192 20700 18256 20704
rect 18192 20644 18196 20700
rect 18196 20644 18252 20700
rect 18252 20644 18256 20700
rect 18192 20640 18256 20644
rect 27952 20700 28016 20704
rect 27952 20644 27956 20700
rect 27956 20644 28012 20700
rect 28012 20644 28016 20700
rect 27952 20640 28016 20644
rect 28032 20700 28096 20704
rect 28032 20644 28036 20700
rect 28036 20644 28092 20700
rect 28092 20644 28096 20700
rect 28032 20640 28096 20644
rect 28112 20700 28176 20704
rect 28112 20644 28116 20700
rect 28116 20644 28172 20700
rect 28172 20644 28176 20700
rect 28112 20640 28176 20644
rect 28192 20700 28256 20704
rect 28192 20644 28196 20700
rect 28196 20644 28252 20700
rect 28252 20644 28256 20700
rect 28192 20640 28256 20644
rect 37952 20700 38016 20704
rect 37952 20644 37956 20700
rect 37956 20644 38012 20700
rect 38012 20644 38016 20700
rect 37952 20640 38016 20644
rect 38032 20700 38096 20704
rect 38032 20644 38036 20700
rect 38036 20644 38092 20700
rect 38092 20644 38096 20700
rect 38032 20640 38096 20644
rect 38112 20700 38176 20704
rect 38112 20644 38116 20700
rect 38116 20644 38172 20700
rect 38172 20644 38176 20700
rect 38112 20640 38176 20644
rect 38192 20700 38256 20704
rect 38192 20644 38196 20700
rect 38196 20644 38252 20700
rect 38252 20644 38256 20700
rect 38192 20640 38256 20644
rect 47952 20700 48016 20704
rect 47952 20644 47956 20700
rect 47956 20644 48012 20700
rect 48012 20644 48016 20700
rect 47952 20640 48016 20644
rect 48032 20700 48096 20704
rect 48032 20644 48036 20700
rect 48036 20644 48092 20700
rect 48092 20644 48096 20700
rect 48032 20640 48096 20644
rect 48112 20700 48176 20704
rect 48112 20644 48116 20700
rect 48116 20644 48172 20700
rect 48172 20644 48176 20700
rect 48112 20640 48176 20644
rect 48192 20700 48256 20704
rect 48192 20644 48196 20700
rect 48196 20644 48252 20700
rect 48252 20644 48256 20700
rect 48192 20640 48256 20644
rect 30420 20632 30484 20636
rect 30420 20576 30470 20632
rect 30470 20576 30484 20632
rect 30420 20572 30484 20576
rect 35204 20632 35268 20636
rect 35204 20576 35218 20632
rect 35218 20576 35268 20632
rect 35204 20572 35268 20576
rect 2952 20156 3016 20160
rect 2952 20100 2956 20156
rect 2956 20100 3012 20156
rect 3012 20100 3016 20156
rect 2952 20096 3016 20100
rect 3032 20156 3096 20160
rect 3032 20100 3036 20156
rect 3036 20100 3092 20156
rect 3092 20100 3096 20156
rect 3032 20096 3096 20100
rect 3112 20156 3176 20160
rect 3112 20100 3116 20156
rect 3116 20100 3172 20156
rect 3172 20100 3176 20156
rect 3112 20096 3176 20100
rect 3192 20156 3256 20160
rect 3192 20100 3196 20156
rect 3196 20100 3252 20156
rect 3252 20100 3256 20156
rect 3192 20096 3256 20100
rect 12952 20156 13016 20160
rect 12952 20100 12956 20156
rect 12956 20100 13012 20156
rect 13012 20100 13016 20156
rect 12952 20096 13016 20100
rect 13032 20156 13096 20160
rect 13032 20100 13036 20156
rect 13036 20100 13092 20156
rect 13092 20100 13096 20156
rect 13032 20096 13096 20100
rect 13112 20156 13176 20160
rect 13112 20100 13116 20156
rect 13116 20100 13172 20156
rect 13172 20100 13176 20156
rect 13112 20096 13176 20100
rect 13192 20156 13256 20160
rect 13192 20100 13196 20156
rect 13196 20100 13252 20156
rect 13252 20100 13256 20156
rect 13192 20096 13256 20100
rect 22952 20156 23016 20160
rect 22952 20100 22956 20156
rect 22956 20100 23012 20156
rect 23012 20100 23016 20156
rect 22952 20096 23016 20100
rect 23032 20156 23096 20160
rect 23032 20100 23036 20156
rect 23036 20100 23092 20156
rect 23092 20100 23096 20156
rect 23032 20096 23096 20100
rect 23112 20156 23176 20160
rect 23112 20100 23116 20156
rect 23116 20100 23172 20156
rect 23172 20100 23176 20156
rect 23112 20096 23176 20100
rect 23192 20156 23256 20160
rect 23192 20100 23196 20156
rect 23196 20100 23252 20156
rect 23252 20100 23256 20156
rect 23192 20096 23256 20100
rect 32952 20156 33016 20160
rect 32952 20100 32956 20156
rect 32956 20100 33012 20156
rect 33012 20100 33016 20156
rect 32952 20096 33016 20100
rect 33032 20156 33096 20160
rect 33032 20100 33036 20156
rect 33036 20100 33092 20156
rect 33092 20100 33096 20156
rect 33032 20096 33096 20100
rect 33112 20156 33176 20160
rect 33112 20100 33116 20156
rect 33116 20100 33172 20156
rect 33172 20100 33176 20156
rect 33112 20096 33176 20100
rect 33192 20156 33256 20160
rect 33192 20100 33196 20156
rect 33196 20100 33252 20156
rect 33252 20100 33256 20156
rect 33192 20096 33256 20100
rect 42952 20156 43016 20160
rect 42952 20100 42956 20156
rect 42956 20100 43012 20156
rect 43012 20100 43016 20156
rect 42952 20096 43016 20100
rect 43032 20156 43096 20160
rect 43032 20100 43036 20156
rect 43036 20100 43092 20156
rect 43092 20100 43096 20156
rect 43032 20096 43096 20100
rect 43112 20156 43176 20160
rect 43112 20100 43116 20156
rect 43116 20100 43172 20156
rect 43172 20100 43176 20156
rect 43112 20096 43176 20100
rect 43192 20156 43256 20160
rect 43192 20100 43196 20156
rect 43196 20100 43252 20156
rect 43252 20100 43256 20156
rect 43192 20096 43256 20100
rect 7952 19612 8016 19616
rect 7952 19556 7956 19612
rect 7956 19556 8012 19612
rect 8012 19556 8016 19612
rect 7952 19552 8016 19556
rect 8032 19612 8096 19616
rect 8032 19556 8036 19612
rect 8036 19556 8092 19612
rect 8092 19556 8096 19612
rect 8032 19552 8096 19556
rect 8112 19612 8176 19616
rect 8112 19556 8116 19612
rect 8116 19556 8172 19612
rect 8172 19556 8176 19612
rect 8112 19552 8176 19556
rect 8192 19612 8256 19616
rect 8192 19556 8196 19612
rect 8196 19556 8252 19612
rect 8252 19556 8256 19612
rect 8192 19552 8256 19556
rect 17952 19612 18016 19616
rect 17952 19556 17956 19612
rect 17956 19556 18012 19612
rect 18012 19556 18016 19612
rect 17952 19552 18016 19556
rect 18032 19612 18096 19616
rect 18032 19556 18036 19612
rect 18036 19556 18092 19612
rect 18092 19556 18096 19612
rect 18032 19552 18096 19556
rect 18112 19612 18176 19616
rect 18112 19556 18116 19612
rect 18116 19556 18172 19612
rect 18172 19556 18176 19612
rect 18112 19552 18176 19556
rect 18192 19612 18256 19616
rect 18192 19556 18196 19612
rect 18196 19556 18252 19612
rect 18252 19556 18256 19612
rect 18192 19552 18256 19556
rect 27952 19612 28016 19616
rect 27952 19556 27956 19612
rect 27956 19556 28012 19612
rect 28012 19556 28016 19612
rect 27952 19552 28016 19556
rect 28032 19612 28096 19616
rect 28032 19556 28036 19612
rect 28036 19556 28092 19612
rect 28092 19556 28096 19612
rect 28032 19552 28096 19556
rect 28112 19612 28176 19616
rect 28112 19556 28116 19612
rect 28116 19556 28172 19612
rect 28172 19556 28176 19612
rect 28112 19552 28176 19556
rect 28192 19612 28256 19616
rect 28192 19556 28196 19612
rect 28196 19556 28252 19612
rect 28252 19556 28256 19612
rect 28192 19552 28256 19556
rect 37952 19612 38016 19616
rect 37952 19556 37956 19612
rect 37956 19556 38012 19612
rect 38012 19556 38016 19612
rect 37952 19552 38016 19556
rect 38032 19612 38096 19616
rect 38032 19556 38036 19612
rect 38036 19556 38092 19612
rect 38092 19556 38096 19612
rect 38032 19552 38096 19556
rect 38112 19612 38176 19616
rect 38112 19556 38116 19612
rect 38116 19556 38172 19612
rect 38172 19556 38176 19612
rect 38112 19552 38176 19556
rect 38192 19612 38256 19616
rect 38192 19556 38196 19612
rect 38196 19556 38252 19612
rect 38252 19556 38256 19612
rect 38192 19552 38256 19556
rect 47952 19612 48016 19616
rect 47952 19556 47956 19612
rect 47956 19556 48012 19612
rect 48012 19556 48016 19612
rect 47952 19552 48016 19556
rect 48032 19612 48096 19616
rect 48032 19556 48036 19612
rect 48036 19556 48092 19612
rect 48092 19556 48096 19612
rect 48032 19552 48096 19556
rect 48112 19612 48176 19616
rect 48112 19556 48116 19612
rect 48116 19556 48172 19612
rect 48172 19556 48176 19612
rect 48112 19552 48176 19556
rect 48192 19612 48256 19616
rect 48192 19556 48196 19612
rect 48196 19556 48252 19612
rect 48252 19556 48256 19612
rect 48192 19552 48256 19556
rect 32812 19212 32876 19276
rect 38516 19212 38580 19276
rect 2952 19068 3016 19072
rect 2952 19012 2956 19068
rect 2956 19012 3012 19068
rect 3012 19012 3016 19068
rect 2952 19008 3016 19012
rect 3032 19068 3096 19072
rect 3032 19012 3036 19068
rect 3036 19012 3092 19068
rect 3092 19012 3096 19068
rect 3032 19008 3096 19012
rect 3112 19068 3176 19072
rect 3112 19012 3116 19068
rect 3116 19012 3172 19068
rect 3172 19012 3176 19068
rect 3112 19008 3176 19012
rect 3192 19068 3256 19072
rect 3192 19012 3196 19068
rect 3196 19012 3252 19068
rect 3252 19012 3256 19068
rect 3192 19008 3256 19012
rect 12952 19068 13016 19072
rect 12952 19012 12956 19068
rect 12956 19012 13012 19068
rect 13012 19012 13016 19068
rect 12952 19008 13016 19012
rect 13032 19068 13096 19072
rect 13032 19012 13036 19068
rect 13036 19012 13092 19068
rect 13092 19012 13096 19068
rect 13032 19008 13096 19012
rect 13112 19068 13176 19072
rect 13112 19012 13116 19068
rect 13116 19012 13172 19068
rect 13172 19012 13176 19068
rect 13112 19008 13176 19012
rect 13192 19068 13256 19072
rect 13192 19012 13196 19068
rect 13196 19012 13252 19068
rect 13252 19012 13256 19068
rect 13192 19008 13256 19012
rect 22952 19068 23016 19072
rect 22952 19012 22956 19068
rect 22956 19012 23012 19068
rect 23012 19012 23016 19068
rect 22952 19008 23016 19012
rect 23032 19068 23096 19072
rect 23032 19012 23036 19068
rect 23036 19012 23092 19068
rect 23092 19012 23096 19068
rect 23032 19008 23096 19012
rect 23112 19068 23176 19072
rect 23112 19012 23116 19068
rect 23116 19012 23172 19068
rect 23172 19012 23176 19068
rect 23112 19008 23176 19012
rect 23192 19068 23256 19072
rect 23192 19012 23196 19068
rect 23196 19012 23252 19068
rect 23252 19012 23256 19068
rect 23192 19008 23256 19012
rect 32952 19068 33016 19072
rect 32952 19012 32956 19068
rect 32956 19012 33012 19068
rect 33012 19012 33016 19068
rect 32952 19008 33016 19012
rect 33032 19068 33096 19072
rect 33032 19012 33036 19068
rect 33036 19012 33092 19068
rect 33092 19012 33096 19068
rect 33032 19008 33096 19012
rect 33112 19068 33176 19072
rect 33112 19012 33116 19068
rect 33116 19012 33172 19068
rect 33172 19012 33176 19068
rect 33112 19008 33176 19012
rect 33192 19068 33256 19072
rect 33192 19012 33196 19068
rect 33196 19012 33252 19068
rect 33252 19012 33256 19068
rect 33192 19008 33256 19012
rect 42952 19068 43016 19072
rect 42952 19012 42956 19068
rect 42956 19012 43012 19068
rect 43012 19012 43016 19068
rect 42952 19008 43016 19012
rect 43032 19068 43096 19072
rect 43032 19012 43036 19068
rect 43036 19012 43092 19068
rect 43092 19012 43096 19068
rect 43032 19008 43096 19012
rect 43112 19068 43176 19072
rect 43112 19012 43116 19068
rect 43116 19012 43172 19068
rect 43172 19012 43176 19068
rect 43112 19008 43176 19012
rect 43192 19068 43256 19072
rect 43192 19012 43196 19068
rect 43196 19012 43252 19068
rect 43252 19012 43256 19068
rect 43192 19008 43256 19012
rect 22692 18804 22756 18868
rect 7952 18524 8016 18528
rect 7952 18468 7956 18524
rect 7956 18468 8012 18524
rect 8012 18468 8016 18524
rect 7952 18464 8016 18468
rect 8032 18524 8096 18528
rect 8032 18468 8036 18524
rect 8036 18468 8092 18524
rect 8092 18468 8096 18524
rect 8032 18464 8096 18468
rect 8112 18524 8176 18528
rect 8112 18468 8116 18524
rect 8116 18468 8172 18524
rect 8172 18468 8176 18524
rect 8112 18464 8176 18468
rect 8192 18524 8256 18528
rect 8192 18468 8196 18524
rect 8196 18468 8252 18524
rect 8252 18468 8256 18524
rect 8192 18464 8256 18468
rect 17952 18524 18016 18528
rect 17952 18468 17956 18524
rect 17956 18468 18012 18524
rect 18012 18468 18016 18524
rect 17952 18464 18016 18468
rect 18032 18524 18096 18528
rect 18032 18468 18036 18524
rect 18036 18468 18092 18524
rect 18092 18468 18096 18524
rect 18032 18464 18096 18468
rect 18112 18524 18176 18528
rect 18112 18468 18116 18524
rect 18116 18468 18172 18524
rect 18172 18468 18176 18524
rect 18112 18464 18176 18468
rect 18192 18524 18256 18528
rect 18192 18468 18196 18524
rect 18196 18468 18252 18524
rect 18252 18468 18256 18524
rect 18192 18464 18256 18468
rect 27952 18524 28016 18528
rect 27952 18468 27956 18524
rect 27956 18468 28012 18524
rect 28012 18468 28016 18524
rect 27952 18464 28016 18468
rect 28032 18524 28096 18528
rect 28032 18468 28036 18524
rect 28036 18468 28092 18524
rect 28092 18468 28096 18524
rect 28032 18464 28096 18468
rect 28112 18524 28176 18528
rect 28112 18468 28116 18524
rect 28116 18468 28172 18524
rect 28172 18468 28176 18524
rect 28112 18464 28176 18468
rect 28192 18524 28256 18528
rect 28192 18468 28196 18524
rect 28196 18468 28252 18524
rect 28252 18468 28256 18524
rect 28192 18464 28256 18468
rect 37952 18524 38016 18528
rect 37952 18468 37956 18524
rect 37956 18468 38012 18524
rect 38012 18468 38016 18524
rect 37952 18464 38016 18468
rect 38032 18524 38096 18528
rect 38032 18468 38036 18524
rect 38036 18468 38092 18524
rect 38092 18468 38096 18524
rect 38032 18464 38096 18468
rect 38112 18524 38176 18528
rect 38112 18468 38116 18524
rect 38116 18468 38172 18524
rect 38172 18468 38176 18524
rect 38112 18464 38176 18468
rect 38192 18524 38256 18528
rect 38192 18468 38196 18524
rect 38196 18468 38252 18524
rect 38252 18468 38256 18524
rect 38192 18464 38256 18468
rect 47952 18524 48016 18528
rect 47952 18468 47956 18524
rect 47956 18468 48012 18524
rect 48012 18468 48016 18524
rect 47952 18464 48016 18468
rect 48032 18524 48096 18528
rect 48032 18468 48036 18524
rect 48036 18468 48092 18524
rect 48092 18468 48096 18524
rect 48032 18464 48096 18468
rect 48112 18524 48176 18528
rect 48112 18468 48116 18524
rect 48116 18468 48172 18524
rect 48172 18468 48176 18524
rect 48112 18464 48176 18468
rect 48192 18524 48256 18528
rect 48192 18468 48196 18524
rect 48196 18468 48252 18524
rect 48252 18468 48256 18524
rect 48192 18464 48256 18468
rect 30972 17988 31036 18052
rect 2952 17980 3016 17984
rect 2952 17924 2956 17980
rect 2956 17924 3012 17980
rect 3012 17924 3016 17980
rect 2952 17920 3016 17924
rect 3032 17980 3096 17984
rect 3032 17924 3036 17980
rect 3036 17924 3092 17980
rect 3092 17924 3096 17980
rect 3032 17920 3096 17924
rect 3112 17980 3176 17984
rect 3112 17924 3116 17980
rect 3116 17924 3172 17980
rect 3172 17924 3176 17980
rect 3112 17920 3176 17924
rect 3192 17980 3256 17984
rect 3192 17924 3196 17980
rect 3196 17924 3252 17980
rect 3252 17924 3256 17980
rect 3192 17920 3256 17924
rect 12952 17980 13016 17984
rect 12952 17924 12956 17980
rect 12956 17924 13012 17980
rect 13012 17924 13016 17980
rect 12952 17920 13016 17924
rect 13032 17980 13096 17984
rect 13032 17924 13036 17980
rect 13036 17924 13092 17980
rect 13092 17924 13096 17980
rect 13032 17920 13096 17924
rect 13112 17980 13176 17984
rect 13112 17924 13116 17980
rect 13116 17924 13172 17980
rect 13172 17924 13176 17980
rect 13112 17920 13176 17924
rect 13192 17980 13256 17984
rect 13192 17924 13196 17980
rect 13196 17924 13252 17980
rect 13252 17924 13256 17980
rect 13192 17920 13256 17924
rect 22952 17980 23016 17984
rect 22952 17924 22956 17980
rect 22956 17924 23012 17980
rect 23012 17924 23016 17980
rect 22952 17920 23016 17924
rect 23032 17980 23096 17984
rect 23032 17924 23036 17980
rect 23036 17924 23092 17980
rect 23092 17924 23096 17980
rect 23032 17920 23096 17924
rect 23112 17980 23176 17984
rect 23112 17924 23116 17980
rect 23116 17924 23172 17980
rect 23172 17924 23176 17980
rect 23112 17920 23176 17924
rect 23192 17980 23256 17984
rect 23192 17924 23196 17980
rect 23196 17924 23252 17980
rect 23252 17924 23256 17980
rect 23192 17920 23256 17924
rect 32952 17980 33016 17984
rect 32952 17924 32956 17980
rect 32956 17924 33012 17980
rect 33012 17924 33016 17980
rect 32952 17920 33016 17924
rect 33032 17980 33096 17984
rect 33032 17924 33036 17980
rect 33036 17924 33092 17980
rect 33092 17924 33096 17980
rect 33032 17920 33096 17924
rect 33112 17980 33176 17984
rect 33112 17924 33116 17980
rect 33116 17924 33172 17980
rect 33172 17924 33176 17980
rect 33112 17920 33176 17924
rect 33192 17980 33256 17984
rect 33192 17924 33196 17980
rect 33196 17924 33252 17980
rect 33252 17924 33256 17980
rect 33192 17920 33256 17924
rect 42952 17980 43016 17984
rect 42952 17924 42956 17980
rect 42956 17924 43012 17980
rect 43012 17924 43016 17980
rect 42952 17920 43016 17924
rect 43032 17980 43096 17984
rect 43032 17924 43036 17980
rect 43036 17924 43092 17980
rect 43092 17924 43096 17980
rect 43032 17920 43096 17924
rect 43112 17980 43176 17984
rect 43112 17924 43116 17980
rect 43116 17924 43172 17980
rect 43172 17924 43176 17980
rect 43112 17920 43176 17924
rect 43192 17980 43256 17984
rect 43192 17924 43196 17980
rect 43196 17924 43252 17980
rect 43252 17924 43256 17980
rect 43192 17920 43256 17924
rect 7952 17436 8016 17440
rect 7952 17380 7956 17436
rect 7956 17380 8012 17436
rect 8012 17380 8016 17436
rect 7952 17376 8016 17380
rect 8032 17436 8096 17440
rect 8032 17380 8036 17436
rect 8036 17380 8092 17436
rect 8092 17380 8096 17436
rect 8032 17376 8096 17380
rect 8112 17436 8176 17440
rect 8112 17380 8116 17436
rect 8116 17380 8172 17436
rect 8172 17380 8176 17436
rect 8112 17376 8176 17380
rect 8192 17436 8256 17440
rect 8192 17380 8196 17436
rect 8196 17380 8252 17436
rect 8252 17380 8256 17436
rect 8192 17376 8256 17380
rect 17952 17436 18016 17440
rect 17952 17380 17956 17436
rect 17956 17380 18012 17436
rect 18012 17380 18016 17436
rect 17952 17376 18016 17380
rect 18032 17436 18096 17440
rect 18032 17380 18036 17436
rect 18036 17380 18092 17436
rect 18092 17380 18096 17436
rect 18032 17376 18096 17380
rect 18112 17436 18176 17440
rect 18112 17380 18116 17436
rect 18116 17380 18172 17436
rect 18172 17380 18176 17436
rect 18112 17376 18176 17380
rect 18192 17436 18256 17440
rect 18192 17380 18196 17436
rect 18196 17380 18252 17436
rect 18252 17380 18256 17436
rect 18192 17376 18256 17380
rect 27952 17436 28016 17440
rect 27952 17380 27956 17436
rect 27956 17380 28012 17436
rect 28012 17380 28016 17436
rect 27952 17376 28016 17380
rect 28032 17436 28096 17440
rect 28032 17380 28036 17436
rect 28036 17380 28092 17436
rect 28092 17380 28096 17436
rect 28032 17376 28096 17380
rect 28112 17436 28176 17440
rect 28112 17380 28116 17436
rect 28116 17380 28172 17436
rect 28172 17380 28176 17436
rect 28112 17376 28176 17380
rect 28192 17436 28256 17440
rect 28192 17380 28196 17436
rect 28196 17380 28252 17436
rect 28252 17380 28256 17436
rect 28192 17376 28256 17380
rect 37952 17436 38016 17440
rect 37952 17380 37956 17436
rect 37956 17380 38012 17436
rect 38012 17380 38016 17436
rect 37952 17376 38016 17380
rect 38032 17436 38096 17440
rect 38032 17380 38036 17436
rect 38036 17380 38092 17436
rect 38092 17380 38096 17436
rect 38032 17376 38096 17380
rect 38112 17436 38176 17440
rect 38112 17380 38116 17436
rect 38116 17380 38172 17436
rect 38172 17380 38176 17436
rect 38112 17376 38176 17380
rect 38192 17436 38256 17440
rect 38192 17380 38196 17436
rect 38196 17380 38252 17436
rect 38252 17380 38256 17436
rect 38192 17376 38256 17380
rect 47952 17436 48016 17440
rect 47952 17380 47956 17436
rect 47956 17380 48012 17436
rect 48012 17380 48016 17436
rect 47952 17376 48016 17380
rect 48032 17436 48096 17440
rect 48032 17380 48036 17436
rect 48036 17380 48092 17436
rect 48092 17380 48096 17436
rect 48032 17376 48096 17380
rect 48112 17436 48176 17440
rect 48112 17380 48116 17436
rect 48116 17380 48172 17436
rect 48172 17380 48176 17436
rect 48112 17376 48176 17380
rect 48192 17436 48256 17440
rect 48192 17380 48196 17436
rect 48196 17380 48252 17436
rect 48252 17380 48256 17436
rect 48192 17376 48256 17380
rect 32812 17308 32876 17372
rect 2952 16892 3016 16896
rect 2952 16836 2956 16892
rect 2956 16836 3012 16892
rect 3012 16836 3016 16892
rect 2952 16832 3016 16836
rect 3032 16892 3096 16896
rect 3032 16836 3036 16892
rect 3036 16836 3092 16892
rect 3092 16836 3096 16892
rect 3032 16832 3096 16836
rect 3112 16892 3176 16896
rect 3112 16836 3116 16892
rect 3116 16836 3172 16892
rect 3172 16836 3176 16892
rect 3112 16832 3176 16836
rect 3192 16892 3256 16896
rect 3192 16836 3196 16892
rect 3196 16836 3252 16892
rect 3252 16836 3256 16892
rect 3192 16832 3256 16836
rect 12952 16892 13016 16896
rect 12952 16836 12956 16892
rect 12956 16836 13012 16892
rect 13012 16836 13016 16892
rect 12952 16832 13016 16836
rect 13032 16892 13096 16896
rect 13032 16836 13036 16892
rect 13036 16836 13092 16892
rect 13092 16836 13096 16892
rect 13032 16832 13096 16836
rect 13112 16892 13176 16896
rect 13112 16836 13116 16892
rect 13116 16836 13172 16892
rect 13172 16836 13176 16892
rect 13112 16832 13176 16836
rect 13192 16892 13256 16896
rect 13192 16836 13196 16892
rect 13196 16836 13252 16892
rect 13252 16836 13256 16892
rect 13192 16832 13256 16836
rect 22952 16892 23016 16896
rect 22952 16836 22956 16892
rect 22956 16836 23012 16892
rect 23012 16836 23016 16892
rect 22952 16832 23016 16836
rect 23032 16892 23096 16896
rect 23032 16836 23036 16892
rect 23036 16836 23092 16892
rect 23092 16836 23096 16892
rect 23032 16832 23096 16836
rect 23112 16892 23176 16896
rect 23112 16836 23116 16892
rect 23116 16836 23172 16892
rect 23172 16836 23176 16892
rect 23112 16832 23176 16836
rect 23192 16892 23256 16896
rect 23192 16836 23196 16892
rect 23196 16836 23252 16892
rect 23252 16836 23256 16892
rect 23192 16832 23256 16836
rect 32952 16892 33016 16896
rect 32952 16836 32956 16892
rect 32956 16836 33012 16892
rect 33012 16836 33016 16892
rect 32952 16832 33016 16836
rect 33032 16892 33096 16896
rect 33032 16836 33036 16892
rect 33036 16836 33092 16892
rect 33092 16836 33096 16892
rect 33032 16832 33096 16836
rect 33112 16892 33176 16896
rect 33112 16836 33116 16892
rect 33116 16836 33172 16892
rect 33172 16836 33176 16892
rect 33112 16832 33176 16836
rect 33192 16892 33256 16896
rect 33192 16836 33196 16892
rect 33196 16836 33252 16892
rect 33252 16836 33256 16892
rect 33192 16832 33256 16836
rect 42952 16892 43016 16896
rect 42952 16836 42956 16892
rect 42956 16836 43012 16892
rect 43012 16836 43016 16892
rect 42952 16832 43016 16836
rect 43032 16892 43096 16896
rect 43032 16836 43036 16892
rect 43036 16836 43092 16892
rect 43092 16836 43096 16892
rect 43032 16832 43096 16836
rect 43112 16892 43176 16896
rect 43112 16836 43116 16892
rect 43116 16836 43172 16892
rect 43172 16836 43176 16892
rect 43112 16832 43176 16836
rect 43192 16892 43256 16896
rect 43192 16836 43196 16892
rect 43196 16836 43252 16892
rect 43252 16836 43256 16892
rect 43192 16832 43256 16836
rect 32628 16628 32692 16692
rect 7952 16348 8016 16352
rect 7952 16292 7956 16348
rect 7956 16292 8012 16348
rect 8012 16292 8016 16348
rect 7952 16288 8016 16292
rect 8032 16348 8096 16352
rect 8032 16292 8036 16348
rect 8036 16292 8092 16348
rect 8092 16292 8096 16348
rect 8032 16288 8096 16292
rect 8112 16348 8176 16352
rect 8112 16292 8116 16348
rect 8116 16292 8172 16348
rect 8172 16292 8176 16348
rect 8112 16288 8176 16292
rect 8192 16348 8256 16352
rect 8192 16292 8196 16348
rect 8196 16292 8252 16348
rect 8252 16292 8256 16348
rect 8192 16288 8256 16292
rect 17952 16348 18016 16352
rect 17952 16292 17956 16348
rect 17956 16292 18012 16348
rect 18012 16292 18016 16348
rect 17952 16288 18016 16292
rect 18032 16348 18096 16352
rect 18032 16292 18036 16348
rect 18036 16292 18092 16348
rect 18092 16292 18096 16348
rect 18032 16288 18096 16292
rect 18112 16348 18176 16352
rect 18112 16292 18116 16348
rect 18116 16292 18172 16348
rect 18172 16292 18176 16348
rect 18112 16288 18176 16292
rect 18192 16348 18256 16352
rect 18192 16292 18196 16348
rect 18196 16292 18252 16348
rect 18252 16292 18256 16348
rect 18192 16288 18256 16292
rect 27952 16348 28016 16352
rect 27952 16292 27956 16348
rect 27956 16292 28012 16348
rect 28012 16292 28016 16348
rect 27952 16288 28016 16292
rect 28032 16348 28096 16352
rect 28032 16292 28036 16348
rect 28036 16292 28092 16348
rect 28092 16292 28096 16348
rect 28032 16288 28096 16292
rect 28112 16348 28176 16352
rect 28112 16292 28116 16348
rect 28116 16292 28172 16348
rect 28172 16292 28176 16348
rect 28112 16288 28176 16292
rect 28192 16348 28256 16352
rect 28192 16292 28196 16348
rect 28196 16292 28252 16348
rect 28252 16292 28256 16348
rect 28192 16288 28256 16292
rect 37952 16348 38016 16352
rect 37952 16292 37956 16348
rect 37956 16292 38012 16348
rect 38012 16292 38016 16348
rect 37952 16288 38016 16292
rect 38032 16348 38096 16352
rect 38032 16292 38036 16348
rect 38036 16292 38092 16348
rect 38092 16292 38096 16348
rect 38032 16288 38096 16292
rect 38112 16348 38176 16352
rect 38112 16292 38116 16348
rect 38116 16292 38172 16348
rect 38172 16292 38176 16348
rect 38112 16288 38176 16292
rect 38192 16348 38256 16352
rect 38192 16292 38196 16348
rect 38196 16292 38252 16348
rect 38252 16292 38256 16348
rect 38192 16288 38256 16292
rect 47952 16348 48016 16352
rect 47952 16292 47956 16348
rect 47956 16292 48012 16348
rect 48012 16292 48016 16348
rect 47952 16288 48016 16292
rect 48032 16348 48096 16352
rect 48032 16292 48036 16348
rect 48036 16292 48092 16348
rect 48092 16292 48096 16348
rect 48032 16288 48096 16292
rect 48112 16348 48176 16352
rect 48112 16292 48116 16348
rect 48116 16292 48172 16348
rect 48172 16292 48176 16348
rect 48112 16288 48176 16292
rect 48192 16348 48256 16352
rect 48192 16292 48196 16348
rect 48196 16292 48252 16348
rect 48252 16292 48256 16348
rect 48192 16288 48256 16292
rect 2952 15804 3016 15808
rect 2952 15748 2956 15804
rect 2956 15748 3012 15804
rect 3012 15748 3016 15804
rect 2952 15744 3016 15748
rect 3032 15804 3096 15808
rect 3032 15748 3036 15804
rect 3036 15748 3092 15804
rect 3092 15748 3096 15804
rect 3032 15744 3096 15748
rect 3112 15804 3176 15808
rect 3112 15748 3116 15804
rect 3116 15748 3172 15804
rect 3172 15748 3176 15804
rect 3112 15744 3176 15748
rect 3192 15804 3256 15808
rect 3192 15748 3196 15804
rect 3196 15748 3252 15804
rect 3252 15748 3256 15804
rect 3192 15744 3256 15748
rect 12952 15804 13016 15808
rect 12952 15748 12956 15804
rect 12956 15748 13012 15804
rect 13012 15748 13016 15804
rect 12952 15744 13016 15748
rect 13032 15804 13096 15808
rect 13032 15748 13036 15804
rect 13036 15748 13092 15804
rect 13092 15748 13096 15804
rect 13032 15744 13096 15748
rect 13112 15804 13176 15808
rect 13112 15748 13116 15804
rect 13116 15748 13172 15804
rect 13172 15748 13176 15804
rect 13112 15744 13176 15748
rect 13192 15804 13256 15808
rect 13192 15748 13196 15804
rect 13196 15748 13252 15804
rect 13252 15748 13256 15804
rect 13192 15744 13256 15748
rect 22952 15804 23016 15808
rect 22952 15748 22956 15804
rect 22956 15748 23012 15804
rect 23012 15748 23016 15804
rect 22952 15744 23016 15748
rect 23032 15804 23096 15808
rect 23032 15748 23036 15804
rect 23036 15748 23092 15804
rect 23092 15748 23096 15804
rect 23032 15744 23096 15748
rect 23112 15804 23176 15808
rect 23112 15748 23116 15804
rect 23116 15748 23172 15804
rect 23172 15748 23176 15804
rect 23112 15744 23176 15748
rect 23192 15804 23256 15808
rect 23192 15748 23196 15804
rect 23196 15748 23252 15804
rect 23252 15748 23256 15804
rect 23192 15744 23256 15748
rect 32952 15804 33016 15808
rect 32952 15748 32956 15804
rect 32956 15748 33012 15804
rect 33012 15748 33016 15804
rect 32952 15744 33016 15748
rect 33032 15804 33096 15808
rect 33032 15748 33036 15804
rect 33036 15748 33092 15804
rect 33092 15748 33096 15804
rect 33032 15744 33096 15748
rect 33112 15804 33176 15808
rect 33112 15748 33116 15804
rect 33116 15748 33172 15804
rect 33172 15748 33176 15804
rect 33112 15744 33176 15748
rect 33192 15804 33256 15808
rect 33192 15748 33196 15804
rect 33196 15748 33252 15804
rect 33252 15748 33256 15804
rect 33192 15744 33256 15748
rect 42952 15804 43016 15808
rect 42952 15748 42956 15804
rect 42956 15748 43012 15804
rect 43012 15748 43016 15804
rect 42952 15744 43016 15748
rect 43032 15804 43096 15808
rect 43032 15748 43036 15804
rect 43036 15748 43092 15804
rect 43092 15748 43096 15804
rect 43032 15744 43096 15748
rect 43112 15804 43176 15808
rect 43112 15748 43116 15804
rect 43116 15748 43172 15804
rect 43172 15748 43176 15804
rect 43112 15744 43176 15748
rect 43192 15804 43256 15808
rect 43192 15748 43196 15804
rect 43196 15748 43252 15804
rect 43252 15748 43256 15804
rect 43192 15744 43256 15748
rect 7952 15260 8016 15264
rect 7952 15204 7956 15260
rect 7956 15204 8012 15260
rect 8012 15204 8016 15260
rect 7952 15200 8016 15204
rect 8032 15260 8096 15264
rect 8032 15204 8036 15260
rect 8036 15204 8092 15260
rect 8092 15204 8096 15260
rect 8032 15200 8096 15204
rect 8112 15260 8176 15264
rect 8112 15204 8116 15260
rect 8116 15204 8172 15260
rect 8172 15204 8176 15260
rect 8112 15200 8176 15204
rect 8192 15260 8256 15264
rect 8192 15204 8196 15260
rect 8196 15204 8252 15260
rect 8252 15204 8256 15260
rect 8192 15200 8256 15204
rect 17952 15260 18016 15264
rect 17952 15204 17956 15260
rect 17956 15204 18012 15260
rect 18012 15204 18016 15260
rect 17952 15200 18016 15204
rect 18032 15260 18096 15264
rect 18032 15204 18036 15260
rect 18036 15204 18092 15260
rect 18092 15204 18096 15260
rect 18032 15200 18096 15204
rect 18112 15260 18176 15264
rect 18112 15204 18116 15260
rect 18116 15204 18172 15260
rect 18172 15204 18176 15260
rect 18112 15200 18176 15204
rect 18192 15260 18256 15264
rect 18192 15204 18196 15260
rect 18196 15204 18252 15260
rect 18252 15204 18256 15260
rect 18192 15200 18256 15204
rect 27952 15260 28016 15264
rect 27952 15204 27956 15260
rect 27956 15204 28012 15260
rect 28012 15204 28016 15260
rect 27952 15200 28016 15204
rect 28032 15260 28096 15264
rect 28032 15204 28036 15260
rect 28036 15204 28092 15260
rect 28092 15204 28096 15260
rect 28032 15200 28096 15204
rect 28112 15260 28176 15264
rect 28112 15204 28116 15260
rect 28116 15204 28172 15260
rect 28172 15204 28176 15260
rect 28112 15200 28176 15204
rect 28192 15260 28256 15264
rect 28192 15204 28196 15260
rect 28196 15204 28252 15260
rect 28252 15204 28256 15260
rect 28192 15200 28256 15204
rect 37952 15260 38016 15264
rect 37952 15204 37956 15260
rect 37956 15204 38012 15260
rect 38012 15204 38016 15260
rect 37952 15200 38016 15204
rect 38032 15260 38096 15264
rect 38032 15204 38036 15260
rect 38036 15204 38092 15260
rect 38092 15204 38096 15260
rect 38032 15200 38096 15204
rect 38112 15260 38176 15264
rect 38112 15204 38116 15260
rect 38116 15204 38172 15260
rect 38172 15204 38176 15260
rect 38112 15200 38176 15204
rect 38192 15260 38256 15264
rect 38192 15204 38196 15260
rect 38196 15204 38252 15260
rect 38252 15204 38256 15260
rect 38192 15200 38256 15204
rect 47952 15260 48016 15264
rect 47952 15204 47956 15260
rect 47956 15204 48012 15260
rect 48012 15204 48016 15260
rect 47952 15200 48016 15204
rect 48032 15260 48096 15264
rect 48032 15204 48036 15260
rect 48036 15204 48092 15260
rect 48092 15204 48096 15260
rect 48032 15200 48096 15204
rect 48112 15260 48176 15264
rect 48112 15204 48116 15260
rect 48116 15204 48172 15260
rect 48172 15204 48176 15260
rect 48112 15200 48176 15204
rect 48192 15260 48256 15264
rect 48192 15204 48196 15260
rect 48196 15204 48252 15260
rect 48252 15204 48256 15260
rect 48192 15200 48256 15204
rect 2952 14716 3016 14720
rect 2952 14660 2956 14716
rect 2956 14660 3012 14716
rect 3012 14660 3016 14716
rect 2952 14656 3016 14660
rect 3032 14716 3096 14720
rect 3032 14660 3036 14716
rect 3036 14660 3092 14716
rect 3092 14660 3096 14716
rect 3032 14656 3096 14660
rect 3112 14716 3176 14720
rect 3112 14660 3116 14716
rect 3116 14660 3172 14716
rect 3172 14660 3176 14716
rect 3112 14656 3176 14660
rect 3192 14716 3256 14720
rect 3192 14660 3196 14716
rect 3196 14660 3252 14716
rect 3252 14660 3256 14716
rect 3192 14656 3256 14660
rect 12952 14716 13016 14720
rect 12952 14660 12956 14716
rect 12956 14660 13012 14716
rect 13012 14660 13016 14716
rect 12952 14656 13016 14660
rect 13032 14716 13096 14720
rect 13032 14660 13036 14716
rect 13036 14660 13092 14716
rect 13092 14660 13096 14716
rect 13032 14656 13096 14660
rect 13112 14716 13176 14720
rect 13112 14660 13116 14716
rect 13116 14660 13172 14716
rect 13172 14660 13176 14716
rect 13112 14656 13176 14660
rect 13192 14716 13256 14720
rect 13192 14660 13196 14716
rect 13196 14660 13252 14716
rect 13252 14660 13256 14716
rect 13192 14656 13256 14660
rect 22952 14716 23016 14720
rect 22952 14660 22956 14716
rect 22956 14660 23012 14716
rect 23012 14660 23016 14716
rect 22952 14656 23016 14660
rect 23032 14716 23096 14720
rect 23032 14660 23036 14716
rect 23036 14660 23092 14716
rect 23092 14660 23096 14716
rect 23032 14656 23096 14660
rect 23112 14716 23176 14720
rect 23112 14660 23116 14716
rect 23116 14660 23172 14716
rect 23172 14660 23176 14716
rect 23112 14656 23176 14660
rect 23192 14716 23256 14720
rect 23192 14660 23196 14716
rect 23196 14660 23252 14716
rect 23252 14660 23256 14716
rect 23192 14656 23256 14660
rect 32952 14716 33016 14720
rect 32952 14660 32956 14716
rect 32956 14660 33012 14716
rect 33012 14660 33016 14716
rect 32952 14656 33016 14660
rect 33032 14716 33096 14720
rect 33032 14660 33036 14716
rect 33036 14660 33092 14716
rect 33092 14660 33096 14716
rect 33032 14656 33096 14660
rect 33112 14716 33176 14720
rect 33112 14660 33116 14716
rect 33116 14660 33172 14716
rect 33172 14660 33176 14716
rect 33112 14656 33176 14660
rect 33192 14716 33256 14720
rect 33192 14660 33196 14716
rect 33196 14660 33252 14716
rect 33252 14660 33256 14716
rect 33192 14656 33256 14660
rect 42952 14716 43016 14720
rect 42952 14660 42956 14716
rect 42956 14660 43012 14716
rect 43012 14660 43016 14716
rect 42952 14656 43016 14660
rect 43032 14716 43096 14720
rect 43032 14660 43036 14716
rect 43036 14660 43092 14716
rect 43092 14660 43096 14716
rect 43032 14656 43096 14660
rect 43112 14716 43176 14720
rect 43112 14660 43116 14716
rect 43116 14660 43172 14716
rect 43172 14660 43176 14716
rect 43112 14656 43176 14660
rect 43192 14716 43256 14720
rect 43192 14660 43196 14716
rect 43196 14660 43252 14716
rect 43252 14660 43256 14716
rect 43192 14656 43256 14660
rect 7952 14172 8016 14176
rect 7952 14116 7956 14172
rect 7956 14116 8012 14172
rect 8012 14116 8016 14172
rect 7952 14112 8016 14116
rect 8032 14172 8096 14176
rect 8032 14116 8036 14172
rect 8036 14116 8092 14172
rect 8092 14116 8096 14172
rect 8032 14112 8096 14116
rect 8112 14172 8176 14176
rect 8112 14116 8116 14172
rect 8116 14116 8172 14172
rect 8172 14116 8176 14172
rect 8112 14112 8176 14116
rect 8192 14172 8256 14176
rect 8192 14116 8196 14172
rect 8196 14116 8252 14172
rect 8252 14116 8256 14172
rect 8192 14112 8256 14116
rect 17952 14172 18016 14176
rect 17952 14116 17956 14172
rect 17956 14116 18012 14172
rect 18012 14116 18016 14172
rect 17952 14112 18016 14116
rect 18032 14172 18096 14176
rect 18032 14116 18036 14172
rect 18036 14116 18092 14172
rect 18092 14116 18096 14172
rect 18032 14112 18096 14116
rect 18112 14172 18176 14176
rect 18112 14116 18116 14172
rect 18116 14116 18172 14172
rect 18172 14116 18176 14172
rect 18112 14112 18176 14116
rect 18192 14172 18256 14176
rect 18192 14116 18196 14172
rect 18196 14116 18252 14172
rect 18252 14116 18256 14172
rect 18192 14112 18256 14116
rect 27952 14172 28016 14176
rect 27952 14116 27956 14172
rect 27956 14116 28012 14172
rect 28012 14116 28016 14172
rect 27952 14112 28016 14116
rect 28032 14172 28096 14176
rect 28032 14116 28036 14172
rect 28036 14116 28092 14172
rect 28092 14116 28096 14172
rect 28032 14112 28096 14116
rect 28112 14172 28176 14176
rect 28112 14116 28116 14172
rect 28116 14116 28172 14172
rect 28172 14116 28176 14172
rect 28112 14112 28176 14116
rect 28192 14172 28256 14176
rect 28192 14116 28196 14172
rect 28196 14116 28252 14172
rect 28252 14116 28256 14172
rect 28192 14112 28256 14116
rect 37952 14172 38016 14176
rect 37952 14116 37956 14172
rect 37956 14116 38012 14172
rect 38012 14116 38016 14172
rect 37952 14112 38016 14116
rect 38032 14172 38096 14176
rect 38032 14116 38036 14172
rect 38036 14116 38092 14172
rect 38092 14116 38096 14172
rect 38032 14112 38096 14116
rect 38112 14172 38176 14176
rect 38112 14116 38116 14172
rect 38116 14116 38172 14172
rect 38172 14116 38176 14172
rect 38112 14112 38176 14116
rect 38192 14172 38256 14176
rect 38192 14116 38196 14172
rect 38196 14116 38252 14172
rect 38252 14116 38256 14172
rect 38192 14112 38256 14116
rect 47952 14172 48016 14176
rect 47952 14116 47956 14172
rect 47956 14116 48012 14172
rect 48012 14116 48016 14172
rect 47952 14112 48016 14116
rect 48032 14172 48096 14176
rect 48032 14116 48036 14172
rect 48036 14116 48092 14172
rect 48092 14116 48096 14172
rect 48032 14112 48096 14116
rect 48112 14172 48176 14176
rect 48112 14116 48116 14172
rect 48116 14116 48172 14172
rect 48172 14116 48176 14172
rect 48112 14112 48176 14116
rect 48192 14172 48256 14176
rect 48192 14116 48196 14172
rect 48196 14116 48252 14172
rect 48252 14116 48256 14172
rect 48192 14112 48256 14116
rect 2952 13628 3016 13632
rect 2952 13572 2956 13628
rect 2956 13572 3012 13628
rect 3012 13572 3016 13628
rect 2952 13568 3016 13572
rect 3032 13628 3096 13632
rect 3032 13572 3036 13628
rect 3036 13572 3092 13628
rect 3092 13572 3096 13628
rect 3032 13568 3096 13572
rect 3112 13628 3176 13632
rect 3112 13572 3116 13628
rect 3116 13572 3172 13628
rect 3172 13572 3176 13628
rect 3112 13568 3176 13572
rect 3192 13628 3256 13632
rect 3192 13572 3196 13628
rect 3196 13572 3252 13628
rect 3252 13572 3256 13628
rect 3192 13568 3256 13572
rect 12952 13628 13016 13632
rect 12952 13572 12956 13628
rect 12956 13572 13012 13628
rect 13012 13572 13016 13628
rect 12952 13568 13016 13572
rect 13032 13628 13096 13632
rect 13032 13572 13036 13628
rect 13036 13572 13092 13628
rect 13092 13572 13096 13628
rect 13032 13568 13096 13572
rect 13112 13628 13176 13632
rect 13112 13572 13116 13628
rect 13116 13572 13172 13628
rect 13172 13572 13176 13628
rect 13112 13568 13176 13572
rect 13192 13628 13256 13632
rect 13192 13572 13196 13628
rect 13196 13572 13252 13628
rect 13252 13572 13256 13628
rect 13192 13568 13256 13572
rect 22952 13628 23016 13632
rect 22952 13572 22956 13628
rect 22956 13572 23012 13628
rect 23012 13572 23016 13628
rect 22952 13568 23016 13572
rect 23032 13628 23096 13632
rect 23032 13572 23036 13628
rect 23036 13572 23092 13628
rect 23092 13572 23096 13628
rect 23032 13568 23096 13572
rect 23112 13628 23176 13632
rect 23112 13572 23116 13628
rect 23116 13572 23172 13628
rect 23172 13572 23176 13628
rect 23112 13568 23176 13572
rect 23192 13628 23256 13632
rect 23192 13572 23196 13628
rect 23196 13572 23252 13628
rect 23252 13572 23256 13628
rect 23192 13568 23256 13572
rect 32952 13628 33016 13632
rect 32952 13572 32956 13628
rect 32956 13572 33012 13628
rect 33012 13572 33016 13628
rect 32952 13568 33016 13572
rect 33032 13628 33096 13632
rect 33032 13572 33036 13628
rect 33036 13572 33092 13628
rect 33092 13572 33096 13628
rect 33032 13568 33096 13572
rect 33112 13628 33176 13632
rect 33112 13572 33116 13628
rect 33116 13572 33172 13628
rect 33172 13572 33176 13628
rect 33112 13568 33176 13572
rect 33192 13628 33256 13632
rect 33192 13572 33196 13628
rect 33196 13572 33252 13628
rect 33252 13572 33256 13628
rect 33192 13568 33256 13572
rect 42952 13628 43016 13632
rect 42952 13572 42956 13628
rect 42956 13572 43012 13628
rect 43012 13572 43016 13628
rect 42952 13568 43016 13572
rect 43032 13628 43096 13632
rect 43032 13572 43036 13628
rect 43036 13572 43092 13628
rect 43092 13572 43096 13628
rect 43032 13568 43096 13572
rect 43112 13628 43176 13632
rect 43112 13572 43116 13628
rect 43116 13572 43172 13628
rect 43172 13572 43176 13628
rect 43112 13568 43176 13572
rect 43192 13628 43256 13632
rect 43192 13572 43196 13628
rect 43196 13572 43252 13628
rect 43252 13572 43256 13628
rect 43192 13568 43256 13572
rect 7952 13084 8016 13088
rect 7952 13028 7956 13084
rect 7956 13028 8012 13084
rect 8012 13028 8016 13084
rect 7952 13024 8016 13028
rect 8032 13084 8096 13088
rect 8032 13028 8036 13084
rect 8036 13028 8092 13084
rect 8092 13028 8096 13084
rect 8032 13024 8096 13028
rect 8112 13084 8176 13088
rect 8112 13028 8116 13084
rect 8116 13028 8172 13084
rect 8172 13028 8176 13084
rect 8112 13024 8176 13028
rect 8192 13084 8256 13088
rect 8192 13028 8196 13084
rect 8196 13028 8252 13084
rect 8252 13028 8256 13084
rect 8192 13024 8256 13028
rect 17952 13084 18016 13088
rect 17952 13028 17956 13084
rect 17956 13028 18012 13084
rect 18012 13028 18016 13084
rect 17952 13024 18016 13028
rect 18032 13084 18096 13088
rect 18032 13028 18036 13084
rect 18036 13028 18092 13084
rect 18092 13028 18096 13084
rect 18032 13024 18096 13028
rect 18112 13084 18176 13088
rect 18112 13028 18116 13084
rect 18116 13028 18172 13084
rect 18172 13028 18176 13084
rect 18112 13024 18176 13028
rect 18192 13084 18256 13088
rect 18192 13028 18196 13084
rect 18196 13028 18252 13084
rect 18252 13028 18256 13084
rect 18192 13024 18256 13028
rect 27952 13084 28016 13088
rect 27952 13028 27956 13084
rect 27956 13028 28012 13084
rect 28012 13028 28016 13084
rect 27952 13024 28016 13028
rect 28032 13084 28096 13088
rect 28032 13028 28036 13084
rect 28036 13028 28092 13084
rect 28092 13028 28096 13084
rect 28032 13024 28096 13028
rect 28112 13084 28176 13088
rect 28112 13028 28116 13084
rect 28116 13028 28172 13084
rect 28172 13028 28176 13084
rect 28112 13024 28176 13028
rect 28192 13084 28256 13088
rect 28192 13028 28196 13084
rect 28196 13028 28252 13084
rect 28252 13028 28256 13084
rect 28192 13024 28256 13028
rect 37952 13084 38016 13088
rect 37952 13028 37956 13084
rect 37956 13028 38012 13084
rect 38012 13028 38016 13084
rect 37952 13024 38016 13028
rect 38032 13084 38096 13088
rect 38032 13028 38036 13084
rect 38036 13028 38092 13084
rect 38092 13028 38096 13084
rect 38032 13024 38096 13028
rect 38112 13084 38176 13088
rect 38112 13028 38116 13084
rect 38116 13028 38172 13084
rect 38172 13028 38176 13084
rect 38112 13024 38176 13028
rect 38192 13084 38256 13088
rect 38192 13028 38196 13084
rect 38196 13028 38252 13084
rect 38252 13028 38256 13084
rect 38192 13024 38256 13028
rect 47952 13084 48016 13088
rect 47952 13028 47956 13084
rect 47956 13028 48012 13084
rect 48012 13028 48016 13084
rect 47952 13024 48016 13028
rect 48032 13084 48096 13088
rect 48032 13028 48036 13084
rect 48036 13028 48092 13084
rect 48092 13028 48096 13084
rect 48032 13024 48096 13028
rect 48112 13084 48176 13088
rect 48112 13028 48116 13084
rect 48116 13028 48172 13084
rect 48172 13028 48176 13084
rect 48112 13024 48176 13028
rect 48192 13084 48256 13088
rect 48192 13028 48196 13084
rect 48196 13028 48252 13084
rect 48252 13028 48256 13084
rect 48192 13024 48256 13028
rect 2952 12540 3016 12544
rect 2952 12484 2956 12540
rect 2956 12484 3012 12540
rect 3012 12484 3016 12540
rect 2952 12480 3016 12484
rect 3032 12540 3096 12544
rect 3032 12484 3036 12540
rect 3036 12484 3092 12540
rect 3092 12484 3096 12540
rect 3032 12480 3096 12484
rect 3112 12540 3176 12544
rect 3112 12484 3116 12540
rect 3116 12484 3172 12540
rect 3172 12484 3176 12540
rect 3112 12480 3176 12484
rect 3192 12540 3256 12544
rect 3192 12484 3196 12540
rect 3196 12484 3252 12540
rect 3252 12484 3256 12540
rect 3192 12480 3256 12484
rect 12952 12540 13016 12544
rect 12952 12484 12956 12540
rect 12956 12484 13012 12540
rect 13012 12484 13016 12540
rect 12952 12480 13016 12484
rect 13032 12540 13096 12544
rect 13032 12484 13036 12540
rect 13036 12484 13092 12540
rect 13092 12484 13096 12540
rect 13032 12480 13096 12484
rect 13112 12540 13176 12544
rect 13112 12484 13116 12540
rect 13116 12484 13172 12540
rect 13172 12484 13176 12540
rect 13112 12480 13176 12484
rect 13192 12540 13256 12544
rect 13192 12484 13196 12540
rect 13196 12484 13252 12540
rect 13252 12484 13256 12540
rect 13192 12480 13256 12484
rect 22952 12540 23016 12544
rect 22952 12484 22956 12540
rect 22956 12484 23012 12540
rect 23012 12484 23016 12540
rect 22952 12480 23016 12484
rect 23032 12540 23096 12544
rect 23032 12484 23036 12540
rect 23036 12484 23092 12540
rect 23092 12484 23096 12540
rect 23032 12480 23096 12484
rect 23112 12540 23176 12544
rect 23112 12484 23116 12540
rect 23116 12484 23172 12540
rect 23172 12484 23176 12540
rect 23112 12480 23176 12484
rect 23192 12540 23256 12544
rect 23192 12484 23196 12540
rect 23196 12484 23252 12540
rect 23252 12484 23256 12540
rect 23192 12480 23256 12484
rect 32952 12540 33016 12544
rect 32952 12484 32956 12540
rect 32956 12484 33012 12540
rect 33012 12484 33016 12540
rect 32952 12480 33016 12484
rect 33032 12540 33096 12544
rect 33032 12484 33036 12540
rect 33036 12484 33092 12540
rect 33092 12484 33096 12540
rect 33032 12480 33096 12484
rect 33112 12540 33176 12544
rect 33112 12484 33116 12540
rect 33116 12484 33172 12540
rect 33172 12484 33176 12540
rect 33112 12480 33176 12484
rect 33192 12540 33256 12544
rect 33192 12484 33196 12540
rect 33196 12484 33252 12540
rect 33252 12484 33256 12540
rect 33192 12480 33256 12484
rect 42952 12540 43016 12544
rect 42952 12484 42956 12540
rect 42956 12484 43012 12540
rect 43012 12484 43016 12540
rect 42952 12480 43016 12484
rect 43032 12540 43096 12544
rect 43032 12484 43036 12540
rect 43036 12484 43092 12540
rect 43092 12484 43096 12540
rect 43032 12480 43096 12484
rect 43112 12540 43176 12544
rect 43112 12484 43116 12540
rect 43116 12484 43172 12540
rect 43172 12484 43176 12540
rect 43112 12480 43176 12484
rect 43192 12540 43256 12544
rect 43192 12484 43196 12540
rect 43196 12484 43252 12540
rect 43252 12484 43256 12540
rect 43192 12480 43256 12484
rect 38516 12276 38580 12340
rect 7952 11996 8016 12000
rect 7952 11940 7956 11996
rect 7956 11940 8012 11996
rect 8012 11940 8016 11996
rect 7952 11936 8016 11940
rect 8032 11996 8096 12000
rect 8032 11940 8036 11996
rect 8036 11940 8092 11996
rect 8092 11940 8096 11996
rect 8032 11936 8096 11940
rect 8112 11996 8176 12000
rect 8112 11940 8116 11996
rect 8116 11940 8172 11996
rect 8172 11940 8176 11996
rect 8112 11936 8176 11940
rect 8192 11996 8256 12000
rect 8192 11940 8196 11996
rect 8196 11940 8252 11996
rect 8252 11940 8256 11996
rect 8192 11936 8256 11940
rect 17952 11996 18016 12000
rect 17952 11940 17956 11996
rect 17956 11940 18012 11996
rect 18012 11940 18016 11996
rect 17952 11936 18016 11940
rect 18032 11996 18096 12000
rect 18032 11940 18036 11996
rect 18036 11940 18092 11996
rect 18092 11940 18096 11996
rect 18032 11936 18096 11940
rect 18112 11996 18176 12000
rect 18112 11940 18116 11996
rect 18116 11940 18172 11996
rect 18172 11940 18176 11996
rect 18112 11936 18176 11940
rect 18192 11996 18256 12000
rect 18192 11940 18196 11996
rect 18196 11940 18252 11996
rect 18252 11940 18256 11996
rect 18192 11936 18256 11940
rect 27952 11996 28016 12000
rect 27952 11940 27956 11996
rect 27956 11940 28012 11996
rect 28012 11940 28016 11996
rect 27952 11936 28016 11940
rect 28032 11996 28096 12000
rect 28032 11940 28036 11996
rect 28036 11940 28092 11996
rect 28092 11940 28096 11996
rect 28032 11936 28096 11940
rect 28112 11996 28176 12000
rect 28112 11940 28116 11996
rect 28116 11940 28172 11996
rect 28172 11940 28176 11996
rect 28112 11936 28176 11940
rect 28192 11996 28256 12000
rect 28192 11940 28196 11996
rect 28196 11940 28252 11996
rect 28252 11940 28256 11996
rect 28192 11936 28256 11940
rect 37952 11996 38016 12000
rect 37952 11940 37956 11996
rect 37956 11940 38012 11996
rect 38012 11940 38016 11996
rect 37952 11936 38016 11940
rect 38032 11996 38096 12000
rect 38032 11940 38036 11996
rect 38036 11940 38092 11996
rect 38092 11940 38096 11996
rect 38032 11936 38096 11940
rect 38112 11996 38176 12000
rect 38112 11940 38116 11996
rect 38116 11940 38172 11996
rect 38172 11940 38176 11996
rect 38112 11936 38176 11940
rect 38192 11996 38256 12000
rect 38192 11940 38196 11996
rect 38196 11940 38252 11996
rect 38252 11940 38256 11996
rect 38192 11936 38256 11940
rect 47952 11996 48016 12000
rect 47952 11940 47956 11996
rect 47956 11940 48012 11996
rect 48012 11940 48016 11996
rect 47952 11936 48016 11940
rect 48032 11996 48096 12000
rect 48032 11940 48036 11996
rect 48036 11940 48092 11996
rect 48092 11940 48096 11996
rect 48032 11936 48096 11940
rect 48112 11996 48176 12000
rect 48112 11940 48116 11996
rect 48116 11940 48172 11996
rect 48172 11940 48176 11996
rect 48112 11936 48176 11940
rect 48192 11996 48256 12000
rect 48192 11940 48196 11996
rect 48196 11940 48252 11996
rect 48252 11940 48256 11996
rect 48192 11936 48256 11940
rect 2952 11452 3016 11456
rect 2952 11396 2956 11452
rect 2956 11396 3012 11452
rect 3012 11396 3016 11452
rect 2952 11392 3016 11396
rect 3032 11452 3096 11456
rect 3032 11396 3036 11452
rect 3036 11396 3092 11452
rect 3092 11396 3096 11452
rect 3032 11392 3096 11396
rect 3112 11452 3176 11456
rect 3112 11396 3116 11452
rect 3116 11396 3172 11452
rect 3172 11396 3176 11452
rect 3112 11392 3176 11396
rect 3192 11452 3256 11456
rect 3192 11396 3196 11452
rect 3196 11396 3252 11452
rect 3252 11396 3256 11452
rect 3192 11392 3256 11396
rect 12952 11452 13016 11456
rect 12952 11396 12956 11452
rect 12956 11396 13012 11452
rect 13012 11396 13016 11452
rect 12952 11392 13016 11396
rect 13032 11452 13096 11456
rect 13032 11396 13036 11452
rect 13036 11396 13092 11452
rect 13092 11396 13096 11452
rect 13032 11392 13096 11396
rect 13112 11452 13176 11456
rect 13112 11396 13116 11452
rect 13116 11396 13172 11452
rect 13172 11396 13176 11452
rect 13112 11392 13176 11396
rect 13192 11452 13256 11456
rect 13192 11396 13196 11452
rect 13196 11396 13252 11452
rect 13252 11396 13256 11452
rect 13192 11392 13256 11396
rect 22952 11452 23016 11456
rect 22952 11396 22956 11452
rect 22956 11396 23012 11452
rect 23012 11396 23016 11452
rect 22952 11392 23016 11396
rect 23032 11452 23096 11456
rect 23032 11396 23036 11452
rect 23036 11396 23092 11452
rect 23092 11396 23096 11452
rect 23032 11392 23096 11396
rect 23112 11452 23176 11456
rect 23112 11396 23116 11452
rect 23116 11396 23172 11452
rect 23172 11396 23176 11452
rect 23112 11392 23176 11396
rect 23192 11452 23256 11456
rect 23192 11396 23196 11452
rect 23196 11396 23252 11452
rect 23252 11396 23256 11452
rect 23192 11392 23256 11396
rect 32952 11452 33016 11456
rect 32952 11396 32956 11452
rect 32956 11396 33012 11452
rect 33012 11396 33016 11452
rect 32952 11392 33016 11396
rect 33032 11452 33096 11456
rect 33032 11396 33036 11452
rect 33036 11396 33092 11452
rect 33092 11396 33096 11452
rect 33032 11392 33096 11396
rect 33112 11452 33176 11456
rect 33112 11396 33116 11452
rect 33116 11396 33172 11452
rect 33172 11396 33176 11452
rect 33112 11392 33176 11396
rect 33192 11452 33256 11456
rect 33192 11396 33196 11452
rect 33196 11396 33252 11452
rect 33252 11396 33256 11452
rect 33192 11392 33256 11396
rect 42952 11452 43016 11456
rect 42952 11396 42956 11452
rect 42956 11396 43012 11452
rect 43012 11396 43016 11452
rect 42952 11392 43016 11396
rect 43032 11452 43096 11456
rect 43032 11396 43036 11452
rect 43036 11396 43092 11452
rect 43092 11396 43096 11452
rect 43032 11392 43096 11396
rect 43112 11452 43176 11456
rect 43112 11396 43116 11452
rect 43116 11396 43172 11452
rect 43172 11396 43176 11452
rect 43112 11392 43176 11396
rect 43192 11452 43256 11456
rect 43192 11396 43196 11452
rect 43196 11396 43252 11452
rect 43252 11396 43256 11452
rect 43192 11392 43256 11396
rect 7952 10908 8016 10912
rect 7952 10852 7956 10908
rect 7956 10852 8012 10908
rect 8012 10852 8016 10908
rect 7952 10848 8016 10852
rect 8032 10908 8096 10912
rect 8032 10852 8036 10908
rect 8036 10852 8092 10908
rect 8092 10852 8096 10908
rect 8032 10848 8096 10852
rect 8112 10908 8176 10912
rect 8112 10852 8116 10908
rect 8116 10852 8172 10908
rect 8172 10852 8176 10908
rect 8112 10848 8176 10852
rect 8192 10908 8256 10912
rect 8192 10852 8196 10908
rect 8196 10852 8252 10908
rect 8252 10852 8256 10908
rect 8192 10848 8256 10852
rect 17952 10908 18016 10912
rect 17952 10852 17956 10908
rect 17956 10852 18012 10908
rect 18012 10852 18016 10908
rect 17952 10848 18016 10852
rect 18032 10908 18096 10912
rect 18032 10852 18036 10908
rect 18036 10852 18092 10908
rect 18092 10852 18096 10908
rect 18032 10848 18096 10852
rect 18112 10908 18176 10912
rect 18112 10852 18116 10908
rect 18116 10852 18172 10908
rect 18172 10852 18176 10908
rect 18112 10848 18176 10852
rect 18192 10908 18256 10912
rect 18192 10852 18196 10908
rect 18196 10852 18252 10908
rect 18252 10852 18256 10908
rect 18192 10848 18256 10852
rect 27952 10908 28016 10912
rect 27952 10852 27956 10908
rect 27956 10852 28012 10908
rect 28012 10852 28016 10908
rect 27952 10848 28016 10852
rect 28032 10908 28096 10912
rect 28032 10852 28036 10908
rect 28036 10852 28092 10908
rect 28092 10852 28096 10908
rect 28032 10848 28096 10852
rect 28112 10908 28176 10912
rect 28112 10852 28116 10908
rect 28116 10852 28172 10908
rect 28172 10852 28176 10908
rect 28112 10848 28176 10852
rect 28192 10908 28256 10912
rect 28192 10852 28196 10908
rect 28196 10852 28252 10908
rect 28252 10852 28256 10908
rect 28192 10848 28256 10852
rect 37952 10908 38016 10912
rect 37952 10852 37956 10908
rect 37956 10852 38012 10908
rect 38012 10852 38016 10908
rect 37952 10848 38016 10852
rect 38032 10908 38096 10912
rect 38032 10852 38036 10908
rect 38036 10852 38092 10908
rect 38092 10852 38096 10908
rect 38032 10848 38096 10852
rect 38112 10908 38176 10912
rect 38112 10852 38116 10908
rect 38116 10852 38172 10908
rect 38172 10852 38176 10908
rect 38112 10848 38176 10852
rect 38192 10908 38256 10912
rect 38192 10852 38196 10908
rect 38196 10852 38252 10908
rect 38252 10852 38256 10908
rect 38192 10848 38256 10852
rect 47952 10908 48016 10912
rect 47952 10852 47956 10908
rect 47956 10852 48012 10908
rect 48012 10852 48016 10908
rect 47952 10848 48016 10852
rect 48032 10908 48096 10912
rect 48032 10852 48036 10908
rect 48036 10852 48092 10908
rect 48092 10852 48096 10908
rect 48032 10848 48096 10852
rect 48112 10908 48176 10912
rect 48112 10852 48116 10908
rect 48116 10852 48172 10908
rect 48172 10852 48176 10908
rect 48112 10848 48176 10852
rect 48192 10908 48256 10912
rect 48192 10852 48196 10908
rect 48196 10852 48252 10908
rect 48252 10852 48256 10908
rect 48192 10848 48256 10852
rect 2952 10364 3016 10368
rect 2952 10308 2956 10364
rect 2956 10308 3012 10364
rect 3012 10308 3016 10364
rect 2952 10304 3016 10308
rect 3032 10364 3096 10368
rect 3032 10308 3036 10364
rect 3036 10308 3092 10364
rect 3092 10308 3096 10364
rect 3032 10304 3096 10308
rect 3112 10364 3176 10368
rect 3112 10308 3116 10364
rect 3116 10308 3172 10364
rect 3172 10308 3176 10364
rect 3112 10304 3176 10308
rect 3192 10364 3256 10368
rect 3192 10308 3196 10364
rect 3196 10308 3252 10364
rect 3252 10308 3256 10364
rect 3192 10304 3256 10308
rect 12952 10364 13016 10368
rect 12952 10308 12956 10364
rect 12956 10308 13012 10364
rect 13012 10308 13016 10364
rect 12952 10304 13016 10308
rect 13032 10364 13096 10368
rect 13032 10308 13036 10364
rect 13036 10308 13092 10364
rect 13092 10308 13096 10364
rect 13032 10304 13096 10308
rect 13112 10364 13176 10368
rect 13112 10308 13116 10364
rect 13116 10308 13172 10364
rect 13172 10308 13176 10364
rect 13112 10304 13176 10308
rect 13192 10364 13256 10368
rect 13192 10308 13196 10364
rect 13196 10308 13252 10364
rect 13252 10308 13256 10364
rect 13192 10304 13256 10308
rect 22952 10364 23016 10368
rect 22952 10308 22956 10364
rect 22956 10308 23012 10364
rect 23012 10308 23016 10364
rect 22952 10304 23016 10308
rect 23032 10364 23096 10368
rect 23032 10308 23036 10364
rect 23036 10308 23092 10364
rect 23092 10308 23096 10364
rect 23032 10304 23096 10308
rect 23112 10364 23176 10368
rect 23112 10308 23116 10364
rect 23116 10308 23172 10364
rect 23172 10308 23176 10364
rect 23112 10304 23176 10308
rect 23192 10364 23256 10368
rect 23192 10308 23196 10364
rect 23196 10308 23252 10364
rect 23252 10308 23256 10364
rect 23192 10304 23256 10308
rect 32952 10364 33016 10368
rect 32952 10308 32956 10364
rect 32956 10308 33012 10364
rect 33012 10308 33016 10364
rect 32952 10304 33016 10308
rect 33032 10364 33096 10368
rect 33032 10308 33036 10364
rect 33036 10308 33092 10364
rect 33092 10308 33096 10364
rect 33032 10304 33096 10308
rect 33112 10364 33176 10368
rect 33112 10308 33116 10364
rect 33116 10308 33172 10364
rect 33172 10308 33176 10364
rect 33112 10304 33176 10308
rect 33192 10364 33256 10368
rect 33192 10308 33196 10364
rect 33196 10308 33252 10364
rect 33252 10308 33256 10364
rect 33192 10304 33256 10308
rect 42952 10364 43016 10368
rect 42952 10308 42956 10364
rect 42956 10308 43012 10364
rect 43012 10308 43016 10364
rect 42952 10304 43016 10308
rect 43032 10364 43096 10368
rect 43032 10308 43036 10364
rect 43036 10308 43092 10364
rect 43092 10308 43096 10364
rect 43032 10304 43096 10308
rect 43112 10364 43176 10368
rect 43112 10308 43116 10364
rect 43116 10308 43172 10364
rect 43172 10308 43176 10364
rect 43112 10304 43176 10308
rect 43192 10364 43256 10368
rect 43192 10308 43196 10364
rect 43196 10308 43252 10364
rect 43252 10308 43256 10364
rect 43192 10304 43256 10308
rect 7952 9820 8016 9824
rect 7952 9764 7956 9820
rect 7956 9764 8012 9820
rect 8012 9764 8016 9820
rect 7952 9760 8016 9764
rect 8032 9820 8096 9824
rect 8032 9764 8036 9820
rect 8036 9764 8092 9820
rect 8092 9764 8096 9820
rect 8032 9760 8096 9764
rect 8112 9820 8176 9824
rect 8112 9764 8116 9820
rect 8116 9764 8172 9820
rect 8172 9764 8176 9820
rect 8112 9760 8176 9764
rect 8192 9820 8256 9824
rect 8192 9764 8196 9820
rect 8196 9764 8252 9820
rect 8252 9764 8256 9820
rect 8192 9760 8256 9764
rect 17952 9820 18016 9824
rect 17952 9764 17956 9820
rect 17956 9764 18012 9820
rect 18012 9764 18016 9820
rect 17952 9760 18016 9764
rect 18032 9820 18096 9824
rect 18032 9764 18036 9820
rect 18036 9764 18092 9820
rect 18092 9764 18096 9820
rect 18032 9760 18096 9764
rect 18112 9820 18176 9824
rect 18112 9764 18116 9820
rect 18116 9764 18172 9820
rect 18172 9764 18176 9820
rect 18112 9760 18176 9764
rect 18192 9820 18256 9824
rect 18192 9764 18196 9820
rect 18196 9764 18252 9820
rect 18252 9764 18256 9820
rect 18192 9760 18256 9764
rect 27952 9820 28016 9824
rect 27952 9764 27956 9820
rect 27956 9764 28012 9820
rect 28012 9764 28016 9820
rect 27952 9760 28016 9764
rect 28032 9820 28096 9824
rect 28032 9764 28036 9820
rect 28036 9764 28092 9820
rect 28092 9764 28096 9820
rect 28032 9760 28096 9764
rect 28112 9820 28176 9824
rect 28112 9764 28116 9820
rect 28116 9764 28172 9820
rect 28172 9764 28176 9820
rect 28112 9760 28176 9764
rect 28192 9820 28256 9824
rect 28192 9764 28196 9820
rect 28196 9764 28252 9820
rect 28252 9764 28256 9820
rect 28192 9760 28256 9764
rect 37952 9820 38016 9824
rect 37952 9764 37956 9820
rect 37956 9764 38012 9820
rect 38012 9764 38016 9820
rect 37952 9760 38016 9764
rect 38032 9820 38096 9824
rect 38032 9764 38036 9820
rect 38036 9764 38092 9820
rect 38092 9764 38096 9820
rect 38032 9760 38096 9764
rect 38112 9820 38176 9824
rect 38112 9764 38116 9820
rect 38116 9764 38172 9820
rect 38172 9764 38176 9820
rect 38112 9760 38176 9764
rect 38192 9820 38256 9824
rect 38192 9764 38196 9820
rect 38196 9764 38252 9820
rect 38252 9764 38256 9820
rect 38192 9760 38256 9764
rect 47952 9820 48016 9824
rect 47952 9764 47956 9820
rect 47956 9764 48012 9820
rect 48012 9764 48016 9820
rect 47952 9760 48016 9764
rect 48032 9820 48096 9824
rect 48032 9764 48036 9820
rect 48036 9764 48092 9820
rect 48092 9764 48096 9820
rect 48032 9760 48096 9764
rect 48112 9820 48176 9824
rect 48112 9764 48116 9820
rect 48116 9764 48172 9820
rect 48172 9764 48176 9820
rect 48112 9760 48176 9764
rect 48192 9820 48256 9824
rect 48192 9764 48196 9820
rect 48196 9764 48252 9820
rect 48252 9764 48256 9820
rect 48192 9760 48256 9764
rect 2952 9276 3016 9280
rect 2952 9220 2956 9276
rect 2956 9220 3012 9276
rect 3012 9220 3016 9276
rect 2952 9216 3016 9220
rect 3032 9276 3096 9280
rect 3032 9220 3036 9276
rect 3036 9220 3092 9276
rect 3092 9220 3096 9276
rect 3032 9216 3096 9220
rect 3112 9276 3176 9280
rect 3112 9220 3116 9276
rect 3116 9220 3172 9276
rect 3172 9220 3176 9276
rect 3112 9216 3176 9220
rect 3192 9276 3256 9280
rect 3192 9220 3196 9276
rect 3196 9220 3252 9276
rect 3252 9220 3256 9276
rect 3192 9216 3256 9220
rect 12952 9276 13016 9280
rect 12952 9220 12956 9276
rect 12956 9220 13012 9276
rect 13012 9220 13016 9276
rect 12952 9216 13016 9220
rect 13032 9276 13096 9280
rect 13032 9220 13036 9276
rect 13036 9220 13092 9276
rect 13092 9220 13096 9276
rect 13032 9216 13096 9220
rect 13112 9276 13176 9280
rect 13112 9220 13116 9276
rect 13116 9220 13172 9276
rect 13172 9220 13176 9276
rect 13112 9216 13176 9220
rect 13192 9276 13256 9280
rect 13192 9220 13196 9276
rect 13196 9220 13252 9276
rect 13252 9220 13256 9276
rect 13192 9216 13256 9220
rect 22952 9276 23016 9280
rect 22952 9220 22956 9276
rect 22956 9220 23012 9276
rect 23012 9220 23016 9276
rect 22952 9216 23016 9220
rect 23032 9276 23096 9280
rect 23032 9220 23036 9276
rect 23036 9220 23092 9276
rect 23092 9220 23096 9276
rect 23032 9216 23096 9220
rect 23112 9276 23176 9280
rect 23112 9220 23116 9276
rect 23116 9220 23172 9276
rect 23172 9220 23176 9276
rect 23112 9216 23176 9220
rect 23192 9276 23256 9280
rect 23192 9220 23196 9276
rect 23196 9220 23252 9276
rect 23252 9220 23256 9276
rect 23192 9216 23256 9220
rect 32952 9276 33016 9280
rect 32952 9220 32956 9276
rect 32956 9220 33012 9276
rect 33012 9220 33016 9276
rect 32952 9216 33016 9220
rect 33032 9276 33096 9280
rect 33032 9220 33036 9276
rect 33036 9220 33092 9276
rect 33092 9220 33096 9276
rect 33032 9216 33096 9220
rect 33112 9276 33176 9280
rect 33112 9220 33116 9276
rect 33116 9220 33172 9276
rect 33172 9220 33176 9276
rect 33112 9216 33176 9220
rect 33192 9276 33256 9280
rect 33192 9220 33196 9276
rect 33196 9220 33252 9276
rect 33252 9220 33256 9276
rect 33192 9216 33256 9220
rect 42952 9276 43016 9280
rect 42952 9220 42956 9276
rect 42956 9220 43012 9276
rect 43012 9220 43016 9276
rect 42952 9216 43016 9220
rect 43032 9276 43096 9280
rect 43032 9220 43036 9276
rect 43036 9220 43092 9276
rect 43092 9220 43096 9276
rect 43032 9216 43096 9220
rect 43112 9276 43176 9280
rect 43112 9220 43116 9276
rect 43116 9220 43172 9276
rect 43172 9220 43176 9276
rect 43112 9216 43176 9220
rect 43192 9276 43256 9280
rect 43192 9220 43196 9276
rect 43196 9220 43252 9276
rect 43252 9220 43256 9276
rect 43192 9216 43256 9220
rect 7952 8732 8016 8736
rect 7952 8676 7956 8732
rect 7956 8676 8012 8732
rect 8012 8676 8016 8732
rect 7952 8672 8016 8676
rect 8032 8732 8096 8736
rect 8032 8676 8036 8732
rect 8036 8676 8092 8732
rect 8092 8676 8096 8732
rect 8032 8672 8096 8676
rect 8112 8732 8176 8736
rect 8112 8676 8116 8732
rect 8116 8676 8172 8732
rect 8172 8676 8176 8732
rect 8112 8672 8176 8676
rect 8192 8732 8256 8736
rect 8192 8676 8196 8732
rect 8196 8676 8252 8732
rect 8252 8676 8256 8732
rect 8192 8672 8256 8676
rect 17952 8732 18016 8736
rect 17952 8676 17956 8732
rect 17956 8676 18012 8732
rect 18012 8676 18016 8732
rect 17952 8672 18016 8676
rect 18032 8732 18096 8736
rect 18032 8676 18036 8732
rect 18036 8676 18092 8732
rect 18092 8676 18096 8732
rect 18032 8672 18096 8676
rect 18112 8732 18176 8736
rect 18112 8676 18116 8732
rect 18116 8676 18172 8732
rect 18172 8676 18176 8732
rect 18112 8672 18176 8676
rect 18192 8732 18256 8736
rect 18192 8676 18196 8732
rect 18196 8676 18252 8732
rect 18252 8676 18256 8732
rect 18192 8672 18256 8676
rect 27952 8732 28016 8736
rect 27952 8676 27956 8732
rect 27956 8676 28012 8732
rect 28012 8676 28016 8732
rect 27952 8672 28016 8676
rect 28032 8732 28096 8736
rect 28032 8676 28036 8732
rect 28036 8676 28092 8732
rect 28092 8676 28096 8732
rect 28032 8672 28096 8676
rect 28112 8732 28176 8736
rect 28112 8676 28116 8732
rect 28116 8676 28172 8732
rect 28172 8676 28176 8732
rect 28112 8672 28176 8676
rect 28192 8732 28256 8736
rect 28192 8676 28196 8732
rect 28196 8676 28252 8732
rect 28252 8676 28256 8732
rect 28192 8672 28256 8676
rect 37952 8732 38016 8736
rect 37952 8676 37956 8732
rect 37956 8676 38012 8732
rect 38012 8676 38016 8732
rect 37952 8672 38016 8676
rect 38032 8732 38096 8736
rect 38032 8676 38036 8732
rect 38036 8676 38092 8732
rect 38092 8676 38096 8732
rect 38032 8672 38096 8676
rect 38112 8732 38176 8736
rect 38112 8676 38116 8732
rect 38116 8676 38172 8732
rect 38172 8676 38176 8732
rect 38112 8672 38176 8676
rect 38192 8732 38256 8736
rect 38192 8676 38196 8732
rect 38196 8676 38252 8732
rect 38252 8676 38256 8732
rect 38192 8672 38256 8676
rect 47952 8732 48016 8736
rect 47952 8676 47956 8732
rect 47956 8676 48012 8732
rect 48012 8676 48016 8732
rect 47952 8672 48016 8676
rect 48032 8732 48096 8736
rect 48032 8676 48036 8732
rect 48036 8676 48092 8732
rect 48092 8676 48096 8732
rect 48032 8672 48096 8676
rect 48112 8732 48176 8736
rect 48112 8676 48116 8732
rect 48116 8676 48172 8732
rect 48172 8676 48176 8732
rect 48112 8672 48176 8676
rect 48192 8732 48256 8736
rect 48192 8676 48196 8732
rect 48196 8676 48252 8732
rect 48252 8676 48256 8732
rect 48192 8672 48256 8676
rect 2952 8188 3016 8192
rect 2952 8132 2956 8188
rect 2956 8132 3012 8188
rect 3012 8132 3016 8188
rect 2952 8128 3016 8132
rect 3032 8188 3096 8192
rect 3032 8132 3036 8188
rect 3036 8132 3092 8188
rect 3092 8132 3096 8188
rect 3032 8128 3096 8132
rect 3112 8188 3176 8192
rect 3112 8132 3116 8188
rect 3116 8132 3172 8188
rect 3172 8132 3176 8188
rect 3112 8128 3176 8132
rect 3192 8188 3256 8192
rect 3192 8132 3196 8188
rect 3196 8132 3252 8188
rect 3252 8132 3256 8188
rect 3192 8128 3256 8132
rect 12952 8188 13016 8192
rect 12952 8132 12956 8188
rect 12956 8132 13012 8188
rect 13012 8132 13016 8188
rect 12952 8128 13016 8132
rect 13032 8188 13096 8192
rect 13032 8132 13036 8188
rect 13036 8132 13092 8188
rect 13092 8132 13096 8188
rect 13032 8128 13096 8132
rect 13112 8188 13176 8192
rect 13112 8132 13116 8188
rect 13116 8132 13172 8188
rect 13172 8132 13176 8188
rect 13112 8128 13176 8132
rect 13192 8188 13256 8192
rect 13192 8132 13196 8188
rect 13196 8132 13252 8188
rect 13252 8132 13256 8188
rect 13192 8128 13256 8132
rect 22952 8188 23016 8192
rect 22952 8132 22956 8188
rect 22956 8132 23012 8188
rect 23012 8132 23016 8188
rect 22952 8128 23016 8132
rect 23032 8188 23096 8192
rect 23032 8132 23036 8188
rect 23036 8132 23092 8188
rect 23092 8132 23096 8188
rect 23032 8128 23096 8132
rect 23112 8188 23176 8192
rect 23112 8132 23116 8188
rect 23116 8132 23172 8188
rect 23172 8132 23176 8188
rect 23112 8128 23176 8132
rect 23192 8188 23256 8192
rect 23192 8132 23196 8188
rect 23196 8132 23252 8188
rect 23252 8132 23256 8188
rect 23192 8128 23256 8132
rect 32952 8188 33016 8192
rect 32952 8132 32956 8188
rect 32956 8132 33012 8188
rect 33012 8132 33016 8188
rect 32952 8128 33016 8132
rect 33032 8188 33096 8192
rect 33032 8132 33036 8188
rect 33036 8132 33092 8188
rect 33092 8132 33096 8188
rect 33032 8128 33096 8132
rect 33112 8188 33176 8192
rect 33112 8132 33116 8188
rect 33116 8132 33172 8188
rect 33172 8132 33176 8188
rect 33112 8128 33176 8132
rect 33192 8188 33256 8192
rect 33192 8132 33196 8188
rect 33196 8132 33252 8188
rect 33252 8132 33256 8188
rect 33192 8128 33256 8132
rect 42952 8188 43016 8192
rect 42952 8132 42956 8188
rect 42956 8132 43012 8188
rect 43012 8132 43016 8188
rect 42952 8128 43016 8132
rect 43032 8188 43096 8192
rect 43032 8132 43036 8188
rect 43036 8132 43092 8188
rect 43092 8132 43096 8188
rect 43032 8128 43096 8132
rect 43112 8188 43176 8192
rect 43112 8132 43116 8188
rect 43116 8132 43172 8188
rect 43172 8132 43176 8188
rect 43112 8128 43176 8132
rect 43192 8188 43256 8192
rect 43192 8132 43196 8188
rect 43196 8132 43252 8188
rect 43252 8132 43256 8188
rect 43192 8128 43256 8132
rect 7952 7644 8016 7648
rect 7952 7588 7956 7644
rect 7956 7588 8012 7644
rect 8012 7588 8016 7644
rect 7952 7584 8016 7588
rect 8032 7644 8096 7648
rect 8032 7588 8036 7644
rect 8036 7588 8092 7644
rect 8092 7588 8096 7644
rect 8032 7584 8096 7588
rect 8112 7644 8176 7648
rect 8112 7588 8116 7644
rect 8116 7588 8172 7644
rect 8172 7588 8176 7644
rect 8112 7584 8176 7588
rect 8192 7644 8256 7648
rect 8192 7588 8196 7644
rect 8196 7588 8252 7644
rect 8252 7588 8256 7644
rect 8192 7584 8256 7588
rect 17952 7644 18016 7648
rect 17952 7588 17956 7644
rect 17956 7588 18012 7644
rect 18012 7588 18016 7644
rect 17952 7584 18016 7588
rect 18032 7644 18096 7648
rect 18032 7588 18036 7644
rect 18036 7588 18092 7644
rect 18092 7588 18096 7644
rect 18032 7584 18096 7588
rect 18112 7644 18176 7648
rect 18112 7588 18116 7644
rect 18116 7588 18172 7644
rect 18172 7588 18176 7644
rect 18112 7584 18176 7588
rect 18192 7644 18256 7648
rect 18192 7588 18196 7644
rect 18196 7588 18252 7644
rect 18252 7588 18256 7644
rect 18192 7584 18256 7588
rect 27952 7644 28016 7648
rect 27952 7588 27956 7644
rect 27956 7588 28012 7644
rect 28012 7588 28016 7644
rect 27952 7584 28016 7588
rect 28032 7644 28096 7648
rect 28032 7588 28036 7644
rect 28036 7588 28092 7644
rect 28092 7588 28096 7644
rect 28032 7584 28096 7588
rect 28112 7644 28176 7648
rect 28112 7588 28116 7644
rect 28116 7588 28172 7644
rect 28172 7588 28176 7644
rect 28112 7584 28176 7588
rect 28192 7644 28256 7648
rect 28192 7588 28196 7644
rect 28196 7588 28252 7644
rect 28252 7588 28256 7644
rect 28192 7584 28256 7588
rect 37952 7644 38016 7648
rect 37952 7588 37956 7644
rect 37956 7588 38012 7644
rect 38012 7588 38016 7644
rect 37952 7584 38016 7588
rect 38032 7644 38096 7648
rect 38032 7588 38036 7644
rect 38036 7588 38092 7644
rect 38092 7588 38096 7644
rect 38032 7584 38096 7588
rect 38112 7644 38176 7648
rect 38112 7588 38116 7644
rect 38116 7588 38172 7644
rect 38172 7588 38176 7644
rect 38112 7584 38176 7588
rect 38192 7644 38256 7648
rect 38192 7588 38196 7644
rect 38196 7588 38252 7644
rect 38252 7588 38256 7644
rect 38192 7584 38256 7588
rect 47952 7644 48016 7648
rect 47952 7588 47956 7644
rect 47956 7588 48012 7644
rect 48012 7588 48016 7644
rect 47952 7584 48016 7588
rect 48032 7644 48096 7648
rect 48032 7588 48036 7644
rect 48036 7588 48092 7644
rect 48092 7588 48096 7644
rect 48032 7584 48096 7588
rect 48112 7644 48176 7648
rect 48112 7588 48116 7644
rect 48116 7588 48172 7644
rect 48172 7588 48176 7644
rect 48112 7584 48176 7588
rect 48192 7644 48256 7648
rect 48192 7588 48196 7644
rect 48196 7588 48252 7644
rect 48252 7588 48256 7644
rect 48192 7584 48256 7588
rect 2952 7100 3016 7104
rect 2952 7044 2956 7100
rect 2956 7044 3012 7100
rect 3012 7044 3016 7100
rect 2952 7040 3016 7044
rect 3032 7100 3096 7104
rect 3032 7044 3036 7100
rect 3036 7044 3092 7100
rect 3092 7044 3096 7100
rect 3032 7040 3096 7044
rect 3112 7100 3176 7104
rect 3112 7044 3116 7100
rect 3116 7044 3172 7100
rect 3172 7044 3176 7100
rect 3112 7040 3176 7044
rect 3192 7100 3256 7104
rect 3192 7044 3196 7100
rect 3196 7044 3252 7100
rect 3252 7044 3256 7100
rect 3192 7040 3256 7044
rect 12952 7100 13016 7104
rect 12952 7044 12956 7100
rect 12956 7044 13012 7100
rect 13012 7044 13016 7100
rect 12952 7040 13016 7044
rect 13032 7100 13096 7104
rect 13032 7044 13036 7100
rect 13036 7044 13092 7100
rect 13092 7044 13096 7100
rect 13032 7040 13096 7044
rect 13112 7100 13176 7104
rect 13112 7044 13116 7100
rect 13116 7044 13172 7100
rect 13172 7044 13176 7100
rect 13112 7040 13176 7044
rect 13192 7100 13256 7104
rect 13192 7044 13196 7100
rect 13196 7044 13252 7100
rect 13252 7044 13256 7100
rect 13192 7040 13256 7044
rect 22952 7100 23016 7104
rect 22952 7044 22956 7100
rect 22956 7044 23012 7100
rect 23012 7044 23016 7100
rect 22952 7040 23016 7044
rect 23032 7100 23096 7104
rect 23032 7044 23036 7100
rect 23036 7044 23092 7100
rect 23092 7044 23096 7100
rect 23032 7040 23096 7044
rect 23112 7100 23176 7104
rect 23112 7044 23116 7100
rect 23116 7044 23172 7100
rect 23172 7044 23176 7100
rect 23112 7040 23176 7044
rect 23192 7100 23256 7104
rect 23192 7044 23196 7100
rect 23196 7044 23252 7100
rect 23252 7044 23256 7100
rect 23192 7040 23256 7044
rect 32952 7100 33016 7104
rect 32952 7044 32956 7100
rect 32956 7044 33012 7100
rect 33012 7044 33016 7100
rect 32952 7040 33016 7044
rect 33032 7100 33096 7104
rect 33032 7044 33036 7100
rect 33036 7044 33092 7100
rect 33092 7044 33096 7100
rect 33032 7040 33096 7044
rect 33112 7100 33176 7104
rect 33112 7044 33116 7100
rect 33116 7044 33172 7100
rect 33172 7044 33176 7100
rect 33112 7040 33176 7044
rect 33192 7100 33256 7104
rect 33192 7044 33196 7100
rect 33196 7044 33252 7100
rect 33252 7044 33256 7100
rect 33192 7040 33256 7044
rect 42952 7100 43016 7104
rect 42952 7044 42956 7100
rect 42956 7044 43012 7100
rect 43012 7044 43016 7100
rect 42952 7040 43016 7044
rect 43032 7100 43096 7104
rect 43032 7044 43036 7100
rect 43036 7044 43092 7100
rect 43092 7044 43096 7100
rect 43032 7040 43096 7044
rect 43112 7100 43176 7104
rect 43112 7044 43116 7100
rect 43116 7044 43172 7100
rect 43172 7044 43176 7100
rect 43112 7040 43176 7044
rect 43192 7100 43256 7104
rect 43192 7044 43196 7100
rect 43196 7044 43252 7100
rect 43252 7044 43256 7100
rect 43192 7040 43256 7044
rect 7952 6556 8016 6560
rect 7952 6500 7956 6556
rect 7956 6500 8012 6556
rect 8012 6500 8016 6556
rect 7952 6496 8016 6500
rect 8032 6556 8096 6560
rect 8032 6500 8036 6556
rect 8036 6500 8092 6556
rect 8092 6500 8096 6556
rect 8032 6496 8096 6500
rect 8112 6556 8176 6560
rect 8112 6500 8116 6556
rect 8116 6500 8172 6556
rect 8172 6500 8176 6556
rect 8112 6496 8176 6500
rect 8192 6556 8256 6560
rect 8192 6500 8196 6556
rect 8196 6500 8252 6556
rect 8252 6500 8256 6556
rect 8192 6496 8256 6500
rect 17952 6556 18016 6560
rect 17952 6500 17956 6556
rect 17956 6500 18012 6556
rect 18012 6500 18016 6556
rect 17952 6496 18016 6500
rect 18032 6556 18096 6560
rect 18032 6500 18036 6556
rect 18036 6500 18092 6556
rect 18092 6500 18096 6556
rect 18032 6496 18096 6500
rect 18112 6556 18176 6560
rect 18112 6500 18116 6556
rect 18116 6500 18172 6556
rect 18172 6500 18176 6556
rect 18112 6496 18176 6500
rect 18192 6556 18256 6560
rect 18192 6500 18196 6556
rect 18196 6500 18252 6556
rect 18252 6500 18256 6556
rect 18192 6496 18256 6500
rect 27952 6556 28016 6560
rect 27952 6500 27956 6556
rect 27956 6500 28012 6556
rect 28012 6500 28016 6556
rect 27952 6496 28016 6500
rect 28032 6556 28096 6560
rect 28032 6500 28036 6556
rect 28036 6500 28092 6556
rect 28092 6500 28096 6556
rect 28032 6496 28096 6500
rect 28112 6556 28176 6560
rect 28112 6500 28116 6556
rect 28116 6500 28172 6556
rect 28172 6500 28176 6556
rect 28112 6496 28176 6500
rect 28192 6556 28256 6560
rect 28192 6500 28196 6556
rect 28196 6500 28252 6556
rect 28252 6500 28256 6556
rect 28192 6496 28256 6500
rect 37952 6556 38016 6560
rect 37952 6500 37956 6556
rect 37956 6500 38012 6556
rect 38012 6500 38016 6556
rect 37952 6496 38016 6500
rect 38032 6556 38096 6560
rect 38032 6500 38036 6556
rect 38036 6500 38092 6556
rect 38092 6500 38096 6556
rect 38032 6496 38096 6500
rect 38112 6556 38176 6560
rect 38112 6500 38116 6556
rect 38116 6500 38172 6556
rect 38172 6500 38176 6556
rect 38112 6496 38176 6500
rect 38192 6556 38256 6560
rect 38192 6500 38196 6556
rect 38196 6500 38252 6556
rect 38252 6500 38256 6556
rect 38192 6496 38256 6500
rect 47952 6556 48016 6560
rect 47952 6500 47956 6556
rect 47956 6500 48012 6556
rect 48012 6500 48016 6556
rect 47952 6496 48016 6500
rect 48032 6556 48096 6560
rect 48032 6500 48036 6556
rect 48036 6500 48092 6556
rect 48092 6500 48096 6556
rect 48032 6496 48096 6500
rect 48112 6556 48176 6560
rect 48112 6500 48116 6556
rect 48116 6500 48172 6556
rect 48172 6500 48176 6556
rect 48112 6496 48176 6500
rect 48192 6556 48256 6560
rect 48192 6500 48196 6556
rect 48196 6500 48252 6556
rect 48252 6500 48256 6556
rect 48192 6496 48256 6500
rect 2952 6012 3016 6016
rect 2952 5956 2956 6012
rect 2956 5956 3012 6012
rect 3012 5956 3016 6012
rect 2952 5952 3016 5956
rect 3032 6012 3096 6016
rect 3032 5956 3036 6012
rect 3036 5956 3092 6012
rect 3092 5956 3096 6012
rect 3032 5952 3096 5956
rect 3112 6012 3176 6016
rect 3112 5956 3116 6012
rect 3116 5956 3172 6012
rect 3172 5956 3176 6012
rect 3112 5952 3176 5956
rect 3192 6012 3256 6016
rect 3192 5956 3196 6012
rect 3196 5956 3252 6012
rect 3252 5956 3256 6012
rect 3192 5952 3256 5956
rect 12952 6012 13016 6016
rect 12952 5956 12956 6012
rect 12956 5956 13012 6012
rect 13012 5956 13016 6012
rect 12952 5952 13016 5956
rect 13032 6012 13096 6016
rect 13032 5956 13036 6012
rect 13036 5956 13092 6012
rect 13092 5956 13096 6012
rect 13032 5952 13096 5956
rect 13112 6012 13176 6016
rect 13112 5956 13116 6012
rect 13116 5956 13172 6012
rect 13172 5956 13176 6012
rect 13112 5952 13176 5956
rect 13192 6012 13256 6016
rect 13192 5956 13196 6012
rect 13196 5956 13252 6012
rect 13252 5956 13256 6012
rect 13192 5952 13256 5956
rect 22952 6012 23016 6016
rect 22952 5956 22956 6012
rect 22956 5956 23012 6012
rect 23012 5956 23016 6012
rect 22952 5952 23016 5956
rect 23032 6012 23096 6016
rect 23032 5956 23036 6012
rect 23036 5956 23092 6012
rect 23092 5956 23096 6012
rect 23032 5952 23096 5956
rect 23112 6012 23176 6016
rect 23112 5956 23116 6012
rect 23116 5956 23172 6012
rect 23172 5956 23176 6012
rect 23112 5952 23176 5956
rect 23192 6012 23256 6016
rect 23192 5956 23196 6012
rect 23196 5956 23252 6012
rect 23252 5956 23256 6012
rect 23192 5952 23256 5956
rect 32952 6012 33016 6016
rect 32952 5956 32956 6012
rect 32956 5956 33012 6012
rect 33012 5956 33016 6012
rect 32952 5952 33016 5956
rect 33032 6012 33096 6016
rect 33032 5956 33036 6012
rect 33036 5956 33092 6012
rect 33092 5956 33096 6012
rect 33032 5952 33096 5956
rect 33112 6012 33176 6016
rect 33112 5956 33116 6012
rect 33116 5956 33172 6012
rect 33172 5956 33176 6012
rect 33112 5952 33176 5956
rect 33192 6012 33256 6016
rect 33192 5956 33196 6012
rect 33196 5956 33252 6012
rect 33252 5956 33256 6012
rect 33192 5952 33256 5956
rect 42952 6012 43016 6016
rect 42952 5956 42956 6012
rect 42956 5956 43012 6012
rect 43012 5956 43016 6012
rect 42952 5952 43016 5956
rect 43032 6012 43096 6016
rect 43032 5956 43036 6012
rect 43036 5956 43092 6012
rect 43092 5956 43096 6012
rect 43032 5952 43096 5956
rect 43112 6012 43176 6016
rect 43112 5956 43116 6012
rect 43116 5956 43172 6012
rect 43172 5956 43176 6012
rect 43112 5952 43176 5956
rect 43192 6012 43256 6016
rect 43192 5956 43196 6012
rect 43196 5956 43252 6012
rect 43252 5956 43256 6012
rect 43192 5952 43256 5956
rect 7952 5468 8016 5472
rect 7952 5412 7956 5468
rect 7956 5412 8012 5468
rect 8012 5412 8016 5468
rect 7952 5408 8016 5412
rect 8032 5468 8096 5472
rect 8032 5412 8036 5468
rect 8036 5412 8092 5468
rect 8092 5412 8096 5468
rect 8032 5408 8096 5412
rect 8112 5468 8176 5472
rect 8112 5412 8116 5468
rect 8116 5412 8172 5468
rect 8172 5412 8176 5468
rect 8112 5408 8176 5412
rect 8192 5468 8256 5472
rect 8192 5412 8196 5468
rect 8196 5412 8252 5468
rect 8252 5412 8256 5468
rect 8192 5408 8256 5412
rect 17952 5468 18016 5472
rect 17952 5412 17956 5468
rect 17956 5412 18012 5468
rect 18012 5412 18016 5468
rect 17952 5408 18016 5412
rect 18032 5468 18096 5472
rect 18032 5412 18036 5468
rect 18036 5412 18092 5468
rect 18092 5412 18096 5468
rect 18032 5408 18096 5412
rect 18112 5468 18176 5472
rect 18112 5412 18116 5468
rect 18116 5412 18172 5468
rect 18172 5412 18176 5468
rect 18112 5408 18176 5412
rect 18192 5468 18256 5472
rect 18192 5412 18196 5468
rect 18196 5412 18252 5468
rect 18252 5412 18256 5468
rect 18192 5408 18256 5412
rect 27952 5468 28016 5472
rect 27952 5412 27956 5468
rect 27956 5412 28012 5468
rect 28012 5412 28016 5468
rect 27952 5408 28016 5412
rect 28032 5468 28096 5472
rect 28032 5412 28036 5468
rect 28036 5412 28092 5468
rect 28092 5412 28096 5468
rect 28032 5408 28096 5412
rect 28112 5468 28176 5472
rect 28112 5412 28116 5468
rect 28116 5412 28172 5468
rect 28172 5412 28176 5468
rect 28112 5408 28176 5412
rect 28192 5468 28256 5472
rect 28192 5412 28196 5468
rect 28196 5412 28252 5468
rect 28252 5412 28256 5468
rect 28192 5408 28256 5412
rect 37952 5468 38016 5472
rect 37952 5412 37956 5468
rect 37956 5412 38012 5468
rect 38012 5412 38016 5468
rect 37952 5408 38016 5412
rect 38032 5468 38096 5472
rect 38032 5412 38036 5468
rect 38036 5412 38092 5468
rect 38092 5412 38096 5468
rect 38032 5408 38096 5412
rect 38112 5468 38176 5472
rect 38112 5412 38116 5468
rect 38116 5412 38172 5468
rect 38172 5412 38176 5468
rect 38112 5408 38176 5412
rect 38192 5468 38256 5472
rect 38192 5412 38196 5468
rect 38196 5412 38252 5468
rect 38252 5412 38256 5468
rect 38192 5408 38256 5412
rect 47952 5468 48016 5472
rect 47952 5412 47956 5468
rect 47956 5412 48012 5468
rect 48012 5412 48016 5468
rect 47952 5408 48016 5412
rect 48032 5468 48096 5472
rect 48032 5412 48036 5468
rect 48036 5412 48092 5468
rect 48092 5412 48096 5468
rect 48032 5408 48096 5412
rect 48112 5468 48176 5472
rect 48112 5412 48116 5468
rect 48116 5412 48172 5468
rect 48172 5412 48176 5468
rect 48112 5408 48176 5412
rect 48192 5468 48256 5472
rect 48192 5412 48196 5468
rect 48196 5412 48252 5468
rect 48252 5412 48256 5468
rect 48192 5408 48256 5412
rect 2952 4924 3016 4928
rect 2952 4868 2956 4924
rect 2956 4868 3012 4924
rect 3012 4868 3016 4924
rect 2952 4864 3016 4868
rect 3032 4924 3096 4928
rect 3032 4868 3036 4924
rect 3036 4868 3092 4924
rect 3092 4868 3096 4924
rect 3032 4864 3096 4868
rect 3112 4924 3176 4928
rect 3112 4868 3116 4924
rect 3116 4868 3172 4924
rect 3172 4868 3176 4924
rect 3112 4864 3176 4868
rect 3192 4924 3256 4928
rect 3192 4868 3196 4924
rect 3196 4868 3252 4924
rect 3252 4868 3256 4924
rect 3192 4864 3256 4868
rect 12952 4924 13016 4928
rect 12952 4868 12956 4924
rect 12956 4868 13012 4924
rect 13012 4868 13016 4924
rect 12952 4864 13016 4868
rect 13032 4924 13096 4928
rect 13032 4868 13036 4924
rect 13036 4868 13092 4924
rect 13092 4868 13096 4924
rect 13032 4864 13096 4868
rect 13112 4924 13176 4928
rect 13112 4868 13116 4924
rect 13116 4868 13172 4924
rect 13172 4868 13176 4924
rect 13112 4864 13176 4868
rect 13192 4924 13256 4928
rect 13192 4868 13196 4924
rect 13196 4868 13252 4924
rect 13252 4868 13256 4924
rect 13192 4864 13256 4868
rect 22952 4924 23016 4928
rect 22952 4868 22956 4924
rect 22956 4868 23012 4924
rect 23012 4868 23016 4924
rect 22952 4864 23016 4868
rect 23032 4924 23096 4928
rect 23032 4868 23036 4924
rect 23036 4868 23092 4924
rect 23092 4868 23096 4924
rect 23032 4864 23096 4868
rect 23112 4924 23176 4928
rect 23112 4868 23116 4924
rect 23116 4868 23172 4924
rect 23172 4868 23176 4924
rect 23112 4864 23176 4868
rect 23192 4924 23256 4928
rect 23192 4868 23196 4924
rect 23196 4868 23252 4924
rect 23252 4868 23256 4924
rect 23192 4864 23256 4868
rect 32952 4924 33016 4928
rect 32952 4868 32956 4924
rect 32956 4868 33012 4924
rect 33012 4868 33016 4924
rect 32952 4864 33016 4868
rect 33032 4924 33096 4928
rect 33032 4868 33036 4924
rect 33036 4868 33092 4924
rect 33092 4868 33096 4924
rect 33032 4864 33096 4868
rect 33112 4924 33176 4928
rect 33112 4868 33116 4924
rect 33116 4868 33172 4924
rect 33172 4868 33176 4924
rect 33112 4864 33176 4868
rect 33192 4924 33256 4928
rect 33192 4868 33196 4924
rect 33196 4868 33252 4924
rect 33252 4868 33256 4924
rect 33192 4864 33256 4868
rect 42952 4924 43016 4928
rect 42952 4868 42956 4924
rect 42956 4868 43012 4924
rect 43012 4868 43016 4924
rect 42952 4864 43016 4868
rect 43032 4924 43096 4928
rect 43032 4868 43036 4924
rect 43036 4868 43092 4924
rect 43092 4868 43096 4924
rect 43032 4864 43096 4868
rect 43112 4924 43176 4928
rect 43112 4868 43116 4924
rect 43116 4868 43172 4924
rect 43172 4868 43176 4924
rect 43112 4864 43176 4868
rect 43192 4924 43256 4928
rect 43192 4868 43196 4924
rect 43196 4868 43252 4924
rect 43252 4868 43256 4924
rect 43192 4864 43256 4868
rect 7952 4380 8016 4384
rect 7952 4324 7956 4380
rect 7956 4324 8012 4380
rect 8012 4324 8016 4380
rect 7952 4320 8016 4324
rect 8032 4380 8096 4384
rect 8032 4324 8036 4380
rect 8036 4324 8092 4380
rect 8092 4324 8096 4380
rect 8032 4320 8096 4324
rect 8112 4380 8176 4384
rect 8112 4324 8116 4380
rect 8116 4324 8172 4380
rect 8172 4324 8176 4380
rect 8112 4320 8176 4324
rect 8192 4380 8256 4384
rect 8192 4324 8196 4380
rect 8196 4324 8252 4380
rect 8252 4324 8256 4380
rect 8192 4320 8256 4324
rect 17952 4380 18016 4384
rect 17952 4324 17956 4380
rect 17956 4324 18012 4380
rect 18012 4324 18016 4380
rect 17952 4320 18016 4324
rect 18032 4380 18096 4384
rect 18032 4324 18036 4380
rect 18036 4324 18092 4380
rect 18092 4324 18096 4380
rect 18032 4320 18096 4324
rect 18112 4380 18176 4384
rect 18112 4324 18116 4380
rect 18116 4324 18172 4380
rect 18172 4324 18176 4380
rect 18112 4320 18176 4324
rect 18192 4380 18256 4384
rect 18192 4324 18196 4380
rect 18196 4324 18252 4380
rect 18252 4324 18256 4380
rect 18192 4320 18256 4324
rect 27952 4380 28016 4384
rect 27952 4324 27956 4380
rect 27956 4324 28012 4380
rect 28012 4324 28016 4380
rect 27952 4320 28016 4324
rect 28032 4380 28096 4384
rect 28032 4324 28036 4380
rect 28036 4324 28092 4380
rect 28092 4324 28096 4380
rect 28032 4320 28096 4324
rect 28112 4380 28176 4384
rect 28112 4324 28116 4380
rect 28116 4324 28172 4380
rect 28172 4324 28176 4380
rect 28112 4320 28176 4324
rect 28192 4380 28256 4384
rect 28192 4324 28196 4380
rect 28196 4324 28252 4380
rect 28252 4324 28256 4380
rect 28192 4320 28256 4324
rect 37952 4380 38016 4384
rect 37952 4324 37956 4380
rect 37956 4324 38012 4380
rect 38012 4324 38016 4380
rect 37952 4320 38016 4324
rect 38032 4380 38096 4384
rect 38032 4324 38036 4380
rect 38036 4324 38092 4380
rect 38092 4324 38096 4380
rect 38032 4320 38096 4324
rect 38112 4380 38176 4384
rect 38112 4324 38116 4380
rect 38116 4324 38172 4380
rect 38172 4324 38176 4380
rect 38112 4320 38176 4324
rect 38192 4380 38256 4384
rect 38192 4324 38196 4380
rect 38196 4324 38252 4380
rect 38252 4324 38256 4380
rect 38192 4320 38256 4324
rect 47952 4380 48016 4384
rect 47952 4324 47956 4380
rect 47956 4324 48012 4380
rect 48012 4324 48016 4380
rect 47952 4320 48016 4324
rect 48032 4380 48096 4384
rect 48032 4324 48036 4380
rect 48036 4324 48092 4380
rect 48092 4324 48096 4380
rect 48032 4320 48096 4324
rect 48112 4380 48176 4384
rect 48112 4324 48116 4380
rect 48116 4324 48172 4380
rect 48172 4324 48176 4380
rect 48112 4320 48176 4324
rect 48192 4380 48256 4384
rect 48192 4324 48196 4380
rect 48196 4324 48252 4380
rect 48252 4324 48256 4380
rect 48192 4320 48256 4324
rect 2952 3836 3016 3840
rect 2952 3780 2956 3836
rect 2956 3780 3012 3836
rect 3012 3780 3016 3836
rect 2952 3776 3016 3780
rect 3032 3836 3096 3840
rect 3032 3780 3036 3836
rect 3036 3780 3092 3836
rect 3092 3780 3096 3836
rect 3032 3776 3096 3780
rect 3112 3836 3176 3840
rect 3112 3780 3116 3836
rect 3116 3780 3172 3836
rect 3172 3780 3176 3836
rect 3112 3776 3176 3780
rect 3192 3836 3256 3840
rect 3192 3780 3196 3836
rect 3196 3780 3252 3836
rect 3252 3780 3256 3836
rect 3192 3776 3256 3780
rect 12952 3836 13016 3840
rect 12952 3780 12956 3836
rect 12956 3780 13012 3836
rect 13012 3780 13016 3836
rect 12952 3776 13016 3780
rect 13032 3836 13096 3840
rect 13032 3780 13036 3836
rect 13036 3780 13092 3836
rect 13092 3780 13096 3836
rect 13032 3776 13096 3780
rect 13112 3836 13176 3840
rect 13112 3780 13116 3836
rect 13116 3780 13172 3836
rect 13172 3780 13176 3836
rect 13112 3776 13176 3780
rect 13192 3836 13256 3840
rect 13192 3780 13196 3836
rect 13196 3780 13252 3836
rect 13252 3780 13256 3836
rect 13192 3776 13256 3780
rect 22952 3836 23016 3840
rect 22952 3780 22956 3836
rect 22956 3780 23012 3836
rect 23012 3780 23016 3836
rect 22952 3776 23016 3780
rect 23032 3836 23096 3840
rect 23032 3780 23036 3836
rect 23036 3780 23092 3836
rect 23092 3780 23096 3836
rect 23032 3776 23096 3780
rect 23112 3836 23176 3840
rect 23112 3780 23116 3836
rect 23116 3780 23172 3836
rect 23172 3780 23176 3836
rect 23112 3776 23176 3780
rect 23192 3836 23256 3840
rect 23192 3780 23196 3836
rect 23196 3780 23252 3836
rect 23252 3780 23256 3836
rect 23192 3776 23256 3780
rect 32952 3836 33016 3840
rect 32952 3780 32956 3836
rect 32956 3780 33012 3836
rect 33012 3780 33016 3836
rect 32952 3776 33016 3780
rect 33032 3836 33096 3840
rect 33032 3780 33036 3836
rect 33036 3780 33092 3836
rect 33092 3780 33096 3836
rect 33032 3776 33096 3780
rect 33112 3836 33176 3840
rect 33112 3780 33116 3836
rect 33116 3780 33172 3836
rect 33172 3780 33176 3836
rect 33112 3776 33176 3780
rect 33192 3836 33256 3840
rect 33192 3780 33196 3836
rect 33196 3780 33252 3836
rect 33252 3780 33256 3836
rect 33192 3776 33256 3780
rect 42952 3836 43016 3840
rect 42952 3780 42956 3836
rect 42956 3780 43012 3836
rect 43012 3780 43016 3836
rect 42952 3776 43016 3780
rect 43032 3836 43096 3840
rect 43032 3780 43036 3836
rect 43036 3780 43092 3836
rect 43092 3780 43096 3836
rect 43032 3776 43096 3780
rect 43112 3836 43176 3840
rect 43112 3780 43116 3836
rect 43116 3780 43172 3836
rect 43172 3780 43176 3836
rect 43112 3776 43176 3780
rect 43192 3836 43256 3840
rect 43192 3780 43196 3836
rect 43196 3780 43252 3836
rect 43252 3780 43256 3836
rect 43192 3776 43256 3780
rect 27108 3436 27172 3500
rect 7952 3292 8016 3296
rect 7952 3236 7956 3292
rect 7956 3236 8012 3292
rect 8012 3236 8016 3292
rect 7952 3232 8016 3236
rect 8032 3292 8096 3296
rect 8032 3236 8036 3292
rect 8036 3236 8092 3292
rect 8092 3236 8096 3292
rect 8032 3232 8096 3236
rect 8112 3292 8176 3296
rect 8112 3236 8116 3292
rect 8116 3236 8172 3292
rect 8172 3236 8176 3292
rect 8112 3232 8176 3236
rect 8192 3292 8256 3296
rect 8192 3236 8196 3292
rect 8196 3236 8252 3292
rect 8252 3236 8256 3292
rect 8192 3232 8256 3236
rect 17952 3292 18016 3296
rect 17952 3236 17956 3292
rect 17956 3236 18012 3292
rect 18012 3236 18016 3292
rect 17952 3232 18016 3236
rect 18032 3292 18096 3296
rect 18032 3236 18036 3292
rect 18036 3236 18092 3292
rect 18092 3236 18096 3292
rect 18032 3232 18096 3236
rect 18112 3292 18176 3296
rect 18112 3236 18116 3292
rect 18116 3236 18172 3292
rect 18172 3236 18176 3292
rect 18112 3232 18176 3236
rect 18192 3292 18256 3296
rect 18192 3236 18196 3292
rect 18196 3236 18252 3292
rect 18252 3236 18256 3292
rect 18192 3232 18256 3236
rect 27952 3292 28016 3296
rect 27952 3236 27956 3292
rect 27956 3236 28012 3292
rect 28012 3236 28016 3292
rect 27952 3232 28016 3236
rect 28032 3292 28096 3296
rect 28032 3236 28036 3292
rect 28036 3236 28092 3292
rect 28092 3236 28096 3292
rect 28032 3232 28096 3236
rect 28112 3292 28176 3296
rect 28112 3236 28116 3292
rect 28116 3236 28172 3292
rect 28172 3236 28176 3292
rect 28112 3232 28176 3236
rect 28192 3292 28256 3296
rect 28192 3236 28196 3292
rect 28196 3236 28252 3292
rect 28252 3236 28256 3292
rect 28192 3232 28256 3236
rect 37952 3292 38016 3296
rect 37952 3236 37956 3292
rect 37956 3236 38012 3292
rect 38012 3236 38016 3292
rect 37952 3232 38016 3236
rect 38032 3292 38096 3296
rect 38032 3236 38036 3292
rect 38036 3236 38092 3292
rect 38092 3236 38096 3292
rect 38032 3232 38096 3236
rect 38112 3292 38176 3296
rect 38112 3236 38116 3292
rect 38116 3236 38172 3292
rect 38172 3236 38176 3292
rect 38112 3232 38176 3236
rect 38192 3292 38256 3296
rect 38192 3236 38196 3292
rect 38196 3236 38252 3292
rect 38252 3236 38256 3292
rect 38192 3232 38256 3236
rect 47952 3292 48016 3296
rect 47952 3236 47956 3292
rect 47956 3236 48012 3292
rect 48012 3236 48016 3292
rect 47952 3232 48016 3236
rect 48032 3292 48096 3296
rect 48032 3236 48036 3292
rect 48036 3236 48092 3292
rect 48092 3236 48096 3292
rect 48032 3232 48096 3236
rect 48112 3292 48176 3296
rect 48112 3236 48116 3292
rect 48116 3236 48172 3292
rect 48172 3236 48176 3292
rect 48112 3232 48176 3236
rect 48192 3292 48256 3296
rect 48192 3236 48196 3292
rect 48196 3236 48252 3292
rect 48252 3236 48256 3292
rect 48192 3232 48256 3236
rect 22508 2892 22572 2956
rect 2952 2748 3016 2752
rect 2952 2692 2956 2748
rect 2956 2692 3012 2748
rect 3012 2692 3016 2748
rect 2952 2688 3016 2692
rect 3032 2748 3096 2752
rect 3032 2692 3036 2748
rect 3036 2692 3092 2748
rect 3092 2692 3096 2748
rect 3032 2688 3096 2692
rect 3112 2748 3176 2752
rect 3112 2692 3116 2748
rect 3116 2692 3172 2748
rect 3172 2692 3176 2748
rect 3112 2688 3176 2692
rect 3192 2748 3256 2752
rect 3192 2692 3196 2748
rect 3196 2692 3252 2748
rect 3252 2692 3256 2748
rect 3192 2688 3256 2692
rect 12952 2748 13016 2752
rect 12952 2692 12956 2748
rect 12956 2692 13012 2748
rect 13012 2692 13016 2748
rect 12952 2688 13016 2692
rect 13032 2748 13096 2752
rect 13032 2692 13036 2748
rect 13036 2692 13092 2748
rect 13092 2692 13096 2748
rect 13032 2688 13096 2692
rect 13112 2748 13176 2752
rect 13112 2692 13116 2748
rect 13116 2692 13172 2748
rect 13172 2692 13176 2748
rect 13112 2688 13176 2692
rect 13192 2748 13256 2752
rect 13192 2692 13196 2748
rect 13196 2692 13252 2748
rect 13252 2692 13256 2748
rect 13192 2688 13256 2692
rect 22952 2748 23016 2752
rect 22952 2692 22956 2748
rect 22956 2692 23012 2748
rect 23012 2692 23016 2748
rect 22952 2688 23016 2692
rect 23032 2748 23096 2752
rect 23032 2692 23036 2748
rect 23036 2692 23092 2748
rect 23092 2692 23096 2748
rect 23032 2688 23096 2692
rect 23112 2748 23176 2752
rect 23112 2692 23116 2748
rect 23116 2692 23172 2748
rect 23172 2692 23176 2748
rect 23112 2688 23176 2692
rect 23192 2748 23256 2752
rect 23192 2692 23196 2748
rect 23196 2692 23252 2748
rect 23252 2692 23256 2748
rect 23192 2688 23256 2692
rect 32952 2748 33016 2752
rect 32952 2692 32956 2748
rect 32956 2692 33012 2748
rect 33012 2692 33016 2748
rect 32952 2688 33016 2692
rect 33032 2748 33096 2752
rect 33032 2692 33036 2748
rect 33036 2692 33092 2748
rect 33092 2692 33096 2748
rect 33032 2688 33096 2692
rect 33112 2748 33176 2752
rect 33112 2692 33116 2748
rect 33116 2692 33172 2748
rect 33172 2692 33176 2748
rect 33112 2688 33176 2692
rect 33192 2748 33256 2752
rect 33192 2692 33196 2748
rect 33196 2692 33252 2748
rect 33252 2692 33256 2748
rect 33192 2688 33256 2692
rect 42952 2748 43016 2752
rect 42952 2692 42956 2748
rect 42956 2692 43012 2748
rect 43012 2692 43016 2748
rect 42952 2688 43016 2692
rect 43032 2748 43096 2752
rect 43032 2692 43036 2748
rect 43036 2692 43092 2748
rect 43092 2692 43096 2748
rect 43032 2688 43096 2692
rect 43112 2748 43176 2752
rect 43112 2692 43116 2748
rect 43116 2692 43172 2748
rect 43172 2692 43176 2748
rect 43112 2688 43176 2692
rect 43192 2748 43256 2752
rect 43192 2692 43196 2748
rect 43196 2692 43252 2748
rect 43252 2692 43256 2748
rect 43192 2688 43256 2692
rect 22140 2620 22204 2684
rect 22692 2484 22756 2548
rect 7952 2204 8016 2208
rect 7952 2148 7956 2204
rect 7956 2148 8012 2204
rect 8012 2148 8016 2204
rect 7952 2144 8016 2148
rect 8032 2204 8096 2208
rect 8032 2148 8036 2204
rect 8036 2148 8092 2204
rect 8092 2148 8096 2204
rect 8032 2144 8096 2148
rect 8112 2204 8176 2208
rect 8112 2148 8116 2204
rect 8116 2148 8172 2204
rect 8172 2148 8176 2204
rect 8112 2144 8176 2148
rect 8192 2204 8256 2208
rect 8192 2148 8196 2204
rect 8196 2148 8252 2204
rect 8252 2148 8256 2204
rect 8192 2144 8256 2148
rect 17952 2204 18016 2208
rect 17952 2148 17956 2204
rect 17956 2148 18012 2204
rect 18012 2148 18016 2204
rect 17952 2144 18016 2148
rect 18032 2204 18096 2208
rect 18032 2148 18036 2204
rect 18036 2148 18092 2204
rect 18092 2148 18096 2204
rect 18032 2144 18096 2148
rect 18112 2204 18176 2208
rect 18112 2148 18116 2204
rect 18116 2148 18172 2204
rect 18172 2148 18176 2204
rect 18112 2144 18176 2148
rect 18192 2204 18256 2208
rect 18192 2148 18196 2204
rect 18196 2148 18252 2204
rect 18252 2148 18256 2204
rect 18192 2144 18256 2148
rect 27952 2204 28016 2208
rect 27952 2148 27956 2204
rect 27956 2148 28012 2204
rect 28012 2148 28016 2204
rect 27952 2144 28016 2148
rect 28032 2204 28096 2208
rect 28032 2148 28036 2204
rect 28036 2148 28092 2204
rect 28092 2148 28096 2204
rect 28032 2144 28096 2148
rect 28112 2204 28176 2208
rect 28112 2148 28116 2204
rect 28116 2148 28172 2204
rect 28172 2148 28176 2204
rect 28112 2144 28176 2148
rect 28192 2204 28256 2208
rect 28192 2148 28196 2204
rect 28196 2148 28252 2204
rect 28252 2148 28256 2204
rect 28192 2144 28256 2148
rect 37952 2204 38016 2208
rect 37952 2148 37956 2204
rect 37956 2148 38012 2204
rect 38012 2148 38016 2204
rect 37952 2144 38016 2148
rect 38032 2204 38096 2208
rect 38032 2148 38036 2204
rect 38036 2148 38092 2204
rect 38092 2148 38096 2204
rect 38032 2144 38096 2148
rect 38112 2204 38176 2208
rect 38112 2148 38116 2204
rect 38116 2148 38172 2204
rect 38172 2148 38176 2204
rect 38112 2144 38176 2148
rect 38192 2204 38256 2208
rect 38192 2148 38196 2204
rect 38196 2148 38252 2204
rect 38252 2148 38256 2204
rect 38192 2144 38256 2148
rect 47952 2204 48016 2208
rect 47952 2148 47956 2204
rect 47956 2148 48012 2204
rect 48012 2148 48016 2204
rect 47952 2144 48016 2148
rect 48032 2204 48096 2208
rect 48032 2148 48036 2204
rect 48036 2148 48092 2204
rect 48092 2148 48096 2204
rect 48032 2144 48096 2148
rect 48112 2204 48176 2208
rect 48112 2148 48116 2204
rect 48116 2148 48172 2204
rect 48172 2148 48176 2204
rect 48112 2144 48176 2148
rect 48192 2204 48256 2208
rect 48192 2148 48196 2204
rect 48196 2148 48252 2204
rect 48252 2148 48256 2204
rect 48192 2144 48256 2148
<< metal4 >>
rect 2944 53888 3264 54448
rect 2944 53824 2952 53888
rect 3016 53824 3032 53888
rect 3096 53824 3112 53888
rect 3176 53824 3192 53888
rect 3256 53824 3264 53888
rect 2944 52800 3264 53824
rect 2944 52736 2952 52800
rect 3016 52736 3032 52800
rect 3096 52736 3112 52800
rect 3176 52736 3192 52800
rect 3256 52736 3264 52800
rect 2944 51712 3264 52736
rect 2944 51648 2952 51712
rect 3016 51648 3032 51712
rect 3096 51648 3112 51712
rect 3176 51648 3192 51712
rect 3256 51648 3264 51712
rect 2944 50624 3264 51648
rect 2944 50560 2952 50624
rect 3016 50560 3032 50624
rect 3096 50560 3112 50624
rect 3176 50560 3192 50624
rect 3256 50560 3264 50624
rect 2944 49536 3264 50560
rect 2944 49472 2952 49536
rect 3016 49472 3032 49536
rect 3096 49472 3112 49536
rect 3176 49472 3192 49536
rect 3256 49472 3264 49536
rect 2944 48448 3264 49472
rect 2944 48384 2952 48448
rect 3016 48384 3032 48448
rect 3096 48384 3112 48448
rect 3176 48384 3192 48448
rect 3256 48384 3264 48448
rect 2944 47360 3264 48384
rect 2944 47296 2952 47360
rect 3016 47296 3032 47360
rect 3096 47296 3112 47360
rect 3176 47296 3192 47360
rect 3256 47296 3264 47360
rect 2944 46272 3264 47296
rect 2944 46208 2952 46272
rect 3016 46208 3032 46272
rect 3096 46208 3112 46272
rect 3176 46208 3192 46272
rect 3256 46208 3264 46272
rect 2944 45184 3264 46208
rect 2944 45120 2952 45184
rect 3016 45120 3032 45184
rect 3096 45120 3112 45184
rect 3176 45120 3192 45184
rect 3256 45120 3264 45184
rect 2944 44096 3264 45120
rect 2944 44032 2952 44096
rect 3016 44032 3032 44096
rect 3096 44032 3112 44096
rect 3176 44032 3192 44096
rect 3256 44032 3264 44096
rect 2944 43008 3264 44032
rect 2944 42944 2952 43008
rect 3016 42944 3032 43008
rect 3096 42944 3112 43008
rect 3176 42944 3192 43008
rect 3256 42944 3264 43008
rect 2944 41920 3264 42944
rect 2944 41856 2952 41920
rect 3016 41856 3032 41920
rect 3096 41856 3112 41920
rect 3176 41856 3192 41920
rect 3256 41856 3264 41920
rect 2944 40832 3264 41856
rect 2944 40768 2952 40832
rect 3016 40768 3032 40832
rect 3096 40768 3112 40832
rect 3176 40768 3192 40832
rect 3256 40768 3264 40832
rect 2944 39744 3264 40768
rect 2944 39680 2952 39744
rect 3016 39680 3032 39744
rect 3096 39680 3112 39744
rect 3176 39680 3192 39744
rect 3256 39680 3264 39744
rect 2944 38656 3264 39680
rect 2944 38592 2952 38656
rect 3016 38592 3032 38656
rect 3096 38592 3112 38656
rect 3176 38592 3192 38656
rect 3256 38592 3264 38656
rect 2944 37568 3264 38592
rect 2944 37504 2952 37568
rect 3016 37504 3032 37568
rect 3096 37504 3112 37568
rect 3176 37504 3192 37568
rect 3256 37504 3264 37568
rect 2944 36480 3264 37504
rect 2944 36416 2952 36480
rect 3016 36416 3032 36480
rect 3096 36416 3112 36480
rect 3176 36416 3192 36480
rect 3256 36416 3264 36480
rect 2944 35392 3264 36416
rect 2944 35328 2952 35392
rect 3016 35328 3032 35392
rect 3096 35328 3112 35392
rect 3176 35328 3192 35392
rect 3256 35328 3264 35392
rect 2944 34304 3264 35328
rect 2944 34240 2952 34304
rect 3016 34240 3032 34304
rect 3096 34240 3112 34304
rect 3176 34240 3192 34304
rect 3256 34240 3264 34304
rect 2944 33216 3264 34240
rect 2944 33152 2952 33216
rect 3016 33152 3032 33216
rect 3096 33152 3112 33216
rect 3176 33152 3192 33216
rect 3256 33152 3264 33216
rect 2944 32128 3264 33152
rect 2944 32064 2952 32128
rect 3016 32064 3032 32128
rect 3096 32064 3112 32128
rect 3176 32064 3192 32128
rect 3256 32064 3264 32128
rect 2944 31040 3264 32064
rect 2944 30976 2952 31040
rect 3016 30976 3032 31040
rect 3096 30976 3112 31040
rect 3176 30976 3192 31040
rect 3256 30976 3264 31040
rect 2944 29952 3264 30976
rect 2944 29888 2952 29952
rect 3016 29888 3032 29952
rect 3096 29888 3112 29952
rect 3176 29888 3192 29952
rect 3256 29888 3264 29952
rect 2944 28864 3264 29888
rect 2944 28800 2952 28864
rect 3016 28800 3032 28864
rect 3096 28800 3112 28864
rect 3176 28800 3192 28864
rect 3256 28800 3264 28864
rect 2944 27776 3264 28800
rect 2944 27712 2952 27776
rect 3016 27712 3032 27776
rect 3096 27712 3112 27776
rect 3176 27712 3192 27776
rect 3256 27712 3264 27776
rect 2944 26688 3264 27712
rect 2944 26624 2952 26688
rect 3016 26624 3032 26688
rect 3096 26624 3112 26688
rect 3176 26624 3192 26688
rect 3256 26624 3264 26688
rect 2944 25600 3264 26624
rect 2944 25536 2952 25600
rect 3016 25536 3032 25600
rect 3096 25536 3112 25600
rect 3176 25536 3192 25600
rect 3256 25536 3264 25600
rect 2944 24512 3264 25536
rect 2944 24448 2952 24512
rect 3016 24448 3032 24512
rect 3096 24448 3112 24512
rect 3176 24448 3192 24512
rect 3256 24448 3264 24512
rect 2944 23424 3264 24448
rect 2944 23360 2952 23424
rect 3016 23360 3032 23424
rect 3096 23360 3112 23424
rect 3176 23360 3192 23424
rect 3256 23360 3264 23424
rect 2944 22336 3264 23360
rect 2944 22272 2952 22336
rect 3016 22272 3032 22336
rect 3096 22272 3112 22336
rect 3176 22272 3192 22336
rect 3256 22272 3264 22336
rect 2944 21248 3264 22272
rect 2944 21184 2952 21248
rect 3016 21184 3032 21248
rect 3096 21184 3112 21248
rect 3176 21184 3192 21248
rect 3256 21184 3264 21248
rect 2944 20160 3264 21184
rect 2944 20096 2952 20160
rect 3016 20096 3032 20160
rect 3096 20096 3112 20160
rect 3176 20096 3192 20160
rect 3256 20096 3264 20160
rect 2944 19072 3264 20096
rect 2944 19008 2952 19072
rect 3016 19008 3032 19072
rect 3096 19008 3112 19072
rect 3176 19008 3192 19072
rect 3256 19008 3264 19072
rect 2944 17984 3264 19008
rect 2944 17920 2952 17984
rect 3016 17920 3032 17984
rect 3096 17920 3112 17984
rect 3176 17920 3192 17984
rect 3256 17920 3264 17984
rect 2944 16896 3264 17920
rect 2944 16832 2952 16896
rect 3016 16832 3032 16896
rect 3096 16832 3112 16896
rect 3176 16832 3192 16896
rect 3256 16832 3264 16896
rect 2944 15808 3264 16832
rect 2944 15744 2952 15808
rect 3016 15744 3032 15808
rect 3096 15744 3112 15808
rect 3176 15744 3192 15808
rect 3256 15744 3264 15808
rect 2944 14720 3264 15744
rect 2944 14656 2952 14720
rect 3016 14656 3032 14720
rect 3096 14656 3112 14720
rect 3176 14656 3192 14720
rect 3256 14656 3264 14720
rect 2944 13632 3264 14656
rect 2944 13568 2952 13632
rect 3016 13568 3032 13632
rect 3096 13568 3112 13632
rect 3176 13568 3192 13632
rect 3256 13568 3264 13632
rect 2944 12544 3264 13568
rect 2944 12480 2952 12544
rect 3016 12480 3032 12544
rect 3096 12480 3112 12544
rect 3176 12480 3192 12544
rect 3256 12480 3264 12544
rect 2944 11456 3264 12480
rect 2944 11392 2952 11456
rect 3016 11392 3032 11456
rect 3096 11392 3112 11456
rect 3176 11392 3192 11456
rect 3256 11392 3264 11456
rect 2944 10368 3264 11392
rect 2944 10304 2952 10368
rect 3016 10304 3032 10368
rect 3096 10304 3112 10368
rect 3176 10304 3192 10368
rect 3256 10304 3264 10368
rect 2944 9280 3264 10304
rect 2944 9216 2952 9280
rect 3016 9216 3032 9280
rect 3096 9216 3112 9280
rect 3176 9216 3192 9280
rect 3256 9216 3264 9280
rect 2944 8192 3264 9216
rect 2944 8128 2952 8192
rect 3016 8128 3032 8192
rect 3096 8128 3112 8192
rect 3176 8128 3192 8192
rect 3256 8128 3264 8192
rect 2944 7104 3264 8128
rect 2944 7040 2952 7104
rect 3016 7040 3032 7104
rect 3096 7040 3112 7104
rect 3176 7040 3192 7104
rect 3256 7040 3264 7104
rect 2944 6016 3264 7040
rect 2944 5952 2952 6016
rect 3016 5952 3032 6016
rect 3096 5952 3112 6016
rect 3176 5952 3192 6016
rect 3256 5952 3264 6016
rect 2944 4928 3264 5952
rect 2944 4864 2952 4928
rect 3016 4864 3032 4928
rect 3096 4864 3112 4928
rect 3176 4864 3192 4928
rect 3256 4864 3264 4928
rect 2944 3840 3264 4864
rect 2944 3776 2952 3840
rect 3016 3776 3032 3840
rect 3096 3776 3112 3840
rect 3176 3776 3192 3840
rect 3256 3776 3264 3840
rect 2944 2752 3264 3776
rect 2944 2688 2952 2752
rect 3016 2688 3032 2752
rect 3096 2688 3112 2752
rect 3176 2688 3192 2752
rect 3256 2688 3264 2752
rect 2944 2128 3264 2688
rect 7944 54432 8264 54448
rect 7944 54368 7952 54432
rect 8016 54368 8032 54432
rect 8096 54368 8112 54432
rect 8176 54368 8192 54432
rect 8256 54368 8264 54432
rect 7944 53344 8264 54368
rect 7944 53280 7952 53344
rect 8016 53280 8032 53344
rect 8096 53280 8112 53344
rect 8176 53280 8192 53344
rect 8256 53280 8264 53344
rect 7944 52256 8264 53280
rect 7944 52192 7952 52256
rect 8016 52192 8032 52256
rect 8096 52192 8112 52256
rect 8176 52192 8192 52256
rect 8256 52192 8264 52256
rect 7944 51168 8264 52192
rect 7944 51104 7952 51168
rect 8016 51104 8032 51168
rect 8096 51104 8112 51168
rect 8176 51104 8192 51168
rect 8256 51104 8264 51168
rect 7944 50080 8264 51104
rect 7944 50016 7952 50080
rect 8016 50016 8032 50080
rect 8096 50016 8112 50080
rect 8176 50016 8192 50080
rect 8256 50016 8264 50080
rect 7944 48992 8264 50016
rect 7944 48928 7952 48992
rect 8016 48928 8032 48992
rect 8096 48928 8112 48992
rect 8176 48928 8192 48992
rect 8256 48928 8264 48992
rect 7944 47904 8264 48928
rect 7944 47840 7952 47904
rect 8016 47840 8032 47904
rect 8096 47840 8112 47904
rect 8176 47840 8192 47904
rect 8256 47840 8264 47904
rect 7944 46816 8264 47840
rect 7944 46752 7952 46816
rect 8016 46752 8032 46816
rect 8096 46752 8112 46816
rect 8176 46752 8192 46816
rect 8256 46752 8264 46816
rect 7944 45728 8264 46752
rect 7944 45664 7952 45728
rect 8016 45664 8032 45728
rect 8096 45664 8112 45728
rect 8176 45664 8192 45728
rect 8256 45664 8264 45728
rect 7944 44640 8264 45664
rect 7944 44576 7952 44640
rect 8016 44576 8032 44640
rect 8096 44576 8112 44640
rect 8176 44576 8192 44640
rect 8256 44576 8264 44640
rect 7944 43552 8264 44576
rect 7944 43488 7952 43552
rect 8016 43488 8032 43552
rect 8096 43488 8112 43552
rect 8176 43488 8192 43552
rect 8256 43488 8264 43552
rect 7944 42464 8264 43488
rect 7944 42400 7952 42464
rect 8016 42400 8032 42464
rect 8096 42400 8112 42464
rect 8176 42400 8192 42464
rect 8256 42400 8264 42464
rect 7944 41376 8264 42400
rect 7944 41312 7952 41376
rect 8016 41312 8032 41376
rect 8096 41312 8112 41376
rect 8176 41312 8192 41376
rect 8256 41312 8264 41376
rect 7944 40288 8264 41312
rect 7944 40224 7952 40288
rect 8016 40224 8032 40288
rect 8096 40224 8112 40288
rect 8176 40224 8192 40288
rect 8256 40224 8264 40288
rect 7944 39200 8264 40224
rect 7944 39136 7952 39200
rect 8016 39136 8032 39200
rect 8096 39136 8112 39200
rect 8176 39136 8192 39200
rect 8256 39136 8264 39200
rect 7944 38112 8264 39136
rect 7944 38048 7952 38112
rect 8016 38048 8032 38112
rect 8096 38048 8112 38112
rect 8176 38048 8192 38112
rect 8256 38048 8264 38112
rect 7944 37024 8264 38048
rect 7944 36960 7952 37024
rect 8016 36960 8032 37024
rect 8096 36960 8112 37024
rect 8176 36960 8192 37024
rect 8256 36960 8264 37024
rect 7944 35936 8264 36960
rect 7944 35872 7952 35936
rect 8016 35872 8032 35936
rect 8096 35872 8112 35936
rect 8176 35872 8192 35936
rect 8256 35872 8264 35936
rect 7944 34848 8264 35872
rect 7944 34784 7952 34848
rect 8016 34784 8032 34848
rect 8096 34784 8112 34848
rect 8176 34784 8192 34848
rect 8256 34784 8264 34848
rect 7944 33760 8264 34784
rect 7944 33696 7952 33760
rect 8016 33696 8032 33760
rect 8096 33696 8112 33760
rect 8176 33696 8192 33760
rect 8256 33696 8264 33760
rect 7944 32672 8264 33696
rect 7944 32608 7952 32672
rect 8016 32608 8032 32672
rect 8096 32608 8112 32672
rect 8176 32608 8192 32672
rect 8256 32608 8264 32672
rect 7944 31584 8264 32608
rect 7944 31520 7952 31584
rect 8016 31520 8032 31584
rect 8096 31520 8112 31584
rect 8176 31520 8192 31584
rect 8256 31520 8264 31584
rect 7944 30496 8264 31520
rect 7944 30432 7952 30496
rect 8016 30432 8032 30496
rect 8096 30432 8112 30496
rect 8176 30432 8192 30496
rect 8256 30432 8264 30496
rect 7944 29408 8264 30432
rect 7944 29344 7952 29408
rect 8016 29344 8032 29408
rect 8096 29344 8112 29408
rect 8176 29344 8192 29408
rect 8256 29344 8264 29408
rect 7944 28320 8264 29344
rect 7944 28256 7952 28320
rect 8016 28256 8032 28320
rect 8096 28256 8112 28320
rect 8176 28256 8192 28320
rect 8256 28256 8264 28320
rect 7944 27232 8264 28256
rect 7944 27168 7952 27232
rect 8016 27168 8032 27232
rect 8096 27168 8112 27232
rect 8176 27168 8192 27232
rect 8256 27168 8264 27232
rect 7944 26144 8264 27168
rect 7944 26080 7952 26144
rect 8016 26080 8032 26144
rect 8096 26080 8112 26144
rect 8176 26080 8192 26144
rect 8256 26080 8264 26144
rect 7944 25056 8264 26080
rect 7944 24992 7952 25056
rect 8016 24992 8032 25056
rect 8096 24992 8112 25056
rect 8176 24992 8192 25056
rect 8256 24992 8264 25056
rect 7944 23968 8264 24992
rect 7944 23904 7952 23968
rect 8016 23904 8032 23968
rect 8096 23904 8112 23968
rect 8176 23904 8192 23968
rect 8256 23904 8264 23968
rect 7944 22880 8264 23904
rect 7944 22816 7952 22880
rect 8016 22816 8032 22880
rect 8096 22816 8112 22880
rect 8176 22816 8192 22880
rect 8256 22816 8264 22880
rect 7944 21792 8264 22816
rect 7944 21728 7952 21792
rect 8016 21728 8032 21792
rect 8096 21728 8112 21792
rect 8176 21728 8192 21792
rect 8256 21728 8264 21792
rect 7944 20704 8264 21728
rect 7944 20640 7952 20704
rect 8016 20640 8032 20704
rect 8096 20640 8112 20704
rect 8176 20640 8192 20704
rect 8256 20640 8264 20704
rect 7944 19616 8264 20640
rect 7944 19552 7952 19616
rect 8016 19552 8032 19616
rect 8096 19552 8112 19616
rect 8176 19552 8192 19616
rect 8256 19552 8264 19616
rect 7944 18528 8264 19552
rect 7944 18464 7952 18528
rect 8016 18464 8032 18528
rect 8096 18464 8112 18528
rect 8176 18464 8192 18528
rect 8256 18464 8264 18528
rect 7944 17440 8264 18464
rect 7944 17376 7952 17440
rect 8016 17376 8032 17440
rect 8096 17376 8112 17440
rect 8176 17376 8192 17440
rect 8256 17376 8264 17440
rect 7944 16352 8264 17376
rect 7944 16288 7952 16352
rect 8016 16288 8032 16352
rect 8096 16288 8112 16352
rect 8176 16288 8192 16352
rect 8256 16288 8264 16352
rect 7944 15264 8264 16288
rect 7944 15200 7952 15264
rect 8016 15200 8032 15264
rect 8096 15200 8112 15264
rect 8176 15200 8192 15264
rect 8256 15200 8264 15264
rect 7944 14176 8264 15200
rect 7944 14112 7952 14176
rect 8016 14112 8032 14176
rect 8096 14112 8112 14176
rect 8176 14112 8192 14176
rect 8256 14112 8264 14176
rect 7944 13088 8264 14112
rect 7944 13024 7952 13088
rect 8016 13024 8032 13088
rect 8096 13024 8112 13088
rect 8176 13024 8192 13088
rect 8256 13024 8264 13088
rect 7944 12000 8264 13024
rect 7944 11936 7952 12000
rect 8016 11936 8032 12000
rect 8096 11936 8112 12000
rect 8176 11936 8192 12000
rect 8256 11936 8264 12000
rect 7944 10912 8264 11936
rect 7944 10848 7952 10912
rect 8016 10848 8032 10912
rect 8096 10848 8112 10912
rect 8176 10848 8192 10912
rect 8256 10848 8264 10912
rect 7944 9824 8264 10848
rect 7944 9760 7952 9824
rect 8016 9760 8032 9824
rect 8096 9760 8112 9824
rect 8176 9760 8192 9824
rect 8256 9760 8264 9824
rect 7944 8736 8264 9760
rect 7944 8672 7952 8736
rect 8016 8672 8032 8736
rect 8096 8672 8112 8736
rect 8176 8672 8192 8736
rect 8256 8672 8264 8736
rect 7944 7648 8264 8672
rect 7944 7584 7952 7648
rect 8016 7584 8032 7648
rect 8096 7584 8112 7648
rect 8176 7584 8192 7648
rect 8256 7584 8264 7648
rect 7944 6560 8264 7584
rect 7944 6496 7952 6560
rect 8016 6496 8032 6560
rect 8096 6496 8112 6560
rect 8176 6496 8192 6560
rect 8256 6496 8264 6560
rect 7944 5472 8264 6496
rect 7944 5408 7952 5472
rect 8016 5408 8032 5472
rect 8096 5408 8112 5472
rect 8176 5408 8192 5472
rect 8256 5408 8264 5472
rect 7944 4384 8264 5408
rect 7944 4320 7952 4384
rect 8016 4320 8032 4384
rect 8096 4320 8112 4384
rect 8176 4320 8192 4384
rect 8256 4320 8264 4384
rect 7944 3296 8264 4320
rect 7944 3232 7952 3296
rect 8016 3232 8032 3296
rect 8096 3232 8112 3296
rect 8176 3232 8192 3296
rect 8256 3232 8264 3296
rect 7944 2208 8264 3232
rect 7944 2144 7952 2208
rect 8016 2144 8032 2208
rect 8096 2144 8112 2208
rect 8176 2144 8192 2208
rect 8256 2144 8264 2208
rect 7944 2128 8264 2144
rect 12944 53888 13264 54448
rect 12944 53824 12952 53888
rect 13016 53824 13032 53888
rect 13096 53824 13112 53888
rect 13176 53824 13192 53888
rect 13256 53824 13264 53888
rect 12944 52800 13264 53824
rect 12944 52736 12952 52800
rect 13016 52736 13032 52800
rect 13096 52736 13112 52800
rect 13176 52736 13192 52800
rect 13256 52736 13264 52800
rect 12944 51712 13264 52736
rect 12944 51648 12952 51712
rect 13016 51648 13032 51712
rect 13096 51648 13112 51712
rect 13176 51648 13192 51712
rect 13256 51648 13264 51712
rect 12944 50624 13264 51648
rect 12944 50560 12952 50624
rect 13016 50560 13032 50624
rect 13096 50560 13112 50624
rect 13176 50560 13192 50624
rect 13256 50560 13264 50624
rect 12944 49536 13264 50560
rect 12944 49472 12952 49536
rect 13016 49472 13032 49536
rect 13096 49472 13112 49536
rect 13176 49472 13192 49536
rect 13256 49472 13264 49536
rect 12944 48448 13264 49472
rect 12944 48384 12952 48448
rect 13016 48384 13032 48448
rect 13096 48384 13112 48448
rect 13176 48384 13192 48448
rect 13256 48384 13264 48448
rect 12944 47360 13264 48384
rect 12944 47296 12952 47360
rect 13016 47296 13032 47360
rect 13096 47296 13112 47360
rect 13176 47296 13192 47360
rect 13256 47296 13264 47360
rect 12944 46272 13264 47296
rect 12944 46208 12952 46272
rect 13016 46208 13032 46272
rect 13096 46208 13112 46272
rect 13176 46208 13192 46272
rect 13256 46208 13264 46272
rect 12944 45184 13264 46208
rect 12944 45120 12952 45184
rect 13016 45120 13032 45184
rect 13096 45120 13112 45184
rect 13176 45120 13192 45184
rect 13256 45120 13264 45184
rect 12944 44096 13264 45120
rect 12944 44032 12952 44096
rect 13016 44032 13032 44096
rect 13096 44032 13112 44096
rect 13176 44032 13192 44096
rect 13256 44032 13264 44096
rect 12944 43008 13264 44032
rect 12944 42944 12952 43008
rect 13016 42944 13032 43008
rect 13096 42944 13112 43008
rect 13176 42944 13192 43008
rect 13256 42944 13264 43008
rect 12944 41920 13264 42944
rect 12944 41856 12952 41920
rect 13016 41856 13032 41920
rect 13096 41856 13112 41920
rect 13176 41856 13192 41920
rect 13256 41856 13264 41920
rect 12944 40832 13264 41856
rect 12944 40768 12952 40832
rect 13016 40768 13032 40832
rect 13096 40768 13112 40832
rect 13176 40768 13192 40832
rect 13256 40768 13264 40832
rect 12944 39744 13264 40768
rect 12944 39680 12952 39744
rect 13016 39680 13032 39744
rect 13096 39680 13112 39744
rect 13176 39680 13192 39744
rect 13256 39680 13264 39744
rect 12944 38656 13264 39680
rect 12944 38592 12952 38656
rect 13016 38592 13032 38656
rect 13096 38592 13112 38656
rect 13176 38592 13192 38656
rect 13256 38592 13264 38656
rect 12944 37568 13264 38592
rect 12944 37504 12952 37568
rect 13016 37504 13032 37568
rect 13096 37504 13112 37568
rect 13176 37504 13192 37568
rect 13256 37504 13264 37568
rect 12944 36480 13264 37504
rect 12944 36416 12952 36480
rect 13016 36416 13032 36480
rect 13096 36416 13112 36480
rect 13176 36416 13192 36480
rect 13256 36416 13264 36480
rect 12944 35392 13264 36416
rect 12944 35328 12952 35392
rect 13016 35328 13032 35392
rect 13096 35328 13112 35392
rect 13176 35328 13192 35392
rect 13256 35328 13264 35392
rect 12944 34304 13264 35328
rect 12944 34240 12952 34304
rect 13016 34240 13032 34304
rect 13096 34240 13112 34304
rect 13176 34240 13192 34304
rect 13256 34240 13264 34304
rect 12944 33216 13264 34240
rect 12944 33152 12952 33216
rect 13016 33152 13032 33216
rect 13096 33152 13112 33216
rect 13176 33152 13192 33216
rect 13256 33152 13264 33216
rect 12944 32128 13264 33152
rect 12944 32064 12952 32128
rect 13016 32064 13032 32128
rect 13096 32064 13112 32128
rect 13176 32064 13192 32128
rect 13256 32064 13264 32128
rect 12944 31040 13264 32064
rect 12944 30976 12952 31040
rect 13016 30976 13032 31040
rect 13096 30976 13112 31040
rect 13176 30976 13192 31040
rect 13256 30976 13264 31040
rect 12944 29952 13264 30976
rect 12944 29888 12952 29952
rect 13016 29888 13032 29952
rect 13096 29888 13112 29952
rect 13176 29888 13192 29952
rect 13256 29888 13264 29952
rect 12944 28864 13264 29888
rect 12944 28800 12952 28864
rect 13016 28800 13032 28864
rect 13096 28800 13112 28864
rect 13176 28800 13192 28864
rect 13256 28800 13264 28864
rect 12944 27776 13264 28800
rect 12944 27712 12952 27776
rect 13016 27712 13032 27776
rect 13096 27712 13112 27776
rect 13176 27712 13192 27776
rect 13256 27712 13264 27776
rect 12944 26688 13264 27712
rect 12944 26624 12952 26688
rect 13016 26624 13032 26688
rect 13096 26624 13112 26688
rect 13176 26624 13192 26688
rect 13256 26624 13264 26688
rect 12944 25600 13264 26624
rect 12944 25536 12952 25600
rect 13016 25536 13032 25600
rect 13096 25536 13112 25600
rect 13176 25536 13192 25600
rect 13256 25536 13264 25600
rect 12944 24512 13264 25536
rect 12944 24448 12952 24512
rect 13016 24448 13032 24512
rect 13096 24448 13112 24512
rect 13176 24448 13192 24512
rect 13256 24448 13264 24512
rect 12944 23424 13264 24448
rect 12944 23360 12952 23424
rect 13016 23360 13032 23424
rect 13096 23360 13112 23424
rect 13176 23360 13192 23424
rect 13256 23360 13264 23424
rect 12944 22336 13264 23360
rect 12944 22272 12952 22336
rect 13016 22272 13032 22336
rect 13096 22272 13112 22336
rect 13176 22272 13192 22336
rect 13256 22272 13264 22336
rect 12944 21248 13264 22272
rect 12944 21184 12952 21248
rect 13016 21184 13032 21248
rect 13096 21184 13112 21248
rect 13176 21184 13192 21248
rect 13256 21184 13264 21248
rect 12944 20160 13264 21184
rect 12944 20096 12952 20160
rect 13016 20096 13032 20160
rect 13096 20096 13112 20160
rect 13176 20096 13192 20160
rect 13256 20096 13264 20160
rect 12944 19072 13264 20096
rect 12944 19008 12952 19072
rect 13016 19008 13032 19072
rect 13096 19008 13112 19072
rect 13176 19008 13192 19072
rect 13256 19008 13264 19072
rect 12944 17984 13264 19008
rect 12944 17920 12952 17984
rect 13016 17920 13032 17984
rect 13096 17920 13112 17984
rect 13176 17920 13192 17984
rect 13256 17920 13264 17984
rect 12944 16896 13264 17920
rect 12944 16832 12952 16896
rect 13016 16832 13032 16896
rect 13096 16832 13112 16896
rect 13176 16832 13192 16896
rect 13256 16832 13264 16896
rect 12944 15808 13264 16832
rect 12944 15744 12952 15808
rect 13016 15744 13032 15808
rect 13096 15744 13112 15808
rect 13176 15744 13192 15808
rect 13256 15744 13264 15808
rect 12944 14720 13264 15744
rect 12944 14656 12952 14720
rect 13016 14656 13032 14720
rect 13096 14656 13112 14720
rect 13176 14656 13192 14720
rect 13256 14656 13264 14720
rect 12944 13632 13264 14656
rect 12944 13568 12952 13632
rect 13016 13568 13032 13632
rect 13096 13568 13112 13632
rect 13176 13568 13192 13632
rect 13256 13568 13264 13632
rect 12944 12544 13264 13568
rect 12944 12480 12952 12544
rect 13016 12480 13032 12544
rect 13096 12480 13112 12544
rect 13176 12480 13192 12544
rect 13256 12480 13264 12544
rect 12944 11456 13264 12480
rect 12944 11392 12952 11456
rect 13016 11392 13032 11456
rect 13096 11392 13112 11456
rect 13176 11392 13192 11456
rect 13256 11392 13264 11456
rect 12944 10368 13264 11392
rect 12944 10304 12952 10368
rect 13016 10304 13032 10368
rect 13096 10304 13112 10368
rect 13176 10304 13192 10368
rect 13256 10304 13264 10368
rect 12944 9280 13264 10304
rect 12944 9216 12952 9280
rect 13016 9216 13032 9280
rect 13096 9216 13112 9280
rect 13176 9216 13192 9280
rect 13256 9216 13264 9280
rect 12944 8192 13264 9216
rect 12944 8128 12952 8192
rect 13016 8128 13032 8192
rect 13096 8128 13112 8192
rect 13176 8128 13192 8192
rect 13256 8128 13264 8192
rect 12944 7104 13264 8128
rect 12944 7040 12952 7104
rect 13016 7040 13032 7104
rect 13096 7040 13112 7104
rect 13176 7040 13192 7104
rect 13256 7040 13264 7104
rect 12944 6016 13264 7040
rect 12944 5952 12952 6016
rect 13016 5952 13032 6016
rect 13096 5952 13112 6016
rect 13176 5952 13192 6016
rect 13256 5952 13264 6016
rect 12944 4928 13264 5952
rect 12944 4864 12952 4928
rect 13016 4864 13032 4928
rect 13096 4864 13112 4928
rect 13176 4864 13192 4928
rect 13256 4864 13264 4928
rect 12944 3840 13264 4864
rect 12944 3776 12952 3840
rect 13016 3776 13032 3840
rect 13096 3776 13112 3840
rect 13176 3776 13192 3840
rect 13256 3776 13264 3840
rect 12944 2752 13264 3776
rect 12944 2688 12952 2752
rect 13016 2688 13032 2752
rect 13096 2688 13112 2752
rect 13176 2688 13192 2752
rect 13256 2688 13264 2752
rect 12944 2128 13264 2688
rect 17944 54432 18264 54448
rect 17944 54368 17952 54432
rect 18016 54368 18032 54432
rect 18096 54368 18112 54432
rect 18176 54368 18192 54432
rect 18256 54368 18264 54432
rect 17944 53344 18264 54368
rect 17944 53280 17952 53344
rect 18016 53280 18032 53344
rect 18096 53280 18112 53344
rect 18176 53280 18192 53344
rect 18256 53280 18264 53344
rect 17944 52256 18264 53280
rect 17944 52192 17952 52256
rect 18016 52192 18032 52256
rect 18096 52192 18112 52256
rect 18176 52192 18192 52256
rect 18256 52192 18264 52256
rect 17944 51168 18264 52192
rect 17944 51104 17952 51168
rect 18016 51104 18032 51168
rect 18096 51104 18112 51168
rect 18176 51104 18192 51168
rect 18256 51104 18264 51168
rect 17944 50080 18264 51104
rect 17944 50016 17952 50080
rect 18016 50016 18032 50080
rect 18096 50016 18112 50080
rect 18176 50016 18192 50080
rect 18256 50016 18264 50080
rect 17944 48992 18264 50016
rect 17944 48928 17952 48992
rect 18016 48928 18032 48992
rect 18096 48928 18112 48992
rect 18176 48928 18192 48992
rect 18256 48928 18264 48992
rect 17944 47904 18264 48928
rect 17944 47840 17952 47904
rect 18016 47840 18032 47904
rect 18096 47840 18112 47904
rect 18176 47840 18192 47904
rect 18256 47840 18264 47904
rect 17944 46816 18264 47840
rect 17944 46752 17952 46816
rect 18016 46752 18032 46816
rect 18096 46752 18112 46816
rect 18176 46752 18192 46816
rect 18256 46752 18264 46816
rect 17944 45728 18264 46752
rect 17944 45664 17952 45728
rect 18016 45664 18032 45728
rect 18096 45664 18112 45728
rect 18176 45664 18192 45728
rect 18256 45664 18264 45728
rect 17944 44640 18264 45664
rect 17944 44576 17952 44640
rect 18016 44576 18032 44640
rect 18096 44576 18112 44640
rect 18176 44576 18192 44640
rect 18256 44576 18264 44640
rect 17944 43552 18264 44576
rect 17944 43488 17952 43552
rect 18016 43488 18032 43552
rect 18096 43488 18112 43552
rect 18176 43488 18192 43552
rect 18256 43488 18264 43552
rect 17944 42464 18264 43488
rect 17944 42400 17952 42464
rect 18016 42400 18032 42464
rect 18096 42400 18112 42464
rect 18176 42400 18192 42464
rect 18256 42400 18264 42464
rect 17944 41376 18264 42400
rect 17944 41312 17952 41376
rect 18016 41312 18032 41376
rect 18096 41312 18112 41376
rect 18176 41312 18192 41376
rect 18256 41312 18264 41376
rect 17944 40288 18264 41312
rect 17944 40224 17952 40288
rect 18016 40224 18032 40288
rect 18096 40224 18112 40288
rect 18176 40224 18192 40288
rect 18256 40224 18264 40288
rect 17944 39200 18264 40224
rect 17944 39136 17952 39200
rect 18016 39136 18032 39200
rect 18096 39136 18112 39200
rect 18176 39136 18192 39200
rect 18256 39136 18264 39200
rect 17944 38112 18264 39136
rect 17944 38048 17952 38112
rect 18016 38048 18032 38112
rect 18096 38048 18112 38112
rect 18176 38048 18192 38112
rect 18256 38048 18264 38112
rect 17944 37024 18264 38048
rect 17944 36960 17952 37024
rect 18016 36960 18032 37024
rect 18096 36960 18112 37024
rect 18176 36960 18192 37024
rect 18256 36960 18264 37024
rect 17944 35936 18264 36960
rect 17944 35872 17952 35936
rect 18016 35872 18032 35936
rect 18096 35872 18112 35936
rect 18176 35872 18192 35936
rect 18256 35872 18264 35936
rect 17944 34848 18264 35872
rect 17944 34784 17952 34848
rect 18016 34784 18032 34848
rect 18096 34784 18112 34848
rect 18176 34784 18192 34848
rect 18256 34784 18264 34848
rect 17944 33760 18264 34784
rect 17944 33696 17952 33760
rect 18016 33696 18032 33760
rect 18096 33696 18112 33760
rect 18176 33696 18192 33760
rect 18256 33696 18264 33760
rect 17944 32672 18264 33696
rect 17944 32608 17952 32672
rect 18016 32608 18032 32672
rect 18096 32608 18112 32672
rect 18176 32608 18192 32672
rect 18256 32608 18264 32672
rect 17944 31584 18264 32608
rect 17944 31520 17952 31584
rect 18016 31520 18032 31584
rect 18096 31520 18112 31584
rect 18176 31520 18192 31584
rect 18256 31520 18264 31584
rect 17944 30496 18264 31520
rect 22944 53888 23264 54448
rect 27944 54432 28264 54448
rect 27944 54368 27952 54432
rect 28016 54368 28032 54432
rect 28096 54368 28112 54432
rect 28176 54368 28192 54432
rect 28256 54368 28264 54432
rect 25083 53956 25149 53957
rect 25083 53892 25084 53956
rect 25148 53892 25149 53956
rect 25083 53891 25149 53892
rect 22944 53824 22952 53888
rect 23016 53824 23032 53888
rect 23096 53824 23112 53888
rect 23176 53824 23192 53888
rect 23256 53824 23264 53888
rect 22944 52800 23264 53824
rect 22944 52736 22952 52800
rect 23016 52736 23032 52800
rect 23096 52736 23112 52800
rect 23176 52736 23192 52800
rect 23256 52736 23264 52800
rect 22944 51712 23264 52736
rect 22944 51648 22952 51712
rect 23016 51648 23032 51712
rect 23096 51648 23112 51712
rect 23176 51648 23192 51712
rect 23256 51648 23264 51712
rect 22944 50624 23264 51648
rect 22944 50560 22952 50624
rect 23016 50560 23032 50624
rect 23096 50560 23112 50624
rect 23176 50560 23192 50624
rect 23256 50560 23264 50624
rect 22944 49536 23264 50560
rect 22944 49472 22952 49536
rect 23016 49472 23032 49536
rect 23096 49472 23112 49536
rect 23176 49472 23192 49536
rect 23256 49472 23264 49536
rect 22944 48448 23264 49472
rect 22944 48384 22952 48448
rect 23016 48384 23032 48448
rect 23096 48384 23112 48448
rect 23176 48384 23192 48448
rect 23256 48384 23264 48448
rect 22944 47360 23264 48384
rect 22944 47296 22952 47360
rect 23016 47296 23032 47360
rect 23096 47296 23112 47360
rect 23176 47296 23192 47360
rect 23256 47296 23264 47360
rect 22944 46272 23264 47296
rect 22944 46208 22952 46272
rect 23016 46208 23032 46272
rect 23096 46208 23112 46272
rect 23176 46208 23192 46272
rect 23256 46208 23264 46272
rect 22944 45184 23264 46208
rect 22944 45120 22952 45184
rect 23016 45120 23032 45184
rect 23096 45120 23112 45184
rect 23176 45120 23192 45184
rect 23256 45120 23264 45184
rect 22944 44096 23264 45120
rect 22944 44032 22952 44096
rect 23016 44032 23032 44096
rect 23096 44032 23112 44096
rect 23176 44032 23192 44096
rect 23256 44032 23264 44096
rect 22944 43008 23264 44032
rect 22944 42944 22952 43008
rect 23016 42944 23032 43008
rect 23096 42944 23112 43008
rect 23176 42944 23192 43008
rect 23256 42944 23264 43008
rect 22944 41920 23264 42944
rect 22944 41856 22952 41920
rect 23016 41856 23032 41920
rect 23096 41856 23112 41920
rect 23176 41856 23192 41920
rect 23256 41856 23264 41920
rect 22944 40832 23264 41856
rect 22944 40768 22952 40832
rect 23016 40768 23032 40832
rect 23096 40768 23112 40832
rect 23176 40768 23192 40832
rect 23256 40768 23264 40832
rect 22944 39744 23264 40768
rect 22944 39680 22952 39744
rect 23016 39680 23032 39744
rect 23096 39680 23112 39744
rect 23176 39680 23192 39744
rect 23256 39680 23264 39744
rect 22944 38656 23264 39680
rect 22944 38592 22952 38656
rect 23016 38592 23032 38656
rect 23096 38592 23112 38656
rect 23176 38592 23192 38656
rect 23256 38592 23264 38656
rect 22944 37568 23264 38592
rect 22944 37504 22952 37568
rect 23016 37504 23032 37568
rect 23096 37504 23112 37568
rect 23176 37504 23192 37568
rect 23256 37504 23264 37568
rect 22944 36480 23264 37504
rect 22944 36416 22952 36480
rect 23016 36416 23032 36480
rect 23096 36416 23112 36480
rect 23176 36416 23192 36480
rect 23256 36416 23264 36480
rect 22944 35392 23264 36416
rect 22944 35328 22952 35392
rect 23016 35328 23032 35392
rect 23096 35328 23112 35392
rect 23176 35328 23192 35392
rect 23256 35328 23264 35392
rect 22944 34304 23264 35328
rect 22944 34240 22952 34304
rect 23016 34240 23032 34304
rect 23096 34240 23112 34304
rect 23176 34240 23192 34304
rect 23256 34240 23264 34304
rect 22944 33216 23264 34240
rect 22944 33152 22952 33216
rect 23016 33152 23032 33216
rect 23096 33152 23112 33216
rect 23176 33152 23192 33216
rect 23256 33152 23264 33216
rect 22944 32128 23264 33152
rect 22944 32064 22952 32128
rect 23016 32064 23032 32128
rect 23096 32064 23112 32128
rect 23176 32064 23192 32128
rect 23256 32064 23264 32128
rect 22507 31244 22573 31245
rect 22507 31180 22508 31244
rect 22572 31180 22573 31244
rect 22507 31179 22573 31180
rect 17944 30432 17952 30496
rect 18016 30432 18032 30496
rect 18096 30432 18112 30496
rect 18176 30432 18192 30496
rect 18256 30432 18264 30496
rect 17944 29408 18264 30432
rect 17944 29344 17952 29408
rect 18016 29344 18032 29408
rect 18096 29344 18112 29408
rect 18176 29344 18192 29408
rect 18256 29344 18264 29408
rect 17944 28320 18264 29344
rect 17944 28256 17952 28320
rect 18016 28256 18032 28320
rect 18096 28256 18112 28320
rect 18176 28256 18192 28320
rect 18256 28256 18264 28320
rect 17944 27232 18264 28256
rect 17944 27168 17952 27232
rect 18016 27168 18032 27232
rect 18096 27168 18112 27232
rect 18176 27168 18192 27232
rect 18256 27168 18264 27232
rect 17944 26144 18264 27168
rect 17944 26080 17952 26144
rect 18016 26080 18032 26144
rect 18096 26080 18112 26144
rect 18176 26080 18192 26144
rect 18256 26080 18264 26144
rect 17944 25056 18264 26080
rect 17944 24992 17952 25056
rect 18016 24992 18032 25056
rect 18096 24992 18112 25056
rect 18176 24992 18192 25056
rect 18256 24992 18264 25056
rect 17944 23968 18264 24992
rect 17944 23904 17952 23968
rect 18016 23904 18032 23968
rect 18096 23904 18112 23968
rect 18176 23904 18192 23968
rect 18256 23904 18264 23968
rect 17944 22880 18264 23904
rect 22139 23628 22205 23629
rect 22139 23564 22140 23628
rect 22204 23564 22205 23628
rect 22139 23563 22205 23564
rect 17944 22816 17952 22880
rect 18016 22816 18032 22880
rect 18096 22816 18112 22880
rect 18176 22816 18192 22880
rect 18256 22816 18264 22880
rect 17944 21792 18264 22816
rect 17944 21728 17952 21792
rect 18016 21728 18032 21792
rect 18096 21728 18112 21792
rect 18176 21728 18192 21792
rect 18256 21728 18264 21792
rect 17944 20704 18264 21728
rect 17944 20640 17952 20704
rect 18016 20640 18032 20704
rect 18096 20640 18112 20704
rect 18176 20640 18192 20704
rect 18256 20640 18264 20704
rect 17944 19616 18264 20640
rect 17944 19552 17952 19616
rect 18016 19552 18032 19616
rect 18096 19552 18112 19616
rect 18176 19552 18192 19616
rect 18256 19552 18264 19616
rect 17944 18528 18264 19552
rect 17944 18464 17952 18528
rect 18016 18464 18032 18528
rect 18096 18464 18112 18528
rect 18176 18464 18192 18528
rect 18256 18464 18264 18528
rect 17944 17440 18264 18464
rect 17944 17376 17952 17440
rect 18016 17376 18032 17440
rect 18096 17376 18112 17440
rect 18176 17376 18192 17440
rect 18256 17376 18264 17440
rect 17944 16352 18264 17376
rect 17944 16288 17952 16352
rect 18016 16288 18032 16352
rect 18096 16288 18112 16352
rect 18176 16288 18192 16352
rect 18256 16288 18264 16352
rect 17944 15264 18264 16288
rect 17944 15200 17952 15264
rect 18016 15200 18032 15264
rect 18096 15200 18112 15264
rect 18176 15200 18192 15264
rect 18256 15200 18264 15264
rect 17944 14176 18264 15200
rect 17944 14112 17952 14176
rect 18016 14112 18032 14176
rect 18096 14112 18112 14176
rect 18176 14112 18192 14176
rect 18256 14112 18264 14176
rect 17944 13088 18264 14112
rect 17944 13024 17952 13088
rect 18016 13024 18032 13088
rect 18096 13024 18112 13088
rect 18176 13024 18192 13088
rect 18256 13024 18264 13088
rect 17944 12000 18264 13024
rect 17944 11936 17952 12000
rect 18016 11936 18032 12000
rect 18096 11936 18112 12000
rect 18176 11936 18192 12000
rect 18256 11936 18264 12000
rect 17944 10912 18264 11936
rect 17944 10848 17952 10912
rect 18016 10848 18032 10912
rect 18096 10848 18112 10912
rect 18176 10848 18192 10912
rect 18256 10848 18264 10912
rect 17944 9824 18264 10848
rect 17944 9760 17952 9824
rect 18016 9760 18032 9824
rect 18096 9760 18112 9824
rect 18176 9760 18192 9824
rect 18256 9760 18264 9824
rect 17944 8736 18264 9760
rect 17944 8672 17952 8736
rect 18016 8672 18032 8736
rect 18096 8672 18112 8736
rect 18176 8672 18192 8736
rect 18256 8672 18264 8736
rect 17944 7648 18264 8672
rect 17944 7584 17952 7648
rect 18016 7584 18032 7648
rect 18096 7584 18112 7648
rect 18176 7584 18192 7648
rect 18256 7584 18264 7648
rect 17944 6560 18264 7584
rect 17944 6496 17952 6560
rect 18016 6496 18032 6560
rect 18096 6496 18112 6560
rect 18176 6496 18192 6560
rect 18256 6496 18264 6560
rect 17944 5472 18264 6496
rect 17944 5408 17952 5472
rect 18016 5408 18032 5472
rect 18096 5408 18112 5472
rect 18176 5408 18192 5472
rect 18256 5408 18264 5472
rect 17944 4384 18264 5408
rect 17944 4320 17952 4384
rect 18016 4320 18032 4384
rect 18096 4320 18112 4384
rect 18176 4320 18192 4384
rect 18256 4320 18264 4384
rect 17944 3296 18264 4320
rect 17944 3232 17952 3296
rect 18016 3232 18032 3296
rect 18096 3232 18112 3296
rect 18176 3232 18192 3296
rect 18256 3232 18264 3296
rect 17944 2208 18264 3232
rect 22142 2685 22202 23563
rect 22510 22949 22570 31179
rect 22944 31040 23264 32064
rect 22944 30976 22952 31040
rect 23016 30976 23032 31040
rect 23096 30976 23112 31040
rect 23176 30976 23192 31040
rect 23256 30976 23264 31040
rect 22944 29952 23264 30976
rect 25086 30429 25146 53891
rect 27944 53344 28264 54368
rect 27944 53280 27952 53344
rect 28016 53280 28032 53344
rect 28096 53280 28112 53344
rect 28176 53280 28192 53344
rect 28256 53280 28264 53344
rect 27944 52256 28264 53280
rect 27944 52192 27952 52256
rect 28016 52192 28032 52256
rect 28096 52192 28112 52256
rect 28176 52192 28192 52256
rect 28256 52192 28264 52256
rect 27944 51168 28264 52192
rect 27944 51104 27952 51168
rect 28016 51104 28032 51168
rect 28096 51104 28112 51168
rect 28176 51104 28192 51168
rect 28256 51104 28264 51168
rect 27944 50080 28264 51104
rect 27944 50016 27952 50080
rect 28016 50016 28032 50080
rect 28096 50016 28112 50080
rect 28176 50016 28192 50080
rect 28256 50016 28264 50080
rect 27944 48992 28264 50016
rect 27944 48928 27952 48992
rect 28016 48928 28032 48992
rect 28096 48928 28112 48992
rect 28176 48928 28192 48992
rect 28256 48928 28264 48992
rect 27944 47904 28264 48928
rect 27944 47840 27952 47904
rect 28016 47840 28032 47904
rect 28096 47840 28112 47904
rect 28176 47840 28192 47904
rect 28256 47840 28264 47904
rect 27944 46816 28264 47840
rect 27944 46752 27952 46816
rect 28016 46752 28032 46816
rect 28096 46752 28112 46816
rect 28176 46752 28192 46816
rect 28256 46752 28264 46816
rect 27944 45728 28264 46752
rect 27944 45664 27952 45728
rect 28016 45664 28032 45728
rect 28096 45664 28112 45728
rect 28176 45664 28192 45728
rect 28256 45664 28264 45728
rect 27944 44640 28264 45664
rect 27944 44576 27952 44640
rect 28016 44576 28032 44640
rect 28096 44576 28112 44640
rect 28176 44576 28192 44640
rect 28256 44576 28264 44640
rect 27944 43552 28264 44576
rect 27944 43488 27952 43552
rect 28016 43488 28032 43552
rect 28096 43488 28112 43552
rect 28176 43488 28192 43552
rect 28256 43488 28264 43552
rect 27944 42464 28264 43488
rect 27944 42400 27952 42464
rect 28016 42400 28032 42464
rect 28096 42400 28112 42464
rect 28176 42400 28192 42464
rect 28256 42400 28264 42464
rect 27944 41376 28264 42400
rect 27944 41312 27952 41376
rect 28016 41312 28032 41376
rect 28096 41312 28112 41376
rect 28176 41312 28192 41376
rect 28256 41312 28264 41376
rect 27944 40288 28264 41312
rect 27944 40224 27952 40288
rect 28016 40224 28032 40288
rect 28096 40224 28112 40288
rect 28176 40224 28192 40288
rect 28256 40224 28264 40288
rect 27944 39200 28264 40224
rect 32944 53888 33264 54448
rect 32944 53824 32952 53888
rect 33016 53824 33032 53888
rect 33096 53824 33112 53888
rect 33176 53824 33192 53888
rect 33256 53824 33264 53888
rect 32944 52800 33264 53824
rect 32944 52736 32952 52800
rect 33016 52736 33032 52800
rect 33096 52736 33112 52800
rect 33176 52736 33192 52800
rect 33256 52736 33264 52800
rect 32944 51712 33264 52736
rect 32944 51648 32952 51712
rect 33016 51648 33032 51712
rect 33096 51648 33112 51712
rect 33176 51648 33192 51712
rect 33256 51648 33264 51712
rect 32944 50624 33264 51648
rect 32944 50560 32952 50624
rect 33016 50560 33032 50624
rect 33096 50560 33112 50624
rect 33176 50560 33192 50624
rect 33256 50560 33264 50624
rect 32944 49536 33264 50560
rect 32944 49472 32952 49536
rect 33016 49472 33032 49536
rect 33096 49472 33112 49536
rect 33176 49472 33192 49536
rect 33256 49472 33264 49536
rect 32944 48448 33264 49472
rect 32944 48384 32952 48448
rect 33016 48384 33032 48448
rect 33096 48384 33112 48448
rect 33176 48384 33192 48448
rect 33256 48384 33264 48448
rect 32944 47360 33264 48384
rect 32944 47296 32952 47360
rect 33016 47296 33032 47360
rect 33096 47296 33112 47360
rect 33176 47296 33192 47360
rect 33256 47296 33264 47360
rect 32944 46272 33264 47296
rect 32944 46208 32952 46272
rect 33016 46208 33032 46272
rect 33096 46208 33112 46272
rect 33176 46208 33192 46272
rect 33256 46208 33264 46272
rect 32944 45184 33264 46208
rect 32944 45120 32952 45184
rect 33016 45120 33032 45184
rect 33096 45120 33112 45184
rect 33176 45120 33192 45184
rect 33256 45120 33264 45184
rect 32944 44096 33264 45120
rect 32944 44032 32952 44096
rect 33016 44032 33032 44096
rect 33096 44032 33112 44096
rect 33176 44032 33192 44096
rect 33256 44032 33264 44096
rect 32944 43008 33264 44032
rect 32944 42944 32952 43008
rect 33016 42944 33032 43008
rect 33096 42944 33112 43008
rect 33176 42944 33192 43008
rect 33256 42944 33264 43008
rect 32944 41920 33264 42944
rect 32944 41856 32952 41920
rect 33016 41856 33032 41920
rect 33096 41856 33112 41920
rect 33176 41856 33192 41920
rect 33256 41856 33264 41920
rect 32944 40832 33264 41856
rect 32944 40768 32952 40832
rect 33016 40768 33032 40832
rect 33096 40768 33112 40832
rect 33176 40768 33192 40832
rect 33256 40768 33264 40832
rect 30419 40084 30485 40085
rect 30419 40020 30420 40084
rect 30484 40020 30485 40084
rect 30419 40019 30485 40020
rect 27944 39136 27952 39200
rect 28016 39136 28032 39200
rect 28096 39136 28112 39200
rect 28176 39136 28192 39200
rect 28256 39136 28264 39200
rect 27944 38112 28264 39136
rect 27944 38048 27952 38112
rect 28016 38048 28032 38112
rect 28096 38048 28112 38112
rect 28176 38048 28192 38112
rect 28256 38048 28264 38112
rect 27944 37024 28264 38048
rect 27944 36960 27952 37024
rect 28016 36960 28032 37024
rect 28096 36960 28112 37024
rect 28176 36960 28192 37024
rect 28256 36960 28264 37024
rect 25635 36004 25701 36005
rect 25635 35940 25636 36004
rect 25700 35940 25701 36004
rect 25635 35939 25701 35940
rect 25083 30428 25149 30429
rect 25083 30364 25084 30428
rect 25148 30364 25149 30428
rect 25083 30363 25149 30364
rect 22944 29888 22952 29952
rect 23016 29888 23032 29952
rect 23096 29888 23112 29952
rect 23176 29888 23192 29952
rect 23256 29888 23264 29952
rect 22944 28864 23264 29888
rect 22944 28800 22952 28864
rect 23016 28800 23032 28864
rect 23096 28800 23112 28864
rect 23176 28800 23192 28864
rect 23256 28800 23264 28864
rect 22944 27776 23264 28800
rect 22944 27712 22952 27776
rect 23016 27712 23032 27776
rect 23096 27712 23112 27776
rect 23176 27712 23192 27776
rect 23256 27712 23264 27776
rect 22944 26688 23264 27712
rect 22944 26624 22952 26688
rect 23016 26624 23032 26688
rect 23096 26624 23112 26688
rect 23176 26624 23192 26688
rect 23256 26624 23264 26688
rect 22944 25600 23264 26624
rect 22944 25536 22952 25600
rect 23016 25536 23032 25600
rect 23096 25536 23112 25600
rect 23176 25536 23192 25600
rect 23256 25536 23264 25600
rect 22944 24512 23264 25536
rect 22944 24448 22952 24512
rect 23016 24448 23032 24512
rect 23096 24448 23112 24512
rect 23176 24448 23192 24512
rect 23256 24448 23264 24512
rect 22944 23424 23264 24448
rect 25638 24309 25698 35939
rect 27944 35936 28264 36960
rect 27944 35872 27952 35936
rect 28016 35872 28032 35936
rect 28096 35872 28112 35936
rect 28176 35872 28192 35936
rect 28256 35872 28264 35936
rect 27944 34848 28264 35872
rect 28763 35732 28829 35733
rect 28763 35668 28764 35732
rect 28828 35668 28829 35732
rect 28763 35667 28829 35668
rect 28579 35052 28645 35053
rect 28579 34988 28580 35052
rect 28644 34988 28645 35052
rect 28579 34987 28645 34988
rect 27944 34784 27952 34848
rect 28016 34784 28032 34848
rect 28096 34784 28112 34848
rect 28176 34784 28192 34848
rect 28256 34784 28264 34848
rect 27944 33760 28264 34784
rect 27944 33696 27952 33760
rect 28016 33696 28032 33760
rect 28096 33696 28112 33760
rect 28176 33696 28192 33760
rect 28256 33696 28264 33760
rect 27944 32672 28264 33696
rect 27944 32608 27952 32672
rect 28016 32608 28032 32672
rect 28096 32608 28112 32672
rect 28176 32608 28192 32672
rect 28256 32608 28264 32672
rect 27944 31584 28264 32608
rect 28582 32197 28642 34987
rect 28579 32196 28645 32197
rect 28579 32132 28580 32196
rect 28644 32132 28645 32196
rect 28579 32131 28645 32132
rect 27944 31520 27952 31584
rect 28016 31520 28032 31584
rect 28096 31520 28112 31584
rect 28176 31520 28192 31584
rect 28256 31520 28264 31584
rect 27944 30496 28264 31520
rect 27944 30432 27952 30496
rect 28016 30432 28032 30496
rect 28096 30432 28112 30496
rect 28176 30432 28192 30496
rect 28256 30432 28264 30496
rect 27944 29408 28264 30432
rect 28766 30157 28826 35667
rect 28763 30156 28829 30157
rect 28763 30092 28764 30156
rect 28828 30092 28829 30156
rect 28763 30091 28829 30092
rect 27944 29344 27952 29408
rect 28016 29344 28032 29408
rect 28096 29344 28112 29408
rect 28176 29344 28192 29408
rect 28256 29344 28264 29408
rect 27944 28320 28264 29344
rect 27944 28256 27952 28320
rect 28016 28256 28032 28320
rect 28096 28256 28112 28320
rect 28176 28256 28192 28320
rect 28256 28256 28264 28320
rect 27659 28252 27725 28253
rect 27659 28188 27660 28252
rect 27724 28188 27725 28252
rect 27659 28187 27725 28188
rect 27107 27708 27173 27709
rect 27107 27644 27108 27708
rect 27172 27644 27173 27708
rect 27107 27643 27173 27644
rect 25635 24308 25701 24309
rect 25635 24244 25636 24308
rect 25700 24244 25701 24308
rect 25635 24243 25701 24244
rect 22944 23360 22952 23424
rect 23016 23360 23032 23424
rect 23096 23360 23112 23424
rect 23176 23360 23192 23424
rect 23256 23360 23264 23424
rect 22507 22948 22573 22949
rect 22507 22884 22508 22948
rect 22572 22884 22573 22948
rect 22507 22883 22573 22884
rect 22510 2957 22570 22883
rect 22944 22336 23264 23360
rect 22944 22272 22952 22336
rect 23016 22272 23032 22336
rect 23096 22272 23112 22336
rect 23176 22272 23192 22336
rect 23256 22272 23264 22336
rect 22944 21248 23264 22272
rect 22944 21184 22952 21248
rect 23016 21184 23032 21248
rect 23096 21184 23112 21248
rect 23176 21184 23192 21248
rect 23256 21184 23264 21248
rect 22944 20160 23264 21184
rect 22944 20096 22952 20160
rect 23016 20096 23032 20160
rect 23096 20096 23112 20160
rect 23176 20096 23192 20160
rect 23256 20096 23264 20160
rect 22944 19072 23264 20096
rect 22944 19008 22952 19072
rect 23016 19008 23032 19072
rect 23096 19008 23112 19072
rect 23176 19008 23192 19072
rect 23256 19008 23264 19072
rect 22691 18868 22757 18869
rect 22691 18804 22692 18868
rect 22756 18804 22757 18868
rect 22691 18803 22757 18804
rect 22507 2956 22573 2957
rect 22507 2892 22508 2956
rect 22572 2892 22573 2956
rect 22507 2891 22573 2892
rect 22139 2684 22205 2685
rect 22139 2620 22140 2684
rect 22204 2620 22205 2684
rect 22139 2619 22205 2620
rect 22694 2549 22754 18803
rect 22944 17984 23264 19008
rect 22944 17920 22952 17984
rect 23016 17920 23032 17984
rect 23096 17920 23112 17984
rect 23176 17920 23192 17984
rect 23256 17920 23264 17984
rect 22944 16896 23264 17920
rect 22944 16832 22952 16896
rect 23016 16832 23032 16896
rect 23096 16832 23112 16896
rect 23176 16832 23192 16896
rect 23256 16832 23264 16896
rect 22944 15808 23264 16832
rect 22944 15744 22952 15808
rect 23016 15744 23032 15808
rect 23096 15744 23112 15808
rect 23176 15744 23192 15808
rect 23256 15744 23264 15808
rect 22944 14720 23264 15744
rect 22944 14656 22952 14720
rect 23016 14656 23032 14720
rect 23096 14656 23112 14720
rect 23176 14656 23192 14720
rect 23256 14656 23264 14720
rect 22944 13632 23264 14656
rect 22944 13568 22952 13632
rect 23016 13568 23032 13632
rect 23096 13568 23112 13632
rect 23176 13568 23192 13632
rect 23256 13568 23264 13632
rect 22944 12544 23264 13568
rect 22944 12480 22952 12544
rect 23016 12480 23032 12544
rect 23096 12480 23112 12544
rect 23176 12480 23192 12544
rect 23256 12480 23264 12544
rect 22944 11456 23264 12480
rect 22944 11392 22952 11456
rect 23016 11392 23032 11456
rect 23096 11392 23112 11456
rect 23176 11392 23192 11456
rect 23256 11392 23264 11456
rect 22944 10368 23264 11392
rect 22944 10304 22952 10368
rect 23016 10304 23032 10368
rect 23096 10304 23112 10368
rect 23176 10304 23192 10368
rect 23256 10304 23264 10368
rect 22944 9280 23264 10304
rect 22944 9216 22952 9280
rect 23016 9216 23032 9280
rect 23096 9216 23112 9280
rect 23176 9216 23192 9280
rect 23256 9216 23264 9280
rect 22944 8192 23264 9216
rect 22944 8128 22952 8192
rect 23016 8128 23032 8192
rect 23096 8128 23112 8192
rect 23176 8128 23192 8192
rect 23256 8128 23264 8192
rect 22944 7104 23264 8128
rect 22944 7040 22952 7104
rect 23016 7040 23032 7104
rect 23096 7040 23112 7104
rect 23176 7040 23192 7104
rect 23256 7040 23264 7104
rect 22944 6016 23264 7040
rect 22944 5952 22952 6016
rect 23016 5952 23032 6016
rect 23096 5952 23112 6016
rect 23176 5952 23192 6016
rect 23256 5952 23264 6016
rect 22944 4928 23264 5952
rect 22944 4864 22952 4928
rect 23016 4864 23032 4928
rect 23096 4864 23112 4928
rect 23176 4864 23192 4928
rect 23256 4864 23264 4928
rect 22944 3840 23264 4864
rect 22944 3776 22952 3840
rect 23016 3776 23032 3840
rect 23096 3776 23112 3840
rect 23176 3776 23192 3840
rect 23256 3776 23264 3840
rect 22944 2752 23264 3776
rect 27110 3501 27170 27643
rect 27662 24173 27722 28187
rect 27944 27232 28264 28256
rect 30422 27301 30482 40019
rect 32944 39744 33264 40768
rect 32944 39680 32952 39744
rect 33016 39680 33032 39744
rect 33096 39680 33112 39744
rect 33176 39680 33192 39744
rect 33256 39680 33264 39744
rect 32944 38656 33264 39680
rect 32944 38592 32952 38656
rect 33016 38592 33032 38656
rect 33096 38592 33112 38656
rect 33176 38592 33192 38656
rect 33256 38592 33264 38656
rect 32944 37568 33264 38592
rect 37944 54432 38264 54448
rect 37944 54368 37952 54432
rect 38016 54368 38032 54432
rect 38096 54368 38112 54432
rect 38176 54368 38192 54432
rect 38256 54368 38264 54432
rect 37944 53344 38264 54368
rect 37944 53280 37952 53344
rect 38016 53280 38032 53344
rect 38096 53280 38112 53344
rect 38176 53280 38192 53344
rect 38256 53280 38264 53344
rect 37944 52256 38264 53280
rect 37944 52192 37952 52256
rect 38016 52192 38032 52256
rect 38096 52192 38112 52256
rect 38176 52192 38192 52256
rect 38256 52192 38264 52256
rect 37944 51168 38264 52192
rect 37944 51104 37952 51168
rect 38016 51104 38032 51168
rect 38096 51104 38112 51168
rect 38176 51104 38192 51168
rect 38256 51104 38264 51168
rect 37944 50080 38264 51104
rect 37944 50016 37952 50080
rect 38016 50016 38032 50080
rect 38096 50016 38112 50080
rect 38176 50016 38192 50080
rect 38256 50016 38264 50080
rect 37944 48992 38264 50016
rect 37944 48928 37952 48992
rect 38016 48928 38032 48992
rect 38096 48928 38112 48992
rect 38176 48928 38192 48992
rect 38256 48928 38264 48992
rect 37944 47904 38264 48928
rect 37944 47840 37952 47904
rect 38016 47840 38032 47904
rect 38096 47840 38112 47904
rect 38176 47840 38192 47904
rect 38256 47840 38264 47904
rect 37944 46816 38264 47840
rect 37944 46752 37952 46816
rect 38016 46752 38032 46816
rect 38096 46752 38112 46816
rect 38176 46752 38192 46816
rect 38256 46752 38264 46816
rect 37944 45728 38264 46752
rect 37944 45664 37952 45728
rect 38016 45664 38032 45728
rect 38096 45664 38112 45728
rect 38176 45664 38192 45728
rect 38256 45664 38264 45728
rect 37944 44640 38264 45664
rect 37944 44576 37952 44640
rect 38016 44576 38032 44640
rect 38096 44576 38112 44640
rect 38176 44576 38192 44640
rect 38256 44576 38264 44640
rect 37944 43552 38264 44576
rect 37944 43488 37952 43552
rect 38016 43488 38032 43552
rect 38096 43488 38112 43552
rect 38176 43488 38192 43552
rect 38256 43488 38264 43552
rect 37944 42464 38264 43488
rect 37944 42400 37952 42464
rect 38016 42400 38032 42464
rect 38096 42400 38112 42464
rect 38176 42400 38192 42464
rect 38256 42400 38264 42464
rect 37944 41376 38264 42400
rect 42944 53888 43264 54448
rect 42944 53824 42952 53888
rect 43016 53824 43032 53888
rect 43096 53824 43112 53888
rect 43176 53824 43192 53888
rect 43256 53824 43264 53888
rect 42944 52800 43264 53824
rect 42944 52736 42952 52800
rect 43016 52736 43032 52800
rect 43096 52736 43112 52800
rect 43176 52736 43192 52800
rect 43256 52736 43264 52800
rect 42944 51712 43264 52736
rect 42944 51648 42952 51712
rect 43016 51648 43032 51712
rect 43096 51648 43112 51712
rect 43176 51648 43192 51712
rect 43256 51648 43264 51712
rect 42944 50624 43264 51648
rect 42944 50560 42952 50624
rect 43016 50560 43032 50624
rect 43096 50560 43112 50624
rect 43176 50560 43192 50624
rect 43256 50560 43264 50624
rect 42944 49536 43264 50560
rect 42944 49472 42952 49536
rect 43016 49472 43032 49536
rect 43096 49472 43112 49536
rect 43176 49472 43192 49536
rect 43256 49472 43264 49536
rect 42944 48448 43264 49472
rect 42944 48384 42952 48448
rect 43016 48384 43032 48448
rect 43096 48384 43112 48448
rect 43176 48384 43192 48448
rect 43256 48384 43264 48448
rect 42944 47360 43264 48384
rect 42944 47296 42952 47360
rect 43016 47296 43032 47360
rect 43096 47296 43112 47360
rect 43176 47296 43192 47360
rect 43256 47296 43264 47360
rect 42944 46272 43264 47296
rect 42944 46208 42952 46272
rect 43016 46208 43032 46272
rect 43096 46208 43112 46272
rect 43176 46208 43192 46272
rect 43256 46208 43264 46272
rect 42944 45184 43264 46208
rect 42944 45120 42952 45184
rect 43016 45120 43032 45184
rect 43096 45120 43112 45184
rect 43176 45120 43192 45184
rect 43256 45120 43264 45184
rect 42944 44096 43264 45120
rect 42944 44032 42952 44096
rect 43016 44032 43032 44096
rect 43096 44032 43112 44096
rect 43176 44032 43192 44096
rect 43256 44032 43264 44096
rect 42944 43008 43264 44032
rect 42944 42944 42952 43008
rect 43016 42944 43032 43008
rect 43096 42944 43112 43008
rect 43176 42944 43192 43008
rect 43256 42944 43264 43008
rect 39987 42124 40053 42125
rect 39987 42060 39988 42124
rect 40052 42060 40053 42124
rect 39987 42059 40053 42060
rect 37944 41312 37952 41376
rect 38016 41312 38032 41376
rect 38096 41312 38112 41376
rect 38176 41312 38192 41376
rect 38256 41312 38264 41376
rect 37944 40288 38264 41312
rect 37944 40224 37952 40288
rect 38016 40224 38032 40288
rect 38096 40224 38112 40288
rect 38176 40224 38192 40288
rect 38256 40224 38264 40288
rect 37944 39200 38264 40224
rect 37944 39136 37952 39200
rect 38016 39136 38032 39200
rect 38096 39136 38112 39200
rect 38176 39136 38192 39200
rect 38256 39136 38264 39200
rect 37944 38112 38264 39136
rect 37944 38048 37952 38112
rect 38016 38048 38032 38112
rect 38096 38048 38112 38112
rect 38176 38048 38192 38112
rect 38256 38048 38264 38112
rect 37595 37772 37661 37773
rect 37595 37708 37596 37772
rect 37660 37708 37661 37772
rect 37595 37707 37661 37708
rect 32944 37504 32952 37568
rect 33016 37504 33032 37568
rect 33096 37504 33112 37568
rect 33176 37504 33192 37568
rect 33256 37504 33264 37568
rect 32944 36480 33264 37504
rect 32944 36416 32952 36480
rect 33016 36416 33032 36480
rect 33096 36416 33112 36480
rect 33176 36416 33192 36480
rect 33256 36416 33264 36480
rect 32944 35392 33264 36416
rect 32944 35328 32952 35392
rect 33016 35328 33032 35392
rect 33096 35328 33112 35392
rect 33176 35328 33192 35392
rect 33256 35328 33264 35392
rect 32944 34304 33264 35328
rect 32944 34240 32952 34304
rect 33016 34240 33032 34304
rect 33096 34240 33112 34304
rect 33176 34240 33192 34304
rect 33256 34240 33264 34304
rect 32944 33216 33264 34240
rect 32944 33152 32952 33216
rect 33016 33152 33032 33216
rect 33096 33152 33112 33216
rect 33176 33152 33192 33216
rect 33256 33152 33264 33216
rect 32944 32128 33264 33152
rect 32944 32064 32952 32128
rect 33016 32064 33032 32128
rect 33096 32064 33112 32128
rect 33176 32064 33192 32128
rect 33256 32064 33264 32128
rect 32944 31040 33264 32064
rect 37411 31924 37477 31925
rect 37411 31860 37412 31924
rect 37476 31860 37477 31924
rect 37411 31859 37477 31860
rect 32944 30976 32952 31040
rect 33016 30976 33032 31040
rect 33096 30976 33112 31040
rect 33176 30976 33192 31040
rect 33256 30976 33264 31040
rect 30787 30156 30853 30157
rect 30787 30092 30788 30156
rect 30852 30092 30853 30156
rect 30787 30091 30853 30092
rect 30419 27300 30485 27301
rect 30419 27236 30420 27300
rect 30484 27236 30485 27300
rect 30419 27235 30485 27236
rect 27944 27168 27952 27232
rect 28016 27168 28032 27232
rect 28096 27168 28112 27232
rect 28176 27168 28192 27232
rect 28256 27168 28264 27232
rect 27944 26144 28264 27168
rect 27944 26080 27952 26144
rect 28016 26080 28032 26144
rect 28096 26080 28112 26144
rect 28176 26080 28192 26144
rect 28256 26080 28264 26144
rect 27944 25056 28264 26080
rect 30419 25260 30485 25261
rect 30419 25196 30420 25260
rect 30484 25196 30485 25260
rect 30419 25195 30485 25196
rect 27944 24992 27952 25056
rect 28016 24992 28032 25056
rect 28096 24992 28112 25056
rect 28176 24992 28192 25056
rect 28256 24992 28264 25056
rect 27659 24172 27725 24173
rect 27659 24108 27660 24172
rect 27724 24108 27725 24172
rect 27659 24107 27725 24108
rect 27944 23968 28264 24992
rect 27944 23904 27952 23968
rect 28016 23904 28032 23968
rect 28096 23904 28112 23968
rect 28176 23904 28192 23968
rect 28256 23904 28264 23968
rect 27944 22880 28264 23904
rect 27944 22816 27952 22880
rect 28016 22816 28032 22880
rect 28096 22816 28112 22880
rect 28176 22816 28192 22880
rect 28256 22816 28264 22880
rect 27944 21792 28264 22816
rect 27944 21728 27952 21792
rect 28016 21728 28032 21792
rect 28096 21728 28112 21792
rect 28176 21728 28192 21792
rect 28256 21728 28264 21792
rect 27944 20704 28264 21728
rect 27944 20640 27952 20704
rect 28016 20640 28032 20704
rect 28096 20640 28112 20704
rect 28176 20640 28192 20704
rect 28256 20640 28264 20704
rect 27944 19616 28264 20640
rect 30422 20637 30482 25195
rect 30790 21997 30850 30091
rect 32944 29952 33264 30976
rect 32944 29888 32952 29952
rect 33016 29888 33032 29952
rect 33096 29888 33112 29952
rect 33176 29888 33192 29952
rect 33256 29888 33264 29952
rect 32944 28864 33264 29888
rect 32944 28800 32952 28864
rect 33016 28800 33032 28864
rect 33096 28800 33112 28864
rect 33176 28800 33192 28864
rect 33256 28800 33264 28864
rect 32944 27776 33264 28800
rect 35203 28388 35269 28389
rect 35203 28324 35204 28388
rect 35268 28324 35269 28388
rect 35203 28323 35269 28324
rect 32944 27712 32952 27776
rect 33016 27712 33032 27776
rect 33096 27712 33112 27776
rect 33176 27712 33192 27776
rect 33256 27712 33264 27776
rect 30971 27028 31037 27029
rect 30971 26964 30972 27028
rect 31036 26964 31037 27028
rect 30971 26963 31037 26964
rect 30787 21996 30853 21997
rect 30787 21932 30788 21996
rect 30852 21932 30853 21996
rect 30787 21931 30853 21932
rect 30419 20636 30485 20637
rect 30419 20572 30420 20636
rect 30484 20572 30485 20636
rect 30419 20571 30485 20572
rect 27944 19552 27952 19616
rect 28016 19552 28032 19616
rect 28096 19552 28112 19616
rect 28176 19552 28192 19616
rect 28256 19552 28264 19616
rect 27944 18528 28264 19552
rect 27944 18464 27952 18528
rect 28016 18464 28032 18528
rect 28096 18464 28112 18528
rect 28176 18464 28192 18528
rect 28256 18464 28264 18528
rect 27944 17440 28264 18464
rect 30974 18053 31034 26963
rect 32944 26688 33264 27712
rect 32944 26624 32952 26688
rect 33016 26624 33032 26688
rect 33096 26624 33112 26688
rect 33176 26624 33192 26688
rect 33256 26624 33264 26688
rect 32627 26348 32693 26349
rect 32627 26284 32628 26348
rect 32692 26284 32693 26348
rect 32627 26283 32693 26284
rect 30971 18052 31037 18053
rect 30971 17988 30972 18052
rect 31036 17988 31037 18052
rect 30971 17987 31037 17988
rect 27944 17376 27952 17440
rect 28016 17376 28032 17440
rect 28096 17376 28112 17440
rect 28176 17376 28192 17440
rect 28256 17376 28264 17440
rect 27944 16352 28264 17376
rect 32630 16693 32690 26283
rect 32944 25600 33264 26624
rect 32944 25536 32952 25600
rect 33016 25536 33032 25600
rect 33096 25536 33112 25600
rect 33176 25536 33192 25600
rect 33256 25536 33264 25600
rect 32944 24512 33264 25536
rect 32944 24448 32952 24512
rect 33016 24448 33032 24512
rect 33096 24448 33112 24512
rect 33176 24448 33192 24512
rect 33256 24448 33264 24512
rect 32944 23424 33264 24448
rect 32944 23360 32952 23424
rect 33016 23360 33032 23424
rect 33096 23360 33112 23424
rect 33176 23360 33192 23424
rect 33256 23360 33264 23424
rect 32944 22336 33264 23360
rect 32944 22272 32952 22336
rect 33016 22272 33032 22336
rect 33096 22272 33112 22336
rect 33176 22272 33192 22336
rect 33256 22272 33264 22336
rect 32944 21248 33264 22272
rect 32944 21184 32952 21248
rect 33016 21184 33032 21248
rect 33096 21184 33112 21248
rect 33176 21184 33192 21248
rect 33256 21184 33264 21248
rect 32944 20160 33264 21184
rect 35206 20637 35266 28323
rect 37414 27029 37474 31859
rect 37598 29069 37658 37707
rect 37944 37024 38264 38048
rect 37944 36960 37952 37024
rect 38016 36960 38032 37024
rect 38096 36960 38112 37024
rect 38176 36960 38192 37024
rect 38256 36960 38264 37024
rect 37779 36820 37845 36821
rect 37779 36756 37780 36820
rect 37844 36756 37845 36820
rect 37779 36755 37845 36756
rect 37782 36141 37842 36755
rect 37779 36140 37845 36141
rect 37779 36076 37780 36140
rect 37844 36076 37845 36140
rect 37779 36075 37845 36076
rect 37782 30293 37842 36075
rect 37944 35936 38264 36960
rect 37944 35872 37952 35936
rect 38016 35872 38032 35936
rect 38096 35872 38112 35936
rect 38176 35872 38192 35936
rect 38256 35872 38264 35936
rect 37944 34848 38264 35872
rect 38883 34916 38949 34917
rect 38883 34852 38884 34916
rect 38948 34852 38949 34916
rect 38883 34851 38949 34852
rect 37944 34784 37952 34848
rect 38016 34784 38032 34848
rect 38096 34784 38112 34848
rect 38176 34784 38192 34848
rect 38256 34784 38264 34848
rect 37944 33760 38264 34784
rect 37944 33696 37952 33760
rect 38016 33696 38032 33760
rect 38096 33696 38112 33760
rect 38176 33696 38192 33760
rect 38256 33696 38264 33760
rect 37944 32672 38264 33696
rect 38886 33557 38946 34851
rect 38883 33556 38949 33557
rect 38883 33492 38884 33556
rect 38948 33492 38949 33556
rect 38883 33491 38949 33492
rect 37944 32608 37952 32672
rect 38016 32608 38032 32672
rect 38096 32608 38112 32672
rect 38176 32608 38192 32672
rect 38256 32608 38264 32672
rect 37944 31584 38264 32608
rect 37944 31520 37952 31584
rect 38016 31520 38032 31584
rect 38096 31520 38112 31584
rect 38176 31520 38192 31584
rect 38256 31520 38264 31584
rect 37944 30496 38264 31520
rect 37944 30432 37952 30496
rect 38016 30432 38032 30496
rect 38096 30432 38112 30496
rect 38176 30432 38192 30496
rect 38256 30432 38264 30496
rect 37779 30292 37845 30293
rect 37779 30228 37780 30292
rect 37844 30228 37845 30292
rect 37779 30227 37845 30228
rect 37944 29408 38264 30432
rect 37944 29344 37952 29408
rect 38016 29344 38032 29408
rect 38096 29344 38112 29408
rect 38176 29344 38192 29408
rect 38256 29344 38264 29408
rect 37595 29068 37661 29069
rect 37595 29004 37596 29068
rect 37660 29004 37661 29068
rect 37595 29003 37661 29004
rect 37944 28320 38264 29344
rect 37944 28256 37952 28320
rect 38016 28256 38032 28320
rect 38096 28256 38112 28320
rect 38176 28256 38192 28320
rect 38256 28256 38264 28320
rect 37944 27232 38264 28256
rect 37944 27168 37952 27232
rect 38016 27168 38032 27232
rect 38096 27168 38112 27232
rect 38176 27168 38192 27232
rect 38256 27168 38264 27232
rect 37411 27028 37477 27029
rect 37411 26964 37412 27028
rect 37476 26964 37477 27028
rect 37411 26963 37477 26964
rect 37944 26144 38264 27168
rect 38515 27028 38581 27029
rect 38515 26964 38516 27028
rect 38580 26964 38581 27028
rect 38515 26963 38581 26964
rect 37944 26080 37952 26144
rect 38016 26080 38032 26144
rect 38096 26080 38112 26144
rect 38176 26080 38192 26144
rect 38256 26080 38264 26144
rect 37944 25056 38264 26080
rect 37944 24992 37952 25056
rect 38016 24992 38032 25056
rect 38096 24992 38112 25056
rect 38176 24992 38192 25056
rect 38256 24992 38264 25056
rect 37944 23968 38264 24992
rect 37944 23904 37952 23968
rect 38016 23904 38032 23968
rect 38096 23904 38112 23968
rect 38176 23904 38192 23968
rect 38256 23904 38264 23968
rect 37944 22880 38264 23904
rect 37944 22816 37952 22880
rect 38016 22816 38032 22880
rect 38096 22816 38112 22880
rect 38176 22816 38192 22880
rect 38256 22816 38264 22880
rect 37944 21792 38264 22816
rect 37944 21728 37952 21792
rect 38016 21728 38032 21792
rect 38096 21728 38112 21792
rect 38176 21728 38192 21792
rect 38256 21728 38264 21792
rect 37944 20704 38264 21728
rect 37944 20640 37952 20704
rect 38016 20640 38032 20704
rect 38096 20640 38112 20704
rect 38176 20640 38192 20704
rect 38256 20640 38264 20704
rect 35203 20636 35269 20637
rect 35203 20572 35204 20636
rect 35268 20572 35269 20636
rect 35203 20571 35269 20572
rect 32944 20096 32952 20160
rect 33016 20096 33032 20160
rect 33096 20096 33112 20160
rect 33176 20096 33192 20160
rect 33256 20096 33264 20160
rect 32811 19276 32877 19277
rect 32811 19212 32812 19276
rect 32876 19212 32877 19276
rect 32811 19211 32877 19212
rect 32814 17373 32874 19211
rect 32944 19072 33264 20096
rect 32944 19008 32952 19072
rect 33016 19008 33032 19072
rect 33096 19008 33112 19072
rect 33176 19008 33192 19072
rect 33256 19008 33264 19072
rect 32944 17984 33264 19008
rect 32944 17920 32952 17984
rect 33016 17920 33032 17984
rect 33096 17920 33112 17984
rect 33176 17920 33192 17984
rect 33256 17920 33264 17984
rect 32811 17372 32877 17373
rect 32811 17308 32812 17372
rect 32876 17308 32877 17372
rect 32811 17307 32877 17308
rect 32944 16896 33264 17920
rect 32944 16832 32952 16896
rect 33016 16832 33032 16896
rect 33096 16832 33112 16896
rect 33176 16832 33192 16896
rect 33256 16832 33264 16896
rect 32627 16692 32693 16693
rect 32627 16628 32628 16692
rect 32692 16628 32693 16692
rect 32627 16627 32693 16628
rect 27944 16288 27952 16352
rect 28016 16288 28032 16352
rect 28096 16288 28112 16352
rect 28176 16288 28192 16352
rect 28256 16288 28264 16352
rect 27944 15264 28264 16288
rect 27944 15200 27952 15264
rect 28016 15200 28032 15264
rect 28096 15200 28112 15264
rect 28176 15200 28192 15264
rect 28256 15200 28264 15264
rect 27944 14176 28264 15200
rect 27944 14112 27952 14176
rect 28016 14112 28032 14176
rect 28096 14112 28112 14176
rect 28176 14112 28192 14176
rect 28256 14112 28264 14176
rect 27944 13088 28264 14112
rect 27944 13024 27952 13088
rect 28016 13024 28032 13088
rect 28096 13024 28112 13088
rect 28176 13024 28192 13088
rect 28256 13024 28264 13088
rect 27944 12000 28264 13024
rect 27944 11936 27952 12000
rect 28016 11936 28032 12000
rect 28096 11936 28112 12000
rect 28176 11936 28192 12000
rect 28256 11936 28264 12000
rect 27944 10912 28264 11936
rect 27944 10848 27952 10912
rect 28016 10848 28032 10912
rect 28096 10848 28112 10912
rect 28176 10848 28192 10912
rect 28256 10848 28264 10912
rect 27944 9824 28264 10848
rect 27944 9760 27952 9824
rect 28016 9760 28032 9824
rect 28096 9760 28112 9824
rect 28176 9760 28192 9824
rect 28256 9760 28264 9824
rect 27944 8736 28264 9760
rect 27944 8672 27952 8736
rect 28016 8672 28032 8736
rect 28096 8672 28112 8736
rect 28176 8672 28192 8736
rect 28256 8672 28264 8736
rect 27944 7648 28264 8672
rect 27944 7584 27952 7648
rect 28016 7584 28032 7648
rect 28096 7584 28112 7648
rect 28176 7584 28192 7648
rect 28256 7584 28264 7648
rect 27944 6560 28264 7584
rect 27944 6496 27952 6560
rect 28016 6496 28032 6560
rect 28096 6496 28112 6560
rect 28176 6496 28192 6560
rect 28256 6496 28264 6560
rect 27944 5472 28264 6496
rect 27944 5408 27952 5472
rect 28016 5408 28032 5472
rect 28096 5408 28112 5472
rect 28176 5408 28192 5472
rect 28256 5408 28264 5472
rect 27944 4384 28264 5408
rect 27944 4320 27952 4384
rect 28016 4320 28032 4384
rect 28096 4320 28112 4384
rect 28176 4320 28192 4384
rect 28256 4320 28264 4384
rect 27107 3500 27173 3501
rect 27107 3436 27108 3500
rect 27172 3436 27173 3500
rect 27107 3435 27173 3436
rect 22944 2688 22952 2752
rect 23016 2688 23032 2752
rect 23096 2688 23112 2752
rect 23176 2688 23192 2752
rect 23256 2688 23264 2752
rect 22691 2548 22757 2549
rect 22691 2484 22692 2548
rect 22756 2484 22757 2548
rect 22691 2483 22757 2484
rect 17944 2144 17952 2208
rect 18016 2144 18032 2208
rect 18096 2144 18112 2208
rect 18176 2144 18192 2208
rect 18256 2144 18264 2208
rect 17944 2128 18264 2144
rect 22944 2128 23264 2688
rect 27944 3296 28264 4320
rect 27944 3232 27952 3296
rect 28016 3232 28032 3296
rect 28096 3232 28112 3296
rect 28176 3232 28192 3296
rect 28256 3232 28264 3296
rect 27944 2208 28264 3232
rect 27944 2144 27952 2208
rect 28016 2144 28032 2208
rect 28096 2144 28112 2208
rect 28176 2144 28192 2208
rect 28256 2144 28264 2208
rect 27944 2128 28264 2144
rect 32944 15808 33264 16832
rect 32944 15744 32952 15808
rect 33016 15744 33032 15808
rect 33096 15744 33112 15808
rect 33176 15744 33192 15808
rect 33256 15744 33264 15808
rect 32944 14720 33264 15744
rect 32944 14656 32952 14720
rect 33016 14656 33032 14720
rect 33096 14656 33112 14720
rect 33176 14656 33192 14720
rect 33256 14656 33264 14720
rect 32944 13632 33264 14656
rect 32944 13568 32952 13632
rect 33016 13568 33032 13632
rect 33096 13568 33112 13632
rect 33176 13568 33192 13632
rect 33256 13568 33264 13632
rect 32944 12544 33264 13568
rect 32944 12480 32952 12544
rect 33016 12480 33032 12544
rect 33096 12480 33112 12544
rect 33176 12480 33192 12544
rect 33256 12480 33264 12544
rect 32944 11456 33264 12480
rect 32944 11392 32952 11456
rect 33016 11392 33032 11456
rect 33096 11392 33112 11456
rect 33176 11392 33192 11456
rect 33256 11392 33264 11456
rect 32944 10368 33264 11392
rect 32944 10304 32952 10368
rect 33016 10304 33032 10368
rect 33096 10304 33112 10368
rect 33176 10304 33192 10368
rect 33256 10304 33264 10368
rect 32944 9280 33264 10304
rect 32944 9216 32952 9280
rect 33016 9216 33032 9280
rect 33096 9216 33112 9280
rect 33176 9216 33192 9280
rect 33256 9216 33264 9280
rect 32944 8192 33264 9216
rect 32944 8128 32952 8192
rect 33016 8128 33032 8192
rect 33096 8128 33112 8192
rect 33176 8128 33192 8192
rect 33256 8128 33264 8192
rect 32944 7104 33264 8128
rect 32944 7040 32952 7104
rect 33016 7040 33032 7104
rect 33096 7040 33112 7104
rect 33176 7040 33192 7104
rect 33256 7040 33264 7104
rect 32944 6016 33264 7040
rect 32944 5952 32952 6016
rect 33016 5952 33032 6016
rect 33096 5952 33112 6016
rect 33176 5952 33192 6016
rect 33256 5952 33264 6016
rect 32944 4928 33264 5952
rect 32944 4864 32952 4928
rect 33016 4864 33032 4928
rect 33096 4864 33112 4928
rect 33176 4864 33192 4928
rect 33256 4864 33264 4928
rect 32944 3840 33264 4864
rect 32944 3776 32952 3840
rect 33016 3776 33032 3840
rect 33096 3776 33112 3840
rect 33176 3776 33192 3840
rect 33256 3776 33264 3840
rect 32944 2752 33264 3776
rect 32944 2688 32952 2752
rect 33016 2688 33032 2752
rect 33096 2688 33112 2752
rect 33176 2688 33192 2752
rect 33256 2688 33264 2752
rect 32944 2128 33264 2688
rect 37944 19616 38264 20640
rect 37944 19552 37952 19616
rect 38016 19552 38032 19616
rect 38096 19552 38112 19616
rect 38176 19552 38192 19616
rect 38256 19552 38264 19616
rect 37944 18528 38264 19552
rect 38518 19277 38578 26963
rect 39990 26349 40050 42059
rect 42944 41920 43264 42944
rect 42944 41856 42952 41920
rect 43016 41856 43032 41920
rect 43096 41856 43112 41920
rect 43176 41856 43192 41920
rect 43256 41856 43264 41920
rect 40539 41716 40605 41717
rect 40539 41652 40540 41716
rect 40604 41652 40605 41716
rect 40539 41651 40605 41652
rect 40542 28525 40602 41651
rect 42944 40832 43264 41856
rect 42944 40768 42952 40832
rect 43016 40768 43032 40832
rect 43096 40768 43112 40832
rect 43176 40768 43192 40832
rect 43256 40768 43264 40832
rect 41275 40628 41341 40629
rect 41275 40564 41276 40628
rect 41340 40564 41341 40628
rect 41275 40563 41341 40564
rect 41278 35869 41338 40563
rect 42944 39744 43264 40768
rect 42944 39680 42952 39744
rect 43016 39680 43032 39744
rect 43096 39680 43112 39744
rect 43176 39680 43192 39744
rect 43256 39680 43264 39744
rect 42944 38656 43264 39680
rect 42944 38592 42952 38656
rect 43016 38592 43032 38656
rect 43096 38592 43112 38656
rect 43176 38592 43192 38656
rect 43256 38592 43264 38656
rect 42944 37568 43264 38592
rect 42944 37504 42952 37568
rect 43016 37504 43032 37568
rect 43096 37504 43112 37568
rect 43176 37504 43192 37568
rect 43256 37504 43264 37568
rect 42944 36480 43264 37504
rect 42944 36416 42952 36480
rect 43016 36416 43032 36480
rect 43096 36416 43112 36480
rect 43176 36416 43192 36480
rect 43256 36416 43264 36480
rect 41275 35868 41341 35869
rect 41275 35804 41276 35868
rect 41340 35804 41341 35868
rect 41275 35803 41341 35804
rect 42944 35392 43264 36416
rect 42944 35328 42952 35392
rect 43016 35328 43032 35392
rect 43096 35328 43112 35392
rect 43176 35328 43192 35392
rect 43256 35328 43264 35392
rect 42944 34304 43264 35328
rect 42944 34240 42952 34304
rect 43016 34240 43032 34304
rect 43096 34240 43112 34304
rect 43176 34240 43192 34304
rect 43256 34240 43264 34304
rect 42944 33216 43264 34240
rect 42944 33152 42952 33216
rect 43016 33152 43032 33216
rect 43096 33152 43112 33216
rect 43176 33152 43192 33216
rect 43256 33152 43264 33216
rect 42944 32128 43264 33152
rect 42944 32064 42952 32128
rect 43016 32064 43032 32128
rect 43096 32064 43112 32128
rect 43176 32064 43192 32128
rect 43256 32064 43264 32128
rect 42944 31040 43264 32064
rect 42944 30976 42952 31040
rect 43016 30976 43032 31040
rect 43096 30976 43112 31040
rect 43176 30976 43192 31040
rect 43256 30976 43264 31040
rect 42944 29952 43264 30976
rect 42944 29888 42952 29952
rect 43016 29888 43032 29952
rect 43096 29888 43112 29952
rect 43176 29888 43192 29952
rect 43256 29888 43264 29952
rect 42944 28864 43264 29888
rect 42944 28800 42952 28864
rect 43016 28800 43032 28864
rect 43096 28800 43112 28864
rect 43176 28800 43192 28864
rect 43256 28800 43264 28864
rect 40539 28524 40605 28525
rect 40539 28460 40540 28524
rect 40604 28460 40605 28524
rect 40539 28459 40605 28460
rect 42944 27776 43264 28800
rect 42944 27712 42952 27776
rect 43016 27712 43032 27776
rect 43096 27712 43112 27776
rect 43176 27712 43192 27776
rect 43256 27712 43264 27776
rect 42944 26688 43264 27712
rect 42944 26624 42952 26688
rect 43016 26624 43032 26688
rect 43096 26624 43112 26688
rect 43176 26624 43192 26688
rect 43256 26624 43264 26688
rect 39987 26348 40053 26349
rect 39987 26284 39988 26348
rect 40052 26284 40053 26348
rect 39987 26283 40053 26284
rect 42944 25600 43264 26624
rect 42944 25536 42952 25600
rect 43016 25536 43032 25600
rect 43096 25536 43112 25600
rect 43176 25536 43192 25600
rect 43256 25536 43264 25600
rect 42944 24512 43264 25536
rect 42944 24448 42952 24512
rect 43016 24448 43032 24512
rect 43096 24448 43112 24512
rect 43176 24448 43192 24512
rect 43256 24448 43264 24512
rect 42944 23424 43264 24448
rect 42944 23360 42952 23424
rect 43016 23360 43032 23424
rect 43096 23360 43112 23424
rect 43176 23360 43192 23424
rect 43256 23360 43264 23424
rect 42944 22336 43264 23360
rect 42944 22272 42952 22336
rect 43016 22272 43032 22336
rect 43096 22272 43112 22336
rect 43176 22272 43192 22336
rect 43256 22272 43264 22336
rect 42944 21248 43264 22272
rect 42944 21184 42952 21248
rect 43016 21184 43032 21248
rect 43096 21184 43112 21248
rect 43176 21184 43192 21248
rect 43256 21184 43264 21248
rect 42944 20160 43264 21184
rect 42944 20096 42952 20160
rect 43016 20096 43032 20160
rect 43096 20096 43112 20160
rect 43176 20096 43192 20160
rect 43256 20096 43264 20160
rect 38515 19276 38581 19277
rect 38515 19212 38516 19276
rect 38580 19212 38581 19276
rect 38515 19211 38581 19212
rect 37944 18464 37952 18528
rect 38016 18464 38032 18528
rect 38096 18464 38112 18528
rect 38176 18464 38192 18528
rect 38256 18464 38264 18528
rect 37944 17440 38264 18464
rect 37944 17376 37952 17440
rect 38016 17376 38032 17440
rect 38096 17376 38112 17440
rect 38176 17376 38192 17440
rect 38256 17376 38264 17440
rect 37944 16352 38264 17376
rect 37944 16288 37952 16352
rect 38016 16288 38032 16352
rect 38096 16288 38112 16352
rect 38176 16288 38192 16352
rect 38256 16288 38264 16352
rect 37944 15264 38264 16288
rect 37944 15200 37952 15264
rect 38016 15200 38032 15264
rect 38096 15200 38112 15264
rect 38176 15200 38192 15264
rect 38256 15200 38264 15264
rect 37944 14176 38264 15200
rect 37944 14112 37952 14176
rect 38016 14112 38032 14176
rect 38096 14112 38112 14176
rect 38176 14112 38192 14176
rect 38256 14112 38264 14176
rect 37944 13088 38264 14112
rect 37944 13024 37952 13088
rect 38016 13024 38032 13088
rect 38096 13024 38112 13088
rect 38176 13024 38192 13088
rect 38256 13024 38264 13088
rect 37944 12000 38264 13024
rect 38518 12341 38578 19211
rect 42944 19072 43264 20096
rect 42944 19008 42952 19072
rect 43016 19008 43032 19072
rect 43096 19008 43112 19072
rect 43176 19008 43192 19072
rect 43256 19008 43264 19072
rect 42944 17984 43264 19008
rect 42944 17920 42952 17984
rect 43016 17920 43032 17984
rect 43096 17920 43112 17984
rect 43176 17920 43192 17984
rect 43256 17920 43264 17984
rect 42944 16896 43264 17920
rect 42944 16832 42952 16896
rect 43016 16832 43032 16896
rect 43096 16832 43112 16896
rect 43176 16832 43192 16896
rect 43256 16832 43264 16896
rect 42944 15808 43264 16832
rect 42944 15744 42952 15808
rect 43016 15744 43032 15808
rect 43096 15744 43112 15808
rect 43176 15744 43192 15808
rect 43256 15744 43264 15808
rect 42944 14720 43264 15744
rect 42944 14656 42952 14720
rect 43016 14656 43032 14720
rect 43096 14656 43112 14720
rect 43176 14656 43192 14720
rect 43256 14656 43264 14720
rect 42944 13632 43264 14656
rect 42944 13568 42952 13632
rect 43016 13568 43032 13632
rect 43096 13568 43112 13632
rect 43176 13568 43192 13632
rect 43256 13568 43264 13632
rect 42944 12544 43264 13568
rect 42944 12480 42952 12544
rect 43016 12480 43032 12544
rect 43096 12480 43112 12544
rect 43176 12480 43192 12544
rect 43256 12480 43264 12544
rect 38515 12340 38581 12341
rect 38515 12276 38516 12340
rect 38580 12276 38581 12340
rect 38515 12275 38581 12276
rect 37944 11936 37952 12000
rect 38016 11936 38032 12000
rect 38096 11936 38112 12000
rect 38176 11936 38192 12000
rect 38256 11936 38264 12000
rect 37944 10912 38264 11936
rect 37944 10848 37952 10912
rect 38016 10848 38032 10912
rect 38096 10848 38112 10912
rect 38176 10848 38192 10912
rect 38256 10848 38264 10912
rect 37944 9824 38264 10848
rect 37944 9760 37952 9824
rect 38016 9760 38032 9824
rect 38096 9760 38112 9824
rect 38176 9760 38192 9824
rect 38256 9760 38264 9824
rect 37944 8736 38264 9760
rect 37944 8672 37952 8736
rect 38016 8672 38032 8736
rect 38096 8672 38112 8736
rect 38176 8672 38192 8736
rect 38256 8672 38264 8736
rect 37944 7648 38264 8672
rect 37944 7584 37952 7648
rect 38016 7584 38032 7648
rect 38096 7584 38112 7648
rect 38176 7584 38192 7648
rect 38256 7584 38264 7648
rect 37944 6560 38264 7584
rect 37944 6496 37952 6560
rect 38016 6496 38032 6560
rect 38096 6496 38112 6560
rect 38176 6496 38192 6560
rect 38256 6496 38264 6560
rect 37944 5472 38264 6496
rect 37944 5408 37952 5472
rect 38016 5408 38032 5472
rect 38096 5408 38112 5472
rect 38176 5408 38192 5472
rect 38256 5408 38264 5472
rect 37944 4384 38264 5408
rect 37944 4320 37952 4384
rect 38016 4320 38032 4384
rect 38096 4320 38112 4384
rect 38176 4320 38192 4384
rect 38256 4320 38264 4384
rect 37944 3296 38264 4320
rect 37944 3232 37952 3296
rect 38016 3232 38032 3296
rect 38096 3232 38112 3296
rect 38176 3232 38192 3296
rect 38256 3232 38264 3296
rect 37944 2208 38264 3232
rect 37944 2144 37952 2208
rect 38016 2144 38032 2208
rect 38096 2144 38112 2208
rect 38176 2144 38192 2208
rect 38256 2144 38264 2208
rect 37944 2128 38264 2144
rect 42944 11456 43264 12480
rect 42944 11392 42952 11456
rect 43016 11392 43032 11456
rect 43096 11392 43112 11456
rect 43176 11392 43192 11456
rect 43256 11392 43264 11456
rect 42944 10368 43264 11392
rect 42944 10304 42952 10368
rect 43016 10304 43032 10368
rect 43096 10304 43112 10368
rect 43176 10304 43192 10368
rect 43256 10304 43264 10368
rect 42944 9280 43264 10304
rect 42944 9216 42952 9280
rect 43016 9216 43032 9280
rect 43096 9216 43112 9280
rect 43176 9216 43192 9280
rect 43256 9216 43264 9280
rect 42944 8192 43264 9216
rect 42944 8128 42952 8192
rect 43016 8128 43032 8192
rect 43096 8128 43112 8192
rect 43176 8128 43192 8192
rect 43256 8128 43264 8192
rect 42944 7104 43264 8128
rect 42944 7040 42952 7104
rect 43016 7040 43032 7104
rect 43096 7040 43112 7104
rect 43176 7040 43192 7104
rect 43256 7040 43264 7104
rect 42944 6016 43264 7040
rect 42944 5952 42952 6016
rect 43016 5952 43032 6016
rect 43096 5952 43112 6016
rect 43176 5952 43192 6016
rect 43256 5952 43264 6016
rect 42944 4928 43264 5952
rect 42944 4864 42952 4928
rect 43016 4864 43032 4928
rect 43096 4864 43112 4928
rect 43176 4864 43192 4928
rect 43256 4864 43264 4928
rect 42944 3840 43264 4864
rect 42944 3776 42952 3840
rect 43016 3776 43032 3840
rect 43096 3776 43112 3840
rect 43176 3776 43192 3840
rect 43256 3776 43264 3840
rect 42944 2752 43264 3776
rect 42944 2688 42952 2752
rect 43016 2688 43032 2752
rect 43096 2688 43112 2752
rect 43176 2688 43192 2752
rect 43256 2688 43264 2752
rect 42944 2128 43264 2688
rect 47944 54432 48264 54448
rect 47944 54368 47952 54432
rect 48016 54368 48032 54432
rect 48096 54368 48112 54432
rect 48176 54368 48192 54432
rect 48256 54368 48264 54432
rect 47944 53344 48264 54368
rect 47944 53280 47952 53344
rect 48016 53280 48032 53344
rect 48096 53280 48112 53344
rect 48176 53280 48192 53344
rect 48256 53280 48264 53344
rect 47944 52256 48264 53280
rect 47944 52192 47952 52256
rect 48016 52192 48032 52256
rect 48096 52192 48112 52256
rect 48176 52192 48192 52256
rect 48256 52192 48264 52256
rect 47944 51168 48264 52192
rect 47944 51104 47952 51168
rect 48016 51104 48032 51168
rect 48096 51104 48112 51168
rect 48176 51104 48192 51168
rect 48256 51104 48264 51168
rect 47944 50080 48264 51104
rect 47944 50016 47952 50080
rect 48016 50016 48032 50080
rect 48096 50016 48112 50080
rect 48176 50016 48192 50080
rect 48256 50016 48264 50080
rect 47944 48992 48264 50016
rect 47944 48928 47952 48992
rect 48016 48928 48032 48992
rect 48096 48928 48112 48992
rect 48176 48928 48192 48992
rect 48256 48928 48264 48992
rect 47944 47904 48264 48928
rect 47944 47840 47952 47904
rect 48016 47840 48032 47904
rect 48096 47840 48112 47904
rect 48176 47840 48192 47904
rect 48256 47840 48264 47904
rect 47944 46816 48264 47840
rect 47944 46752 47952 46816
rect 48016 46752 48032 46816
rect 48096 46752 48112 46816
rect 48176 46752 48192 46816
rect 48256 46752 48264 46816
rect 47944 45728 48264 46752
rect 47944 45664 47952 45728
rect 48016 45664 48032 45728
rect 48096 45664 48112 45728
rect 48176 45664 48192 45728
rect 48256 45664 48264 45728
rect 47944 44640 48264 45664
rect 47944 44576 47952 44640
rect 48016 44576 48032 44640
rect 48096 44576 48112 44640
rect 48176 44576 48192 44640
rect 48256 44576 48264 44640
rect 47944 43552 48264 44576
rect 47944 43488 47952 43552
rect 48016 43488 48032 43552
rect 48096 43488 48112 43552
rect 48176 43488 48192 43552
rect 48256 43488 48264 43552
rect 47944 42464 48264 43488
rect 47944 42400 47952 42464
rect 48016 42400 48032 42464
rect 48096 42400 48112 42464
rect 48176 42400 48192 42464
rect 48256 42400 48264 42464
rect 47944 41376 48264 42400
rect 47944 41312 47952 41376
rect 48016 41312 48032 41376
rect 48096 41312 48112 41376
rect 48176 41312 48192 41376
rect 48256 41312 48264 41376
rect 47944 40288 48264 41312
rect 47944 40224 47952 40288
rect 48016 40224 48032 40288
rect 48096 40224 48112 40288
rect 48176 40224 48192 40288
rect 48256 40224 48264 40288
rect 47944 39200 48264 40224
rect 47944 39136 47952 39200
rect 48016 39136 48032 39200
rect 48096 39136 48112 39200
rect 48176 39136 48192 39200
rect 48256 39136 48264 39200
rect 47944 38112 48264 39136
rect 47944 38048 47952 38112
rect 48016 38048 48032 38112
rect 48096 38048 48112 38112
rect 48176 38048 48192 38112
rect 48256 38048 48264 38112
rect 47944 37024 48264 38048
rect 47944 36960 47952 37024
rect 48016 36960 48032 37024
rect 48096 36960 48112 37024
rect 48176 36960 48192 37024
rect 48256 36960 48264 37024
rect 47944 35936 48264 36960
rect 47944 35872 47952 35936
rect 48016 35872 48032 35936
rect 48096 35872 48112 35936
rect 48176 35872 48192 35936
rect 48256 35872 48264 35936
rect 47944 34848 48264 35872
rect 47944 34784 47952 34848
rect 48016 34784 48032 34848
rect 48096 34784 48112 34848
rect 48176 34784 48192 34848
rect 48256 34784 48264 34848
rect 47944 33760 48264 34784
rect 47944 33696 47952 33760
rect 48016 33696 48032 33760
rect 48096 33696 48112 33760
rect 48176 33696 48192 33760
rect 48256 33696 48264 33760
rect 47944 32672 48264 33696
rect 47944 32608 47952 32672
rect 48016 32608 48032 32672
rect 48096 32608 48112 32672
rect 48176 32608 48192 32672
rect 48256 32608 48264 32672
rect 47944 31584 48264 32608
rect 47944 31520 47952 31584
rect 48016 31520 48032 31584
rect 48096 31520 48112 31584
rect 48176 31520 48192 31584
rect 48256 31520 48264 31584
rect 47944 30496 48264 31520
rect 47944 30432 47952 30496
rect 48016 30432 48032 30496
rect 48096 30432 48112 30496
rect 48176 30432 48192 30496
rect 48256 30432 48264 30496
rect 47944 29408 48264 30432
rect 47944 29344 47952 29408
rect 48016 29344 48032 29408
rect 48096 29344 48112 29408
rect 48176 29344 48192 29408
rect 48256 29344 48264 29408
rect 47944 28320 48264 29344
rect 47944 28256 47952 28320
rect 48016 28256 48032 28320
rect 48096 28256 48112 28320
rect 48176 28256 48192 28320
rect 48256 28256 48264 28320
rect 47944 27232 48264 28256
rect 47944 27168 47952 27232
rect 48016 27168 48032 27232
rect 48096 27168 48112 27232
rect 48176 27168 48192 27232
rect 48256 27168 48264 27232
rect 47944 26144 48264 27168
rect 47944 26080 47952 26144
rect 48016 26080 48032 26144
rect 48096 26080 48112 26144
rect 48176 26080 48192 26144
rect 48256 26080 48264 26144
rect 47944 25056 48264 26080
rect 47944 24992 47952 25056
rect 48016 24992 48032 25056
rect 48096 24992 48112 25056
rect 48176 24992 48192 25056
rect 48256 24992 48264 25056
rect 47944 23968 48264 24992
rect 47944 23904 47952 23968
rect 48016 23904 48032 23968
rect 48096 23904 48112 23968
rect 48176 23904 48192 23968
rect 48256 23904 48264 23968
rect 47944 22880 48264 23904
rect 47944 22816 47952 22880
rect 48016 22816 48032 22880
rect 48096 22816 48112 22880
rect 48176 22816 48192 22880
rect 48256 22816 48264 22880
rect 47944 21792 48264 22816
rect 47944 21728 47952 21792
rect 48016 21728 48032 21792
rect 48096 21728 48112 21792
rect 48176 21728 48192 21792
rect 48256 21728 48264 21792
rect 47944 20704 48264 21728
rect 47944 20640 47952 20704
rect 48016 20640 48032 20704
rect 48096 20640 48112 20704
rect 48176 20640 48192 20704
rect 48256 20640 48264 20704
rect 47944 19616 48264 20640
rect 47944 19552 47952 19616
rect 48016 19552 48032 19616
rect 48096 19552 48112 19616
rect 48176 19552 48192 19616
rect 48256 19552 48264 19616
rect 47944 18528 48264 19552
rect 47944 18464 47952 18528
rect 48016 18464 48032 18528
rect 48096 18464 48112 18528
rect 48176 18464 48192 18528
rect 48256 18464 48264 18528
rect 47944 17440 48264 18464
rect 47944 17376 47952 17440
rect 48016 17376 48032 17440
rect 48096 17376 48112 17440
rect 48176 17376 48192 17440
rect 48256 17376 48264 17440
rect 47944 16352 48264 17376
rect 47944 16288 47952 16352
rect 48016 16288 48032 16352
rect 48096 16288 48112 16352
rect 48176 16288 48192 16352
rect 48256 16288 48264 16352
rect 47944 15264 48264 16288
rect 47944 15200 47952 15264
rect 48016 15200 48032 15264
rect 48096 15200 48112 15264
rect 48176 15200 48192 15264
rect 48256 15200 48264 15264
rect 47944 14176 48264 15200
rect 47944 14112 47952 14176
rect 48016 14112 48032 14176
rect 48096 14112 48112 14176
rect 48176 14112 48192 14176
rect 48256 14112 48264 14176
rect 47944 13088 48264 14112
rect 47944 13024 47952 13088
rect 48016 13024 48032 13088
rect 48096 13024 48112 13088
rect 48176 13024 48192 13088
rect 48256 13024 48264 13088
rect 47944 12000 48264 13024
rect 47944 11936 47952 12000
rect 48016 11936 48032 12000
rect 48096 11936 48112 12000
rect 48176 11936 48192 12000
rect 48256 11936 48264 12000
rect 47944 10912 48264 11936
rect 47944 10848 47952 10912
rect 48016 10848 48032 10912
rect 48096 10848 48112 10912
rect 48176 10848 48192 10912
rect 48256 10848 48264 10912
rect 47944 9824 48264 10848
rect 47944 9760 47952 9824
rect 48016 9760 48032 9824
rect 48096 9760 48112 9824
rect 48176 9760 48192 9824
rect 48256 9760 48264 9824
rect 47944 8736 48264 9760
rect 47944 8672 47952 8736
rect 48016 8672 48032 8736
rect 48096 8672 48112 8736
rect 48176 8672 48192 8736
rect 48256 8672 48264 8736
rect 47944 7648 48264 8672
rect 47944 7584 47952 7648
rect 48016 7584 48032 7648
rect 48096 7584 48112 7648
rect 48176 7584 48192 7648
rect 48256 7584 48264 7648
rect 47944 6560 48264 7584
rect 47944 6496 47952 6560
rect 48016 6496 48032 6560
rect 48096 6496 48112 6560
rect 48176 6496 48192 6560
rect 48256 6496 48264 6560
rect 47944 5472 48264 6496
rect 47944 5408 47952 5472
rect 48016 5408 48032 5472
rect 48096 5408 48112 5472
rect 48176 5408 48192 5472
rect 48256 5408 48264 5472
rect 47944 4384 48264 5408
rect 47944 4320 47952 4384
rect 48016 4320 48032 4384
rect 48096 4320 48112 4384
rect 48176 4320 48192 4384
rect 48256 4320 48264 4384
rect 47944 3296 48264 4320
rect 47944 3232 47952 3296
rect 48016 3232 48032 3296
rect 48096 3232 48112 3296
rect 48176 3232 48192 3296
rect 48256 3232 48264 3296
rect 47944 2208 48264 3232
rect 47944 2144 47952 2208
rect 48016 2144 48032 2208
rect 48096 2144 48112 2208
rect 48176 2144 48192 2208
rect 48256 2144 48264 2208
rect 47944 2128 48264 2144
use sky130_fd_sc_hd__clkbuf_2  _109_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 45908 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _110_
timestamp 1676037725
transform 1 0 45632 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _111_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 46092 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _112_
timestamp 1676037725
transform 1 0 46184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _113_
timestamp 1676037725
transform 1 0 46184 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _114_
timestamp 1676037725
transform 1 0 45448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _115_
timestamp 1676037725
transform 1 0 44712 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _116_
timestamp 1676037725
transform 1 0 29992 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1676037725
transform 1 0 44252 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _118_
timestamp 1676037725
transform 1 0 43608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _119_
timestamp 1676037725
transform 1 0 40480 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _120_
timestamp 1676037725
transform 1 0 42872 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _121_
timestamp 1676037725
transform 1 0 43608 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _122_
timestamp 1676037725
transform 1 0 43608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _123_
timestamp 1676037725
transform 1 0 44344 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1676037725
transform 1 0 44068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _125_
timestamp 1676037725
transform 1 0 43976 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _126_
timestamp 1676037725
transform 1 0 43700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _127_
timestamp 1676037725
transform 1 0 44068 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _128_
timestamp 1676037725
transform 1 0 44252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _129_
timestamp 1676037725
transform 1 0 45172 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _130_
timestamp 1676037725
transform 1 0 45908 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _131_
timestamp 1676037725
transform 1 0 46644 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _132_
timestamp 1676037725
transform 1 0 45908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _133_
timestamp 1676037725
transform 1 0 47104 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _134_
timestamp 1676037725
transform 1 0 47748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1676037725
transform 1 0 46828 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _136_
timestamp 1676037725
transform 1 0 48024 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1676037725
transform 1 0 47196 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _138_
timestamp 1676037725
transform 1 0 24564 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1676037725
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _140_
timestamp 1676037725
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _141_
timestamp 1676037725
transform 1 0 24380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _142_
timestamp 1676037725
transform 1 0 27140 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _143_
timestamp 1676037725
transform 1 0 27876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _144_
timestamp 1676037725
transform 1 0 28888 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _145_
timestamp 1676037725
transform 1 0 31740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _146_
timestamp 1676037725
transform 1 0 28704 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _147_
timestamp 1676037725
transform 1 0 28888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _148_
timestamp 1676037725
transform 1 0 29808 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _149_
timestamp 1676037725
transform 1 0 28612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _150_
timestamp 1676037725
transform 1 0 33028 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1676037725
transform 1 0 33764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _152_
timestamp 1676037725
transform 1 0 31464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _153_
timestamp 1676037725
transform 1 0 32292 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _154_
timestamp 1676037725
transform 1 0 34040 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _155_
timestamp 1676037725
transform 1 0 34868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _156_
timestamp 1676037725
transform 1 0 36156 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _157_
timestamp 1676037725
transform 1 0 37720 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _158_
timestamp 1676037725
transform 1 0 37076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _159_
timestamp 1676037725
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1676037725
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _161_
timestamp 1676037725
transform 1 0 35788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _162_
timestamp 1676037725
transform 1 0 35604 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _163_
timestamp 1676037725
transform 1 0 38824 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _164_
timestamp 1676037725
transform 1 0 36432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _165_
timestamp 1676037725
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _166_
timestamp 1676037725
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _167_
timestamp 1676037725
transform 1 0 37444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _168_
timestamp 1676037725
transform 1 0 5612 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _169_
timestamp 1676037725
transform 1 0 7084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _170_
timestamp 1676037725
transform 1 0 7820 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _171_
timestamp 1676037725
transform 1 0 12144 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _172_
timestamp 1676037725
transform 1 0 9016 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _173_
timestamp 1676037725
transform 1 0 9660 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _174_
timestamp 1676037725
transform 1 0 10580 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _175_
timestamp 1676037725
transform 1 0 12880 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _176_
timestamp 1676037725
transform 1 0 11960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _177_
timestamp 1676037725
transform 1 0 12144 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _178_
timestamp 1676037725
transform 1 0 13340 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _179_
timestamp 1676037725
transform 1 0 14260 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _180_
timestamp 1676037725
transform 1 0 14168 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _181_
timestamp 1676037725
transform 1 0 14812 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _182_
timestamp 1676037725
transform 1 0 16008 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _183_
timestamp 1676037725
transform 1 0 14536 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _184_
timestamp 1676037725
transform 1 0 16744 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _185_
timestamp 1676037725
transform 1 0 17112 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _186_
timestamp 1676037725
transform 1 0 18952 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _187_
timestamp 1676037725
transform 1 0 17848 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _188_
timestamp 1676037725
transform 1 0 20240 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1676037725
transform 1 0 20148 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _190_
timestamp 1676037725
transform 1 0 21068 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _191_
timestamp 1676037725
transform 1 0 20148 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _192_
timestamp 1676037725
transform 1 0 20056 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _193_
timestamp 1676037725
transform 1 0 22632 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _194_
timestamp 1676037725
transform 1 0 21988 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _195_
timestamp 1676037725
transform 1 0 23000 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1676037725
transform 1 0 24656 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _197_
timestamp 1676037725
transform 1 0 23552 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _198_
timestamp 1676037725
transform 1 0 5428 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _199_
timestamp 1676037725
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _200_
timestamp 1676037725
transform 1 0 4048 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _201_
timestamp 1676037725
transform 1 0 4048 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _202_
timestamp 1676037725
transform 1 0 5244 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _203_
timestamp 1676037725
transform 1 0 4968 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1676037725
transform 1 0 4876 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _205_
timestamp 1676037725
transform 1 0 4876 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1676037725
transform 1 0 45816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _207_
timestamp 1676037725
transform 1 0 2024 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _208_
timestamp 1676037725
transform 1 0 48576 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 1676037725
transform 1 0 46828 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1676037725
transform 1 0 46092 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _211_
timestamp 1676037725
transform 1 0 47840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _212_
timestamp 1676037725
transform 1 0 48576 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 1676037725
transform 1 0 48760 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _214_
timestamp 1676037725
transform 1 0 48024 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _215_
timestamp 1676037725
transform 1 0 48576 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1676037725
transform 1 0 47932 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 1676037725
transform 1 0 47932 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _218_
timestamp 1676037725
transform 1 0 48576 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1676037725
transform 1 0 47932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1676037725
transform 1 0 47932 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1676037725
transform 1 0 25024 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1676037725
transform 1 0 26496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1676037725
transform 1 0 30452 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1676037725
transform 1 0 31464 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1676037725
transform 1 0 34776 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1676037725
transform 1 0 37720 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1676037725
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1676037725
transform 1 0 22448 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1676037725
transform 1 0 21896 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1676037725
transform 1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1676037725
transform 1 0 28428 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1676037725
transform 1 0 29440 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1676037725
transform 1 0 26220 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1676037725
transform 1 0 33488 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1676037725
transform 1 0 33488 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1676037725
transform 1 0 23184 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1676037725
transform 1 0 36156 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1676037725
transform 1 0 23828 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1676037725
transform 1 0 38088 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1676037725
transform 1 0 22080 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1676037725
transform 1 0 22356 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1676037725
transform 1 0 21160 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1676037725
transform 1 0 20884 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1676037725
transform 1 0 25576 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1676037725
transform 1 0 26036 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1676037725
transform 1 0 41216 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1676037725
transform 1 0 39192 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1676037725
transform 1 0 23184 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1676037725
transform 1 0 21436 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1676037725
transform 1 0 30912 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1676037725
transform 1 0 22264 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1676037725
transform 1 0 21160 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1676037725
transform 1 0 21160 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1676037725
transform 1 0 27784 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1676037725
transform 1 0 18400 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_39
timestamp 1676037725
transform 1 0 38640 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_40
timestamp 1676037725
transform 1 0 31740 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_41
timestamp 1676037725
transform -1 0 35696 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 -1 8704
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_1_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23000 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_2_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20792 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_0.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19688 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21988 0 -1 23936
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 -1 19584
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21804 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_1.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19596 0 1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23000 0 -1 18496
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24748 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21620 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_2.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 19688 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 20976 0 1 17408
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22448 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.cby_0__1_.mem_right_ipin_3.sky130_fd_sc_hd__dfrtp_1_3_
timestamp 1676037725
transform 1 0 17112 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_0_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 26404 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27324 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 25852 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23368 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25208 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25116 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_2_
timestamp 1676037725
transform 1 0 20700 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3__271 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 23828 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l2_in_3_
timestamp 1676037725
transform 1 0 24564 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 22080 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l3_in_1_
timestamp 1676037725
transform 1 0 20700 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19320 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28796 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28428 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28244 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27140 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23000 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27140 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25760 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_2_
timestamp 1676037725
transform 1 0 18124 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3__272
timestamp 1676037725
transform 1 0 25760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l2_in_3_
timestamp 1676037725
transform 1 0 24564 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l3_in_1_
timestamp 1676037725
transform 1 0 22448 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19872 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29992 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28428 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27232 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l1_in_4_
timestamp 1676037725
transform 1 0 23276 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25944 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_2_
timestamp 1676037725
transform 1 0 20700 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3__273
timestamp 1676037725
transform 1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l2_in_3_
timestamp 1676037725
transform 1 0 22908 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l3_in_1_
timestamp 1676037725
transform 1 0 19320 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.mux_l4_in_0_
timestamp 1676037725
transform 1 0 19412 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 14260 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_2_
timestamp 1676037725
transform 1 0 26680 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_3_
timestamp 1676037725
transform 1 0 25024 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l1_in_4_
timestamp 1676037725
transform 1 0 20240 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_2_
timestamp 1676037725
transform 1 0 19412 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3__274
timestamp 1676037725
transform 1 0 22632 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l2_in_3_
timestamp 1676037725
transform 1 0 22264 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20700 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l3_in_1_
timestamp 1676037725
transform 1 0 19320 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.mux_l4_in_0_
timestamp 1676037725
transform 1 0 17388 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 13432 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7360 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 7636 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10580 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 9108 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14628 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7544 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 10580 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 8740 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 12880 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7820 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 8372 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE
timestamp 1676037725
transform 1 0 12512 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9108 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 14720 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__ebufn_8  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.IN_PROTECT_GATE
timestamp 1676037725
transform 1 0 7636 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.INV_SOC_DIR
timestamp 1676037725
transform 1 0 9108 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.ISOL_EN_GATE pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 17848 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_1  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.OUT_PROTECT_GATE
timestamp 1676037725
transform 1 0 9568 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22724 0 -1 16320
box -38 -48 2154 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 27048 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_prog_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 20516 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_prog_clk
timestamp 1676037725
transform 1 0 21436 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_prog_clk
timestamp 1676037725
transform 1 0 28428 0 -1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_prog_clk
timestamp 1676037725
transform 1 0 28244 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_prog_clk
timestamp 1676037725
transform 1 0 20976 0 1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_prog_clk
timestamp 1676037725
transform 1 0 22448 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_prog_clk
timestamp 1676037725
transform 1 0 27232 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_prog_clk
timestamp 1676037725
transform 1 0 27140 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_prog_clk
timestamp 1676037725
transform 1 0 34868 0 1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_prog_clk
timestamp 1676037725
transform 1 0 32844 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_prog_clk
timestamp 1676037725
transform 1 0 37444 0 -1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_prog_clk
timestamp 1676037725
transform 1 0 37628 0 -1 28288
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_prog_clk
timestamp 1676037725
transform 1 0 31832 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_prog_clk
timestamp 1676037725
transform 1 0 30452 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_prog_clk
timestamp 1676037725
transform 1 0 37076 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_prog_clk
timestamp 1676037725
transform 1 0 35972 0 -1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3772 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43
timestamp 1676037725
transform 1 0 5060 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1676037725
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1676037725
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57
timestamp 1676037725
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1676037725
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72
timestamp 1676037725
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1676037725
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_85
timestamp 1676037725
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93
timestamp 1676037725
transform 1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_100
timestamp 1676037725
transform 1 0 10304 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1676037725
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1676037725
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_123
timestamp 1676037725
transform 1 0 12420 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_131
timestamp 1676037725
transform 1 0 13156 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1676037725
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_141 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_148
timestamp 1676037725
transform 1 0 14720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_156
timestamp 1676037725
transform 1 0 15456 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1676037725
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1676037725
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_179
timestamp 1676037725
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1676037725
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1676037725
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_197
timestamp 1676037725
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_201
timestamp 1676037725
transform 1 0 19596 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_208
timestamp 1676037725
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1676037725
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_225
timestamp 1676037725
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_233
timestamp 1676037725
transform 1 0 22540 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_250
timestamp 1676037725
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_253
timestamp 1676037725
transform 1 0 24380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_261
timestamp 1676037725
transform 1 0 25116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_278
timestamp 1676037725
transform 1 0 26680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_281
timestamp 1676037725
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1676037725
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_307
timestamp 1676037725
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1676037725
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_327
timestamp 1676037725
transform 1 0 31188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1676037725
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_337
timestamp 1676037725
transform 1 0 32108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_355
timestamp 1676037725
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1676037725
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1676037725
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_383
timestamp 1676037725
transform 1 0 36340 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1676037725
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_393
timestamp 1676037725
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_411
timestamp 1676037725
transform 1 0 38916 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_419
timestamp 1676037725
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_421
timestamp 1676037725
transform 1 0 39836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_439
timestamp 1676037725
transform 1 0 41492 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_447
timestamp 1676037725
transform 1 0 42228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_449
timestamp 1676037725
transform 1 0 42412 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_467
timestamp 1676037725
transform 1 0 44068 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1676037725
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_477
timestamp 1676037725
transform 1 0 44988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_481
timestamp 1676037725
transform 1 0 45356 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_502
timestamp 1676037725
transform 1 0 47288 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1676037725
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_523
timestamp 1676037725
transform 1 0 49220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1676037725
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1676037725
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_28
timestamp 1676037725
transform 1 0 3680 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_33
timestamp 1676037725
transform 1 0 4140 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1676037725
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1676037725
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1676037725
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_65
timestamp 1676037725
transform 1 0 7084 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_77
timestamp 1676037725
transform 1 0 8188 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1676037725
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1676037725
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1676037725
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1676037725
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_129
timestamp 1676037725
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_145
timestamp 1676037725
transform 1 0 14444 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_157
timestamp 1676037725
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1676037725
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1676037725
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_187
timestamp 1676037725
transform 1 0 18308 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_195
timestamp 1676037725
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_207
timestamp 1676037725
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_211
timestamp 1676037725
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1676037725
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 1676037725
transform 1 0 21804 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_237
timestamp 1676037725
transform 1 0 22908 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1676037725
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_277
timestamp 1676037725
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_281
timestamp 1676037725
transform 1 0 26956 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1676037725
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_321
timestamp 1676037725
transform 1 0 30636 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_333
timestamp 1676037725
transform 1 0 31740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_337
timestamp 1676037725
transform 1 0 32108 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_355
timestamp 1676037725
transform 1 0 33764 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_375
timestamp 1676037725
transform 1 0 35604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_387
timestamp 1676037725
transform 1 0 36708 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1676037725
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1676037725
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_411
timestamp 1676037725
transform 1 0 38916 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_431
timestamp 1676037725
transform 1 0 40756 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_443
timestamp 1676037725
transform 1 0 41860 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 1676037725
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_449
timestamp 1676037725
transform 1 0 42412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_467
timestamp 1676037725
transform 1 0 44068 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_487
timestamp 1676037725
transform 1 0 45908 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_495
timestamp 1676037725
transform 1 0 46644 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_502
timestamp 1676037725
transform 1 0 47288 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_505
timestamp 1676037725
transform 1 0 47564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_525
timestamp 1676037725
transform 1 0 49404 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_3
timestamp 1676037725
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_8
timestamp 1676037725
transform 1 0 1840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1676037725
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1676037725
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1676037725
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1676037725
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1676037725
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1676037725
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1676037725
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1676037725
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1676037725
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1676037725
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1676037725
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1676037725
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1676037725
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1676037725
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1676037725
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1676037725
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1676037725
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1676037725
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1676037725
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1676037725
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1676037725
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1676037725
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1676037725
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1676037725
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1676037725
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1676037725
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_271
timestamp 1676037725
transform 1 0 26036 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_283
timestamp 1676037725
transform 1 0 27140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_295
timestamp 1676037725
transform 1 0 28244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1676037725
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_309
timestamp 1676037725
transform 1 0 29532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_327
timestamp 1676037725
transform 1 0 31188 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_347
timestamp 1676037725
transform 1 0 33028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_359
timestamp 1676037725
transform 1 0 34132 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1676037725
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_365
timestamp 1676037725
transform 1 0 34684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_383
timestamp 1676037725
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_403
timestamp 1676037725
transform 1 0 38180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_415
timestamp 1676037725
transform 1 0 39284 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_419
timestamp 1676037725
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1676037725
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_439
timestamp 1676037725
transform 1 0 41492 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_459
timestamp 1676037725
transform 1 0 43332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_471
timestamp 1676037725
transform 1 0 44436 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_475
timestamp 1676037725
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_477
timestamp 1676037725
transform 1 0 44988 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_495
timestamp 1676037725
transform 1 0 46644 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_507
timestamp 1676037725
transform 1 0 47748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_525
timestamp 1676037725
transform 1 0 49404 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1676037725
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1676037725
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1676037725
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1676037725
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1676037725
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1676037725
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1676037725
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1676037725
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1676037725
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1676037725
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1676037725
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1676037725
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1676037725
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1676037725
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1676037725
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1676037725
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1676037725
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1676037725
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1676037725
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1676037725
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1676037725
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1676037725
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1676037725
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1676037725
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1676037725
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1676037725
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1676037725
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1676037725
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1676037725
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1676037725
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1676037725
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1676037725
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1676037725
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1676037725
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1676037725
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1676037725
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1676037725
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_349
timestamp 1676037725
transform 1 0 33212 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1676037725
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1676037725
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1676037725
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1676037725
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_405
timestamp 1676037725
transform 1 0 38364 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_429
timestamp 1676037725
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_441
timestamp 1676037725
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1676037725
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1676037725
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_477
timestamp 1676037725
transform 1 0 44988 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_485
timestamp 1676037725
transform 1 0 45724 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_489
timestamp 1676037725
transform 1 0 46092 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_501
timestamp 1676037725
transform 1 0 47196 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_505
timestamp 1676037725
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_521
timestamp 1676037725
transform 1 0 49036 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1676037725
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1676037725
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1676037725
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1676037725
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1676037725
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1676037725
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1676037725
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1676037725
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1676037725
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1676037725
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1676037725
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1676037725
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1676037725
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1676037725
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1676037725
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1676037725
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1676037725
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1676037725
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1676037725
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1676037725
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1676037725
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1676037725
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1676037725
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1676037725
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1676037725
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1676037725
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1676037725
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1676037725
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1676037725
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1676037725
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1676037725
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1676037725
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1676037725
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1676037725
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1676037725
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1676037725
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1676037725
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1676037725
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1676037725
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1676037725
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1676037725
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1676037725
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_401
timestamp 1676037725
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1676037725
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1676037725
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1676037725
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1676037725
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_445
timestamp 1676037725
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_457
timestamp 1676037725
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_469
timestamp 1676037725
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_475
timestamp 1676037725
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_477
timestamp 1676037725
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_489
timestamp 1676037725
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_501
timestamp 1676037725
transform 1 0 47196 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_525
timestamp 1676037725
transform 1 0 49404 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1676037725
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1676037725
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1676037725
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1676037725
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1676037725
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1676037725
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1676037725
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1676037725
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1676037725
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1676037725
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1676037725
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1676037725
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1676037725
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1676037725
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1676037725
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1676037725
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1676037725
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1676037725
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1676037725
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1676037725
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1676037725
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1676037725
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1676037725
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1676037725
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1676037725
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1676037725
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1676037725
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1676037725
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1676037725
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1676037725
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1676037725
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1676037725
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_305
timestamp 1676037725
transform 1 0 29164 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_310
timestamp 1676037725
transform 1 0 29624 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_318
timestamp 1676037725
transform 1 0 30360 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_330
timestamp 1676037725
transform 1 0 31464 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1676037725
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1676037725
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1676037725
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1676037725
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1676037725
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1676037725
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1676037725
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_405
timestamp 1676037725
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_417
timestamp 1676037725
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_429
timestamp 1676037725
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1676037725
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1676037725
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_449
timestamp 1676037725
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_461
timestamp 1676037725
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_473
timestamp 1676037725
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_485
timestamp 1676037725
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_497
timestamp 1676037725
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_503
timestamp 1676037725
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_505
timestamp 1676037725
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_517
timestamp 1676037725
transform 1 0 48668 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_521
timestamp 1676037725
transform 1 0 49036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_525
timestamp 1676037725
transform 1 0 49404 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1676037725
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1676037725
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1676037725
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1676037725
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1676037725
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1676037725
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1676037725
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1676037725
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1676037725
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1676037725
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1676037725
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1676037725
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1676037725
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1676037725
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1676037725
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1676037725
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1676037725
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1676037725
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1676037725
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1676037725
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1676037725
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1676037725
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1676037725
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1676037725
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1676037725
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1676037725
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1676037725
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1676037725
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1676037725
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1676037725
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1676037725
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1676037725
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1676037725
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1676037725
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1676037725
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1676037725
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1676037725
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1676037725
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1676037725
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1676037725
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1676037725
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1676037725
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_401
timestamp 1676037725
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1676037725
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1676037725
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_421
timestamp 1676037725
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1676037725
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1676037725
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_457
timestamp 1676037725
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1676037725
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1676037725
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_477
timestamp 1676037725
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_489
timestamp 1676037725
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_501
timestamp 1676037725
transform 1 0 47196 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_525
timestamp 1676037725
transform 1 0 49404 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1676037725
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1676037725
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1676037725
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1676037725
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1676037725
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1676037725
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1676037725
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1676037725
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1676037725
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1676037725
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1676037725
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1676037725
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1676037725
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1676037725
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1676037725
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1676037725
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1676037725
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1676037725
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1676037725
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1676037725
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1676037725
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1676037725
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1676037725
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1676037725
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1676037725
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1676037725
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1676037725
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1676037725
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1676037725
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1676037725
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1676037725
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1676037725
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1676037725
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1676037725
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1676037725
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1676037725
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1676037725
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1676037725
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1676037725
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1676037725
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1676037725
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1676037725
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1676037725
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1676037725
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1676037725
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1676037725
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1676037725
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1676037725
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_449
timestamp 1676037725
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_461
timestamp 1676037725
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_473
timestamp 1676037725
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_485
timestamp 1676037725
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1676037725
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1676037725
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_505
timestamp 1676037725
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_517
timestamp 1676037725
transform 1 0 48668 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_525
timestamp 1676037725
transform 1 0 49404 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1676037725
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1676037725
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1676037725
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1676037725
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1676037725
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1676037725
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1676037725
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1676037725
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1676037725
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1676037725
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1676037725
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1676037725
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1676037725
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1676037725
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1676037725
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1676037725
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1676037725
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1676037725
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1676037725
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1676037725
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1676037725
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1676037725
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1676037725
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1676037725
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1676037725
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1676037725
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1676037725
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1676037725
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1676037725
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1676037725
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1676037725
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1676037725
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1676037725
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1676037725
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1676037725
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1676037725
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1676037725
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1676037725
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1676037725
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1676037725
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1676037725
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_389
timestamp 1676037725
transform 1 0 36892 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_399
timestamp 1676037725
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_407
timestamp 1676037725
transform 1 0 38548 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1676037725
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_421
timestamp 1676037725
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1676037725
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1676037725
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_457
timestamp 1676037725
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1676037725
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1676037725
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_477
timestamp 1676037725
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_489
timestamp 1676037725
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_501
timestamp 1676037725
transform 1 0 47196 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_525
timestamp 1676037725
transform 1 0 49404 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1676037725
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1676037725
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1676037725
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1676037725
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1676037725
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1676037725
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1676037725
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1676037725
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1676037725
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1676037725
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1676037725
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1676037725
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1676037725
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1676037725
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1676037725
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1676037725
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1676037725
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1676037725
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1676037725
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1676037725
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1676037725
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1676037725
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1676037725
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1676037725
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1676037725
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1676037725
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1676037725
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1676037725
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1676037725
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1676037725
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1676037725
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1676037725
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1676037725
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1676037725
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1676037725
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1676037725
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1676037725
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1676037725
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1676037725
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_373
timestamp 1676037725
transform 1 0 35420 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_379
timestamp 1676037725
transform 1 0 35972 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1676037725
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_393
timestamp 1676037725
transform 1 0 37260 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_399
timestamp 1676037725
transform 1 0 37812 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_411
timestamp 1676037725
transform 1 0 38916 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_423
timestamp 1676037725
transform 1 0 40020 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_435
timestamp 1676037725
transform 1 0 41124 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1676037725
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_449
timestamp 1676037725
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_461
timestamp 1676037725
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_473
timestamp 1676037725
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_485
timestamp 1676037725
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_497
timestamp 1676037725
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_503
timestamp 1676037725
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_505
timestamp 1676037725
transform 1 0 47564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_525
timestamp 1676037725
transform 1 0 49404 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1676037725
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1676037725
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1676037725
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1676037725
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1676037725
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1676037725
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1676037725
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1676037725
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1676037725
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1676037725
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1676037725
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1676037725
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1676037725
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1676037725
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1676037725
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1676037725
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1676037725
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1676037725
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1676037725
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1676037725
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1676037725
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1676037725
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1676037725
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1676037725
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1676037725
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1676037725
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1676037725
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1676037725
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1676037725
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1676037725
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1676037725
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1676037725
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1676037725
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1676037725
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1676037725
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1676037725
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1676037725
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1676037725
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1676037725
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1676037725
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1676037725
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1676037725
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_401
timestamp 1676037725
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1676037725
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1676037725
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_421
timestamp 1676037725
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1676037725
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1676037725
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_457
timestamp 1676037725
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1676037725
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1676037725
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_477
timestamp 1676037725
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_489
timestamp 1676037725
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_501
timestamp 1676037725
transform 1 0 47196 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_525
timestamp 1676037725
transform 1 0 49404 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1676037725
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1676037725
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1676037725
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1676037725
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1676037725
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1676037725
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1676037725
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1676037725
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_81
timestamp 1676037725
transform 1 0 8556 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1676037725
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1676037725
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1676037725
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1676037725
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1676037725
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1676037725
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1676037725
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1676037725
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1676037725
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1676037725
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1676037725
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1676037725
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1676037725
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1676037725
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1676037725
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1676037725
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1676037725
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1676037725
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1676037725
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1676037725
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1676037725
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1676037725
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1676037725
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1676037725
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1676037725
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1676037725
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1676037725
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1676037725
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_373
timestamp 1676037725
transform 1 0 35420 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_381
timestamp 1676037725
transform 1 0 36156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_388
timestamp 1676037725
transform 1 0 36800 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_393
timestamp 1676037725
transform 1 0 37260 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_397
timestamp 1676037725
transform 1 0 37628 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_402
timestamp 1676037725
transform 1 0 38088 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_414
timestamp 1676037725
transform 1 0 39192 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_426
timestamp 1676037725
transform 1 0 40296 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_438
timestamp 1676037725
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_446
timestamp 1676037725
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_449
timestamp 1676037725
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_461
timestamp 1676037725
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_473
timestamp 1676037725
transform 1 0 44620 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_481
timestamp 1676037725
transform 1 0 45356 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_488
timestamp 1676037725
transform 1 0 46000 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_500
timestamp 1676037725
transform 1 0 47104 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_505
timestamp 1676037725
transform 1 0 47564 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_525
timestamp 1676037725
transform 1 0 49404 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1676037725
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1676037725
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1676037725
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1676037725
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1676037725
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1676037725
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1676037725
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1676037725
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1676037725
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1676037725
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1676037725
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1676037725
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1676037725
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1676037725
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1676037725
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1676037725
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1676037725
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1676037725
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1676037725
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1676037725
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1676037725
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1676037725
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1676037725
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1676037725
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1676037725
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1676037725
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1676037725
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1676037725
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1676037725
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1676037725
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1676037725
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1676037725
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1676037725
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1676037725
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1676037725
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1676037725
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1676037725
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1676037725
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1676037725
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1676037725
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1676037725
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1676037725
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1676037725
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1676037725
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1676037725
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_421
timestamp 1676037725
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1676037725
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1676037725
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_457
timestamp 1676037725
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1676037725
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1676037725
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_477
timestamp 1676037725
transform 1 0 44988 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_485
timestamp 1676037725
transform 1 0 45724 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_491
timestamp 1676037725
transform 1 0 46276 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_503
timestamp 1676037725
transform 1 0 47380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1676037725
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1676037725
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_520
timestamp 1676037725
transform 1 0 48944 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_526
timestamp 1676037725
transform 1 0 49496 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1676037725
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1676037725
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1676037725
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1676037725
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1676037725
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1676037725
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1676037725
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1676037725
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1676037725
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1676037725
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1676037725
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1676037725
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1676037725
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1676037725
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1676037725
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1676037725
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1676037725
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1676037725
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1676037725
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1676037725
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1676037725
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1676037725
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1676037725
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1676037725
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1676037725
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1676037725
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1676037725
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1676037725
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1676037725
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1676037725
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1676037725
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1676037725
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1676037725
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1676037725
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1676037725
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1676037725
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_337
timestamp 1676037725
transform 1 0 32108 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_343
timestamp 1676037725
transform 1 0 32660 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_355
timestamp 1676037725
transform 1 0 33764 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_367
timestamp 1676037725
transform 1 0 34868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_375
timestamp 1676037725
transform 1 0 35604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_381
timestamp 1676037725
transform 1 0 36156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_389
timestamp 1676037725
transform 1 0 36892 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1676037725
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1676037725
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1676037725
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1676037725
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1676037725
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1676037725
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_449
timestamp 1676037725
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_461
timestamp 1676037725
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_473
timestamp 1676037725
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_485
timestamp 1676037725
transform 1 0 45724 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_492
timestamp 1676037725
transform 1 0 46368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_505
timestamp 1676037725
transform 1 0 47564 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_525
timestamp 1676037725
transform 1 0 49404 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1676037725
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1676037725
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1676037725
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1676037725
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1676037725
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1676037725
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1676037725
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1676037725
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1676037725
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1676037725
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1676037725
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1676037725
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1676037725
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1676037725
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1676037725
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1676037725
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1676037725
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1676037725
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1676037725
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1676037725
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1676037725
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1676037725
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1676037725
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1676037725
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1676037725
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1676037725
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1676037725
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1676037725
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1676037725
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1676037725
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_289
timestamp 1676037725
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_297
timestamp 1676037725
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1676037725
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1676037725
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1676037725
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1676037725
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_337
timestamp 1676037725
transform 1 0 32108 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_349
timestamp 1676037725
transform 1 0 33212 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 1676037725
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1676037725
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1676037725
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1676037725
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_401
timestamp 1676037725
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1676037725
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1676037725
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1676037725
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1676037725
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_445
timestamp 1676037725
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_457
timestamp 1676037725
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1676037725
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1676037725
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_477
timestamp 1676037725
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_489
timestamp 1676037725
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_501
timestamp 1676037725
transform 1 0 47196 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_525
timestamp 1676037725
transform 1 0 49404 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1676037725
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1676037725
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1676037725
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1676037725
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1676037725
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1676037725
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1676037725
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1676037725
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1676037725
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1676037725
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1676037725
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1676037725
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1676037725
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1676037725
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1676037725
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1676037725
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1676037725
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1676037725
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1676037725
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1676037725
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1676037725
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1676037725
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1676037725
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1676037725
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1676037725
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1676037725
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_249
timestamp 1676037725
transform 1 0 24012 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_257
timestamp 1676037725
transform 1 0 24748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_269
timestamp 1676037725
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_277
timestamp 1676037725
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1676037725
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1676037725
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1676037725
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1676037725
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1676037725
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1676037725
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1676037725
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1676037725
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1676037725
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1676037725
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1676037725
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1676037725
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1676037725
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1676037725
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1676037725
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_432
timestamp 1676037725
transform 1 0 40848 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_444
timestamp 1676037725
transform 1 0 41952 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1676037725
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_461
timestamp 1676037725
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_473
timestamp 1676037725
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_485
timestamp 1676037725
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_497
timestamp 1676037725
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1676037725
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1676037725
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_525
timestamp 1676037725
transform 1 0 49404 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1676037725
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1676037725
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1676037725
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1676037725
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1676037725
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1676037725
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1676037725
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1676037725
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1676037725
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1676037725
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1676037725
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1676037725
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1676037725
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1676037725
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1676037725
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 1676037725
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_146
timestamp 1676037725
transform 1 0 14536 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_158
timestamp 1676037725
transform 1 0 15640 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_170
timestamp 1676037725
transform 1 0 16744 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_182
timestamp 1676037725
transform 1 0 17848 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1676037725
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1676037725
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1676037725
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1676037725
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1676037725
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1676037725
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1676037725
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1676037725
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1676037725
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1676037725
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1676037725
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1676037725
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1676037725
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1676037725
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1676037725
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1676037725
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1676037725
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1676037725
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1676037725
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1676037725
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1676037725
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1676037725
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1676037725
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1676037725
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1676037725
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1676037725
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1676037725
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1676037725
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_457
timestamp 1676037725
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1676037725
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1676037725
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_477
timestamp 1676037725
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_489
timestamp 1676037725
transform 1 0 46092 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_494
timestamp 1676037725
transform 1 0 46552 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_506
timestamp 1676037725
transform 1 0 47656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_525
timestamp 1676037725
transform 1 0 49404 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1676037725
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1676037725
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1676037725
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1676037725
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1676037725
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1676037725
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1676037725
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1676037725
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1676037725
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1676037725
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1676037725
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1676037725
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1676037725
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1676037725
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1676037725
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1676037725
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1676037725
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1676037725
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1676037725
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1676037725
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1676037725
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1676037725
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1676037725
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1676037725
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1676037725
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1676037725
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1676037725
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1676037725
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1676037725
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1676037725
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1676037725
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1676037725
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1676037725
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1676037725
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1676037725
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1676037725
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1676037725
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1676037725
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1676037725
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1676037725
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1676037725
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1676037725
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1676037725
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1676037725
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1676037725
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_429
timestamp 1676037725
transform 1 0 40572 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_437
timestamp 1676037725
transform 1 0 41308 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1676037725
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1676037725
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1676037725
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_461
timestamp 1676037725
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_473
timestamp 1676037725
transform 1 0 44620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_478
timestamp 1676037725
transform 1 0 45080 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_486
timestamp 1676037725
transform 1 0 45816 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_494
timestamp 1676037725
transform 1 0 46552 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_502
timestamp 1676037725
transform 1 0 47288 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_505
timestamp 1676037725
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_517
timestamp 1676037725
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_525
timestamp 1676037725
transform 1 0 49404 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1676037725
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1676037725
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1676037725
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1676037725
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1676037725
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1676037725
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1676037725
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1676037725
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1676037725
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1676037725
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1676037725
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1676037725
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1676037725
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1676037725
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1676037725
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1676037725
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1676037725
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1676037725
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1676037725
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1676037725
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1676037725
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1676037725
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1676037725
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1676037725
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1676037725
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1676037725
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1676037725
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1676037725
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1676037725
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1676037725
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_289
timestamp 1676037725
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_297
timestamp 1676037725
transform 1 0 28428 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1676037725
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1676037725
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1676037725
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1676037725
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1676037725
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1676037725
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1676037725
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1676037725
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1676037725
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1676037725
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_401
timestamp 1676037725
transform 1 0 37996 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_409
timestamp 1676037725
transform 1 0 38732 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_414
timestamp 1676037725
transform 1 0 39192 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1676037725
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_433
timestamp 1676037725
transform 1 0 40940 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_437
timestamp 1676037725
transform 1 0 41308 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_449
timestamp 1676037725
transform 1 0 42412 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_461
timestamp 1676037725
transform 1 0 43516 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_472
timestamp 1676037725
transform 1 0 44528 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_477
timestamp 1676037725
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_489
timestamp 1676037725
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_501
timestamp 1676037725
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_525
timestamp 1676037725
transform 1 0 49404 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1676037725
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1676037725
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1676037725
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1676037725
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1676037725
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1676037725
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1676037725
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1676037725
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1676037725
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1676037725
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1676037725
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1676037725
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1676037725
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1676037725
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1676037725
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1676037725
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1676037725
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1676037725
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1676037725
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1676037725
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1676037725
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1676037725
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1676037725
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1676037725
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1676037725
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1676037725
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1676037725
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1676037725
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1676037725
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1676037725
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_281
timestamp 1676037725
transform 1 0 26956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_287
timestamp 1676037725
transform 1 0 27508 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_295
timestamp 1676037725
transform 1 0 28244 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_310
timestamp 1676037725
transform 1 0 29624 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_323
timestamp 1676037725
transform 1 0 30820 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1676037725
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1676037725
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_349
timestamp 1676037725
transform 1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_353
timestamp 1676037725
transform 1 0 33580 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_374
timestamp 1676037725
transform 1 0 35512 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_387
timestamp 1676037725
transform 1 0 36708 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1676037725
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1676037725
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1676037725
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_417
timestamp 1676037725
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_429
timestamp 1676037725
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_441
timestamp 1676037725
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_447
timestamp 1676037725
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1676037725
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_461
timestamp 1676037725
transform 1 0 43516 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_466
timestamp 1676037725
transform 1 0 43976 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_478
timestamp 1676037725
transform 1 0 45080 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_490
timestamp 1676037725
transform 1 0 46184 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_502
timestamp 1676037725
transform 1 0 47288 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_505
timestamp 1676037725
transform 1 0 47564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_525
timestamp 1676037725
transform 1 0 49404 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1676037725
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1676037725
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1676037725
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1676037725
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1676037725
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1676037725
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1676037725
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1676037725
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1676037725
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1676037725
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1676037725
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1676037725
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1676037725
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1676037725
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1676037725
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1676037725
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1676037725
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1676037725
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1676037725
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1676037725
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1676037725
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1676037725
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1676037725
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1676037725
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1676037725
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1676037725
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1676037725
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1676037725
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_265
timestamp 1676037725
transform 1 0 25484 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_270
timestamp 1676037725
transform 1 0 25944 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_282
timestamp 1676037725
transform 1 0 27048 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_294
timestamp 1676037725
transform 1 0 28152 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_304
timestamp 1676037725
transform 1 0 29072 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1676037725
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1676037725
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1676037725
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1676037725
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_357
timestamp 1676037725
transform 1 0 33948 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_362
timestamp 1676037725
transform 1 0 34408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_365
timestamp 1676037725
transform 1 0 34684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_387
timestamp 1676037725
transform 1 0 36708 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1676037725
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_402
timestamp 1676037725
transform 1 0 38088 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_409
timestamp 1676037725
transform 1 0 38732 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_417
timestamp 1676037725
transform 1 0 39468 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_421
timestamp 1676037725
transform 1 0 39836 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_427
timestamp 1676037725
transform 1 0 40388 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_432
timestamp 1676037725
transform 1 0 40848 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_444
timestamp 1676037725
transform 1 0 41952 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_456
timestamp 1676037725
transform 1 0 43056 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_468
timestamp 1676037725
transform 1 0 44160 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_477
timestamp 1676037725
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_489
timestamp 1676037725
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_501
timestamp 1676037725
transform 1 0 47196 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_525
timestamp 1676037725
transform 1 0 49404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 1676037725
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_21
timestamp 1676037725
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_33
timestamp 1676037725
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_45
timestamp 1676037725
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_53
timestamp 1676037725
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1676037725
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1676037725
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1676037725
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1676037725
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1676037725
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1676037725
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1676037725
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1676037725
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1676037725
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1676037725
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1676037725
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1676037725
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1676037725
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1676037725
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1676037725
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1676037725
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1676037725
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1676037725
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1676037725
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1676037725
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1676037725
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1676037725
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1676037725
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1676037725
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1676037725
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_293
timestamp 1676037725
transform 1 0 28060 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_301
timestamp 1676037725
transform 1 0 28796 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_306
timestamp 1676037725
transform 1 0 29256 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_318
timestamp 1676037725
transform 1 0 30360 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_322
timestamp 1676037725
transform 1 0 30728 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1676037725
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1676037725
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_349
timestamp 1676037725
transform 1 0 33212 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_355
timestamp 1676037725
transform 1 0 33764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_376
timestamp 1676037725
transform 1 0 35696 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_384
timestamp 1676037725
transform 1 0 36432 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1676037725
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_393
timestamp 1676037725
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_399
timestamp 1676037725
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_407
timestamp 1676037725
transform 1 0 38548 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_414
timestamp 1676037725
transform 1 0 39192 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_426
timestamp 1676037725
transform 1 0 40296 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_438
timestamp 1676037725
transform 1 0 41400 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_443
timestamp 1676037725
transform 1 0 41860 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1676037725
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_449
timestamp 1676037725
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_461
timestamp 1676037725
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_473
timestamp 1676037725
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_485
timestamp 1676037725
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_497
timestamp 1676037725
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1676037725
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_505
timestamp 1676037725
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_525
timestamp 1676037725
transform 1 0 49404 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1676037725
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1676037725
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1676037725
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1676037725
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1676037725
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1676037725
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1676037725
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1676037725
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1676037725
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1676037725
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1676037725
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1676037725
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1676037725
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1676037725
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1676037725
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1676037725
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1676037725
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1676037725
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1676037725
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1676037725
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1676037725
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1676037725
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1676037725
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1676037725
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1676037725
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1676037725
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1676037725
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1676037725
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_265
timestamp 1676037725
transform 1 0 25484 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1676037725
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1676037725
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1676037725
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1676037725
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1676037725
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_333
timestamp 1676037725
transform 1 0 31740 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_339
timestamp 1676037725
transform 1 0 32292 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_352
timestamp 1676037725
transform 1 0 33488 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_365
timestamp 1676037725
transform 1 0 34684 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_371
timestamp 1676037725
transform 1 0 35236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_383
timestamp 1676037725
transform 1 0 36340 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_391
timestamp 1676037725
transform 1 0 37076 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_401
timestamp 1676037725
transform 1 0 37996 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_408
timestamp 1676037725
transform 1 0 38640 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1676037725
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_426
timestamp 1676037725
transform 1 0 40296 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_438
timestamp 1676037725
transform 1 0 41400 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_450
timestamp 1676037725
transform 1 0 42504 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_462
timestamp 1676037725
transform 1 0 43608 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_474
timestamp 1676037725
transform 1 0 44712 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_477
timestamp 1676037725
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_489
timestamp 1676037725
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_501
timestamp 1676037725
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_513
timestamp 1676037725
transform 1 0 48300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_525
timestamp 1676037725
transform 1 0 49404 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1676037725
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1676037725
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1676037725
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1676037725
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1676037725
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1676037725
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1676037725
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1676037725
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1676037725
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1676037725
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1676037725
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1676037725
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1676037725
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1676037725
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1676037725
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1676037725
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1676037725
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1676037725
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1676037725
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1676037725
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1676037725
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_205
timestamp 1676037725
transform 1 0 19964 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_209
timestamp 1676037725
transform 1 0 20332 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_219
timestamp 1676037725
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1676037725
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_225
timestamp 1676037725
transform 1 0 21804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_231
timestamp 1676037725
transform 1 0 22356 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_252
timestamp 1676037725
transform 1 0 24288 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1676037725
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_268
timestamp 1676037725
transform 1 0 25760 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1676037725
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_281
timestamp 1676037725
transform 1 0 26956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_287
timestamp 1676037725
transform 1 0 27508 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_308
timestamp 1676037725
transform 1 0 29440 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1676037725
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_323
timestamp 1676037725
transform 1 0 30820 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_329
timestamp 1676037725
transform 1 0 31372 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_334
timestamp 1676037725
transform 1 0 31832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_337
timestamp 1676037725
transform 1 0 32108 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_348
timestamp 1676037725
transform 1 0 33120 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_360
timestamp 1676037725
transform 1 0 34224 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_372
timestamp 1676037725
transform 1 0 35328 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_384
timestamp 1676037725
transform 1 0 36432 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1676037725
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_404
timestamp 1676037725
transform 1 0 38272 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_416
timestamp 1676037725
transform 1 0 39376 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_428
timestamp 1676037725
transform 1 0 40480 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_443
timestamp 1676037725
transform 1 0 41860 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1676037725
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_449
timestamp 1676037725
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_461
timestamp 1676037725
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_473
timestamp 1676037725
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_485
timestamp 1676037725
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_497
timestamp 1676037725
transform 1 0 46828 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_503
timestamp 1676037725
transform 1 0 47380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_505
timestamp 1676037725
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_525
timestamp 1676037725
transform 1 0 49404 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1676037725
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1676037725
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1676037725
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1676037725
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1676037725
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1676037725
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1676037725
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1676037725
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1676037725
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1676037725
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1676037725
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1676037725
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1676037725
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1676037725
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1676037725
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1676037725
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1676037725
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1676037725
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1676037725
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1676037725
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1676037725
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1676037725
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1676037725
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1676037725
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1676037725
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1676037725
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1676037725
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 1676037725
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_259
timestamp 1676037725
transform 1 0 24932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_271
timestamp 1676037725
transform 1 0 26036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_284
timestamp 1676037725
transform 1 0 27232 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_297
timestamp 1676037725
transform 1 0 28428 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_301
timestamp 1676037725
transform 1 0 28796 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_306
timestamp 1676037725
transform 1 0 29256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_309
timestamp 1676037725
transform 1 0 29532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_331
timestamp 1676037725
transform 1 0 31556 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_339
timestamp 1676037725
transform 1 0 32292 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_343
timestamp 1676037725
transform 1 0 32660 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_356
timestamp 1676037725
transform 1 0 33856 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1676037725
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_377
timestamp 1676037725
transform 1 0 35788 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_398
timestamp 1676037725
transform 1 0 37720 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_410
timestamp 1676037725
transform 1 0 38824 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_418
timestamp 1676037725
transform 1 0 39560 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_421
timestamp 1676037725
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_433
timestamp 1676037725
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_445
timestamp 1676037725
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_457
timestamp 1676037725
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1676037725
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1676037725
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_477
timestamp 1676037725
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_489
timestamp 1676037725
transform 1 0 46092 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_501
timestamp 1676037725
transform 1 0 47196 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_525
timestamp 1676037725
transform 1 0 49404 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_3
timestamp 1676037725
transform 1 0 1380 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_21
timestamp 1676037725
transform 1 0 3036 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1676037725
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1676037725
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1676037725
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1676037725
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1676037725
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1676037725
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1676037725
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1676037725
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1676037725
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1676037725
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1676037725
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1676037725
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1676037725
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1676037725
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1676037725
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1676037725
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1676037725
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1676037725
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1676037725
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1676037725
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1676037725
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_225
timestamp 1676037725
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_233
timestamp 1676037725
transform 1 0 22540 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_258
timestamp 1676037725
transform 1 0 24840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_262
timestamp 1676037725
transform 1 0 25208 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1676037725
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1676037725
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_292
timestamp 1676037725
transform 1 0 27968 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_300
timestamp 1676037725
transform 1 0 28704 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_321
timestamp 1676037725
transform 1 0 30636 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_333
timestamp 1676037725
transform 1 0 31740 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_337
timestamp 1676037725
transform 1 0 32108 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_345
timestamp 1676037725
transform 1 0 32844 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_355
timestamp 1676037725
transform 1 0 33764 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_362
timestamp 1676037725
transform 1 0 34408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_369
timestamp 1676037725
transform 1 0 35052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_377
timestamp 1676037725
transform 1 0 35788 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_383
timestamp 1676037725
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1676037725
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1676037725
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_398
timestamp 1676037725
transform 1 0 37720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_406
timestamp 1676037725
transform 1 0 38456 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_411
timestamp 1676037725
transform 1 0 38916 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_423
timestamp 1676037725
transform 1 0 40020 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_435
timestamp 1676037725
transform 1 0 41124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1676037725
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_449
timestamp 1676037725
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_461
timestamp 1676037725
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_473
timestamp 1676037725
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_485
timestamp 1676037725
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1676037725
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1676037725
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_505
timestamp 1676037725
transform 1 0 47564 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_525
timestamp 1676037725
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1676037725
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1676037725
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1676037725
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1676037725
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_41
timestamp 1676037725
transform 1 0 4876 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_51
timestamp 1676037725
transform 1 0 5796 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_63
timestamp 1676037725
transform 1 0 6900 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1676037725
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1676037725
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1676037725
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1676037725
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1676037725
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1676037725
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1676037725
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1676037725
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1676037725
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1676037725
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1676037725
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1676037725
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1676037725
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1676037725
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_197
timestamp 1676037725
transform 1 0 19228 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_219
timestamp 1676037725
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_243
timestamp 1676037725
transform 1 0 23460 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1676037725
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 1676037725
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_264
timestamp 1676037725
transform 1 0 25392 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_270
timestamp 1676037725
transform 1 0 25944 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_275
timestamp 1676037725
transform 1 0 26404 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_292
timestamp 1676037725
transform 1 0 27968 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1676037725
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1676037725
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1676037725
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1676037725
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_345
timestamp 1676037725
transform 1 0 32844 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1676037725
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1676037725
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_387
timestamp 1676037725
transform 1 0 36708 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_26_404
timestamp 1676037725
transform 1 0 38272 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_416
timestamp 1676037725
transform 1 0 39376 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_421
timestamp 1676037725
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_433
timestamp 1676037725
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_445
timestamp 1676037725
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_457
timestamp 1676037725
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1676037725
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1676037725
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_477
timestamp 1676037725
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_489
timestamp 1676037725
transform 1 0 46092 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_501
timestamp 1676037725
transform 1 0 47196 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_525
timestamp 1676037725
transform 1 0 49404 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1676037725
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1676037725
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1676037725
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1676037725
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1676037725
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1676037725
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1676037725
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1676037725
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1676037725
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1676037725
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1676037725
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1676037725
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1676037725
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1676037725
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1676037725
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1676037725
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1676037725
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1676037725
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1676037725
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1676037725
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1676037725
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_201
timestamp 1676037725
transform 1 0 19596 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1676037725
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1676037725
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_246
timestamp 1676037725
transform 1 0 23736 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_254
timestamp 1676037725
transform 1 0 24472 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1676037725
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_281
timestamp 1676037725
transform 1 0 26956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_293
timestamp 1676037725
transform 1 0 28060 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_306
timestamp 1676037725
transform 1 0 29256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_334
timestamp 1676037725
transform 1 0 31832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1676037725
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_342
timestamp 1676037725
transform 1 0 32568 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_350
timestamp 1676037725
transform 1 0 33304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_361
timestamp 1676037725
transform 1 0 34316 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_374
timestamp 1676037725
transform 1 0 35512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_381
timestamp 1676037725
transform 1 0 36156 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1676037725
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_393
timestamp 1676037725
transform 1 0 37260 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_399
timestamp 1676037725
transform 1 0 37812 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_403
timestamp 1676037725
transform 1 0 38180 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_415
timestamp 1676037725
transform 1 0 39284 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_427
timestamp 1676037725
transform 1 0 40388 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_439
timestamp 1676037725
transform 1 0 41492 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1676037725
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_449
timestamp 1676037725
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_461
timestamp 1676037725
transform 1 0 43516 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_466
timestamp 1676037725
transform 1 0 43976 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_478
timestamp 1676037725
transform 1 0 45080 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_490
timestamp 1676037725
transform 1 0 46184 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_502
timestamp 1676037725
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_505
timestamp 1676037725
transform 1 0 47564 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_517
timestamp 1676037725
transform 1 0 48668 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_525
timestamp 1676037725
transform 1 0 49404 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1676037725
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1676037725
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1676037725
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1676037725
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1676037725
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1676037725
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1676037725
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1676037725
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1676037725
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1676037725
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1676037725
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1676037725
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1676037725
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1676037725
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1676037725
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1676037725
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1676037725
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1676037725
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_177
timestamp 1676037725
transform 1 0 17388 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1676037725
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1676037725
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_208
timestamp 1676037725
transform 1 0 20240 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_239
timestamp 1676037725
transform 1 0 23092 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_246
timestamp 1676037725
transform 1 0 23736 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1676037725
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1676037725
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_277
timestamp 1676037725
transform 1 0 26588 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_28_294
timestamp 1676037725
transform 1 0 28152 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_306
timestamp 1676037725
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1676037725
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1676037725
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_341
timestamp 1676037725
transform 1 0 32476 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1676037725
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_28_365
timestamp 1676037725
transform 1 0 34684 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_373
timestamp 1676037725
transform 1 0 35420 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_394
timestamp 1676037725
transform 1 0 37352 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_418
timestamp 1676037725
transform 1 0 39560 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_421
timestamp 1676037725
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_433
timestamp 1676037725
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_445
timestamp 1676037725
transform 1 0 42044 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_453
timestamp 1676037725
transform 1 0 42780 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_458
timestamp 1676037725
transform 1 0 43240 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_466
timestamp 1676037725
transform 1 0 43976 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_474
timestamp 1676037725
transform 1 0 44712 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_477
timestamp 1676037725
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_489
timestamp 1676037725
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_501
timestamp 1676037725
transform 1 0 47196 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_525
timestamp 1676037725
transform 1 0 49404 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_3
timestamp 1676037725
transform 1 0 1380 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_21
timestamp 1676037725
transform 1 0 3036 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_33
timestamp 1676037725
transform 1 0 4140 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_45
timestamp 1676037725
transform 1 0 5244 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_53
timestamp 1676037725
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1676037725
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1676037725
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1676037725
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1676037725
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1676037725
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1676037725
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1676037725
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1676037725
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1676037725
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1676037725
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1676037725
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1676037725
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1676037725
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1676037725
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_193
timestamp 1676037725
transform 1 0 18860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_197
timestamp 1676037725
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_207
timestamp 1676037725
transform 1 0 20148 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_222
timestamp 1676037725
transform 1 0 21528 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1676037725
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_237
timestamp 1676037725
transform 1 0 22908 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1676037725
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1676037725
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1676037725
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_281
timestamp 1676037725
transform 1 0 26956 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_293
timestamp 1676037725
transform 1 0 28060 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_308
timestamp 1676037725
transform 1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_321
timestamp 1676037725
transform 1 0 30636 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_333
timestamp 1676037725
transform 1 0 31740 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_337
timestamp 1676037725
transform 1 0 32108 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_359
timestamp 1676037725
transform 1 0 34132 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_383
timestamp 1676037725
transform 1 0 36340 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1676037725
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1676037725
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_404
timestamp 1676037725
transform 1 0 38272 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_416
timestamp 1676037725
transform 1 0 39376 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_428
timestamp 1676037725
transform 1 0 40480 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_440
timestamp 1676037725
transform 1 0 41584 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_449
timestamp 1676037725
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_461
timestamp 1676037725
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_473
timestamp 1676037725
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_485
timestamp 1676037725
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1676037725
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1676037725
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_505
timestamp 1676037725
transform 1 0 47564 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_525
timestamp 1676037725
transform 1 0 49404 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1676037725
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1676037725
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1676037725
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_29
timestamp 1676037725
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1676037725
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1676037725
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1676037725
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1676037725
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1676037725
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1676037725
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1676037725
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1676037725
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1676037725
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1676037725
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1676037725
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1676037725
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1676037725
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1676037725
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_177
timestamp 1676037725
transform 1 0 17388 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_181
timestamp 1676037725
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1676037725
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1676037725
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1676037725
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_205
timestamp 1676037725
transform 1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_217
timestamp 1676037725
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1676037725
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1676037725
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_264
timestamp 1676037725
transform 1 0 25392 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_279
timestamp 1676037725
transform 1 0 26772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1676037725
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_306
timestamp 1676037725
transform 1 0 29256 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1676037725
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_321
timestamp 1676037725
transform 1 0 30636 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1676037725
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1676037725
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1676037725
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1676037725
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1676037725
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_377
timestamp 1676037725
transform 1 0 35788 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_385
timestamp 1676037725
transform 1 0 36524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_409
timestamp 1676037725
transform 1 0 38732 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_417
timestamp 1676037725
transform 1 0 39468 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_421
timestamp 1676037725
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_433
timestamp 1676037725
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_445
timestamp 1676037725
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_457
timestamp 1676037725
transform 1 0 43148 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_465
timestamp 1676037725
transform 1 0 43884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_471
timestamp 1676037725
transform 1 0 44436 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1676037725
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_477
timestamp 1676037725
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_489
timestamp 1676037725
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_501
timestamp 1676037725
transform 1 0 47196 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_525
timestamp 1676037725
transform 1 0 49404 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1676037725
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1676037725
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1676037725
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1676037725
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1676037725
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1676037725
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1676037725
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1676037725
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1676037725
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1676037725
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1676037725
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1676037725
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1676037725
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1676037725
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1676037725
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1676037725
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1676037725
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1676037725
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1676037725
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1676037725
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_193
timestamp 1676037725
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_201
timestamp 1676037725
transform 1 0 19596 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_213
timestamp 1676037725
transform 1 0 20700 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_221
timestamp 1676037725
transform 1 0 21436 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_225
timestamp 1676037725
transform 1 0 21804 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_233
timestamp 1676037725
transform 1 0 22540 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_238
timestamp 1676037725
transform 1 0 23000 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_251
timestamp 1676037725
transform 1 0 24196 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_278
timestamp 1676037725
transform 1 0 26680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1676037725
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_292
timestamp 1676037725
transform 1 0 27968 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1676037725
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1676037725
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1676037725
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1676037725
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1676037725
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_349
timestamp 1676037725
transform 1 0 33212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_353
timestamp 1676037725
transform 1 0 33580 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_375
timestamp 1676037725
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1676037725
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1676037725
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1676037725
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_415
timestamp 1676037725
transform 1 0 39284 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_427
timestamp 1676037725
transform 1 0 40388 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_439
timestamp 1676037725
transform 1 0 41492 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1676037725
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_449
timestamp 1676037725
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_461
timestamp 1676037725
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_473
timestamp 1676037725
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_485
timestamp 1676037725
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_497
timestamp 1676037725
transform 1 0 46828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1676037725
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_505
timestamp 1676037725
transform 1 0 47564 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_525
timestamp 1676037725
transform 1 0 49404 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1676037725
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1676037725
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1676037725
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1676037725
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1676037725
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1676037725
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1676037725
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1676037725
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1676037725
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1676037725
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1676037725
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1676037725
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1676037725
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1676037725
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1676037725
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_141
timestamp 1676037725
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_146
timestamp 1676037725
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_158
timestamp 1676037725
transform 1 0 15640 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_170
timestamp 1676037725
transform 1 0 16744 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_182
timestamp 1676037725
transform 1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1676037725
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_197
timestamp 1676037725
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_221
timestamp 1676037725
transform 1 0 21436 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1676037725
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1676037725
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_253
timestamp 1676037725
transform 1 0 24380 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_261
timestamp 1676037725
transform 1 0 25116 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_271
timestamp 1676037725
transform 1 0 26036 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_277
timestamp 1676037725
transform 1 0 26588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_287
timestamp 1676037725
transform 1 0 27508 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_299
timestamp 1676037725
transform 1 0 28612 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1676037725
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1676037725
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1676037725
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_333
timestamp 1676037725
transform 1 0 31740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_337
timestamp 1676037725
transform 1 0 32108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_342
timestamp 1676037725
transform 1 0 32568 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_346
timestamp 1676037725
transform 1 0 32936 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_351
timestamp 1676037725
transform 1 0 33396 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1676037725
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1676037725
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1676037725
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_371
timestamp 1676037725
transform 1 0 35236 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_378
timestamp 1676037725
transform 1 0 35880 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_390
timestamp 1676037725
transform 1 0 36984 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_402
timestamp 1676037725
transform 1 0 38088 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_414
timestamp 1676037725
transform 1 0 39192 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_421
timestamp 1676037725
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_433
timestamp 1676037725
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_445
timestamp 1676037725
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_457
timestamp 1676037725
transform 1 0 43148 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_465
timestamp 1676037725
transform 1 0 43884 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_470
timestamp 1676037725
transform 1 0 44344 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_477
timestamp 1676037725
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_489
timestamp 1676037725
transform 1 0 46092 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_501
timestamp 1676037725
transform 1 0 47196 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_513
timestamp 1676037725
transform 1 0 48300 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_525
timestamp 1676037725
transform 1 0 49404 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1676037725
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_21
timestamp 1676037725
transform 1 0 3036 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_33
timestamp 1676037725
transform 1 0 4140 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_45
timestamp 1676037725
transform 1 0 5244 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1676037725
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1676037725
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1676037725
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1676037725
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1676037725
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1676037725
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1676037725
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1676037725
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1676037725
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1676037725
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1676037725
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1676037725
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1676037725
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1676037725
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1676037725
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1676037725
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_205
timestamp 1676037725
transform 1 0 19964 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1676037725
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1676037725
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_237
timestamp 1676037725
transform 1 0 22908 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_259
timestamp 1676037725
transform 1 0 24932 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_267
timestamp 1676037725
transform 1 0 25668 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1676037725
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1676037725
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1676037725
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_305
timestamp 1676037725
transform 1 0 29164 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_313
timestamp 1676037725
transform 1 0 29900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_323
timestamp 1676037725
transform 1 0 30820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1676037725
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_33_337
timestamp 1676037725
transform 1 0 32108 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1676037725
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1676037725
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1676037725
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_385
timestamp 1676037725
transform 1 0 36524 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_390
timestamp 1676037725
transform 1 0 36984 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1676037725
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_405
timestamp 1676037725
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_417
timestamp 1676037725
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_429
timestamp 1676037725
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1676037725
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1676037725
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_449
timestamp 1676037725
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_461
timestamp 1676037725
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_473
timestamp 1676037725
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_485
timestamp 1676037725
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1676037725
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1676037725
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_505
timestamp 1676037725
transform 1 0 47564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_525
timestamp 1676037725
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1676037725
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1676037725
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1676037725
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_34_29
timestamp 1676037725
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_36
timestamp 1676037725
transform 1 0 4416 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_48
timestamp 1676037725
transform 1 0 5520 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_60
timestamp 1676037725
transform 1 0 6624 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_72
timestamp 1676037725
transform 1 0 7728 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_85
timestamp 1676037725
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_95
timestamp 1676037725
transform 1 0 9844 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_107
timestamp 1676037725
transform 1 0 10948 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_119
timestamp 1676037725
transform 1 0 12052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_131
timestamp 1676037725
transform 1 0 13156 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1676037725
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1676037725
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1676037725
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1676037725
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1676037725
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1676037725
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1676037725
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1676037725
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1676037725
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1676037725
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1676037725
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1676037725
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1676037725
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1676037725
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1676037725
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1676037725
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1676037725
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1676037725
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1676037725
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1676037725
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_326
timestamp 1676037725
transform 1 0 31096 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_333
timestamp 1676037725
transform 1 0 31740 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_340
timestamp 1676037725
transform 1 0 32384 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_352
timestamp 1676037725
transform 1 0 33488 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1676037725
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_377
timestamp 1676037725
transform 1 0 35788 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_385
timestamp 1676037725
transform 1 0 36524 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_389
timestamp 1676037725
transform 1 0 36892 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_397
timestamp 1676037725
transform 1 0 37628 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_408
timestamp 1676037725
transform 1 0 38640 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_421
timestamp 1676037725
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_433
timestamp 1676037725
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_445
timestamp 1676037725
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_457
timestamp 1676037725
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1676037725
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1676037725
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_477
timestamp 1676037725
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_489
timestamp 1676037725
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_501
timestamp 1676037725
transform 1 0 47196 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_525
timestamp 1676037725
transform 1 0 49404 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1676037725
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1676037725
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1676037725
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1676037725
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1676037725
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1676037725
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1676037725
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1676037725
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_81
timestamp 1676037725
transform 1 0 8556 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_89
timestamp 1676037725
transform 1 0 9292 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_100
timestamp 1676037725
transform 1 0 10304 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1676037725
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1676037725
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_137
timestamp 1676037725
transform 1 0 13708 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_146
timestamp 1676037725
transform 1 0 14536 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_158
timestamp 1676037725
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_166
timestamp 1676037725
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1676037725
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1676037725
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_193
timestamp 1676037725
transform 1 0 18860 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_208
timestamp 1676037725
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_212
timestamp 1676037725
transform 1 0 20608 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1676037725
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_225
timestamp 1676037725
transform 1 0 21804 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_231
timestamp 1676037725
transform 1 0 22356 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_253
timestamp 1676037725
transform 1 0 24380 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_270
timestamp 1676037725
transform 1 0 25944 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1676037725
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_281
timestamp 1676037725
transform 1 0 26956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_289
timestamp 1676037725
transform 1 0 27692 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_295
timestamp 1676037725
transform 1 0 28244 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_308
timestamp 1676037725
transform 1 0 29440 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1676037725
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_337
timestamp 1676037725
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_361
timestamp 1676037725
transform 1 0 34316 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_369
timestamp 1676037725
transform 1 0 35052 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_373
timestamp 1676037725
transform 1 0 35420 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_380
timestamp 1676037725
transform 1 0 36064 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1676037725
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_405
timestamp 1676037725
transform 1 0 38364 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_426
timestamp 1676037725
transform 1 0 40296 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_438
timestamp 1676037725
transform 1 0 41400 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_446
timestamp 1676037725
transform 1 0 42136 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_449
timestamp 1676037725
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_461
timestamp 1676037725
transform 1 0 43516 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_35_467
timestamp 1676037725
transform 1 0 44068 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_479
timestamp 1676037725
transform 1 0 45172 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_491
timestamp 1676037725
transform 1 0 46276 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1676037725
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1676037725
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_35_525
timestamp 1676037725
transform 1 0 49404 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1676037725
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1676037725
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1676037725
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1676037725
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_41
timestamp 1676037725
transform 1 0 4876 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_49
timestamp 1676037725
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_61
timestamp 1676037725
transform 1 0 6716 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1676037725
transform 1 0 7820 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_81
timestamp 1676037725
transform 1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1676037725
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1676037725
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1676037725
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_121
timestamp 1676037725
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_130
timestamp 1676037725
transform 1 0 13064 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_137
timestamp 1676037725
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_141
timestamp 1676037725
transform 1 0 14076 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_147
timestamp 1676037725
transform 1 0 14628 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_168
timestamp 1676037725
transform 1 0 16560 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_180
timestamp 1676037725
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1676037725
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_197
timestamp 1676037725
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_219
timestamp 1676037725
transform 1 0 21252 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_227
timestamp 1676037725
transform 1 0 21988 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1676037725
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1676037725
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_253
timestamp 1676037725
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_259
timestamp 1676037725
transform 1 0 24932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_262
timestamp 1676037725
transform 1 0 25208 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_275
timestamp 1676037725
transform 1 0 26404 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_287
timestamp 1676037725
transform 1 0 27508 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_295
timestamp 1676037725
transform 1 0 28244 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1676037725
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_309
timestamp 1676037725
transform 1 0 29532 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_314
timestamp 1676037725
transform 1 0 29992 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_326
timestamp 1676037725
transform 1 0 31096 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_338
timestamp 1676037725
transform 1 0 32200 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_350
timestamp 1676037725
transform 1 0 33304 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1676037725
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_365
timestamp 1676037725
transform 1 0 34684 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_371
timestamp 1676037725
transform 1 0 35236 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_393
timestamp 1676037725
transform 1 0 37260 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_400
timestamp 1676037725
transform 1 0 37904 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_412
timestamp 1676037725
transform 1 0 39008 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_421
timestamp 1676037725
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_433
timestamp 1676037725
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_445
timestamp 1676037725
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_457
timestamp 1676037725
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1676037725
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1676037725
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_477
timestamp 1676037725
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_489
timestamp 1676037725
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_501
timestamp 1676037725
transform 1 0 47196 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_525
timestamp 1676037725
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1676037725
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1676037725
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1676037725
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1676037725
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1676037725
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1676037725
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1676037725
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1676037725
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1676037725
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1676037725
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1676037725
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1676037725
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1676037725
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1676037725
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1676037725
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1676037725
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1676037725
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1676037725
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1676037725
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_186
timestamp 1676037725
transform 1 0 18216 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_207
timestamp 1676037725
transform 1 0 20148 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_222
timestamp 1676037725
transform 1 0 21528 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1676037725
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1676037725
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_250
timestamp 1676037725
transform 1 0 24104 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_254
timestamp 1676037725
transform 1 0 24472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_264
timestamp 1676037725
transform 1 0 25392 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_271
timestamp 1676037725
transform 1 0 26036 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1676037725
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_281
timestamp 1676037725
transform 1 0 26956 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_303
timestamp 1676037725
transform 1 0 28980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_309
timestamp 1676037725
transform 1 0 29532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_319
timestamp 1676037725
transform 1 0 30452 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_37_334
timestamp 1676037725
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1676037725
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_342
timestamp 1676037725
transform 1 0 32568 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_363
timestamp 1676037725
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_375
timestamp 1676037725
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1676037725
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1676037725
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_393
timestamp 1676037725
transform 1 0 37260 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_420
timestamp 1676037725
transform 1 0 39744 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_432
timestamp 1676037725
transform 1 0 40848 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_444
timestamp 1676037725
transform 1 0 41952 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_449
timestamp 1676037725
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_461
timestamp 1676037725
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_473
timestamp 1676037725
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_485
timestamp 1676037725
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1676037725
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1676037725
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_505
timestamp 1676037725
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_517
timestamp 1676037725
transform 1 0 48668 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_525
timestamp 1676037725
transform 1 0 49404 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1676037725
transform 1 0 1380 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_21
timestamp 1676037725
transform 1 0 3036 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1676037725
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_38_29
timestamp 1676037725
transform 1 0 3772 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_36
timestamp 1676037725
transform 1 0 4416 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_38_46
timestamp 1676037725
transform 1 0 5336 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_58
timestamp 1676037725
transform 1 0 6440 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_70
timestamp 1676037725
transform 1 0 7544 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_82
timestamp 1676037725
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_85
timestamp 1676037725
transform 1 0 8924 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_90
timestamp 1676037725
transform 1 0 9384 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_102
timestamp 1676037725
transform 1 0 10488 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_114
timestamp 1676037725
transform 1 0 11592 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_126
timestamp 1676037725
transform 1 0 12696 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1676037725
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1676037725
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1676037725
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_165
timestamp 1676037725
transform 1 0 16284 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_173
timestamp 1676037725
transform 1 0 17020 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_194
timestamp 1676037725
transform 1 0 18952 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1676037725
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_219
timestamp 1676037725
transform 1 0 21252 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_231
timestamp 1676037725
transform 1 0 22356 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_234
timestamp 1676037725
transform 1 0 22632 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1676037725
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1676037725
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_253
timestamp 1676037725
transform 1 0 24380 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_264
timestamp 1676037725
transform 1 0 25392 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_276
timestamp 1676037725
transform 1 0 26496 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_282
timestamp 1676037725
transform 1 0 27048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1676037725
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1676037725
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_309
timestamp 1676037725
transform 1 0 29532 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_335
timestamp 1676037725
transform 1 0 31924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_359
timestamp 1676037725
transform 1 0 34132 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1676037725
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1676037725
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_387
timestamp 1676037725
transform 1 0 36708 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_398
timestamp 1676037725
transform 1 0 37720 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_402
timestamp 1676037725
transform 1 0 38088 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_412
timestamp 1676037725
transform 1 0 39008 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_421
timestamp 1676037725
transform 1 0 39836 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_426
timestamp 1676037725
transform 1 0 40296 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_438
timestamp 1676037725
transform 1 0 41400 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_450
timestamp 1676037725
transform 1 0 42504 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_462
timestamp 1676037725
transform 1 0 43608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_466
timestamp 1676037725
transform 1 0 43976 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_471
timestamp 1676037725
transform 1 0 44436 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1676037725
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_477
timestamp 1676037725
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_489
timestamp 1676037725
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_501
timestamp 1676037725
transform 1 0 47196 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_525
timestamp 1676037725
transform 1 0 49404 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1676037725
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1676037725
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1676037725
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1676037725
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1676037725
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1676037725
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1676037725
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1676037725
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_81
timestamp 1676037725
transform 1 0 8556 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_91
timestamp 1676037725
transform 1 0 9476 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_103
timestamp 1676037725
transform 1 0 10580 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1676037725
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1676037725
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_125
timestamp 1676037725
transform 1 0 12604 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_39_148
timestamp 1676037725
transform 1 0 14720 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_160
timestamp 1676037725
transform 1 0 15824 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1676037725
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1676037725
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_193
timestamp 1676037725
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_197
timestamp 1676037725
transform 1 0 19228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_207
timestamp 1676037725
transform 1 0 20148 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1676037725
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1676037725
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_250
timestamp 1676037725
transform 1 0 24104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_254
timestamp 1676037725
transform 1 0 24472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_258
timestamp 1676037725
transform 1 0 24840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_265
timestamp 1676037725
transform 1 0 25484 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_278
timestamp 1676037725
transform 1 0 26680 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1676037725
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_293
timestamp 1676037725
transform 1 0 28060 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_304
timestamp 1676037725
transform 1 0 29072 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_316
timestamp 1676037725
transform 1 0 30176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_328
timestamp 1676037725
transform 1 0 31280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_337
timestamp 1676037725
transform 1 0 32108 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_359
timestamp 1676037725
transform 1 0 34132 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_372
timestamp 1676037725
transform 1 0 35328 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_384
timestamp 1676037725
transform 1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1676037725
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_405
timestamp 1676037725
transform 1 0 38364 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_429
timestamp 1676037725
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1676037725
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1676037725
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_449
timestamp 1676037725
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_461
timestamp 1676037725
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_473
timestamp 1676037725
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_485
timestamp 1676037725
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1676037725
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1676037725
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_505
timestamp 1676037725
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_39_525
timestamp 1676037725
transform 1 0 49404 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1676037725
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1676037725
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1676037725
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1676037725
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1676037725
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1676037725
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1676037725
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1676037725
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1676037725
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1676037725
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_97
timestamp 1676037725
transform 1 0 10028 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1676037725
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1676037725
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1676037725
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1676037725
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_141
timestamp 1676037725
transform 1 0 14076 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_40_167
timestamp 1676037725
transform 1 0 16468 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_179
timestamp 1676037725
transform 1 0 17572 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1676037725
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1676037725
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1676037725
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1676037725
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1676037725
transform 1 0 20700 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_234
timestamp 1676037725
transform 1 0 22632 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_246
timestamp 1676037725
transform 1 0 23736 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_253
timestamp 1676037725
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_259
timestamp 1676037725
transform 1 0 24932 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_269
timestamp 1676037725
transform 1 0 25852 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_284
timestamp 1676037725
transform 1 0 27232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_297
timestamp 1676037725
transform 1 0 28428 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_305
timestamp 1676037725
transform 1 0 29164 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1676037725
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_320
timestamp 1676037725
transform 1 0 30544 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_332
timestamp 1676037725
transform 1 0 31648 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_344
timestamp 1676037725
transform 1 0 32752 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_352
timestamp 1676037725
transform 1 0 33488 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_362
timestamp 1676037725
transform 1 0 34408 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_365
timestamp 1676037725
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_388
timestamp 1676037725
transform 1 0 36800 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_401
timestamp 1676037725
transform 1 0 37996 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_413
timestamp 1676037725
transform 1 0 39100 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_419
timestamp 1676037725
transform 1 0 39652 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_421
timestamp 1676037725
transform 1 0 39836 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_432
timestamp 1676037725
transform 1 0 40848 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_444
timestamp 1676037725
transform 1 0 41952 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_456
timestamp 1676037725
transform 1 0 43056 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_468
timestamp 1676037725
transform 1 0 44160 0 1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_40_477
timestamp 1676037725
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_489
timestamp 1676037725
transform 1 0 46092 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_501
timestamp 1676037725
transform 1 0 47196 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_525
timestamp 1676037725
transform 1 0 49404 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1676037725
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1676037725
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1676037725
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1676037725
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1676037725
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1676037725
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1676037725
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_69
timestamp 1676037725
transform 1 0 7452 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_77
timestamp 1676037725
transform 1 0 8188 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_82
timestamp 1676037725
transform 1 0 8648 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_94
timestamp 1676037725
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1676037725
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1676037725
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1676037725
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1676037725
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1676037725
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1676037725
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1676037725
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1676037725
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1676037725
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_193
timestamp 1676037725
transform 1 0 18860 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_201
timestamp 1676037725
transform 1 0 19596 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_222
timestamp 1676037725
transform 1 0 21528 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1676037725
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1676037725
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1676037725
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_261
timestamp 1676037725
transform 1 0 25116 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_273
timestamp 1676037725
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1676037725
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1676037725
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_303
timestamp 1676037725
transform 1 0 28980 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_327
timestamp 1676037725
transform 1 0 31188 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1676037725
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_337
timestamp 1676037725
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_349
timestamp 1676037725
transform 1 0 33212 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_380
timestamp 1676037725
transform 1 0 36064 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1676037725
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_404
timestamp 1676037725
transform 1 0 38272 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_416
timestamp 1676037725
transform 1 0 39376 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_422
timestamp 1676037725
transform 1 0 39928 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_426
timestamp 1676037725
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_438
timestamp 1676037725
transform 1 0 41400 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_446
timestamp 1676037725
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_449
timestamp 1676037725
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_461
timestamp 1676037725
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_473
timestamp 1676037725
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_485
timestamp 1676037725
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_497
timestamp 1676037725
transform 1 0 46828 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1676037725
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_505
timestamp 1676037725
transform 1 0 47564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_525
timestamp 1676037725
transform 1 0 49404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_3
timestamp 1676037725
transform 1 0 1380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_21
timestamp 1676037725
transform 1 0 3036 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1676037725
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1676037725
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_44
timestamp 1676037725
transform 1 0 5152 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_56
timestamp 1676037725
transform 1 0 6256 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_68
timestamp 1676037725
transform 1 0 7360 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1676037725
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1676037725
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_97
timestamp 1676037725
transform 1 0 10028 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1676037725
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1676037725
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1676037725
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1676037725
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1676037725
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_146
timestamp 1676037725
transform 1 0 14536 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_158
timestamp 1676037725
transform 1 0 15640 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_170
timestamp 1676037725
transform 1 0 16744 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_182
timestamp 1676037725
transform 1 0 17848 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1676037725
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1676037725
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1676037725
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_221
timestamp 1676037725
transform 1 0 21436 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_229
timestamp 1676037725
transform 1 0 22172 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_239
timestamp 1676037725
transform 1 0 23092 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1676037725
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1676037725
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_264
timestamp 1676037725
transform 1 0 25392 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_290
timestamp 1676037725
transform 1 0 27784 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1676037725
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_309
timestamp 1676037725
transform 1 0 29532 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_314
timestamp 1676037725
transform 1 0 29992 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_331
timestamp 1676037725
transform 1 0 31556 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_344
timestamp 1676037725
transform 1 0 32752 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_361
timestamp 1676037725
transform 1 0 34316 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_365
timestamp 1676037725
transform 1 0 34684 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_369
timestamp 1676037725
transform 1 0 35052 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_379
timestamp 1676037725
transform 1 0 35972 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_394
timestamp 1676037725
transform 1 0 37352 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_418
timestamp 1676037725
transform 1 0 39560 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_421
timestamp 1676037725
transform 1 0 39836 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_432
timestamp 1676037725
transform 1 0 40848 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_444
timestamp 1676037725
transform 1 0 41952 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_456
timestamp 1676037725
transform 1 0 43056 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_468
timestamp 1676037725
transform 1 0 44160 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_473
timestamp 1676037725
transform 1 0 44620 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_477
timestamp 1676037725
transform 1 0 44988 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_483
timestamp 1676037725
transform 1 0 45540 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_491
timestamp 1676037725
transform 1 0 46276 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_503
timestamp 1676037725
transform 1 0 47380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_515
timestamp 1676037725
transform 1 0 48484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1676037725
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1676037725
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1676037725
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1676037725
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1676037725
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1676037725
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1676037725
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1676037725
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_92
timestamp 1676037725
transform 1 0 9568 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_104
timestamp 1676037725
transform 1 0 10672 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1676037725
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1676037725
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1676037725
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1676037725
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1676037725
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1676037725
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1676037725
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1676037725
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1676037725
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1676037725
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1676037725
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1676037725
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1676037725
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_233
timestamp 1676037725
transform 1 0 22540 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_237
timestamp 1676037725
transform 1 0 22908 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_245
timestamp 1676037725
transform 1 0 23644 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_255
timestamp 1676037725
transform 1 0 24564 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_262
timestamp 1676037725
transform 1 0 25208 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_271
timestamp 1676037725
transform 1 0 26036 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1676037725
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_281
timestamp 1676037725
transform 1 0 26956 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_292
timestamp 1676037725
transform 1 0 27968 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_316
timestamp 1676037725
transform 1 0 30176 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_333
timestamp 1676037725
transform 1 0 31740 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1676037725
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_348
timestamp 1676037725
transform 1 0 33120 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_360
timestamp 1676037725
transform 1 0 34224 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_366
timestamp 1676037725
transform 1 0 34776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_376
timestamp 1676037725
transform 1 0 35696 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_383
timestamp 1676037725
transform 1 0 36340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1676037725
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1676037725
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_408
timestamp 1676037725
transform 1 0 38640 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_421
timestamp 1676037725
transform 1 0 39836 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_425
timestamp 1676037725
transform 1 0 40204 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1676037725
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_449
timestamp 1676037725
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_461
timestamp 1676037725
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_473
timestamp 1676037725
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_485
timestamp 1676037725
transform 1 0 45724 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_491
timestamp 1676037725
transform 1 0 46276 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_499
timestamp 1676037725
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1676037725
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_505
timestamp 1676037725
transform 1 0 47564 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_517
timestamp 1676037725
transform 1 0 48668 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_521
timestamp 1676037725
transform 1 0 49036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_525
timestamp 1676037725
transform 1 0 49404 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1676037725
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1676037725
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1676037725
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1676037725
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1676037725
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1676037725
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_65
timestamp 1676037725
transform 1 0 7084 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_71
timestamp 1676037725
transform 1 0 7636 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_75
timestamp 1676037725
transform 1 0 8004 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1676037725
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_85
timestamp 1676037725
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_95
timestamp 1676037725
transform 1 0 9844 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_107
timestamp 1676037725
transform 1 0 10948 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_119
timestamp 1676037725
transform 1 0 12052 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_131
timestamp 1676037725
transform 1 0 13156 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1676037725
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1676037725
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1676037725
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1676037725
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1676037725
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1676037725
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1676037725
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1676037725
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1676037725
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_221
timestamp 1676037725
transform 1 0 21436 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_227
timestamp 1676037725
transform 1 0 21988 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1676037725
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_253
timestamp 1676037725
transform 1 0 24380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_44_264
timestamp 1676037725
transform 1 0 25392 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_270
timestamp 1676037725
transform 1 0 25944 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1676037725
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_295
timestamp 1676037725
transform 1 0 28244 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1676037725
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1676037725
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_330
timestamp 1676037725
transform 1 0 31464 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_336
timestamp 1676037725
transform 1 0 32016 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1676037725
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1676037725
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1676037725
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_378
timestamp 1676037725
transform 1 0 35880 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_390
timestamp 1676037725
transform 1 0 36984 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_403
timestamp 1676037725
transform 1 0 38180 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_415
timestamp 1676037725
transform 1 0 39284 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1676037725
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_421
timestamp 1676037725
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_444
timestamp 1676037725
transform 1 0 41952 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_456
timestamp 1676037725
transform 1 0 43056 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_468
timestamp 1676037725
transform 1 0 44160 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_44_477
timestamp 1676037725
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_489
timestamp 1676037725
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_504
timestamp 1676037725
transform 1 0 47472 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_508
timestamp 1676037725
transform 1 0 47840 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_511
timestamp 1676037725
transform 1 0 48116 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_525
timestamp 1676037725
transform 1 0 49404 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1676037725
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1676037725
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1676037725
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1676037725
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1676037725
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1676037725
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1676037725
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1676037725
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_94
timestamp 1676037725
transform 1 0 9752 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_106
timestamp 1676037725
transform 1 0 10856 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1676037725
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1676037725
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1676037725
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1676037725
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1676037725
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1676037725
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1676037725
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1676037725
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1676037725
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1676037725
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1676037725
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1676037725
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1676037725
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1676037725
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_244
timestamp 1676037725
transform 1 0 23552 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_248
timestamp 1676037725
transform 1 0 23920 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1676037725
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_265
timestamp 1676037725
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1676037725
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1676037725
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_294
timestamp 1676037725
transform 1 0 28152 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_318
timestamp 1676037725
transform 1 0 30360 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_331
timestamp 1676037725
transform 1 0 31556 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1676037725
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_337
timestamp 1676037725
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_345
timestamp 1676037725
transform 1 0 32844 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_355
timestamp 1676037725
transform 1 0 33764 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_380
timestamp 1676037725
transform 1 0 36064 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_386
timestamp 1676037725
transform 1 0 36616 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_390
timestamp 1676037725
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1676037725
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_406
timestamp 1676037725
transform 1 0 38456 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_418
timestamp 1676037725
transform 1 0 39560 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1676037725
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_449
timestamp 1676037725
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_461
timestamp 1676037725
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_473
timestamp 1676037725
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_485
timestamp 1676037725
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_500
timestamp 1676037725
transform 1 0 47104 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_505
timestamp 1676037725
transform 1 0 47564 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_511
timestamp 1676037725
transform 1 0 48116 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_525
timestamp 1676037725
transform 1 0 49404 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1676037725
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_21
timestamp 1676037725
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1676037725
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1676037725
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1676037725
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1676037725
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_65
timestamp 1676037725
transform 1 0 7084 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_46_74
timestamp 1676037725
transform 1 0 7912 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_82
timestamp 1676037725
transform 1 0 8648 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1676037725
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1676037725
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1676037725
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1676037725
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1676037725
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1676037725
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1676037725
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1676037725
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1676037725
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1676037725
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1676037725
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1676037725
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1676037725
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1676037725
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1676037725
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_233
timestamp 1676037725
transform 1 0 22540 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_239
timestamp 1676037725
transform 1 0 23092 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_243
timestamp 1676037725
transform 1 0 23460 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1676037725
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_253
timestamp 1676037725
transform 1 0 24380 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_257
timestamp 1676037725
transform 1 0 24748 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_278
timestamp 1676037725
transform 1 0 26680 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_286
timestamp 1676037725
transform 1 0 27416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_298
timestamp 1676037725
transform 1 0 28520 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1676037725
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_309
timestamp 1676037725
transform 1 0 29532 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_315
timestamp 1676037725
transform 1 0 30084 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_325
timestamp 1676037725
transform 1 0 31004 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_331
timestamp 1676037725
transform 1 0 31556 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_341
timestamp 1676037725
transform 1 0 32476 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_356
timestamp 1676037725
transform 1 0 33856 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1676037725
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_376
timestamp 1676037725
transform 1 0 35696 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_388
timestamp 1676037725
transform 1 0 36800 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_409
timestamp 1676037725
transform 1 0 38732 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_417
timestamp 1676037725
transform 1 0 39468 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_421
timestamp 1676037725
transform 1 0 39836 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_46_444
timestamp 1676037725
transform 1 0 41952 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_456
timestamp 1676037725
transform 1 0 43056 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_46_467
timestamp 1676037725
transform 1 0 44068 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1676037725
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_477
timestamp 1676037725
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_489
timestamp 1676037725
transform 1 0 46092 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_497
timestamp 1676037725
transform 1 0 46828 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_504
timestamp 1676037725
transform 1 0 47472 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_512
timestamp 1676037725
transform 1 0 48208 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_525
timestamp 1676037725
transform 1 0 49404 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1676037725
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1676037725
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1676037725
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_39
timestamp 1676037725
transform 1 0 4692 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1676037725
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1676037725
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_69
timestamp 1676037725
transform 1 0 7452 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_91
timestamp 1676037725
transform 1 0 9476 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_103
timestamp 1676037725
transform 1 0 10580 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1676037725
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1676037725
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1676037725
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1676037725
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1676037725
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1676037725
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1676037725
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1676037725
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1676037725
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1676037725
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1676037725
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1676037725
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1676037725
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1676037725
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_251
timestamp 1676037725
transform 1 0 24196 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_275
timestamp 1676037725
transform 1 0 26404 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1676037725
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_281
timestamp 1676037725
transform 1 0 26956 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_289
timestamp 1676037725
transform 1 0 27692 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_311
timestamp 1676037725
transform 1 0 29716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1676037725
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1676037725
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_47_359
timestamp 1676037725
transform 1 0 34132 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_371
timestamp 1676037725
transform 1 0 35236 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1676037725
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_393
timestamp 1676037725
transform 1 0 37260 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_408
timestamp 1676037725
transform 1 0 38640 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_421
timestamp 1676037725
transform 1 0 39836 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_433
timestamp 1676037725
transform 1 0 40940 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_445
timestamp 1676037725
transform 1 0 42044 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_47_449
timestamp 1676037725
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_461
timestamp 1676037725
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_473
timestamp 1676037725
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_485
timestamp 1676037725
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1676037725
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1676037725
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_505
timestamp 1676037725
transform 1 0 47564 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_509
timestamp 1676037725
transform 1 0 47932 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_514
timestamp 1676037725
transform 1 0 48392 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_526
timestamp 1676037725
transform 1 0 49496 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1676037725
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1676037725
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1676037725
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1676037725
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1676037725
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1676037725
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1676037725
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1676037725
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1676037725
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1676037725
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1676037725
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1676037725
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1676037725
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1676037725
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1676037725
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1676037725
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1676037725
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1676037725
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1676037725
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1676037725
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1676037725
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1676037725
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_209
timestamp 1676037725
transform 1 0 20332 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_215
timestamp 1676037725
transform 1 0 20884 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_227
timestamp 1676037725
transform 1 0 21988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_233
timestamp 1676037725
transform 1 0 22540 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_246
timestamp 1676037725
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1676037725
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1676037725
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_277
timestamp 1676037725
transform 1 0 26588 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_281
timestamp 1676037725
transform 1 0 26956 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_302
timestamp 1676037725
transform 1 0 28888 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_309
timestamp 1676037725
transform 1 0 29532 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_314
timestamp 1676037725
transform 1 0 29992 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_320
timestamp 1676037725
transform 1 0 30544 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_330
timestamp 1676037725
transform 1 0 31464 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_342
timestamp 1676037725
transform 1 0 32568 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_350
timestamp 1676037725
transform 1 0 33304 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1676037725
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1676037725
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_376
timestamp 1676037725
transform 1 0 35696 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_398
timestamp 1676037725
transform 1 0 37720 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_404
timestamp 1676037725
transform 1 0 38272 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_417
timestamp 1676037725
transform 1 0 39468 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_421
timestamp 1676037725
transform 1 0 39836 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_432
timestamp 1676037725
transform 1 0 40848 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_444
timestamp 1676037725
transform 1 0 41952 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_456
timestamp 1676037725
transform 1 0 43056 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_468
timestamp 1676037725
transform 1 0 44160 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_48_477
timestamp 1676037725
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_489
timestamp 1676037725
transform 1 0 46092 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_501
timestamp 1676037725
transform 1 0 47196 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_513
timestamp 1676037725
transform 1 0 48300 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_521
timestamp 1676037725
transform 1 0 49036 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_525
timestamp 1676037725
transform 1 0 49404 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1676037725
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1676037725
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1676037725
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1676037725
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1676037725
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1676037725
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1676037725
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1676037725
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1676037725
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1676037725
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1676037725
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1676037725
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1676037725
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1676037725
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1676037725
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1676037725
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1676037725
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1676037725
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1676037725
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1676037725
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1676037725
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1676037725
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_217
timestamp 1676037725
transform 1 0 21068 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_220
timestamp 1676037725
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_225
timestamp 1676037725
transform 1 0 21804 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_236
timestamp 1676037725
transform 1 0 22816 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_242
timestamp 1676037725
transform 1 0 23368 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_254
timestamp 1676037725
transform 1 0 24472 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_266
timestamp 1676037725
transform 1 0 25576 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1676037725
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1676037725
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_309
timestamp 1676037725
transform 1 0 29532 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_322
timestamp 1676037725
transform 1 0 30728 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1676037725
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1676037725
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_349
timestamp 1676037725
transform 1 0 33212 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_377
timestamp 1676037725
transform 1 0 35788 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1676037725
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1676037725
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_405
timestamp 1676037725
transform 1 0 38364 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_409
timestamp 1676037725
transform 1 0 38732 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_424
timestamp 1676037725
transform 1 0 40112 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_430
timestamp 1676037725
transform 1 0 40664 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_440
timestamp 1676037725
transform 1 0 41584 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_449
timestamp 1676037725
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_461
timestamp 1676037725
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_473
timestamp 1676037725
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_485
timestamp 1676037725
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_497
timestamp 1676037725
transform 1 0 46828 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_503
timestamp 1676037725
transform 1 0 47380 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_505
timestamp 1676037725
transform 1 0 47564 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_517
timestamp 1676037725
transform 1 0 48668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_521
timestamp 1676037725
transform 1 0 49036 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_525
timestamp 1676037725
transform 1 0 49404 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_3
timestamp 1676037725
transform 1 0 1380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_21
timestamp 1676037725
transform 1 0 3036 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1676037725
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1676037725
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1676037725
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1676037725
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1676037725
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1676037725
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1676037725
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1676037725
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1676037725
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1676037725
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1676037725
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1676037725
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1676037725
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1676037725
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1676037725
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1676037725
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1676037725
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1676037725
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1676037725
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1676037725
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1676037725
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_221
timestamp 1676037725
transform 1 0 21436 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_229
timestamp 1676037725
transform 1 0 22172 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_243
timestamp 1676037725
transform 1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1676037725
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_253
timestamp 1676037725
transform 1 0 24380 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_261
timestamp 1676037725
transform 1 0 25116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_272
timestamp 1676037725
transform 1 0 26128 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_279
timestamp 1676037725
transform 1 0 26772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_291
timestamp 1676037725
transform 1 0 27876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_303
timestamp 1676037725
transform 1 0 28980 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1676037725
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1676037725
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_320
timestamp 1676037725
transform 1 0 30544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_332
timestamp 1676037725
transform 1 0 31648 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_344
timestamp 1676037725
transform 1 0 32752 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1676037725
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1676037725
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_377
timestamp 1676037725
transform 1 0 35788 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_403
timestamp 1676037725
transform 1 0 38180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_415
timestamp 1676037725
transform 1 0 39284 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1676037725
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_421
timestamp 1676037725
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_453
timestamp 1676037725
transform 1 0 42780 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_465
timestamp 1676037725
transform 1 0 43884 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_473
timestamp 1676037725
transform 1 0 44620 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_477
timestamp 1676037725
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_489
timestamp 1676037725
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_501
timestamp 1676037725
transform 1 0 47196 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_513
timestamp 1676037725
transform 1 0 48300 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_525
timestamp 1676037725
transform 1 0 49404 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1676037725
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1676037725
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1676037725
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1676037725
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1676037725
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1676037725
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_57
timestamp 1676037725
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_65
timestamp 1676037725
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_89
timestamp 1676037725
transform 1 0 9292 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_101
timestamp 1676037725
transform 1 0 10396 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_109
timestamp 1676037725
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1676037725
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1676037725
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1676037725
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1676037725
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1676037725
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1676037725
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1676037725
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1676037725
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1676037725
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1676037725
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1676037725
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1676037725
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1676037725
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_237
timestamp 1676037725
transform 1 0 22908 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_245
timestamp 1676037725
transform 1 0 23644 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_252
timestamp 1676037725
transform 1 0 24288 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_262
timestamp 1676037725
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_268
timestamp 1676037725
transform 1 0 25760 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_281
timestamp 1676037725
transform 1 0 26956 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_289
timestamp 1676037725
transform 1 0 27692 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_292
timestamp 1676037725
transform 1 0 27968 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1676037725
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_317
timestamp 1676037725
transform 1 0 30268 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_327
timestamp 1676037725
transform 1 0 31188 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1676037725
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1676037725
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_349
timestamp 1676037725
transform 1 0 33212 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_353
timestamp 1676037725
transform 1 0 33580 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_363
timestamp 1676037725
transform 1 0 34500 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_371
timestamp 1676037725
transform 1 0 35236 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_383
timestamp 1676037725
transform 1 0 36340 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1676037725
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1676037725
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_404
timestamp 1676037725
transform 1 0 38272 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_428
timestamp 1676037725
transform 1 0 40480 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1676037725
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1676037725
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_449
timestamp 1676037725
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_461
timestamp 1676037725
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_473
timestamp 1676037725
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_485
timestamp 1676037725
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1676037725
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1676037725
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_505
timestamp 1676037725
transform 1 0 47564 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_517
timestamp 1676037725
transform 1 0 48668 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_521
timestamp 1676037725
transform 1 0 49036 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_525
timestamp 1676037725
transform 1 0 49404 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1676037725
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1676037725
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1676037725
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1676037725
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1676037725
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1676037725
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1676037725
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1676037725
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1676037725
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1676037725
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1676037725
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1676037725
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1676037725
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1676037725
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1676037725
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1676037725
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1676037725
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1676037725
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1676037725
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1676037725
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1676037725
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1676037725
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_209
timestamp 1676037725
transform 1 0 20332 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_217
timestamp 1676037725
transform 1 0 21068 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_230
timestamp 1676037725
transform 1 0 22264 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_238
timestamp 1676037725
transform 1 0 23000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1676037725
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_253
timestamp 1676037725
transform 1 0 24380 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_257
timestamp 1676037725
transform 1 0 24748 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_278
timestamp 1676037725
transform 1 0 26680 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_302
timestamp 1676037725
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1676037725
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_320
timestamp 1676037725
transform 1 0 30544 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_348
timestamp 1676037725
transform 1 0 33120 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1676037725
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_365
timestamp 1676037725
transform 1 0 34684 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_377
timestamp 1676037725
transform 1 0 35788 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_390
timestamp 1676037725
transform 1 0 36984 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1676037725
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_407
timestamp 1676037725
transform 1 0 38548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_52_417
timestamp 1676037725
transform 1 0 39468 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_421
timestamp 1676037725
transform 1 0 39836 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_432
timestamp 1676037725
transform 1 0 40848 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_436
timestamp 1676037725
transform 1 0 41216 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_440
timestamp 1676037725
transform 1 0 41584 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_447
timestamp 1676037725
transform 1 0 42228 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_458
timestamp 1676037725
transform 1 0 43240 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_470
timestamp 1676037725
transform 1 0 44344 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_477
timestamp 1676037725
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_489
timestamp 1676037725
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_501
timestamp 1676037725
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_513
timestamp 1676037725
transform 1 0 48300 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_525
timestamp 1676037725
transform 1 0 49404 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1676037725
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1676037725
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1676037725
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1676037725
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1676037725
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1676037725
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1676037725
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1676037725
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1676037725
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1676037725
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1676037725
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1676037725
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1676037725
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1676037725
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1676037725
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1676037725
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1676037725
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1676037725
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1676037725
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1676037725
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1676037725
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1676037725
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_217
timestamp 1676037725
transform 1 0 21068 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1676037725
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1676037725
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_236
timestamp 1676037725
transform 1 0 22816 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_242
timestamp 1676037725
transform 1 0 23368 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_252
timestamp 1676037725
transform 1 0 24288 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_278
timestamp 1676037725
transform 1 0 26680 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1676037725
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1676037725
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1676037725
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1676037725
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1676037725
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1676037725
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_337
timestamp 1676037725
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_345
timestamp 1676037725
transform 1 0 32844 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_355
timestamp 1676037725
transform 1 0 33764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_361
timestamp 1676037725
transform 1 0 34316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_382
timestamp 1676037725
transform 1 0 36248 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1676037725
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_393
timestamp 1676037725
transform 1 0 37260 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_399
timestamp 1676037725
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_412
timestamp 1676037725
transform 1 0 39008 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_424
timestamp 1676037725
transform 1 0 40112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_428
timestamp 1676037725
transform 1 0 40480 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_432
timestamp 1676037725
transform 1 0 40848 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_444
timestamp 1676037725
transform 1 0 41952 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_449
timestamp 1676037725
transform 1 0 42412 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_460
timestamp 1676037725
transform 1 0 43424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_472
timestamp 1676037725
transform 1 0 44528 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_480
timestamp 1676037725
transform 1 0 45264 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_484
timestamp 1676037725
transform 1 0 45632 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_496
timestamp 1676037725
transform 1 0 46736 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1676037725
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_513
timestamp 1676037725
transform 1 0 48300 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_525
timestamp 1676037725
transform 1 0 49404 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1676037725
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1676037725
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1676037725
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1676037725
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1676037725
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1676037725
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1676037725
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1676037725
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1676037725
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1676037725
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1676037725
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1676037725
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1676037725
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1676037725
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1676037725
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1676037725
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1676037725
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1676037725
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1676037725
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1676037725
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1676037725
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1676037725
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1676037725
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_221
timestamp 1676037725
transform 1 0 21436 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1676037725
transform 1 0 21896 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_250
timestamp 1676037725
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1676037725
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_258
timestamp 1676037725
transform 1 0 24840 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_266
timestamp 1676037725
transform 1 0 25576 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_291
timestamp 1676037725
transform 1 0 27876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_306
timestamp 1676037725
transform 1 0 29256 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1676037725
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1676037725
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_335
timestamp 1676037725
transform 1 0 31924 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_348
timestamp 1676037725
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1676037725
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1676037725
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_371
timestamp 1676037725
transform 1 0 35236 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_381
timestamp 1676037725
transform 1 0 36156 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_393
timestamp 1676037725
transform 1 0 37260 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_399
timestamp 1676037725
transform 1 0 37812 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_409
timestamp 1676037725
transform 1 0 38732 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1676037725
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_421
timestamp 1676037725
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_433
timestamp 1676037725
transform 1 0 40940 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_441
timestamp 1676037725
transform 1 0 41676 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_464
timestamp 1676037725
transform 1 0 43792 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_477
timestamp 1676037725
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_489
timestamp 1676037725
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_501
timestamp 1676037725
transform 1 0 47196 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_511
timestamp 1676037725
transform 1 0 48116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_525
timestamp 1676037725
transform 1 0 49404 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_3
timestamp 1676037725
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_8
timestamp 1676037725
transform 1 0 1840 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_20
timestamp 1676037725
transform 1 0 2944 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_32
timestamp 1676037725
transform 1 0 4048 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_44
timestamp 1676037725
transform 1 0 5152 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1676037725
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1676037725
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1676037725
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1676037725
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1676037725
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1676037725
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1676037725
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1676037725
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1676037725
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1676037725
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1676037725
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1676037725
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_169
timestamp 1676037725
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_184
timestamp 1676037725
transform 1 0 18032 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1676037725
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1676037725
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1676037725
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1676037725
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1676037725
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_237
timestamp 1676037725
transform 1 0 22908 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_245
timestamp 1676037725
transform 1 0 23644 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_268
timestamp 1676037725
transform 1 0 25760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_281
timestamp 1676037725
transform 1 0 26956 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_293
timestamp 1676037725
transform 1 0 28060 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_302
timestamp 1676037725
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_314
timestamp 1676037725
transform 1 0 29992 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1676037725
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1676037725
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_337
timestamp 1676037725
transform 1 0 32108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_361
timestamp 1676037725
transform 1 0 34316 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1676037725
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1676037725
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1676037725
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_405
timestamp 1676037725
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_437
timestamp 1676037725
transform 1 0 41308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_445
timestamp 1676037725
transform 1 0 42044 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_449
timestamp 1676037725
transform 1 0 42412 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_454
timestamp 1676037725
transform 1 0 42872 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_466
timestamp 1676037725
transform 1 0 43976 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_472
timestamp 1676037725
transform 1 0 44528 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_476
timestamp 1676037725
transform 1 0 44896 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_488
timestamp 1676037725
transform 1 0 46000 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_500
timestamp 1676037725
transform 1 0 47104 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1676037725
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_513
timestamp 1676037725
transform 1 0 48300 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_525
timestamp 1676037725
transform 1 0 49404 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1676037725
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1676037725
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1676037725
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1676037725
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1676037725
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1676037725
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1676037725
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1676037725
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1676037725
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1676037725
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1676037725
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1676037725
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1676037725
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1676037725
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1676037725
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1676037725
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1676037725
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1676037725
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1676037725
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1676037725
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1676037725
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1676037725
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1676037725
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_221
timestamp 1676037725
transform 1 0 21436 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_229
timestamp 1676037725
transform 1 0 22172 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1676037725
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1676037725
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_265
timestamp 1676037725
transform 1 0 25484 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_273
timestamp 1676037725
transform 1 0 26220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_286
timestamp 1676037725
transform 1 0 27416 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_294
timestamp 1676037725
transform 1 0 28152 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1676037725
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_309
timestamp 1676037725
transform 1 0 29532 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_320
timestamp 1676037725
transform 1 0 30544 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1676037725
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1676037725
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_357
timestamp 1676037725
transform 1 0 33948 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1676037725
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_376
timestamp 1676037725
transform 1 0 35696 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_398
timestamp 1676037725
transform 1 0 37720 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_404
timestamp 1676037725
transform 1 0 38272 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_414
timestamp 1676037725
transform 1 0 39192 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_421
timestamp 1676037725
transform 1 0 39836 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_436
timestamp 1676037725
transform 1 0 41216 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_449
timestamp 1676037725
transform 1 0 42412 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_461
timestamp 1676037725
transform 1 0 43516 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_465
timestamp 1676037725
transform 1 0 43884 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_473
timestamp 1676037725
transform 1 0 44620 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_477
timestamp 1676037725
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_489
timestamp 1676037725
transform 1 0 46092 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_501
timestamp 1676037725
transform 1 0 47196 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_513
timestamp 1676037725
transform 1 0 48300 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_521
timestamp 1676037725
transform 1 0 49036 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_525
timestamp 1676037725
transform 1 0 49404 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1676037725
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1676037725
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1676037725
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1676037725
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1676037725
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1676037725
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1676037725
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1676037725
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1676037725
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1676037725
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1676037725
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1676037725
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1676037725
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1676037725
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1676037725
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1676037725
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1676037725
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1676037725
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1676037725
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1676037725
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1676037725
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1676037725
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1676037725
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1676037725
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1676037725
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1676037725
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_57_254
timestamp 1676037725
transform 1 0 24472 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_266
timestamp 1676037725
transform 1 0 25576 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_278
timestamp 1676037725
transform 1 0 26680 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1676037725
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_293
timestamp 1676037725
transform 1 0 28060 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_299
timestamp 1676037725
transform 1 0 28612 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_309
timestamp 1676037725
transform 1 0 29532 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_322
timestamp 1676037725
transform 1 0 30728 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1676037725
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1676037725
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1676037725
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_349
timestamp 1676037725
transform 1 0 33212 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_377
timestamp 1676037725
transform 1 0 35788 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_383
timestamp 1676037725
transform 1 0 36340 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1676037725
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_393
timestamp 1676037725
transform 1 0 37260 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_404
timestamp 1676037725
transform 1 0 38272 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_419
timestamp 1676037725
transform 1 0 39652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_425
timestamp 1676037725
transform 1 0 40204 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_446
timestamp 1676037725
transform 1 0 42136 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_449
timestamp 1676037725
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_461
timestamp 1676037725
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_473
timestamp 1676037725
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_485
timestamp 1676037725
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1676037725
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1676037725
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_505
timestamp 1676037725
transform 1 0 47564 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_517
timestamp 1676037725
transform 1 0 48668 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_525
timestamp 1676037725
transform 1 0 49404 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1676037725
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1676037725
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1676037725
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1676037725
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1676037725
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1676037725
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1676037725
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1676037725
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1676037725
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1676037725
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1676037725
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1676037725
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1676037725
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1676037725
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1676037725
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1676037725
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1676037725
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1676037725
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1676037725
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1676037725
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1676037725
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1676037725
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp 1676037725
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_237
timestamp 1676037725
transform 1 0 22908 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_250
timestamp 1676037725
transform 1 0 24104 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1676037725
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_264
timestamp 1676037725
transform 1 0 25392 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_272
timestamp 1676037725
transform 1 0 26128 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_293
timestamp 1676037725
transform 1 0 28060 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_305
timestamp 1676037725
transform 1 0 29164 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_309
timestamp 1676037725
transform 1 0 29532 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_314
timestamp 1676037725
transform 1 0 29992 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_58_331
timestamp 1676037725
transform 1 0 31556 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_342
timestamp 1676037725
transform 1 0 32568 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_354
timestamp 1676037725
transform 1 0 33672 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_362
timestamp 1676037725
transform 1 0 34408 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_365
timestamp 1676037725
transform 1 0 34684 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_373
timestamp 1676037725
transform 1 0 35420 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_376
timestamp 1676037725
transform 1 0 35696 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_389
timestamp 1676037725
transform 1 0 36892 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_397
timestamp 1676037725
transform 1 0 37628 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_400
timestamp 1676037725
transform 1 0 37904 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_413
timestamp 1676037725
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_419
timestamp 1676037725
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_421
timestamp 1676037725
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_433
timestamp 1676037725
transform 1 0 40940 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_441
timestamp 1676037725
transform 1 0 41676 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_451
timestamp 1676037725
transform 1 0 42596 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_463
timestamp 1676037725
transform 1 0 43700 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1676037725
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_477
timestamp 1676037725
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_489
timestamp 1676037725
transform 1 0 46092 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_501
timestamp 1676037725
transform 1 0 47196 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_513
timestamp 1676037725
transform 1 0 48300 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_521
timestamp 1676037725
transform 1 0 49036 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_525
timestamp 1676037725
transform 1 0 49404 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_3
timestamp 1676037725
transform 1 0 1380 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_8
timestamp 1676037725
transform 1 0 1840 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_20
timestamp 1676037725
transform 1 0 2944 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_32
timestamp 1676037725
transform 1 0 4048 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_44
timestamp 1676037725
transform 1 0 5152 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1676037725
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1676037725
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1676037725
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1676037725
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1676037725
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1676037725
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1676037725
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1676037725
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1676037725
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1676037725
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1676037725
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1676037725
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1676037725
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1676037725
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1676037725
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1676037725
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1676037725
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1676037725
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1676037725
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_237
timestamp 1676037725
transform 1 0 22908 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_260
timestamp 1676037725
transform 1 0 25024 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1676037725
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1676037725
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1676037725
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_293
timestamp 1676037725
transform 1 0 28060 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_324
timestamp 1676037725
transform 1 0 30912 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_334
timestamp 1676037725
transform 1 0 31832 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_337
timestamp 1676037725
transform 1 0 32108 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_348
timestamp 1676037725
transform 1 0 33120 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_354
timestamp 1676037725
transform 1 0 33672 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_378
timestamp 1676037725
transform 1 0 35880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1676037725
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1676037725
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_405
timestamp 1676037725
transform 1 0 38364 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_411
timestamp 1676037725
transform 1 0 38916 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_421
timestamp 1676037725
transform 1 0 39836 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_434
timestamp 1676037725
transform 1 0 41032 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_445
timestamp 1676037725
transform 1 0 42044 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_59_449
timestamp 1676037725
transform 1 0 42412 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_464
timestamp 1676037725
transform 1 0 43792 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_476
timestamp 1676037725
transform 1 0 44896 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_488
timestamp 1676037725
transform 1 0 46000 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_500
timestamp 1676037725
transform 1 0 47104 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_505
timestamp 1676037725
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_517
timestamp 1676037725
transform 1 0 48668 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_521
timestamp 1676037725
transform 1 0 49036 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_59_525
timestamp 1676037725
transform 1 0 49404 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1676037725
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1676037725
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1676037725
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1676037725
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1676037725
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1676037725
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1676037725
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1676037725
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1676037725
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1676037725
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1676037725
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1676037725
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1676037725
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1676037725
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1676037725
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1676037725
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1676037725
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1676037725
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1676037725
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1676037725
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1676037725
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1676037725
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1676037725
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_221
timestamp 1676037725
transform 1 0 21436 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_244
timestamp 1676037725
transform 1 0 23552 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_253
timestamp 1676037725
transform 1 0 24380 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_264
timestamp 1676037725
transform 1 0 25392 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_270
timestamp 1676037725
transform 1 0 25944 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_280
timestamp 1676037725
transform 1 0 26864 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_304
timestamp 1676037725
transform 1 0 29072 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_309
timestamp 1676037725
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_317
timestamp 1676037725
transform 1 0 30268 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_321
timestamp 1676037725
transform 1 0 30636 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_334
timestamp 1676037725
transform 1 0 31832 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_358
timestamp 1676037725
transform 1 0 34040 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1676037725
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_377
timestamp 1676037725
transform 1 0 35788 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_60_388
timestamp 1676037725
transform 1 0 36800 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_403
timestamp 1676037725
transform 1 0 38180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_416
timestamp 1676037725
transform 1 0 39376 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_421
timestamp 1676037725
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_433
timestamp 1676037725
transform 1 0 40940 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_437
timestamp 1676037725
transform 1 0 41308 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_447
timestamp 1676037725
transform 1 0 42228 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_451
timestamp 1676037725
transform 1 0 42596 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_472
timestamp 1676037725
transform 1 0 44528 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_477
timestamp 1676037725
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_489
timestamp 1676037725
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_501
timestamp 1676037725
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_513
timestamp 1676037725
transform 1 0 48300 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_521
timestamp 1676037725
transform 1 0 49036 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_525
timestamp 1676037725
transform 1 0 49404 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1676037725
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1676037725
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1676037725
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1676037725
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1676037725
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1676037725
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1676037725
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1676037725
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1676037725
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1676037725
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1676037725
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1676037725
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1676037725
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1676037725
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1676037725
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1676037725
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1676037725
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1676037725
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1676037725
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1676037725
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_193
timestamp 1676037725
transform 1 0 18860 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_199
timestamp 1676037725
transform 1 0 19412 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1676037725
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_225
timestamp 1676037725
transform 1 0 21804 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_247
timestamp 1676037725
transform 1 0 23828 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_255
timestamp 1676037725
transform 1 0 24564 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_276
timestamp 1676037725
transform 1 0 26496 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_281
timestamp 1676037725
transform 1 0 26956 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_286
timestamp 1676037725
transform 1 0 27416 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_298
timestamp 1676037725
transform 1 0 28520 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_324
timestamp 1676037725
transform 1 0 30912 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_330
timestamp 1676037725
transform 1 0 31464 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_334
timestamp 1676037725
transform 1 0 31832 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1676037725
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_348
timestamp 1676037725
transform 1 0 33120 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_354
timestamp 1676037725
transform 1 0 33672 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_371
timestamp 1676037725
transform 1 0 35236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_384
timestamp 1676037725
transform 1 0 36432 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_393
timestamp 1676037725
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_401
timestamp 1676037725
transform 1 0 37996 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_423
timestamp 1676037725
transform 1 0 40020 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_436
timestamp 1676037725
transform 1 0 41216 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_449
timestamp 1676037725
transform 1 0 42412 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_471
timestamp 1676037725
transform 1 0 44436 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_483
timestamp 1676037725
transform 1 0 45540 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_495
timestamp 1676037725
transform 1 0 46644 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1676037725
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_505
timestamp 1676037725
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_517
timestamp 1676037725
transform 1 0 48668 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_521
timestamp 1676037725
transform 1 0 49036 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_525
timestamp 1676037725
transform 1 0 49404 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1676037725
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1676037725
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1676037725
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1676037725
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1676037725
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1676037725
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1676037725
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1676037725
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1676037725
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1676037725
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1676037725
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1676037725
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1676037725
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1676037725
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1676037725
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1676037725
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1676037725
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1676037725
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1676037725
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1676037725
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1676037725
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1676037725
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1676037725
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_221
timestamp 1676037725
transform 1 0 21436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_225
timestamp 1676037725
transform 1 0 21804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_228
timestamp 1676037725
transform 1 0 22080 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_241
timestamp 1676037725
transform 1 0 23276 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_249
timestamp 1676037725
transform 1 0 24012 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1676037725
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1676037725
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_277
timestamp 1676037725
transform 1 0 26588 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_62_286
timestamp 1676037725
transform 1 0 27416 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_299
timestamp 1676037725
transform 1 0 28612 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1676037725
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1676037725
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1676037725
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_333
timestamp 1676037725
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1676037725
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1676037725
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1676037725
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_365
timestamp 1676037725
transform 1 0 34684 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_378
timestamp 1676037725
transform 1 0 35880 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_391
timestamp 1676037725
transform 1 0 37076 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_404
timestamp 1676037725
transform 1 0 38272 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_416
timestamp 1676037725
transform 1 0 39376 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_421
timestamp 1676037725
transform 1 0 39836 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_433
timestamp 1676037725
transform 1 0 40940 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_446
timestamp 1676037725
transform 1 0 42136 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_459
timestamp 1676037725
transform 1 0 43332 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_471
timestamp 1676037725
transform 1 0 44436 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1676037725
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_477
timestamp 1676037725
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_489
timestamp 1676037725
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_501
timestamp 1676037725
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_513
timestamp 1676037725
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_525
timestamp 1676037725
transform 1 0 49404 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1676037725
transform 1 0 1380 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_8
timestamp 1676037725
transform 1 0 1840 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_20
timestamp 1676037725
transform 1 0 2944 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_32
timestamp 1676037725
transform 1 0 4048 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_44
timestamp 1676037725
transform 1 0 5152 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1676037725
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1676037725
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1676037725
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1676037725
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1676037725
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1676037725
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1676037725
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1676037725
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1676037725
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1676037725
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1676037725
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1676037725
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1676037725
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1676037725
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_193
timestamp 1676037725
transform 1 0 18860 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_208
timestamp 1676037725
transform 1 0 20240 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1676037725
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_225
timestamp 1676037725
transform 1 0 21804 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_233
timestamp 1676037725
transform 1 0 22540 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_238
timestamp 1676037725
transform 1 0 23000 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_265
timestamp 1676037725
transform 1 0 25484 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_63_278
timestamp 1676037725
transform 1 0 26680 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_281
timestamp 1676037725
transform 1 0 26956 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_292
timestamp 1676037725
transform 1 0 27968 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_304
timestamp 1676037725
transform 1 0 29072 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_312
timestamp 1676037725
transform 1 0 29808 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_322
timestamp 1676037725
transform 1 0 30728 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_330
timestamp 1676037725
transform 1 0 31464 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_334
timestamp 1676037725
transform 1 0 31832 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1676037725
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_348
timestamp 1676037725
transform 1 0 33120 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_360
timestamp 1676037725
transform 1 0 34224 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_381
timestamp 1676037725
transform 1 0 36156 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1676037725
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1676037725
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_404
timestamp 1676037725
transform 1 0 38272 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_416
timestamp 1676037725
transform 1 0 39376 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_440
timestamp 1676037725
transform 1 0 41584 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_449
timestamp 1676037725
transform 1 0 42412 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_460
timestamp 1676037725
transform 1 0 43424 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_472
timestamp 1676037725
transform 1 0 44528 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_484
timestamp 1676037725
transform 1 0 45632 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_496
timestamp 1676037725
transform 1 0 46736 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_63_505
timestamp 1676037725
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_517
timestamp 1676037725
transform 1 0 48668 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_521
timestamp 1676037725
transform 1 0 49036 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_525
timestamp 1676037725
transform 1 0 49404 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1676037725
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1676037725
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1676037725
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1676037725
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1676037725
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1676037725
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1676037725
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1676037725
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1676037725
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1676037725
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1676037725
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_109
timestamp 1676037725
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_121
timestamp 1676037725
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1676037725
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1676037725
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1676037725
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1676037725
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1676037725
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1676037725
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1676037725
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1676037725
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1676037725
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1676037725
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_221
timestamp 1676037725
transform 1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_227
timestamp 1676037725
transform 1 0 21988 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_237
timestamp 1676037725
transform 1 0 22908 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_250
timestamp 1676037725
transform 1 0 24104 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_253
timestamp 1676037725
transform 1 0 24380 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_258
timestamp 1676037725
transform 1 0 24840 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_264
timestamp 1676037725
transform 1 0 25392 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_274
timestamp 1676037725
transform 1 0 26312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_278
timestamp 1676037725
transform 1 0 26680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_299
timestamp 1676037725
transform 1 0 28612 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_306
timestamp 1676037725
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1676037725
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_320
timestamp 1676037725
transform 1 0 30544 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_333
timestamp 1676037725
transform 1 0 31740 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_346
timestamp 1676037725
transform 1 0 32936 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_350
timestamp 1676037725
transform 1 0 33304 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1676037725
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1676037725
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1676037725
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_389
timestamp 1676037725
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_401
timestamp 1676037725
transform 1 0 37996 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_416
timestamp 1676037725
transform 1 0 39376 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_421
timestamp 1676037725
transform 1 0 39836 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_432
timestamp 1676037725
transform 1 0 40848 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_439
timestamp 1676037725
transform 1 0 41492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_445
timestamp 1676037725
transform 1 0 42044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_466
timestamp 1676037725
transform 1 0 43976 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_474
timestamp 1676037725
transform 1 0 44712 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_477
timestamp 1676037725
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_489
timestamp 1676037725
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_501
timestamp 1676037725
transform 1 0 47196 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_511
timestamp 1676037725
transform 1 0 48116 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_64_525
timestamp 1676037725
transform 1 0 49404 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_3
timestamp 1676037725
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_15
timestamp 1676037725
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_27
timestamp 1676037725
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_39
timestamp 1676037725
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_51
timestamp 1676037725
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1676037725
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1676037725
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_69
timestamp 1676037725
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_81
timestamp 1676037725
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_93
timestamp 1676037725
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1676037725
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1676037725
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1676037725
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1676037725
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1676037725
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1676037725
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1676037725
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1676037725
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1676037725
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1676037725
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1676037725
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1676037725
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1676037725
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1676037725
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1676037725
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1676037725
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_235
timestamp 1676037725
transform 1 0 22724 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_259
timestamp 1676037725
transform 1 0 24932 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_271
timestamp 1676037725
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1676037725
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_281
timestamp 1676037725
transform 1 0 26956 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_306
timestamp 1676037725
transform 1 0 29256 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_315
timestamp 1676037725
transform 1 0 30084 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_330
timestamp 1676037725
transform 1 0 31464 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_337
timestamp 1676037725
transform 1 0 32108 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_348
timestamp 1676037725
transform 1 0 33120 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1676037725
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_373
timestamp 1676037725
transform 1 0 35420 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_390
timestamp 1676037725
transform 1 0 36984 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_393
timestamp 1676037725
transform 1 0 37260 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_404
timestamp 1676037725
transform 1 0 38272 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_428
timestamp 1676037725
transform 1 0 40480 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1676037725
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1676037725
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_449
timestamp 1676037725
transform 1 0 42412 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_460
timestamp 1676037725
transform 1 0 43424 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_472
timestamp 1676037725
transform 1 0 44528 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_484
timestamp 1676037725
transform 1 0 45632 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_496
timestamp 1676037725
transform 1 0 46736 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_65_505
timestamp 1676037725
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_517
timestamp 1676037725
transform 1 0 48668 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_521
timestamp 1676037725
transform 1 0 49036 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1676037725
transform 1 0 49404 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_3
timestamp 1676037725
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_15
timestamp 1676037725
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1676037725
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1676037725
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1676037725
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1676037725
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1676037725
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1676037725
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1676037725
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1676037725
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1676037725
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1676037725
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1676037725
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1676037725
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1676037725
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1676037725
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1676037725
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1676037725
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1676037725
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1676037725
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1676037725
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1676037725
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_209
timestamp 1676037725
transform 1 0 20332 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_237
timestamp 1676037725
transform 1 0 22908 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_250
timestamp 1676037725
transform 1 0 24104 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1676037725
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_265
timestamp 1676037725
transform 1 0 25484 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_273
timestamp 1676037725
transform 1 0 26220 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_278
timestamp 1676037725
transform 1 0 26680 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_291
timestamp 1676037725
transform 1 0 27876 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_306
timestamp 1676037725
transform 1 0 29256 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_309
timestamp 1676037725
transform 1 0 29532 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_354
timestamp 1676037725
transform 1 0 33672 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_362
timestamp 1676037725
transform 1 0 34408 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_365
timestamp 1676037725
transform 1 0 34684 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_387
timestamp 1676037725
transform 1 0 36708 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_402
timestamp 1676037725
transform 1 0 38088 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_416
timestamp 1676037725
transform 1 0 39376 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_421
timestamp 1676037725
transform 1 0 39836 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_432
timestamp 1676037725
transform 1 0 40848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_438
timestamp 1676037725
transform 1 0 41400 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_459
timestamp 1676037725
transform 1 0 43332 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_471
timestamp 1676037725
transform 1 0 44436 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1676037725
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_477
timestamp 1676037725
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_489
timestamp 1676037725
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_501
timestamp 1676037725
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_513
timestamp 1676037725
transform 1 0 48300 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_521
timestamp 1676037725
transform 1 0 49036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_525
timestamp 1676037725
transform 1 0 49404 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1676037725
transform 1 0 1380 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_8
timestamp 1676037725
transform 1 0 1840 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_20
timestamp 1676037725
transform 1 0 2944 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_32
timestamp 1676037725
transform 1 0 4048 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_44
timestamp 1676037725
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1676037725
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1676037725
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1676037725
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1676037725
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1676037725
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1676037725
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1676037725
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1676037725
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1676037725
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1676037725
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1676037725
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1676037725
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1676037725
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1676037725
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_193
timestamp 1676037725
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_205
timestamp 1676037725
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1676037725
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1676037725
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_225
timestamp 1676037725
transform 1 0 21804 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_229
timestamp 1676037725
transform 1 0 22172 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_232
timestamp 1676037725
transform 1 0 22448 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_245
timestamp 1676037725
transform 1 0 23644 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_253
timestamp 1676037725
transform 1 0 24380 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_263
timestamp 1676037725
transform 1 0 25300 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1676037725
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_281
timestamp 1676037725
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_294
timestamp 1676037725
transform 1 0 28152 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_307
timestamp 1676037725
transform 1 0 29348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_319
timestamp 1676037725
transform 1 0 30452 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_323
timestamp 1676037725
transform 1 0 30820 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_326
timestamp 1676037725
transform 1 0 31096 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_332
timestamp 1676037725
transform 1 0 31648 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_337
timestamp 1676037725
transform 1 0 32108 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_349
timestamp 1676037725
transform 1 0 33212 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_362
timestamp 1676037725
transform 1 0 34408 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_377
timestamp 1676037725
transform 1 0 35788 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_390
timestamp 1676037725
transform 1 0 36984 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_393
timestamp 1676037725
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_404
timestamp 1676037725
transform 1 0 38272 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_424
timestamp 1676037725
transform 1 0 40112 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_446
timestamp 1676037725
transform 1 0 42136 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_449
timestamp 1676037725
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_461
timestamp 1676037725
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_473
timestamp 1676037725
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_485
timestamp 1676037725
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_497
timestamp 1676037725
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_503
timestamp 1676037725
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_505
timestamp 1676037725
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_517
timestamp 1676037725
transform 1 0 48668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_525
timestamp 1676037725
transform 1 0 49404 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_3
timestamp 1676037725
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_15
timestamp 1676037725
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1676037725
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1676037725
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1676037725
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1676037725
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1676037725
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1676037725
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1676037725
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1676037725
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1676037725
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1676037725
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1676037725
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1676037725
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1676037725
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1676037725
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1676037725
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1676037725
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1676037725
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1676037725
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1676037725
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_197
timestamp 1676037725
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_209
timestamp 1676037725
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_223
timestamp 1676037725
transform 1 0 21620 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_236
timestamp 1676037725
transform 1 0 22816 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_248
timestamp 1676037725
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_253
timestamp 1676037725
transform 1 0 24380 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_68_275
timestamp 1676037725
transform 1 0 26404 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_287
timestamp 1676037725
transform 1 0 27508 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_299
timestamp 1676037725
transform 1 0 28612 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1676037725
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_309
timestamp 1676037725
transform 1 0 29532 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_315
timestamp 1676037725
transform 1 0 30084 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_336
timestamp 1676037725
transform 1 0 32016 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_68_351
timestamp 1676037725
transform 1 0 33396 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1676037725
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1676037725
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_377
timestamp 1676037725
transform 1 0 35788 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_399
timestamp 1676037725
transform 1 0 37812 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_403
timestamp 1676037725
transform 1 0 38180 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_407
timestamp 1676037725
transform 1 0 38548 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1676037725
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_421
timestamp 1676037725
transform 1 0 39836 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_429
timestamp 1676037725
transform 1 0 40572 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_453
timestamp 1676037725
transform 1 0 42780 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_465
timestamp 1676037725
transform 1 0 43884 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_473
timestamp 1676037725
transform 1 0 44620 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_477
timestamp 1676037725
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_489
timestamp 1676037725
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_501
timestamp 1676037725
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_513
timestamp 1676037725
transform 1 0 48300 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_525
timestamp 1676037725
transform 1 0 49404 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_69_3
timestamp 1676037725
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_15
timestamp 1676037725
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_27
timestamp 1676037725
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_39
timestamp 1676037725
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1676037725
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1676037725
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1676037725
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1676037725
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1676037725
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1676037725
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1676037725
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1676037725
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1676037725
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1676037725
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1676037725
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1676037725
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1676037725
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1676037725
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1676037725
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1676037725
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1676037725
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1676037725
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1676037725
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1676037725
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1676037725
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_237
timestamp 1676037725
transform 1 0 22908 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1676037725
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1676037725
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1676037725
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1676037725
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_293
timestamp 1676037725
transform 1 0 28060 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_314
timestamp 1676037725
transform 1 0 29992 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_326
timestamp 1676037725
transform 1 0 31096 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_334
timestamp 1676037725
transform 1 0 31832 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_337
timestamp 1676037725
transform 1 0 32108 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_359
timestamp 1676037725
transform 1 0 34132 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1676037725
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1676037725
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_393
timestamp 1676037725
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_405
timestamp 1676037725
transform 1 0 38364 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_427
timestamp 1676037725
transform 1 0 40388 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_440
timestamp 1676037725
transform 1 0 41584 0 -1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_69_449
timestamp 1676037725
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_461
timestamp 1676037725
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_473
timestamp 1676037725
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_485
timestamp 1676037725
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_497
timestamp 1676037725
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_503
timestamp 1676037725
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_505
timestamp 1676037725
transform 1 0 47564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_513
timestamp 1676037725
transform 1 0 48300 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_525
timestamp 1676037725
transform 1 0 49404 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_3
timestamp 1676037725
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_15
timestamp 1676037725
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1676037725
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1676037725
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1676037725
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1676037725
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1676037725
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1676037725
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1676037725
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1676037725
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1676037725
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1676037725
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1676037725
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1676037725
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1676037725
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1676037725
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1676037725
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1676037725
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1676037725
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1676037725
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1676037725
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1676037725
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1676037725
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1676037725
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_233
timestamp 1676037725
transform 1 0 22540 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_250
timestamp 1676037725
transform 1 0 24104 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1676037725
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_274
timestamp 1676037725
transform 1 0 26312 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_70_287
timestamp 1676037725
transform 1 0 27508 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_299
timestamp 1676037725
transform 1 0 28612 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1676037725
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_309
timestamp 1676037725
transform 1 0 29532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_331
timestamp 1676037725
transform 1 0 31556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_337
timestamp 1676037725
transform 1 0 32108 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_347
timestamp 1676037725
transform 1 0 33028 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_70_362
timestamp 1676037725
transform 1 0 34408 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_365
timestamp 1676037725
transform 1 0 34684 0 1 40256
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_70_380
timestamp 1676037725
transform 1 0 36064 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_392
timestamp 1676037725
transform 1 0 37168 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_404
timestamp 1676037725
transform 1 0 38272 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_408
timestamp 1676037725
transform 1 0 38640 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_418
timestamp 1676037725
transform 1 0 39560 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_70_421
timestamp 1676037725
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_433
timestamp 1676037725
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_445
timestamp 1676037725
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_457
timestamp 1676037725
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1676037725
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1676037725
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_477
timestamp 1676037725
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_489
timestamp 1676037725
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_501
timestamp 1676037725
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_513
timestamp 1676037725
transform 1 0 48300 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_525
timestamp 1676037725
transform 1 0 49404 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_3
timestamp 1676037725
transform 1 0 1380 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_15
timestamp 1676037725
transform 1 0 2484 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_27
timestamp 1676037725
transform 1 0 3588 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_39
timestamp 1676037725
transform 1 0 4692 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_47
timestamp 1676037725
transform 1 0 5428 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_53
timestamp 1676037725
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1676037725
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1676037725
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1676037725
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_97
timestamp 1676037725
transform 1 0 10028 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_107
timestamp 1676037725
transform 1 0 10948 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1676037725
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1676037725
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1676037725
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1676037725
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1676037725
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1676037725
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1676037725
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1676037725
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1676037725
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1676037725
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_205
timestamp 1676037725
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_217
timestamp 1676037725
transform 1 0 21068 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_220
timestamp 1676037725
transform 1 0 21344 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_225
timestamp 1676037725
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_236
timestamp 1676037725
transform 1 0 22816 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_242
timestamp 1676037725
transform 1 0 23368 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_254
timestamp 1676037725
transform 1 0 24472 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_277
timestamp 1676037725
transform 1 0 26588 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_281
timestamp 1676037725
transform 1 0 26956 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_71_304
timestamp 1676037725
transform 1 0 29072 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_317
timestamp 1676037725
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1676037725
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1676037725
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_337
timestamp 1676037725
transform 1 0 32108 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_345
timestamp 1676037725
transform 1 0 32844 0 -1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_71_368
timestamp 1676037725
transform 1 0 34960 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_380
timestamp 1676037725
transform 1 0 36064 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_393
timestamp 1676037725
transform 1 0 37260 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_401
timestamp 1676037725
transform 1 0 37996 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_423
timestamp 1676037725
transform 1 0 40020 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_435
timestamp 1676037725
transform 1 0 41124 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1676037725
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_449
timestamp 1676037725
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_461
timestamp 1676037725
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_473
timestamp 1676037725
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_485
timestamp 1676037725
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_497
timestamp 1676037725
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_503
timestamp 1676037725
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_505
timestamp 1676037725
transform 1 0 47564 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_513
timestamp 1676037725
transform 1 0 48300 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_525
timestamp 1676037725
transform 1 0 49404 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_72_3
timestamp 1676037725
transform 1 0 1380 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_72_9
timestamp 1676037725
transform 1 0 1932 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_21
timestamp 1676037725
transform 1 0 3036 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1676037725
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1676037725
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1676037725
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1676037725
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1676037725
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1676037725
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1676037725
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1676037725
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1676037725
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1676037725
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1676037725
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1676037725
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1676037725
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1676037725
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1676037725
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1676037725
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1676037725
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1676037725
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1676037725
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1676037725
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_209
timestamp 1676037725
transform 1 0 20332 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_217
timestamp 1676037725
transform 1 0 21068 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_220
timestamp 1676037725
transform 1 0 21344 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_247
timestamp 1676037725
transform 1 0 23828 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1676037725
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1676037725
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1676037725
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_277
timestamp 1676037725
transform 1 0 26588 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_290
timestamp 1676037725
transform 1 0 27784 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_302
timestamp 1676037725
transform 1 0 28888 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1676037725
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_321
timestamp 1676037725
transform 1 0 30636 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_72_349
timestamp 1676037725
transform 1 0 33212 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_361
timestamp 1676037725
transform 1 0 34316 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_72_365
timestamp 1676037725
transform 1 0 34684 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_387
timestamp 1676037725
transform 1 0 36708 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_411
timestamp 1676037725
transform 1 0 38916 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1676037725
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_421
timestamp 1676037725
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_433
timestamp 1676037725
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_445
timestamp 1676037725
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_457
timestamp 1676037725
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1676037725
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1676037725
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_477
timestamp 1676037725
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_489
timestamp 1676037725
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_501
timestamp 1676037725
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_513
timestamp 1676037725
transform 1 0 48300 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_519
timestamp 1676037725
transform 1 0 48852 0 1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_3
timestamp 1676037725
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_15
timestamp 1676037725
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_27
timestamp 1676037725
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_39
timestamp 1676037725
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_51
timestamp 1676037725
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1676037725
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_57
timestamp 1676037725
transform 1 0 6348 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_69
timestamp 1676037725
transform 1 0 7452 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_77
timestamp 1676037725
transform 1 0 8188 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_85
timestamp 1676037725
transform 1 0 8924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_90
timestamp 1676037725
transform 1 0 9384 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_102
timestamp 1676037725
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_110
timestamp 1676037725
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1676037725
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1676037725
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1676037725
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1676037725
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1676037725
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1676037725
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_169
timestamp 1676037725
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_173
timestamp 1676037725
transform 1 0 17020 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_178
timestamp 1676037725
transform 1 0 17480 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_190
timestamp 1676037725
transform 1 0 18584 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_202
timestamp 1676037725
transform 1 0 19688 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_210
timestamp 1676037725
transform 1 0 20424 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_215
timestamp 1676037725
transform 1 0 20884 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1676037725
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_225
timestamp 1676037725
transform 1 0 21804 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_232
timestamp 1676037725
transform 1 0 22448 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_244
timestamp 1676037725
transform 1 0 23552 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_73_270
timestamp 1676037725
transform 1 0 25944 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_278
timestamp 1676037725
transform 1 0 26680 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_281
timestamp 1676037725
transform 1 0 26956 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_310
timestamp 1676037725
transform 1 0 29624 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_334
timestamp 1676037725
transform 1 0 31832 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1676037725
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_349
timestamp 1676037725
transform 1 0 33212 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_355
timestamp 1676037725
transform 1 0 33764 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_376
timestamp 1676037725
transform 1 0 35696 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_388
timestamp 1676037725
transform 1 0 36800 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_393
timestamp 1676037725
transform 1 0 37260 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_401
timestamp 1676037725
transform 1 0 37996 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_424
timestamp 1676037725
transform 1 0 40112 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_432
timestamp 1676037725
transform 1 0 40848 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_444
timestamp 1676037725
transform 1 0 41952 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_449
timestamp 1676037725
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_461
timestamp 1676037725
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_473
timestamp 1676037725
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_485
timestamp 1676037725
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1676037725
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1676037725
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_505
timestamp 1676037725
transform 1 0 47564 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_513
timestamp 1676037725
transform 1 0 48300 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_525
timestamp 1676037725
transform 1 0 49404 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_3
timestamp 1676037725
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_15
timestamp 1676037725
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1676037725
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_29
timestamp 1676037725
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_41
timestamp 1676037725
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_53
timestamp 1676037725
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_65
timestamp 1676037725
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1676037725
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1676037725
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1676037725
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1676037725
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1676037725
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1676037725
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1676037725
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1676037725
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1676037725
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1676037725
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1676037725
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1676037725
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1676037725
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1676037725
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1676037725
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1676037725
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1676037725
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1676037725
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1676037725
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1676037725
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1676037725
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_265
timestamp 1676037725
transform 1 0 25484 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_286
timestamp 1676037725
transform 1 0 27416 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_298
timestamp 1676037725
transform 1 0 28520 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_306
timestamp 1676037725
transform 1 0 29256 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1676037725
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1676037725
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1676037725
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1676037725
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1676037725
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1676037725
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_365
timestamp 1676037725
transform 1 0 34684 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_373
timestamp 1676037725
transform 1 0 35420 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_395
timestamp 1676037725
transform 1 0 37444 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_407
timestamp 1676037725
transform 1 0 38548 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1676037725
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_421
timestamp 1676037725
transform 1 0 39836 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_432
timestamp 1676037725
transform 1 0 40848 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_444
timestamp 1676037725
transform 1 0 41952 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_456
timestamp 1676037725
transform 1 0 43056 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_468
timestamp 1676037725
transform 1 0 44160 0 1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_74_477
timestamp 1676037725
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_489
timestamp 1676037725
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_501
timestamp 1676037725
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_513
timestamp 1676037725
transform 1 0 48300 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_525
timestamp 1676037725
transform 1 0 49404 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_3
timestamp 1676037725
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_9
timestamp 1676037725
transform 1 0 1932 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_13
timestamp 1676037725
transform 1 0 2300 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_25
timestamp 1676037725
transform 1 0 3404 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_37
timestamp 1676037725
transform 1 0 4508 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_49
timestamp 1676037725
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1676037725
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1676037725
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1676037725
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1676037725
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1676037725
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1676037725
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1676037725
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_113
timestamp 1676037725
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_117
timestamp 1676037725
transform 1 0 11868 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_122
timestamp 1676037725
transform 1 0 12328 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_134
timestamp 1676037725
transform 1 0 13432 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_146
timestamp 1676037725
transform 1 0 14536 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_158
timestamp 1676037725
transform 1 0 15640 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_166
timestamp 1676037725
transform 1 0 16376 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_169
timestamp 1676037725
transform 1 0 16652 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_174
timestamp 1676037725
transform 1 0 17112 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_186
timestamp 1676037725
transform 1 0 18216 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_75_198
timestamp 1676037725
transform 1 0 19320 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_206
timestamp 1676037725
transform 1 0 20056 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_211
timestamp 1676037725
transform 1 0 20516 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_218
timestamp 1676037725
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1676037725
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1676037725
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1676037725
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_261
timestamp 1676037725
transform 1 0 25116 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1676037725
transform 1 0 26680 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_75_281
timestamp 1676037725
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_293
timestamp 1676037725
transform 1 0 28060 0 -1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_75_321
timestamp 1676037725
transform 1 0 30636 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_333
timestamp 1676037725
transform 1 0 31740 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_337
timestamp 1676037725
transform 1 0 32108 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_359
timestamp 1676037725
transform 1 0 34132 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_75_383
timestamp 1676037725
transform 1 0 36340 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1676037725
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_393
timestamp 1676037725
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_405
timestamp 1676037725
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_417
timestamp 1676037725
transform 1 0 39468 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_430
timestamp 1676037725
transform 1 0 40664 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_442
timestamp 1676037725
transform 1 0 41768 0 -1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_75_449
timestamp 1676037725
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_461
timestamp 1676037725
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_473
timestamp 1676037725
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_485
timestamp 1676037725
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_497
timestamp 1676037725
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_503
timestamp 1676037725
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_505
timestamp 1676037725
transform 1 0 47564 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_513
timestamp 1676037725
transform 1 0 48300 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_525
timestamp 1676037725
transform 1 0 49404 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_3
timestamp 1676037725
transform 1 0 1380 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_8
timestamp 1676037725
transform 1 0 1840 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_20
timestamp 1676037725
transform 1 0 2944 0 1 43520
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1676037725
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1676037725
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1676037725
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1676037725
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1676037725
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1676037725
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1676037725
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1676037725
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_109
timestamp 1676037725
transform 1 0 11132 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_117
timestamp 1676037725
transform 1 0 11868 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_124
timestamp 1676037725
transform 1 0 12512 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_132
timestamp 1676037725
transform 1 0 13248 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_137
timestamp 1676037725
transform 1 0 13708 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1676037725
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_153
timestamp 1676037725
transform 1 0 15180 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_161
timestamp 1676037725
transform 1 0 15916 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_166
timestamp 1676037725
transform 1 0 16376 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_174
timestamp 1676037725
transform 1 0 17112 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_186
timestamp 1676037725
transform 1 0 18216 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_194
timestamp 1676037725
transform 1 0 18952 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_197
timestamp 1676037725
transform 1 0 19228 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_205
timestamp 1676037725
transform 1 0 19964 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_76_212
timestamp 1676037725
transform 1 0 20608 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_216
timestamp 1676037725
transform 1 0 20976 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_221
timestamp 1676037725
transform 1 0 21436 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_227
timestamp 1676037725
transform 1 0 21988 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_233
timestamp 1676037725
transform 1 0 22540 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_238
timestamp 1676037725
transform 1 0 23000 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_250
timestamp 1676037725
transform 1 0 24104 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1676037725
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1676037725
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_277
timestamp 1676037725
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_289
timestamp 1676037725
transform 1 0 27692 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1676037725
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_309
timestamp 1676037725
transform 1 0 29532 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_76_335
timestamp 1676037725
transform 1 0 31924 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_359
timestamp 1676037725
transform 1 0 34132 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1676037725
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_365
timestamp 1676037725
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_377
timestamp 1676037725
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_389
timestamp 1676037725
transform 1 0 36892 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_402
timestamp 1676037725
transform 1 0 38088 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_414
timestamp 1676037725
transform 1 0 39192 0 1 43520
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_76_421
timestamp 1676037725
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_433
timestamp 1676037725
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_445
timestamp 1676037725
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_457
timestamp 1676037725
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1676037725
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1676037725
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_477
timestamp 1676037725
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_489
timestamp 1676037725
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_501
timestamp 1676037725
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_513
timestamp 1676037725
transform 1 0 48300 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_525
timestamp 1676037725
transform 1 0 49404 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_3
timestamp 1676037725
transform 1 0 1380 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_15
timestamp 1676037725
transform 1 0 2484 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_27
timestamp 1676037725
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_39
timestamp 1676037725
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1676037725
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1676037725
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1676037725
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1676037725
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1676037725
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1676037725
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1676037725
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1676037725
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1676037725
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1676037725
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_137
timestamp 1676037725
transform 1 0 13708 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_141
timestamp 1676037725
transform 1 0 14076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_146
timestamp 1676037725
transform 1 0 14536 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_158
timestamp 1676037725
transform 1 0 15640 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_166
timestamp 1676037725
transform 1 0 16376 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1676037725
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1676037725
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1676037725
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1676037725
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1676037725
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1676037725
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_225
timestamp 1676037725
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_237
timestamp 1676037725
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_249
timestamp 1676037725
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_261
timestamp 1676037725
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1676037725
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1676037725
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1676037725
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1676037725
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1676037725
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1676037725
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1676037725
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1676037725
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1676037725
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_349
timestamp 1676037725
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_361
timestamp 1676037725
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_373
timestamp 1676037725
transform 1 0 35420 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_390
timestamp 1676037725
transform 1 0 36984 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_77_393
timestamp 1676037725
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_405
timestamp 1676037725
transform 1 0 38364 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_418
timestamp 1676037725
transform 1 0 39560 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_430
timestamp 1676037725
transform 1 0 40664 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_442
timestamp 1676037725
transform 1 0 41768 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_449
timestamp 1676037725
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_461
timestamp 1676037725
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_473
timestamp 1676037725
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_485
timestamp 1676037725
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_497
timestamp 1676037725
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_503
timestamp 1676037725
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_505
timestamp 1676037725
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_517
timestamp 1676037725
transform 1 0 48668 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_521
timestamp 1676037725
transform 1 0 49036 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_525
timestamp 1676037725
transform 1 0 49404 0 -1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_3
timestamp 1676037725
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_15
timestamp 1676037725
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_27
timestamp 1676037725
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_29
timestamp 1676037725
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_41
timestamp 1676037725
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_53
timestamp 1676037725
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_65
timestamp 1676037725
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1676037725
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1676037725
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1676037725
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1676037725
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1676037725
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1676037725
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1676037725
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1676037725
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1676037725
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_153
timestamp 1676037725
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_165
timestamp 1676037725
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_177
timestamp 1676037725
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1676037725
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1676037725
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1676037725
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1676037725
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1676037725
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_233
timestamp 1676037725
transform 1 0 22540 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_240
timestamp 1676037725
transform 1 0 23184 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_253
timestamp 1676037725
transform 1 0 24380 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_259
timestamp 1676037725
transform 1 0 24932 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_263
timestamp 1676037725
transform 1 0 25300 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_275
timestamp 1676037725
transform 1 0 26404 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_287
timestamp 1676037725
transform 1 0 27508 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_299
timestamp 1676037725
transform 1 0 28612 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1676037725
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1676037725
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1676037725
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1676037725
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_345
timestamp 1676037725
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1676037725
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1676037725
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_78_365
timestamp 1676037725
transform 1 0 34684 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_78_376
timestamp 1676037725
transform 1 0 35696 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_388
timestamp 1676037725
transform 1 0 36800 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_400
timestamp 1676037725
transform 1 0 37904 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_412
timestamp 1676037725
transform 1 0 39008 0 1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_78_421
timestamp 1676037725
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_433
timestamp 1676037725
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_445
timestamp 1676037725
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_457
timestamp 1676037725
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1676037725
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1676037725
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_477
timestamp 1676037725
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_489
timestamp 1676037725
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_501
timestamp 1676037725
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_78_513
timestamp 1676037725
transform 1 0 48300 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_525
timestamp 1676037725
transform 1 0 49404 0 1 44608
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_79_3
timestamp 1676037725
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_15
timestamp 1676037725
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_27
timestamp 1676037725
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_39
timestamp 1676037725
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_51
timestamp 1676037725
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1676037725
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1676037725
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1676037725
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1676037725
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1676037725
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1676037725
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1676037725
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1676037725
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_125
timestamp 1676037725
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_137
timestamp 1676037725
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_153
timestamp 1676037725
transform 1 0 15180 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_165
timestamp 1676037725
transform 1 0 16284 0 -1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_79_169
timestamp 1676037725
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_181
timestamp 1676037725
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_193
timestamp 1676037725
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_205
timestamp 1676037725
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1676037725
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1676037725
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1676037725
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1676037725
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1676037725
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1676037725
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1676037725
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1676037725
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1676037725
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1676037725
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1676037725
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1676037725
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1676037725
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1676037725
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_337
timestamp 1676037725
transform 1 0 32108 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_79_348
timestamp 1676037725
transform 1 0 33120 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_361
timestamp 1676037725
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_373
timestamp 1676037725
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1676037725
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1676037725
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_393
timestamp 1676037725
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_405
timestamp 1676037725
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_417
timestamp 1676037725
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_429
timestamp 1676037725
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1676037725
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1676037725
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_449
timestamp 1676037725
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_461
timestamp 1676037725
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_473
timestamp 1676037725
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_485
timestamp 1676037725
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_497
timestamp 1676037725
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_503
timestamp 1676037725
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_505
timestamp 1676037725
transform 1 0 47564 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_512
timestamp 1676037725
transform 1 0 48208 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_519
timestamp 1676037725
transform 1 0 48852 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1676037725
transform 1 0 1380 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_80_9
timestamp 1676037725
transform 1 0 1932 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_21
timestamp 1676037725
transform 1 0 3036 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1676037725
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_29
timestamp 1676037725
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_41
timestamp 1676037725
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_53
timestamp 1676037725
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_65
timestamp 1676037725
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_77
timestamp 1676037725
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1676037725
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_85
timestamp 1676037725
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_97
timestamp 1676037725
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_109
timestamp 1676037725
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_121
timestamp 1676037725
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1676037725
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1676037725
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_141
timestamp 1676037725
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_153
timestamp 1676037725
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_165
timestamp 1676037725
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_177
timestamp 1676037725
transform 1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_185
timestamp 1676037725
transform 1 0 18124 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_191
timestamp 1676037725
transform 1 0 18676 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1676037725
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_197
timestamp 1676037725
transform 1 0 19228 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_203
timestamp 1676037725
transform 1 0 19780 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_215
timestamp 1676037725
transform 1 0 20884 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_227
timestamp 1676037725
transform 1 0 21988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_239
timestamp 1676037725
transform 1 0 23092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1676037725
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_253
timestamp 1676037725
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_265
timestamp 1676037725
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_80_277
timestamp 1676037725
transform 1 0 26588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_281
timestamp 1676037725
transform 1 0 26956 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_293
timestamp 1676037725
transform 1 0 28060 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_305
timestamp 1676037725
transform 1 0 29164 0 1 45696
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_80_309
timestamp 1676037725
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_321
timestamp 1676037725
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_333
timestamp 1676037725
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_345
timestamp 1676037725
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1676037725
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1676037725
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_365
timestamp 1676037725
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_377
timestamp 1676037725
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_389
timestamp 1676037725
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_401
timestamp 1676037725
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1676037725
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1676037725
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_421
timestamp 1676037725
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_433
timestamp 1676037725
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_445
timestamp 1676037725
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_457
timestamp 1676037725
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_469
timestamp 1676037725
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_475
timestamp 1676037725
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_477
timestamp 1676037725
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_489
timestamp 1676037725
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_501
timestamp 1676037725
transform 1 0 47196 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_525
timestamp 1676037725
transform 1 0 49404 0 1 45696
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_81_3
timestamp 1676037725
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_15
timestamp 1676037725
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_27
timestamp 1676037725
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_39
timestamp 1676037725
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_51
timestamp 1676037725
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1676037725
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_57
timestamp 1676037725
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_69
timestamp 1676037725
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_81
timestamp 1676037725
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_93
timestamp 1676037725
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1676037725
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1676037725
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_113
timestamp 1676037725
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_125
timestamp 1676037725
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_137
timestamp 1676037725
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_149
timestamp 1676037725
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1676037725
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1676037725
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_169
timestamp 1676037725
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_181
timestamp 1676037725
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_193
timestamp 1676037725
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_205
timestamp 1676037725
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1676037725
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1676037725
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_225
timestamp 1676037725
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_237
timestamp 1676037725
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_249
timestamp 1676037725
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_261
timestamp 1676037725
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1676037725
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1676037725
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_281
timestamp 1676037725
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_293
timestamp 1676037725
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_305
timestamp 1676037725
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_317
timestamp 1676037725
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1676037725
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1676037725
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_337
timestamp 1676037725
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_349
timestamp 1676037725
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_361
timestamp 1676037725
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_373
timestamp 1676037725
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1676037725
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1676037725
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_393
timestamp 1676037725
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_405
timestamp 1676037725
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_417
timestamp 1676037725
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_429
timestamp 1676037725
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1676037725
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1676037725
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_449
timestamp 1676037725
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_461
timestamp 1676037725
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_473
timestamp 1676037725
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_81_485
timestamp 1676037725
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_497
timestamp 1676037725
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_503
timestamp 1676037725
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_505
timestamp 1676037725
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_517
timestamp 1676037725
transform 1 0 48668 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_521
timestamp 1676037725
transform 1 0 49036 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_525
timestamp 1676037725
transform 1 0 49404 0 -1 46784
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_82_3
timestamp 1676037725
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_15
timestamp 1676037725
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1676037725
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_29
timestamp 1676037725
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_41
timestamp 1676037725
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_53
timestamp 1676037725
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_65
timestamp 1676037725
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_77
timestamp 1676037725
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1676037725
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_85
timestamp 1676037725
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_97
timestamp 1676037725
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_109
timestamp 1676037725
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_121
timestamp 1676037725
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1676037725
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1676037725
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_141
timestamp 1676037725
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_153
timestamp 1676037725
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_165
timestamp 1676037725
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_177
timestamp 1676037725
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1676037725
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1676037725
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_197
timestamp 1676037725
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_209
timestamp 1676037725
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_221
timestamp 1676037725
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_233
timestamp 1676037725
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_245
timestamp 1676037725
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_251
timestamp 1676037725
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_253
timestamp 1676037725
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_265
timestamp 1676037725
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_277
timestamp 1676037725
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_289
timestamp 1676037725
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1676037725
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1676037725
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_309
timestamp 1676037725
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_321
timestamp 1676037725
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_333
timestamp 1676037725
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_345
timestamp 1676037725
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1676037725
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1676037725
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_365
timestamp 1676037725
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_377
timestamp 1676037725
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_389
timestamp 1676037725
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_401
timestamp 1676037725
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1676037725
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1676037725
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_421
timestamp 1676037725
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_433
timestamp 1676037725
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_445
timestamp 1676037725
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_457
timestamp 1676037725
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_469
timestamp 1676037725
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_475
timestamp 1676037725
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_82_477
timestamp 1676037725
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_82_489
timestamp 1676037725
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_501
timestamp 1676037725
transform 1 0 47196 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_509
timestamp 1676037725
transform 1 0 47932 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_514
timestamp 1676037725
transform 1 0 48392 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_521
timestamp 1676037725
transform 1 0 49036 0 1 46784
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_83_3
timestamp 1676037725
transform 1 0 1380 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_15
timestamp 1676037725
transform 1 0 2484 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_27
timestamp 1676037725
transform 1 0 3588 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_39
timestamp 1676037725
transform 1 0 4692 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_51
timestamp 1676037725
transform 1 0 5796 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_55
timestamp 1676037725
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_57
timestamp 1676037725
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_69
timestamp 1676037725
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_81
timestamp 1676037725
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_93
timestamp 1676037725
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_105
timestamp 1676037725
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_111
timestamp 1676037725
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_113
timestamp 1676037725
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_125
timestamp 1676037725
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_137
timestamp 1676037725
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_149
timestamp 1676037725
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_161
timestamp 1676037725
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_167
timestamp 1676037725
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_169
timestamp 1676037725
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_181
timestamp 1676037725
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_193
timestamp 1676037725
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_205
timestamp 1676037725
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1676037725
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1676037725
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_225
timestamp 1676037725
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_237
timestamp 1676037725
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_249
timestamp 1676037725
transform 1 0 24012 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_255
timestamp 1676037725
transform 1 0 24564 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_259
timestamp 1676037725
transform 1 0 24932 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_271
timestamp 1676037725
transform 1 0 26036 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_279
timestamp 1676037725
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_281
timestamp 1676037725
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_293
timestamp 1676037725
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_305
timestamp 1676037725
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_317
timestamp 1676037725
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_329
timestamp 1676037725
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_335
timestamp 1676037725
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_337
timestamp 1676037725
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_349
timestamp 1676037725
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_361
timestamp 1676037725
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_373
timestamp 1676037725
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_385
timestamp 1676037725
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_391
timestamp 1676037725
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_393
timestamp 1676037725
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_405
timestamp 1676037725
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_417
timestamp 1676037725
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_429
timestamp 1676037725
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_441
timestamp 1676037725
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_447
timestamp 1676037725
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_449
timestamp 1676037725
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_461
timestamp 1676037725
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_473
timestamp 1676037725
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_83_485
timestamp 1676037725
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_497
timestamp 1676037725
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1676037725
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_83_505
timestamp 1676037725
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_517
timestamp 1676037725
transform 1 0 48668 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_525
timestamp 1676037725
transform 1 0 49404 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_3
timestamp 1676037725
transform 1 0 1380 0 1 47872
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_84_9
timestamp 1676037725
transform 1 0 1932 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_21
timestamp 1676037725
transform 1 0 3036 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_27
timestamp 1676037725
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_29
timestamp 1676037725
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_41
timestamp 1676037725
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_53
timestamp 1676037725
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_65
timestamp 1676037725
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1676037725
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1676037725
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_85
timestamp 1676037725
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_84_97
timestamp 1676037725
transform 1 0 10028 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_121
timestamp 1676037725
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_133
timestamp 1676037725
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_139
timestamp 1676037725
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_141
timestamp 1676037725
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_153
timestamp 1676037725
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_165
timestamp 1676037725
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_177
timestamp 1676037725
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_189
timestamp 1676037725
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_195
timestamp 1676037725
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_197
timestamp 1676037725
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_209
timestamp 1676037725
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_221
timestamp 1676037725
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_233
timestamp 1676037725
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_245
timestamp 1676037725
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_251
timestamp 1676037725
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_253
timestamp 1676037725
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_265
timestamp 1676037725
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_277
timestamp 1676037725
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_289
timestamp 1676037725
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_301
timestamp 1676037725
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1676037725
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_309
timestamp 1676037725
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_321
timestamp 1676037725
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_333
timestamp 1676037725
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_345
timestamp 1676037725
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_357
timestamp 1676037725
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_363
timestamp 1676037725
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_365
timestamp 1676037725
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_377
timestamp 1676037725
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_389
timestamp 1676037725
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_401
timestamp 1676037725
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_413
timestamp 1676037725
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_419
timestamp 1676037725
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_421
timestamp 1676037725
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_433
timestamp 1676037725
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_445
timestamp 1676037725
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_457
timestamp 1676037725
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1676037725
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1676037725
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_84_477
timestamp 1676037725
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_84_489
timestamp 1676037725
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_501
timestamp 1676037725
transform 1 0 47196 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_512
timestamp 1676037725
transform 1 0 48208 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_520
timestamp 1676037725
transform 1 0 48944 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_526
timestamp 1676037725
transform 1 0 49496 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_3
timestamp 1676037725
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_15
timestamp 1676037725
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_27
timestamp 1676037725
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_39
timestamp 1676037725
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_51
timestamp 1676037725
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_55
timestamp 1676037725
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_57
timestamp 1676037725
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_69
timestamp 1676037725
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_81
timestamp 1676037725
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_93
timestamp 1676037725
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_105
timestamp 1676037725
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_111
timestamp 1676037725
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_113
timestamp 1676037725
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_125
timestamp 1676037725
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_137
timestamp 1676037725
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_149
timestamp 1676037725
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_161
timestamp 1676037725
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_167
timestamp 1676037725
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_169
timestamp 1676037725
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_181
timestamp 1676037725
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_193
timestamp 1676037725
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_205
timestamp 1676037725
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_217
timestamp 1676037725
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_223
timestamp 1676037725
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_225
timestamp 1676037725
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_237
timestamp 1676037725
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_249
timestamp 1676037725
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_261
timestamp 1676037725
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_273
timestamp 1676037725
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_279
timestamp 1676037725
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_281
timestamp 1676037725
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_293
timestamp 1676037725
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_305
timestamp 1676037725
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_317
timestamp 1676037725
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_329
timestamp 1676037725
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_335
timestamp 1676037725
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_337
timestamp 1676037725
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_349
timestamp 1676037725
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_361
timestamp 1676037725
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_373
timestamp 1676037725
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_385
timestamp 1676037725
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_391
timestamp 1676037725
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_393
timestamp 1676037725
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_405
timestamp 1676037725
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_417
timestamp 1676037725
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_429
timestamp 1676037725
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_441
timestamp 1676037725
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_447
timestamp 1676037725
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_449
timestamp 1676037725
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_461
timestamp 1676037725
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_473
timestamp 1676037725
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_85_485
timestamp 1676037725
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_85_497
timestamp 1676037725
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_503
timestamp 1676037725
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_85_505
timestamp 1676037725
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_517
timestamp 1676037725
transform 1 0 48668 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_525
timestamp 1676037725
transform 1 0 49404 0 -1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_3
timestamp 1676037725
transform 1 0 1380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_15
timestamp 1676037725
transform 1 0 2484 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1676037725
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_29
timestamp 1676037725
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_41
timestamp 1676037725
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_53
timestamp 1676037725
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_65
timestamp 1676037725
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_77
timestamp 1676037725
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_83
timestamp 1676037725
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_85
timestamp 1676037725
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_97
timestamp 1676037725
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_109
timestamp 1676037725
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_121
timestamp 1676037725
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_133
timestamp 1676037725
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_139
timestamp 1676037725
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_141
timestamp 1676037725
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_153
timestamp 1676037725
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_165
timestamp 1676037725
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_177
timestamp 1676037725
transform 1 0 17388 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_181
timestamp 1676037725
transform 1 0 17756 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_186
timestamp 1676037725
transform 1 0 18216 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_194
timestamp 1676037725
transform 1 0 18952 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_197
timestamp 1676037725
transform 1 0 19228 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_205
timestamp 1676037725
transform 1 0 19964 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_86_211
timestamp 1676037725
transform 1 0 20516 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_223
timestamp 1676037725
transform 1 0 21620 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_235
timestamp 1676037725
transform 1 0 22724 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_247
timestamp 1676037725
transform 1 0 23828 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_251
timestamp 1676037725
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_253
timestamp 1676037725
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_265
timestamp 1676037725
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_277
timestamp 1676037725
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_289
timestamp 1676037725
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_301
timestamp 1676037725
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_307
timestamp 1676037725
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_309
timestamp 1676037725
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_321
timestamp 1676037725
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_333
timestamp 1676037725
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_345
timestamp 1676037725
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_357
timestamp 1676037725
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_363
timestamp 1676037725
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_365
timestamp 1676037725
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_377
timestamp 1676037725
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_389
timestamp 1676037725
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_401
timestamp 1676037725
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_413
timestamp 1676037725
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_419
timestamp 1676037725
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_421
timestamp 1676037725
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_433
timestamp 1676037725
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_445
timestamp 1676037725
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_457
timestamp 1676037725
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_86_469
timestamp 1676037725
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_475
timestamp 1676037725
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_86_477
timestamp 1676037725
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_489
timestamp 1676037725
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_86_501
timestamp 1676037725
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_86_513
timestamp 1676037725
transform 1 0 48300 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_525
timestamp 1676037725
transform 1 0 49404 0 1 48960
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_3
timestamp 1676037725
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_15
timestamp 1676037725
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_27
timestamp 1676037725
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_39
timestamp 1676037725
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_51
timestamp 1676037725
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_55
timestamp 1676037725
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_57
timestamp 1676037725
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_69
timestamp 1676037725
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_81
timestamp 1676037725
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_93
timestamp 1676037725
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_105
timestamp 1676037725
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_111
timestamp 1676037725
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_87_113
timestamp 1676037725
transform 1 0 11500 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_119
timestamp 1676037725
transform 1 0 12052 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_124
timestamp 1676037725
transform 1 0 12512 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_136
timestamp 1676037725
transform 1 0 13616 0 -1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_144
timestamp 1676037725
transform 1 0 14352 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_87_150
timestamp 1676037725
transform 1 0 14904 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_162
timestamp 1676037725
transform 1 0 16008 0 -1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_87_169
timestamp 1676037725
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_181
timestamp 1676037725
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_193
timestamp 1676037725
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_205
timestamp 1676037725
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_217
timestamp 1676037725
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_223
timestamp 1676037725
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_225
timestamp 1676037725
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_237
timestamp 1676037725
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_249
timestamp 1676037725
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_261
timestamp 1676037725
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_273
timestamp 1676037725
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_279
timestamp 1676037725
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_281
timestamp 1676037725
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_293
timestamp 1676037725
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_305
timestamp 1676037725
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_317
timestamp 1676037725
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_329
timestamp 1676037725
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_335
timestamp 1676037725
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_337
timestamp 1676037725
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_349
timestamp 1676037725
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_361
timestamp 1676037725
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_373
timestamp 1676037725
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_385
timestamp 1676037725
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_391
timestamp 1676037725
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_393
timestamp 1676037725
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_405
timestamp 1676037725
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_417
timestamp 1676037725
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_429
timestamp 1676037725
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_441
timestamp 1676037725
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_447
timestamp 1676037725
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_449
timestamp 1676037725
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_461
timestamp 1676037725
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_473
timestamp 1676037725
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_87_485
timestamp 1676037725
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_87_497
timestamp 1676037725
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_87_503
timestamp 1676037725
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_87_505
timestamp 1676037725
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_517
timestamp 1676037725
transform 1 0 48668 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_87_525
timestamp 1676037725
transform 1 0 49404 0 -1 50048
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_88_3
timestamp 1676037725
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_15
timestamp 1676037725
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_88_27
timestamp 1676037725
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_29
timestamp 1676037725
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_41
timestamp 1676037725
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_53
timestamp 1676037725
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_65
timestamp 1676037725
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_77
timestamp 1676037725
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_83
timestamp 1676037725
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_85
timestamp 1676037725
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_97
timestamp 1676037725
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_109
timestamp 1676037725
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_121
timestamp 1676037725
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_133
timestamp 1676037725
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_139
timestamp 1676037725
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_141
timestamp 1676037725
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_153
timestamp 1676037725
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_165
timestamp 1676037725
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_177
timestamp 1676037725
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_189
timestamp 1676037725
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_195
timestamp 1676037725
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_197
timestamp 1676037725
transform 1 0 19228 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_205
timestamp 1676037725
transform 1 0 19964 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_210
timestamp 1676037725
transform 1 0 20424 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_222
timestamp 1676037725
transform 1 0 21528 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_234
timestamp 1676037725
transform 1 0 22632 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_246
timestamp 1676037725
transform 1 0 23736 0 1 50048
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_88_253
timestamp 1676037725
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_265
timestamp 1676037725
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_277
timestamp 1676037725
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_289
timestamp 1676037725
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_301
timestamp 1676037725
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_307
timestamp 1676037725
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_309
timestamp 1676037725
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_321
timestamp 1676037725
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_333
timestamp 1676037725
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_345
timestamp 1676037725
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_357
timestamp 1676037725
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_363
timestamp 1676037725
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_365
timestamp 1676037725
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_377
timestamp 1676037725
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_389
timestamp 1676037725
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_401
timestamp 1676037725
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_413
timestamp 1676037725
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_419
timestamp 1676037725
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_421
timestamp 1676037725
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_433
timestamp 1676037725
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_445
timestamp 1676037725
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_457
timestamp 1676037725
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_88_469
timestamp 1676037725
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_88_475
timestamp 1676037725
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_88_477
timestamp 1676037725
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_489
timestamp 1676037725
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_88_501
timestamp 1676037725
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_513
timestamp 1676037725
transform 1 0 48300 0 1 50048
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_525
timestamp 1676037725
transform 1 0 49404 0 1 50048
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_3
timestamp 1676037725
transform 1 0 1380 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_9
timestamp 1676037725
transform 1 0 1932 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_21
timestamp 1676037725
transform 1 0 3036 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_33
timestamp 1676037725
transform 1 0 4140 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_45
timestamp 1676037725
transform 1 0 5244 0 -1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_89_53
timestamp 1676037725
transform 1 0 5980 0 -1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_89_57
timestamp 1676037725
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_69
timestamp 1676037725
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_81
timestamp 1676037725
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_93
timestamp 1676037725
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_105
timestamp 1676037725
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_111
timestamp 1676037725
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_113
timestamp 1676037725
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_125
timestamp 1676037725
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_137
timestamp 1676037725
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_149
timestamp 1676037725
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_161
timestamp 1676037725
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_167
timestamp 1676037725
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_169
timestamp 1676037725
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_181
timestamp 1676037725
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_193
timestamp 1676037725
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_205
timestamp 1676037725
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_217
timestamp 1676037725
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_223
timestamp 1676037725
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_225
timestamp 1676037725
transform 1 0 21804 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_89_231
timestamp 1676037725
transform 1 0 22356 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_237
timestamp 1676037725
transform 1 0 22908 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_242
timestamp 1676037725
transform 1 0 23368 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_254
timestamp 1676037725
transform 1 0 24472 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_266
timestamp 1676037725
transform 1 0 25576 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_278
timestamp 1676037725
transform 1 0 26680 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_89_281
timestamp 1676037725
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_293
timestamp 1676037725
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_305
timestamp 1676037725
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_317
timestamp 1676037725
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_329
timestamp 1676037725
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_335
timestamp 1676037725
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_337
timestamp 1676037725
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_349
timestamp 1676037725
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_361
timestamp 1676037725
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_373
timestamp 1676037725
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_385
timestamp 1676037725
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_391
timestamp 1676037725
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_393
timestamp 1676037725
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_405
timestamp 1676037725
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_417
timestamp 1676037725
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_429
timestamp 1676037725
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_441
timestamp 1676037725
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_447
timestamp 1676037725
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_449
timestamp 1676037725
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_461
timestamp 1676037725
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_473
timestamp 1676037725
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_89_485
timestamp 1676037725
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_89_497
timestamp 1676037725
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_89_503
timestamp 1676037725
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_89_505
timestamp 1676037725
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_517
timestamp 1676037725
transform 1 0 48668 0 -1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_525
timestamp 1676037725
transform 1 0 49404 0 -1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_3
timestamp 1676037725
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_15
timestamp 1676037725
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_27
timestamp 1676037725
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_29
timestamp 1676037725
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_41
timestamp 1676037725
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_53
timestamp 1676037725
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_65
timestamp 1676037725
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_77
timestamp 1676037725
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_83
timestamp 1676037725
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_85
timestamp 1676037725
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_97
timestamp 1676037725
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_109
timestamp 1676037725
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_121
timestamp 1676037725
transform 1 0 12236 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_127
timestamp 1676037725
transform 1 0 12788 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_90_132
timestamp 1676037725
transform 1 0 13248 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_141
timestamp 1676037725
transform 1 0 14076 0 1 51136
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_90_147
timestamp 1676037725
transform 1 0 14628 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_159
timestamp 1676037725
transform 1 0 15732 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_171
timestamp 1676037725
transform 1 0 16836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_183
timestamp 1676037725
transform 1 0 17940 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_195
timestamp 1676037725
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_197
timestamp 1676037725
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_209
timestamp 1676037725
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_221
timestamp 1676037725
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_233
timestamp 1676037725
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_245
timestamp 1676037725
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_251
timestamp 1676037725
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_90_253
timestamp 1676037725
transform 1 0 24380 0 1 51136
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_90_259
timestamp 1676037725
transform 1 0 24932 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_271
timestamp 1676037725
transform 1 0 26036 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_283
timestamp 1676037725
transform 1 0 27140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_295
timestamp 1676037725
transform 1 0 28244 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_90_307
timestamp 1676037725
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_309
timestamp 1676037725
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_321
timestamp 1676037725
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_333
timestamp 1676037725
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_345
timestamp 1676037725
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_357
timestamp 1676037725
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_363
timestamp 1676037725
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_365
timestamp 1676037725
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_377
timestamp 1676037725
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_389
timestamp 1676037725
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_401
timestamp 1676037725
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_413
timestamp 1676037725
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_419
timestamp 1676037725
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_421
timestamp 1676037725
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_433
timestamp 1676037725
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_445
timestamp 1676037725
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_457
timestamp 1676037725
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_90_469
timestamp 1676037725
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_90_475
timestamp 1676037725
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_90_477
timestamp 1676037725
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_489
timestamp 1676037725
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_90_501
timestamp 1676037725
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_513
timestamp 1676037725
transform 1 0 48300 0 1 51136
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_90_525
timestamp 1676037725
transform 1 0 49404 0 1 51136
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1676037725
transform 1 0 1380 0 -1 52224
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_91_21
timestamp 1676037725
transform 1 0 3036 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_33
timestamp 1676037725
transform 1 0 4140 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_45
timestamp 1676037725
transform 1 0 5244 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_91_53
timestamp 1676037725
transform 1 0 5980 0 -1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_91_57
timestamp 1676037725
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_69
timestamp 1676037725
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_81
timestamp 1676037725
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_93
timestamp 1676037725
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_105
timestamp 1676037725
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_111
timestamp 1676037725
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_113
timestamp 1676037725
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_125
timestamp 1676037725
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_137
timestamp 1676037725
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_149
timestamp 1676037725
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_161
timestamp 1676037725
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_167
timestamp 1676037725
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_169
timestamp 1676037725
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_181
timestamp 1676037725
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_193
timestamp 1676037725
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_205
timestamp 1676037725
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_217
timestamp 1676037725
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_223
timestamp 1676037725
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_225
timestamp 1676037725
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_237
timestamp 1676037725
transform 1 0 22908 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_243
timestamp 1676037725
transform 1 0 23460 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_247
timestamp 1676037725
transform 1 0 23828 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_259
timestamp 1676037725
transform 1 0 24932 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_271
timestamp 1676037725
transform 1 0 26036 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_91_279
timestamp 1676037725
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_281
timestamp 1676037725
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_293
timestamp 1676037725
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_305
timestamp 1676037725
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_317
timestamp 1676037725
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_329
timestamp 1676037725
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_335
timestamp 1676037725
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_337
timestamp 1676037725
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_349
timestamp 1676037725
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_361
timestamp 1676037725
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_373
timestamp 1676037725
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_385
timestamp 1676037725
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_391
timestamp 1676037725
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_393
timestamp 1676037725
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_405
timestamp 1676037725
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_417
timestamp 1676037725
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_429
timestamp 1676037725
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_441
timestamp 1676037725
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_447
timestamp 1676037725
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_449
timestamp 1676037725
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_461
timestamp 1676037725
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_473
timestamp 1676037725
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_91_485
timestamp 1676037725
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_497
timestamp 1676037725
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_91_503
timestamp 1676037725
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_91_505
timestamp 1676037725
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_517
timestamp 1676037725
transform 1 0 48668 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_91_525
timestamp 1676037725
transform 1 0 49404 0 -1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_3
timestamp 1676037725
transform 1 0 1380 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_92_21
timestamp 1676037725
transform 1 0 3036 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_27
timestamp 1676037725
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_29
timestamp 1676037725
transform 1 0 3772 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_49
timestamp 1676037725
transform 1 0 5612 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_61
timestamp 1676037725
transform 1 0 6716 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_73
timestamp 1676037725
transform 1 0 7820 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_81
timestamp 1676037725
transform 1 0 8556 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_85
timestamp 1676037725
transform 1 0 8924 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_105
timestamp 1676037725
transform 1 0 10764 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_117
timestamp 1676037725
transform 1 0 11868 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_129
timestamp 1676037725
transform 1 0 12972 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_137
timestamp 1676037725
transform 1 0 13708 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_92_141
timestamp 1676037725
transform 1 0 14076 0 1 52224
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_92_161
timestamp 1676037725
transform 1 0 15916 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_173
timestamp 1676037725
transform 1 0 17020 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_185
timestamp 1676037725
transform 1 0 18124 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_92_193
timestamp 1676037725
transform 1 0 18860 0 1 52224
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_92_197
timestamp 1676037725
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_209
timestamp 1676037725
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_221
timestamp 1676037725
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_233
timestamp 1676037725
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_245
timestamp 1676037725
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_251
timestamp 1676037725
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_253
timestamp 1676037725
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_265
timestamp 1676037725
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_277
timestamp 1676037725
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_289
timestamp 1676037725
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_301
timestamp 1676037725
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_307
timestamp 1676037725
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_309
timestamp 1676037725
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_321
timestamp 1676037725
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_333
timestamp 1676037725
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_345
timestamp 1676037725
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_357
timestamp 1676037725
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_363
timestamp 1676037725
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_365
timestamp 1676037725
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_377
timestamp 1676037725
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_389
timestamp 1676037725
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_401
timestamp 1676037725
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_413
timestamp 1676037725
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_419
timestamp 1676037725
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_421
timestamp 1676037725
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_433
timestamp 1676037725
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_445
timestamp 1676037725
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_457
timestamp 1676037725
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_92_469
timestamp 1676037725
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_92_475
timestamp 1676037725
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_92_477
timestamp 1676037725
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_489
timestamp 1676037725
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_92_501
timestamp 1676037725
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_92_513
timestamp 1676037725
transform 1 0 48300 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_521
timestamp 1676037725
transform 1 0 49036 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_525
timestamp 1676037725
transform 1 0 49404 0 1 52224
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_3
timestamp 1676037725
transform 1 0 1380 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_9
timestamp 1676037725
transform 1 0 1932 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_93_33
timestamp 1676037725
transform 1 0 4140 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_37
timestamp 1676037725
transform 1 0 4508 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_54
timestamp 1676037725
transform 1 0 6072 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_57
timestamp 1676037725
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_69
timestamp 1676037725
transform 1 0 7452 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_89
timestamp 1676037725
transform 1 0 9292 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_93
timestamp 1676037725
transform 1 0 9660 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_110
timestamp 1676037725
transform 1 0 11224 0 -1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_93_113
timestamp 1676037725
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_125
timestamp 1676037725
transform 1 0 12604 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_145
timestamp 1676037725
transform 1 0 14444 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_149
timestamp 1676037725
transform 1 0 14812 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_166
timestamp 1676037725
transform 1 0 16376 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_169
timestamp 1676037725
transform 1 0 16652 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_93_193
timestamp 1676037725
transform 1 0 18860 0 -1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_93_217
timestamp 1676037725
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_223
timestamp 1676037725
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_225
timestamp 1676037725
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_237
timestamp 1676037725
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_249
timestamp 1676037725
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_261
timestamp 1676037725
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_273
timestamp 1676037725
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_279
timestamp 1676037725
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_281
timestamp 1676037725
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_293
timestamp 1676037725
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_305
timestamp 1676037725
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_317
timestamp 1676037725
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_329
timestamp 1676037725
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_335
timestamp 1676037725
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_337
timestamp 1676037725
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_349
timestamp 1676037725
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_361
timestamp 1676037725
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_373
timestamp 1676037725
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_385
timestamp 1676037725
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_391
timestamp 1676037725
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_393
timestamp 1676037725
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_405
timestamp 1676037725
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_417
timestamp 1676037725
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_429
timestamp 1676037725
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_93_441
timestamp 1676037725
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_93_447
timestamp 1676037725
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_93_449
timestamp 1676037725
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_461
timestamp 1676037725
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_93_473
timestamp 1676037725
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_485
timestamp 1676037725
transform 1 0 45724 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_492
timestamp 1676037725
transform 1 0 46368 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_93_496
timestamp 1676037725
transform 1 0 46736 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_93_500
timestamp 1676037725
transform 1 0 47104 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_93_505
timestamp 1676037725
transform 1 0 47564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_93_525
timestamp 1676037725
transform 1 0 49404 0 -1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_94_3
timestamp 1676037725
transform 1 0 1380 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_94_25
timestamp 1676037725
transform 1 0 3404 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_29
timestamp 1676037725
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_41
timestamp 1676037725
transform 1 0 4876 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_61
timestamp 1676037725
transform 1 0 6716 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_81
timestamp 1676037725
transform 1 0 8556 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_85
timestamp 1676037725
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_97
timestamp 1676037725
transform 1 0 10028 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_117
timestamp 1676037725
transform 1 0 11868 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1676037725
transform 1 0 13708 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_141
timestamp 1676037725
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_153
timestamp 1676037725
transform 1 0 15180 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_157
timestamp 1676037725
transform 1 0 15548 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_174
timestamp 1676037725
transform 1 0 17112 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1676037725
transform 1 0 18952 0 1 53312
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_94_197
timestamp 1676037725
transform 1 0 19228 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_94_221
timestamp 1676037725
transform 1 0 21436 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_241
timestamp 1676037725
transform 1 0 23276 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_94_248
timestamp 1676037725
transform 1 0 23920 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_94_253
timestamp 1676037725
transform 1 0 24380 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_259
timestamp 1676037725
transform 1 0 24932 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_271
timestamp 1676037725
transform 1 0 26036 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_283
timestamp 1676037725
transform 1 0 27140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_295
timestamp 1676037725
transform 1 0 28244 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_94_307
timestamp 1676037725
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_309
timestamp 1676037725
transform 1 0 29532 0 1 53312
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_94_314
timestamp 1676037725
transform 1 0 29992 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_326
timestamp 1676037725
transform 1 0 31096 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_334
timestamp 1676037725
transform 1 0 31832 0 1 53312
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_94_340
timestamp 1676037725
transform 1 0 32384 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_352
timestamp 1676037725
transform 1 0 33488 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_365
timestamp 1676037725
transform 1 0 34684 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_372
timestamp 1676037725
transform 1 0 35328 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_384
timestamp 1676037725
transform 1 0 36432 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_396
timestamp 1676037725
transform 1 0 37536 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_94_400
timestamp 1676037725
transform 1 0 37904 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_94_404
timestamp 1676037725
transform 1 0 38272 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_416
timestamp 1676037725
transform 1 0 39376 0 1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_94_421
timestamp 1676037725
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_433
timestamp 1676037725
transform 1 0 40940 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_444
timestamp 1676037725
transform 1 0 41952 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_94_456
timestamp 1676037725
transform 1 0 43056 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_468
timestamp 1676037725
transform 1 0 44160 0 1 53312
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_94_477
timestamp 1676037725
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_489
timestamp 1676037725
transform 1 0 46092 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_94_513
timestamp 1676037725
transform 1 0 48300 0 1 53312
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_524
timestamp 1676037725
transform 1 0 49312 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_95_3
timestamp 1676037725
transform 1 0 1380 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_9
timestamp 1676037725
transform 1 0 1932 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_26
timestamp 1676037725
transform 1 0 3496 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_29
timestamp 1676037725
transform 1 0 3772 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_34
timestamp 1676037725
transform 1 0 4232 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_54
timestamp 1676037725
transform 1 0 6072 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_57
timestamp 1676037725
transform 1 0 6348 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_65
timestamp 1676037725
transform 1 0 7084 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_82
timestamp 1676037725
transform 1 0 8648 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_85
timestamp 1676037725
transform 1 0 8924 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_93
timestamp 1676037725
transform 1 0 9660 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_110
timestamp 1676037725
transform 1 0 11224 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_113
timestamp 1676037725
transform 1 0 11500 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_121
timestamp 1676037725
transform 1 0 12236 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_138
timestamp 1676037725
transform 1 0 13800 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_141
timestamp 1676037725
transform 1 0 14076 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_149
timestamp 1676037725
transform 1 0 14812 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1676037725
transform 1 0 16376 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_169
timestamp 1676037725
transform 1 0 16652 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_177
timestamp 1676037725
transform 1 0 17388 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_194
timestamp 1676037725
transform 1 0 18952 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_197
timestamp 1676037725
transform 1 0 19228 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_205
timestamp 1676037725
transform 1 0 19964 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_222
timestamp 1676037725
transform 1 0 21528 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_225
timestamp 1676037725
transform 1 0 21804 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_249
timestamp 1676037725
transform 1 0 24012 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_95_253
timestamp 1676037725
transform 1 0 24380 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_261
timestamp 1676037725
transform 1 0 25116 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_269
timestamp 1676037725
transform 1 0 25852 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_276
timestamp 1676037725
transform 1 0 26496 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_281
timestamp 1676037725
transform 1 0 26956 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_287
timestamp 1676037725
transform 1 0 27508 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_295
timestamp 1676037725
transform 1 0 28244 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_303
timestamp 1676037725
transform 1 0 28980 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_307
timestamp 1676037725
transform 1 0 29348 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_95_309
timestamp 1676037725
transform 1 0 29532 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_317
timestamp 1676037725
transform 1 0 30268 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_325
timestamp 1676037725
transform 1 0 31004 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_333
timestamp 1676037725
transform 1 0 31740 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_337
timestamp 1676037725
transform 1 0 32108 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_95_349
timestamp 1676037725
transform 1 0 33212 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_357
timestamp 1676037725
transform 1 0 33948 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_363
timestamp 1676037725
transform 1 0 34500 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_365
timestamp 1676037725
transform 1 0 34684 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_371
timestamp 1676037725
transform 1 0 35236 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_95_381
timestamp 1676037725
transform 1 0 36156 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_95_389
timestamp 1676037725
transform 1 0 36892 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_393
timestamp 1676037725
transform 1 0 37260 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_399
timestamp 1676037725
transform 1 0 37812 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_407
timestamp 1676037725
transform 1 0 38548 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_95_413
timestamp 1676037725
transform 1 0 39100 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_95_419
timestamp 1676037725
transform 1 0 39652 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_421
timestamp 1676037725
transform 1 0 39836 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_427
timestamp 1676037725
transform 1 0 40388 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_435
timestamp 1676037725
transform 1 0 41124 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_95_442
timestamp 1676037725
transform 1 0 41768 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_95_449
timestamp 1676037725
transform 1 0 42412 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_457
timestamp 1676037725
transform 1 0 43148 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_464
timestamp 1676037725
transform 1 0 43792 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_95_471
timestamp 1676037725
transform 1 0 44436 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_95_475
timestamp 1676037725
transform 1 0 44804 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_477
timestamp 1676037725
transform 1 0 44988 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_482
timestamp 1676037725
transform 1 0 45448 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_490
timestamp 1676037725
transform 1 0 46184 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_495
timestamp 1676037725
transform 1 0 46644 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_502
timestamp 1676037725
transform 1 0 47288 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_505
timestamp 1676037725
transform 1 0 47564 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_525
timestamp 1676037725
transform 1 0 49404 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1676037725
transform 1 0 3956 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1676037725
transform 1 0 1564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1676037725
transform 1 0 49128 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 48484 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1676037725
transform 1 0 49128 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1676037725
transform 1 0 49128 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1676037725
transform 1 0 49128 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1676037725
transform 1 0 49128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1676037725
transform 1 0 49128 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1676037725
transform 1 0 49128 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1676037725
transform 1 0 48484 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1676037725
transform 1 0 49128 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1676037725
transform 1 0 49128 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1676037725
transform 1 0 48484 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1676037725
transform 1 0 48484 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1676037725
transform 1 0 48484 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1676037725
transform 1 0 48484 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1676037725
transform 1 0 48484 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1676037725
transform 1 0 48484 0 -1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1676037725
transform 1 0 48484 0 1 42432
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1676037725
transform 1 0 48484 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1676037725
transform 1 0 48484 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1676037725
transform 1 0 48484 0 1 44608
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1676037725
transform 1 0 49128 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1676037725
transform 1 0 48484 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1676037725
transform 1 0 48484 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1676037725
transform 1 0 49128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1676037725
transform 1 0 49128 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1676037725
transform 1 0 48484 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1676037725
transform 1 0 49128 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1676037725
transform 1 0 48484 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1676037725
transform 1 0 48484 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1676037725
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input34 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 8096 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input35
timestamp 1676037725
transform 1 0 9108 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1676037725
transform 1 0 10028 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input37 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1676037725
transform 1 0 10672 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input39
timestamp 1676037725
transform 1 0 11868 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1676037725
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input41
timestamp 1676037725
transform 1 0 13248 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input42
timestamp 1676037725
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input43
timestamp 1676037725
transform 1 0 14352 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1676037725
transform 1 0 1564 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1676037725
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1676037725
transform 1 0 15824 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input47
timestamp 1676037725
transform 1 0 17020 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input48
timestamp 1676037725
transform 1 0 17756 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1676037725
transform 1 0 18032 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1676037725
transform 1 0 19228 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 1676037725
transform 1 0 19688 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1676037725
transform 1 0 20608 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1676037725
transform 1 0 20608 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1676037725
transform 1 0 21988 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1676037725
transform 1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1676037725
transform 1 0 2944 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1676037725
transform 1 0 3772 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1676037725
transform 1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input59
timestamp 1676037725
transform 1 0 5244 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input60
timestamp 1676037725
transform 1 0 5520 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1676037725
transform 1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1676037725
transform 1 0 7176 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1676037725
transform 1 0 23644 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input64
timestamp 1676037725
transform 1 0 30636 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1676037725
transform 1 0 31372 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1676037725
transform 1 0 32108 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1676037725
transform 1 0 32844 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1676037725
transform 1 0 33580 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1676037725
transform 1 0 34868 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1676037725
transform 1 0 35052 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input71
timestamp 1676037725
transform 1 0 35788 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1676037725
transform 1 0 36524 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1676037725
transform 1 0 37444 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1676037725
transform 1 0 24564 0 1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1676037725
transform 1 0 37996 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input76
timestamp 1676037725
transform 1 0 38732 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input77
timestamp 1676037725
transform 1 0 40020 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input78
timestamp 1676037725
transform 1 0 40756 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1676037725
transform 1 0 41492 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1676037725
transform 1 0 41676 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input81
timestamp 1676037725
transform 1 0 42596 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1676037725
transform 1 0 43516 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1676037725
transform 1 0 44160 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1676037725
transform 1 0 45172 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input85
timestamp 1676037725
transform 1 0 24748 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1676037725
transform 1 0 25484 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1676037725
transform 1 0 26220 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input88
timestamp 1676037725
transform 1 0 27140 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input89
timestamp 1676037725
transform 1 0 27876 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1676037725
transform 1 0 28612 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1676037725
transform 1 0 29716 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1676037725
transform 1 0 29900 0 -1 54400
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1676037725
transform 1 0 1564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1676037725
transform 1 0 1564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1676037725
transform 1 0 1564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1676037725
transform 1 0 1564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input97
timestamp 1676037725
transform 1 0 1564 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input98
timestamp 1676037725
transform 1 0 45448 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1676037725
transform 1 0 1564 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1676037725
transform 1 0 47012 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input101
timestamp 1676037725
transform 1 0 46920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1676037725
transform 1 0 49128 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1676037725
transform 1 0 49036 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1676037725
transform 1 0 49036 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input105
timestamp 1676037725
transform 1 0 49036 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1676037725
transform 1 0 49036 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input107
timestamp 1676037725
transform 1 0 49036 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1676037725
transform 1 0 49036 0 1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input109
timestamp 1676037725
transform 1 0 48852 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input110
timestamp 1676037725
transform 1 0 49036 0 1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input111
timestamp 1676037725
transform 1 0 49036 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input112
timestamp 1676037725
transform 1 0 48668 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1676037725
transform 1 0 49128 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1676037725
transform 1 0 46368 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1676037725
transform 1 0 1564 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1676037725
transform 1 0 1564 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1676037725
transform 1 0 1564 0 -1 51136
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1676037725
transform 1 0 1564 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  left_tile_270
timestamp 1676037725
transform 1 0 49128 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output119 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 47932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output120
timestamp 1676037725
transform 1 0 1564 0 -1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output121
timestamp 1676037725
transform 1 0 47932 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output122
timestamp 1676037725
transform 1 0 47932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output123
timestamp 1676037725
transform 1 0 47932 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output124
timestamp 1676037725
transform 1 0 47932 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output125
timestamp 1676037725
transform 1 0 47932 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output126
timestamp 1676037725
transform 1 0 47932 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output127
timestamp 1676037725
transform 1 0 47932 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output128
timestamp 1676037725
transform 1 0 47932 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output129
timestamp 1676037725
transform 1 0 47932 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output130
timestamp 1676037725
transform 1 0 47932 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output131
timestamp 1676037725
transform 1 0 47932 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output132
timestamp 1676037725
transform 1 0 47932 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output133
timestamp 1676037725
transform 1 0 47932 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output134
timestamp 1676037725
transform 1 0 47932 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output135
timestamp 1676037725
transform 1 0 47932 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output136
timestamp 1676037725
transform 1 0 47932 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output137
timestamp 1676037725
transform 1 0 47932 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output138
timestamp 1676037725
transform 1 0 47932 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output139
timestamp 1676037725
transform 1 0 47932 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output140
timestamp 1676037725
transform 1 0 47932 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output141
timestamp 1676037725
transform 1 0 47932 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output142
timestamp 1676037725
transform 1 0 47932 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output143
timestamp 1676037725
transform 1 0 47932 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output144
timestamp 1676037725
transform 1 0 47932 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output145
timestamp 1676037725
transform 1 0 47932 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output146
timestamp 1676037725
transform 1 0 47932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output147
timestamp 1676037725
transform 1 0 47932 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output148
timestamp 1676037725
transform 1 0 47932 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output149
timestamp 1676037725
transform 1 0 47932 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output150
timestamp 1676037725
transform 1 0 22632 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output151
timestamp 1676037725
transform 1 0 32292 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output152
timestamp 1676037725
transform 1 0 31556 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output153
timestamp 1676037725
transform 1 0 32292 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output154
timestamp 1676037725
transform 1 0 34132 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output155
timestamp 1676037725
transform 1 0 34868 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output156
timestamp 1676037725
transform 1 0 33948 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output157
timestamp 1676037725
transform 1 0 34868 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output158
timestamp 1676037725
transform 1 0 37444 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output159
timestamp 1676037725
transform 1 0 36708 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output160
timestamp 1676037725
transform 1 0 37444 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output161
timestamp 1676037725
transform 1 0 23276 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output162
timestamp 1676037725
transform 1 0 39284 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output163
timestamp 1676037725
transform 1 0 40020 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output164
timestamp 1676037725
transform 1 0 39100 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output165
timestamp 1676037725
transform 1 0 40020 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output166
timestamp 1676037725
transform 1 0 42596 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output167
timestamp 1676037725
transform 1 0 41860 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output168
timestamp 1676037725
transform 1 0 42596 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output169
timestamp 1676037725
transform 1 0 44436 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output170
timestamp 1676037725
transform 1 0 43516 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output171
timestamp 1676037725
transform 1 0 45172 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output172
timestamp 1676037725
transform 1 0 24564 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output173
timestamp 1676037725
transform 1 0 25116 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output174
timestamp 1676037725
transform 1 0 25208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output175
timestamp 1676037725
transform 1 0 27140 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output176
timestamp 1676037725
transform 1 0 27324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output177
timestamp 1676037725
transform 1 0 29716 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output178
timestamp 1676037725
transform 1 0 29164 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output179
timestamp 1676037725
transform 1 0 29716 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output180
timestamp 1676037725
transform 1 0 1564 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output181
timestamp 1676037725
transform 1 0 7176 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output182
timestamp 1676037725
transform 1 0 9292 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output183
timestamp 1676037725
transform 1 0 9752 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output184
timestamp 1676037725
transform 1 0 10396 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output185
timestamp 1676037725
transform 1 0 9752 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output186
timestamp 1676037725
transform 1 0 12236 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output187
timestamp 1676037725
transform 1 0 12972 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output188
timestamp 1676037725
transform 1 0 12328 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output189
timestamp 1676037725
transform 1 0 14444 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output190
timestamp 1676037725
transform 1 0 14904 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output191
timestamp 1676037725
transform 1 0 1932 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output192
timestamp 1676037725
transform 1 0 15640 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output193
timestamp 1676037725
transform 1 0 14904 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output194
timestamp 1676037725
transform 1 0 17388 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output195
timestamp 1676037725
transform 1 0 17480 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output196
timestamp 1676037725
transform 1 0 17480 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output197
timestamp 1676037725
transform 1 0 19596 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output198
timestamp 1676037725
transform 1 0 19964 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output199
timestamp 1676037725
transform 1 0 20056 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output200
timestamp 1676037725
transform 1 0 21804 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output201
timestamp 1676037725
transform 1 0 22540 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output202
timestamp 1676037725
transform 1 0 2668 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output203
timestamp 1676037725
transform 1 0 2024 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output204
timestamp 1676037725
transform 1 0 4140 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output205
timestamp 1676037725
transform 1 0 4600 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output206
timestamp 1676037725
transform 1 0 5244 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output207
timestamp 1676037725
transform 1 0 4600 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output208
timestamp 1676037725
transform 1 0 7084 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output209
timestamp 1676037725
transform 1 0 7820 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output210
timestamp 1676037725
transform 1 0 1564 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output211
timestamp 1676037725
transform 1 0 1564 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output212
timestamp 1676037725
transform 1 0 1564 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output213
timestamp 1676037725
transform 1 0 1564 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output214
timestamp 1676037725
transform 1 0 1564 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output215
timestamp 1676037725
transform 1 0 1564 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output216
timestamp 1676037725
transform 1 0 1564 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output217
timestamp 1676037725
transform 1 0 1564 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output218
timestamp 1676037725
transform 1 0 47748 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output219
timestamp 1676037725
transform 1 0 47932 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output220
timestamp 1676037725
transform 1 0 46828 0 1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output221
timestamp 1676037725
transform 1 0 47932 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output222
timestamp 1676037725
transform 1 0 47932 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output223
timestamp 1676037725
transform 1 0 47932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output224
timestamp 1676037725
transform 1 0 47932 0 -1 53312
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1676037725
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1676037725
transform -1 0 49864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1676037725
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1676037725
transform -1 0 49864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1676037725
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1676037725
transform -1 0 49864 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1676037725
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1676037725
transform -1 0 49864 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1676037725
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1676037725
transform -1 0 49864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1676037725
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1676037725
transform -1 0 49864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1676037725
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1676037725
transform -1 0 49864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1676037725
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1676037725
transform -1 0 49864 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1676037725
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1676037725
transform -1 0 49864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1676037725
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1676037725
transform -1 0 49864 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1676037725
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1676037725
transform -1 0 49864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1676037725
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1676037725
transform -1 0 49864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1676037725
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1676037725
transform -1 0 49864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1676037725
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1676037725
transform -1 0 49864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1676037725
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1676037725
transform -1 0 49864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1676037725
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1676037725
transform -1 0 49864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1676037725
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1676037725
transform -1 0 49864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1676037725
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1676037725
transform -1 0 49864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1676037725
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1676037725
transform -1 0 49864 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1676037725
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1676037725
transform -1 0 49864 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1676037725
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1676037725
transform -1 0 49864 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1676037725
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1676037725
transform -1 0 49864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1676037725
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1676037725
transform -1 0 49864 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1676037725
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1676037725
transform -1 0 49864 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1676037725
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1676037725
transform -1 0 49864 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1676037725
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1676037725
transform -1 0 49864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1676037725
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1676037725
transform -1 0 49864 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1676037725
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1676037725
transform -1 0 49864 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1676037725
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1676037725
transform -1 0 49864 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1676037725
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1676037725
transform -1 0 49864 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1676037725
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1676037725
transform -1 0 49864 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1676037725
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1676037725
transform -1 0 49864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1676037725
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1676037725
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1676037725
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1676037725
transform -1 0 49864 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1676037725
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1676037725
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1676037725
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1676037725
transform -1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1676037725
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1676037725
transform -1 0 49864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1676037725
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1676037725
transform -1 0 49864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1676037725
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1676037725
transform -1 0 49864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1676037725
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1676037725
transform -1 0 49864 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1676037725
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1676037725
transform -1 0 49864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1676037725
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1676037725
transform -1 0 49864 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1676037725
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1676037725
transform -1 0 49864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1676037725
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1676037725
transform -1 0 49864 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1676037725
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1676037725
transform -1 0 49864 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1676037725
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1676037725
transform -1 0 49864 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1676037725
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1676037725
transform -1 0 49864 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1676037725
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1676037725
transform -1 0 49864 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1676037725
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1676037725
transform -1 0 49864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1676037725
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1676037725
transform -1 0 49864 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1676037725
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1676037725
transform -1 0 49864 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1676037725
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1676037725
transform -1 0 49864 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1676037725
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1676037725
transform -1 0 49864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1676037725
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1676037725
transform -1 0 49864 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1676037725
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1676037725
transform -1 0 49864 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1676037725
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1676037725
transform -1 0 49864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1676037725
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1676037725
transform -1 0 49864 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1676037725
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1676037725
transform -1 0 49864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1676037725
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1676037725
transform -1 0 49864 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1676037725
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1676037725
transform -1 0 49864 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1676037725
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1676037725
transform -1 0 49864 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1676037725
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1676037725
transform -1 0 49864 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1676037725
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1676037725
transform -1 0 49864 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1676037725
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1676037725
transform -1 0 49864 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1676037725
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1676037725
transform -1 0 49864 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1676037725
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1676037725
transform -1 0 49864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1676037725
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1676037725
transform -1 0 49864 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1676037725
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1676037725
transform -1 0 49864 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1676037725
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1676037725
transform -1 0 49864 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1676037725
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1676037725
transform -1 0 49864 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1676037725
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1676037725
transform -1 0 49864 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1676037725
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1676037725
transform -1 0 49864 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1676037725
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1676037725
transform -1 0 49864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1676037725
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1676037725
transform -1 0 49864 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1676037725
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1676037725
transform -1 0 49864 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1676037725
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1676037725
transform -1 0 49864 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1676037725
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1676037725
transform -1 0 49864 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1676037725
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1676037725
transform -1 0 49864 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1676037725
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1676037725
transform -1 0 49864 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1676037725
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1676037725
transform -1 0 49864 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1676037725
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1676037725
transform -1 0 49864 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1676037725
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1676037725
transform -1 0 49864 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1676037725
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1676037725
transform -1 0 49864 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1676037725
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1676037725
transform -1 0 49864 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1676037725
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1676037725
transform -1 0 49864 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1676037725
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1676037725
transform -1 0 49864 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1676037725
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1676037725
transform -1 0 49864 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1676037725
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1676037725
transform -1 0 49864 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1676037725
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1676037725
transform -1 0 49864 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1676037725
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1676037725
transform -1 0 49864 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1676037725
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1676037725
transform -1 0 49864 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1676037725
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1676037725
transform -1 0 49864 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1676037725
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1676037725
transform -1 0 49864 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1676037725
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1676037725
transform -1 0 49864 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1676037725
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1676037725
transform -1 0 49864 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1676037725
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1676037725
transform -1 0 49864 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33672 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30084 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_1.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29808 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_3.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32476 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35328 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38732 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_5.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38456 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37628 0 -1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34960 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_7.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33948 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_11.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32108 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34132 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36892 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_13.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 37720 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_21.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 40296 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40020 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 36340 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_29.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33948 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34408 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32476 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_37.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 31280 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 35880 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_45.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 39468 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34040 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_bottom_track_53.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21712 0 1 41344
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33948 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38640 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 40940 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 41860 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 42596 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 42688 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 42136 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38640 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38180 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 39652 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 40296 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 41492 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 40848 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 38180 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_8.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 38548 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 38272 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35972 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34868 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37076 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35604 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 34684 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34868 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33856 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_14.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 33120 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34500 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_16.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 31372 0 1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30084 0 1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_18.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29992 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28796 0 -1 43520
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28152 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 28244 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27232 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 26220 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_22.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 27048 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27692 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_24.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27876 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 28520 0 -1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_26.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28336 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29348 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_30.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27140 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25944 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_32.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24564 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_34.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 22356 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22080 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 19412 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19412 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22448 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_38.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 25852 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27600 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_40.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 28796 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29992 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 30636 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_46.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 32292 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34500 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_48.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35512 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 36892 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_50.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 37444 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 37720 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 35880 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 34868 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_54.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 33672 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 33856 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_right_track_56.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34868 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 10120 0 1 47872
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24104 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_0.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 25576 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27692 0 -1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 30176 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_2.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 29716 0 1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 29716 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 29072 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_4.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 26772 0 1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 27140 0 -1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24656 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_6.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23092 0 -1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23368 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21712 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_10.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 21988 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 23092 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_12.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23920 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 25760 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24840 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_20.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 22264 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 22264 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 21068 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_28.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 19504 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 21068 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 24564 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_36.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 23276 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 24748 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_44.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 27232 0 -1 41344
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_0_
timestamp 1676037725
transform 1 0 32292 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_1_
timestamp 1676037725
transform 1 0 34316 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  sb_0__1_.mem_top_track_52.sky130_fd_sc_hd__dfrtp_1_2_
timestamp 1676037725
transform 1 0 32200 0 1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31648 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35512 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l1_in_2_
timestamp 1676037725
transform 1 0 25576 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_0_
timestamp 1676037725
transform 1 0 31924 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1__275
timestamp 1676037725
transform 1 0 29716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28612 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_1.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30268 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 29900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32936 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33488 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1__225
timestamp 1676037725
transform 1 0 31464 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29992 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_3.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32384 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32384 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_0_
timestamp 1676037725
transform 1 0 35972 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40848 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37168 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_0_
timestamp 1676037725
transform 1 0 39008 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1__228
timestamp 1676037725
transform 1 0 40020 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38180 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_5.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37812 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38640 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_2_
timestamp 1676037725
transform 1 0 33580 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3__230
timestamp 1676037725
transform 1 0 32292 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l1_in_3_
timestamp 1676037725
transform 1 0 31004 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35144 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34500 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_7.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33672 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32200 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32936 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38364 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_2_
timestamp 1676037725
transform 1 0 32292 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3__276
timestamp 1676037725
transform 1 0 29716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l1_in_3_
timestamp 1676037725
transform 1 0 27600 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_11.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32384 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33672 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40388 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l1_in_2_
timestamp 1676037725
transform 1 0 34868 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36892 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1__277
timestamp 1676037725
transform 1 0 36708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36524 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_13.mux_l3_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 34868 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34960 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_1_
timestamp 1676037725
transform 1 0 41584 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37352 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_21.mux_l2_in_1__278
timestamp 1676037725
transform 1 0 40020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_21.mux_l3_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38640 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40204 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l1_in_2_
timestamp 1676037725
transform 1 0 39008 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35328 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1__279
timestamp 1676037725
transform 1 0 36156 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l2_in_1_
timestamp 1676037725
transform 1 0 36064 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_29.mux_l3_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 32108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38272 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1__226
timestamp 1676037725
transform 1 0 29716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27692 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_37.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30820 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 27968 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l1_in_0_
timestamp 1676037725
transform 1 0 41308 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_0_
timestamp 1676037725
transform 1 0 41768 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1__227
timestamp 1676037725
transform 1 0 42596 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l2_in_1_
timestamp 1676037725
transform 1 0 42596 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_45.mux_l3_in_0_
timestamp 1676037725
transform 1 0 39284 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35604 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1__229
timestamp 1676037725
transform 1 0 31556 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32016 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_bottom_track_53.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24012 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37904 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38180 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_0.mux_l2_in_1__231
timestamp 1676037725
transform 1 0 38456 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38640 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43792 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 41124 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40388 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 37444 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 42504 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_2.mux_l2_in_1__237
timestamp 1676037725
transform 1 0 41768 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 41400 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 42964 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 45356 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38548 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40020 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_4.mux_l2_in_1__248
timestamp 1676037725
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 34868 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 39008 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 42964 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 39836 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 40020 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l1_in_2_
timestamp 1676037725
transform -1 0 36892 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 40756 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_6.mux_l2_in_1__257
timestamp 1676037725
transform 1 0 41216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 40112 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 44620 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_0_
timestamp 1676037725
transform 1 0 38732 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_1_
timestamp 1676037725
transform 1 0 39284 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l1_in_2_
timestamp 1676037725
transform 1 0 34408 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_0_
timestamp 1676037725
transform 1 0 38732 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_8.mux_l2_in_1__258
timestamp 1676037725
transform 1 0 38272 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l2_in_1_
timestamp 1676037725
transform 1 0 38456 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_8.mux_l3_in_0_
timestamp 1676037725
transform 1 0 40848 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 43608 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37260 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30728 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_10.mux_l2_in_1__232
timestamp 1676037725
transform 1 0 31096 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35972 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41308 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 36156 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_12.mux_l2_in_1__233
timestamp 1676037725
transform 1 0 32292 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 36248 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41952 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l1_in_0_
timestamp 1676037725
transform 1 0 34868 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34960 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l2_in_1_
timestamp 1676037725
transform 1 0 32292 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_14.mux_l2_in_1__234
timestamp 1676037725
transform 1 0 31556 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_14.mux_l3_in_0_
timestamp 1676037725
transform 1 0 35052 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40572 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l2_in_1_
timestamp 1676037725
transform 1 0 29716 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_16.mux_l2_in_1__235
timestamp 1676037725
transform 1 0 28980 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_16.mux_l3_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 39284 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32200 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27140 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_18.mux_l2_in_1__236
timestamp 1676037725
transform 1 0 27140 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_18.mux_l3_in_0_
timestamp 1676037725
transform 1 0 32844 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37536 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32108 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_20.mux_l2_in_1__238
timestamp 1676037725
transform 1 0 28612 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 27232 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l1_in_0_
timestamp 1676037725
transform 1 0 26680 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_22.mux_l2_in_1__239
timestamp 1676037725
transform 1 0 26496 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25300 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_22.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30636 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26036 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_24.mux_l1_in_1__240
timestamp 1676037725
transform 1 0 26404 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_24.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30636 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37444 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31924 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_26.mux_l1_in_1__241
timestamp 1676037725
transform 1 0 25760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l1_in_1_
timestamp 1676037725
transform 1 0 25392 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_26.mux_l2_in_0_
timestamp 1676037725
transform 1 0 30728 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 37628 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30728 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_28.mux_l1_in_1__242
timestamp 1676037725
transform 1 0 24564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 24564 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29624 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30176 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l1_in_1_
timestamp 1676037725
transform 1 0 26404 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_30.mux_l1_in_1__243
timestamp 1676037725
transform 1 0 25208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_30.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36616 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_32.mux_l1_in_1__244
timestamp 1676037725
transform 1 0 24932 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23736 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_32.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28336 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35788 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_34.mux_l1_in_1__245
timestamp 1676037725
transform 1 0 23184 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l1_in_1_
timestamp 1676037725
transform 1 0 22724 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_34.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27140 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 35144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 18124 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_36.mux_l2_in_1__246
timestamp 1676037725
transform 1 0 14260 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 20424 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 30452 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l1_in_0_
timestamp 1676037725
transform 1 0 25300 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_38.mux_l2_in_0__247
timestamp 1676037725
transform 1 0 30544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_38.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29808 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 36708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_40.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_40.mux_l2_in_0__249
timestamp 1676037725
transform 1 0 32016 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38456 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 29808 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_44.mux_l2_in_0__250
timestamp 1676037725
transform 1 0 34776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 33028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 38916 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30912 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_46.mux_l2_in_0__251
timestamp 1676037725
transform 1 0 35880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_46.mux_l2_in_0_
timestamp 1676037725
transform 1 0 34684 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33212 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_48.mux_l2_in_0__252
timestamp 1676037725
transform 1 0 37904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_48.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41584 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_0_
timestamp 1676037725
transform 1 0 37812 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_50.mux_l1_in_1__253
timestamp 1676037725
transform 1 0 34132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l1_in_1_
timestamp 1676037725
transform 1 0 32936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_50.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41584 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_52.mux_l2_in_0__254
timestamp 1676037725
transform 1 0 38364 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37168 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41400 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32660 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_54.mux_l2_in_0__255
timestamp 1676037725
transform 1 0 37812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_54.mux_l2_in_0_
timestamp 1676037725
transform 1 0 35880 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 40572 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33488 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_right_track_56.mux_l2_in_0__256
timestamp 1676037725
transform 1 0 37444 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_right_track_56.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37444 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 41032 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35236 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_2_
timestamp 1676037725
transform 1 0 31004 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_0.mux_l1_in_3__259
timestamp 1676037725
transform 1 0 22724 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l1_in_3_
timestamp 1676037725
transform 1 0 22448 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_0_
timestamp 1676037725
transform 1 0 26956 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25852 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_0.mux_l3_in_0_
timestamp 1676037725
transform 1 0 25852 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 24656 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33580 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38548 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l1_in_2_
timestamp 1676037725
transform 1 0 26588 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32568 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_2.mux_l2_in_1__262
timestamp 1676037725
transform 1 0 29808 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l2_in_1_
timestamp 1676037725
transform 1 0 30912 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_2.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29440 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 26680 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_0_
timestamp 1676037725
transform 1 0 32384 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_1_
timestamp 1676037725
transform 1 0 38824 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l1_in_2_
timestamp 1676037725
transform 1 0 24380 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_0_
timestamp 1676037725
transform 1 0 32292 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_4.mux_l2_in_1__266
timestamp 1676037725
transform 1 0 27140 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l2_in_1_
timestamp 1676037725
transform 1 0 26036 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_4.mux_l3_in_0_
timestamp 1676037725
transform 1 0 27324 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 25024 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_0_
timestamp 1676037725
transform 1 0 22816 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37444 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_2_
timestamp 1676037725
transform 1 0 30360 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l1_in_3_
timestamp 1676037725
transform 1 0 21988 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_6.mux_l1_in_3__269
timestamp 1676037725
transform 1 0 21252 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_0_
timestamp 1676037725
transform 1 0 27048 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l2_in_1_
timestamp 1676037725
transform 1 0 25392 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_6.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24472 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22908 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_0_
timestamp 1676037725
transform 1 0 21988 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_1_
timestamp 1676037725
transform 1 0 35604 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_2_
timestamp 1676037725
transform 1 0 28336 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_10.mux_l1_in_3__260
timestamp 1676037725
transform 1 0 21620 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l1_in_3_
timestamp 1676037725
transform 1 0 21436 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25484 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23644 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_10.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22264 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_0_
timestamp 1676037725
transform 1 0 30084 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_1_
timestamp 1676037725
transform 1 0 36156 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l1_in_2_
timestamp 1676037725
transform 1 0 21988 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_12.mux_l2_in_1__261
timestamp 1676037725
transform 1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23460 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_12.mux_l3_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 22172 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_0_
timestamp 1676037725
transform 1 0 31004 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_1_
timestamp 1676037725
transform 1 0 37352 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l1_in_2_
timestamp 1676037725
transform 1 0 22908 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_0_
timestamp 1676037725
transform 1 0 29716 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l2_in_1_
timestamp 1676037725
transform 1 0 23184 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_20.mux_l2_in_1__263
timestamp 1676037725
transform 1 0 24012 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_20.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20608 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_0_
timestamp 1676037725
transform 1 0 27784 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l1_in_1_
timestamp 1676037725
transform 1 0 28428 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_0_
timestamp 1676037725
transform 1 0 24564 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_28.mux_l2_in_1__264
timestamp 1676037725
transform 1 0 18584 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l2_in_1_
timestamp 1676037725
transform 1 0 17204 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_28.mux_l3_in_0_
timestamp 1676037725
transform 1 0 19412 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 16836 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l1_in_0_
timestamp 1676037725
transform 1 0 28520 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_0_
timestamp 1676037725
transform 1 0 28428 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_36.mux_l2_in_1__265
timestamp 1676037725
transform 1 0 22448 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l2_in_1_
timestamp 1676037725
transform 1 0 22080 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_36.mux_l3_in_0_
timestamp 1676037725
transform 1 0 23276 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 18400 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_0_
timestamp 1676037725
transform 1 0 33396 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_44.mux_l1_in_1__267
timestamp 1676037725
transform 1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l1_in_1_
timestamp 1676037725
transform 1 0 23276 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_44.mux_l2_in_0_
timestamp 1676037725
transform 1 0 25484 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 19504 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l1_in_0_
timestamp 1676037725
transform 1 0 42596 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_0_
timestamp 1676037725
transform 1 0 37352 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  sb_0__1_.mux_top_track_52.mux_l2_in_1__268
timestamp 1676037725
transform 1 0 29716 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l2_in_1_
timestamp 1676037725
transform 1 0 28704 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  sb_0__1_.mux_top_track_52.mux_l3_in_0_
timestamp 1676037725
transform 1 0 29900 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__buf_4_0_
timestamp 1676037725
transform 1 0 20884 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1676037725
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1676037725
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1676037725
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1676037725
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1676037725
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1676037725
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1676037725
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1676037725
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1676037725
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1676037725
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1676037725
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1676037725
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1676037725
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1676037725
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1676037725
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1676037725
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1676037725
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1676037725
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1676037725
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1676037725
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1676037725
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1676037725
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1676037725
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1676037725
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1676037725
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1676037725
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1676037725
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1676037725
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1676037725
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1676037725
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1676037725
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1676037725
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1676037725
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1676037725
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1676037725
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1676037725
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1676037725
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1676037725
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1676037725
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1676037725
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1676037725
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1676037725
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1676037725
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1676037725
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1676037725
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1676037725
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1676037725
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1676037725
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1676037725
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1676037725
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1676037725
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1676037725
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1676037725
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1676037725
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1676037725
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1676037725
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1676037725
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1676037725
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1676037725
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1676037725
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1676037725
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1676037725
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1676037725
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1676037725
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1676037725
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1676037725
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1676037725
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1676037725
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1676037725
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1676037725
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1676037725
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1676037725
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1676037725
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1676037725
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1676037725
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1676037725
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1676037725
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1676037725
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1676037725
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1676037725
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1676037725
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1676037725
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1676037725
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1676037725
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1676037725
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1676037725
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1676037725
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1676037725
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1676037725
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1676037725
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1676037725
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1676037725
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1676037725
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1676037725
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1676037725
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1676037725
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1676037725
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1676037725
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1676037725
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1676037725
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1676037725
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1676037725
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1676037725
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1676037725
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1676037725
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1676037725
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1676037725
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1676037725
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1676037725
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1676037725
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1676037725
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1676037725
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1676037725
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1676037725
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1676037725
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1676037725
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1676037725
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1676037725
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1676037725
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1676037725
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1676037725
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1676037725
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1676037725
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1676037725
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1676037725
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1676037725
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1676037725
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1676037725
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1676037725
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1676037725
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1676037725
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1676037725
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1676037725
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1676037725
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1676037725
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1676037725
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1676037725
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1676037725
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1676037725
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1676037725
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1676037725
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1676037725
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1676037725
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1676037725
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1676037725
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1676037725
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1676037725
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1676037725
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1676037725
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1676037725
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1676037725
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1676037725
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1676037725
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1676037725
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1676037725
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1676037725
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1676037725
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1676037725
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1676037725
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1676037725
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1676037725
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1676037725
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1676037725
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1676037725
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1676037725
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1676037725
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1676037725
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1676037725
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1676037725
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1676037725
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1676037725
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1676037725
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1676037725
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1676037725
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1676037725
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1676037725
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1676037725
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1676037725
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1676037725
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1676037725
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1676037725
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1676037725
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1676037725
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1676037725
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1676037725
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1676037725
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1676037725
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1676037725
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1676037725
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1676037725
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1676037725
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1676037725
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1676037725
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1676037725
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1676037725
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1676037725
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1676037725
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1676037725
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1676037725
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1676037725
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1676037725
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1676037725
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1676037725
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1676037725
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1676037725
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1676037725
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1676037725
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1676037725
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1676037725
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1676037725
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1676037725
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1676037725
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1676037725
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1676037725
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1676037725
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1676037725
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1676037725
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1676037725
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1676037725
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1676037725
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1676037725
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1676037725
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1676037725
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1676037725
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1676037725
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1676037725
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1676037725
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1676037725
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1676037725
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1676037725
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1676037725
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1676037725
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1676037725
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1676037725
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1676037725
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1676037725
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1676037725
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1676037725
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1676037725
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1676037725
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1676037725
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1676037725
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1676037725
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1676037725
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1676037725
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1676037725
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1676037725
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1676037725
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1676037725
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1676037725
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1676037725
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1676037725
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1676037725
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1676037725
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1676037725
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1676037725
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1676037725
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1676037725
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1676037725
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1676037725
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1676037725
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1676037725
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1676037725
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1676037725
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1676037725
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1676037725
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1676037725
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1676037725
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1676037725
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1676037725
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1676037725
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1676037725
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1676037725
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1676037725
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1676037725
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1676037725
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1676037725
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1676037725
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1676037725
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1676037725
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1676037725
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1676037725
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1676037725
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1676037725
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1676037725
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1676037725
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1676037725
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1676037725
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1676037725
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1676037725
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1676037725
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1676037725
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1676037725
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1676037725
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1676037725
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1676037725
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1676037725
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1676037725
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1676037725
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1676037725
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1676037725
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1676037725
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1676037725
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1676037725
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1676037725
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1676037725
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1676037725
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1676037725
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1676037725
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1676037725
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1676037725
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1676037725
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1676037725
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1676037725
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1676037725
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1676037725
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1676037725
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1676037725
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1676037725
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1676037725
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1676037725
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1676037725
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1676037725
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1676037725
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1676037725
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1676037725
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1676037725
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1676037725
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1676037725
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1676037725
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1676037725
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1676037725
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1676037725
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1676037725
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1676037725
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1676037725
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1676037725
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1676037725
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1676037725
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1676037725
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1676037725
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1676037725
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1676037725
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1676037725
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1676037725
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1676037725
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1676037725
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1676037725
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1676037725
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1676037725
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1676037725
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1676037725
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1676037725
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1676037725
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1676037725
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1676037725
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1676037725
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1676037725
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1676037725
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1676037725
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1676037725
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1676037725
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1676037725
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1676037725
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1676037725
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1676037725
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1676037725
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1676037725
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1676037725
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1676037725
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1676037725
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1676037725
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1676037725
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1676037725
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1676037725
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1676037725
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1676037725
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1676037725
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1676037725
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1676037725
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1676037725
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1676037725
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1676037725
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1676037725
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1676037725
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1676037725
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1676037725
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1676037725
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1676037725
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1676037725
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1676037725
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1676037725
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1676037725
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1676037725
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1676037725
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1676037725
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1676037725
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1676037725
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1676037725
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1676037725
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1676037725
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1676037725
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1676037725
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1676037725
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1676037725
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1676037725
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1676037725
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1676037725
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1676037725
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1676037725
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1676037725
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1676037725
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1676037725
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1676037725
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1676037725
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1676037725
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1676037725
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1676037725
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1676037725
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1676037725
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1676037725
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1676037725
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1676037725
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1676037725
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1676037725
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1676037725
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1676037725
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1676037725
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1676037725
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1676037725
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1676037725
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1676037725
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1676037725
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1676037725
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1676037725
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1676037725
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1676037725
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1676037725
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1676037725
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1676037725
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1676037725
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1676037725
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1676037725
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1676037725
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1676037725
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1676037725
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1676037725
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1676037725
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1676037725
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1676037725
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1676037725
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1676037725
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1676037725
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1676037725
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1676037725
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1676037725
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1676037725
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1676037725
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1676037725
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1676037725
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1676037725
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1676037725
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1676037725
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1676037725
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1676037725
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1676037725
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1676037725
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1676037725
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1676037725
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1676037725
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1676037725
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1676037725
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1676037725
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1676037725
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1676037725
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1676037725
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1676037725
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1676037725
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1676037725
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1676037725
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1676037725
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1676037725
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1676037725
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1676037725
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1676037725
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1676037725
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1676037725
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1676037725
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1676037725
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1676037725
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1676037725
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1676037725
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1676037725
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1676037725
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1676037725
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1676037725
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1676037725
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1676037725
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1676037725
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1676037725
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1676037725
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1676037725
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1676037725
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1676037725
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1676037725
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1676037725
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1676037725
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1676037725
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1676037725
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1676037725
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1676037725
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1676037725
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1676037725
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1676037725
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1676037725
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1676037725
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1676037725
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1676037725
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1676037725
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1676037725
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1676037725
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1676037725
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1676037725
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1676037725
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1676037725
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1676037725
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1676037725
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1676037725
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1676037725
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1676037725
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1676037725
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1676037725
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1676037725
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1676037725
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1676037725
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1676037725
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1676037725
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1676037725
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1676037725
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1676037725
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1676037725
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1676037725
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1676037725
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1676037725
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1676037725
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1676037725
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1676037725
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1676037725
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1676037725
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1676037725
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1676037725
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1676037725
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1676037725
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1676037725
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1676037725
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1676037725
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1676037725
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1676037725
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1676037725
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1676037725
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1676037725
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1676037725
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1676037725
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1676037725
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1676037725
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1676037725
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1676037725
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1676037725
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1676037725
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1676037725
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1676037725
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1676037725
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1676037725
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1676037725
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1676037725
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1676037725
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1676037725
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1676037725
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1676037725
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1676037725
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1676037725
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1676037725
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1676037725
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1676037725
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1676037725
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1676037725
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1676037725
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1676037725
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1676037725
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1676037725
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1676037725
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1676037725
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1676037725
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1676037725
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1676037725
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1676037725
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1676037725
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1676037725
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1676037725
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1676037725
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1676037725
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1676037725
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1676037725
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1676037725
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1676037725
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1676037725
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1676037725
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1676037725
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1676037725
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1676037725
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1676037725
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1676037725
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1676037725
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1676037725
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1676037725
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1676037725
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1676037725
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1676037725
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1676037725
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1676037725
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1676037725
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1676037725
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1676037725
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1676037725
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1676037725
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1676037725
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1676037725
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1676037725
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1676037725
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1676037725
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1676037725
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1676037725
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1676037725
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1676037725
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1676037725
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1676037725
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1676037725
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1676037725
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1676037725
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1676037725
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1676037725
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1676037725
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1676037725
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1676037725
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1676037725
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1676037725
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1676037725
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1676037725
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1676037725
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1676037725
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1676037725
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1676037725
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1676037725
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1676037725
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1676037725
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1676037725
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1676037725
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1676037725
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1676037725
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1676037725
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1676037725
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1676037725
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1676037725
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1676037725
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1676037725
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1676037725
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1676037725
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1676037725
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1676037725
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1676037725
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1676037725
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1676037725
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1676037725
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1676037725
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1676037725
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1676037725
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1676037725
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1676037725
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1676037725
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1676037725
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1676037725
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1676037725
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1676037725
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1676037725
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1676037725
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1676037725
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1676037725
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1676037725
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1676037725
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1676037725
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1676037725
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1676037725
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1676037725
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1676037725
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1676037725
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1676037725
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1676037725
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1676037725
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1676037725
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1676037725
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1676037725
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1676037725
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1676037725
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1676037725
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1676037725
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1676037725
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1676037725
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1676037725
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1676037725
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1676037725
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1676037725
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1676037725
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1676037725
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1676037725
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1676037725
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1676037725
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1676037725
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1676037725
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1676037725
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1676037725
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1676037725
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1676037725
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1676037725
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1676037725
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1676037725
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1676037725
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1676037725
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1676037725
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1676037725
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1676037725
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1676037725
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1676037725
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1676037725
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1676037725
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1676037725
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1676037725
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1676037725
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1676037725
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1676037725
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1676037725
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1676037725
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1676037725
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1676037725
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1676037725
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1676037725
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1676037725
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1676037725
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1676037725
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1676037725
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1676037725
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1676037725
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1676037725
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1676037725
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1676037725
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1676037725
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1676037725
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1676037725
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1676037725
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1676037725
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1676037725
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1676037725
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1676037725
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1676037725
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1676037725
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1676037725
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1676037725
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1676037725
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1676037725
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1676037725
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1676037725
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1676037725
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1676037725
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1676037725
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1676037725
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1676037725
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1676037725
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1676037725
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1676037725
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1676037725
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1676037725
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1676037725
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1676037725
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1676037725
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1676037725
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1676037725
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1676037725
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1676037725
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1676037725
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1676037725
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1676037725
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1676037725
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1676037725
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1676037725
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1676037725
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1676037725
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1676037725
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1676037725
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1676037725
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1676037725
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1676037725
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1676037725
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1676037725
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1676037725
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1676037725
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1676037725
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1676037725
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1676037725
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1676037725
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1676037725
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1676037725
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1676037725
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1676037725
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1676037725
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1676037725
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1676037725
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1676037725
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1676037725
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1676037725
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1676037725
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1676037725
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1676037725
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1676037725
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1676037725
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1676037725
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1676037725
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1676037725
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1676037725
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1676037725
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1676037725
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1676037725
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1676037725
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1676037725
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1676037725
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1676037725
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1676037725
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1676037725
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1676037725
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1676037725
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1676037725
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1676037725
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1676037725
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1676037725
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1676037725
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1676037725
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1676037725
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1676037725
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1676037725
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1676037725
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1676037725
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1676037725
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1676037725
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1676037725
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1676037725
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1676037725
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1676037725
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1676037725
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1676037725
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1676037725
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1676037725
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1676037725
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1676037725
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1676037725
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1676037725
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1676037725
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1676037725
transform 1 0 3680 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1676037725
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1676037725
transform 1 0 8832 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1676037725
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1676037725
transform 1 0 13984 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1676037725
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1676037725
transform 1 0 19136 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1676037725
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1676037725
transform 1 0 24288 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1676037725
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1676037725
transform 1 0 29440 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1676037725
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1676037725
transform 1 0 34592 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1676037725
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1676037725
transform 1 0 39744 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1676037725
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1676037725
transform 1 0 44896 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1676037725
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
<< labels >>
flabel metal4 s 7944 2128 8264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 17944 2128 18264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 27944 2128 28264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 37944 2128 38264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 47944 2128 48264 54448 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 2944 2128 3264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12944 2128 13264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 22944 2128 23264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 32944 2128 33264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 42944 2128 43264 54448 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 54952 800 55072 0 FreeSans 480 0 0 0 ccff_head
port 2 nsew signal input
flabel metal3 s 0 1776 800 1896 0 FreeSans 480 0 0 0 ccff_head_0
port 3 nsew signal input
flabel metal3 s 50200 4224 51000 4344 0 FreeSans 480 0 0 0 ccff_tail
port 4 nsew signal tristate
flabel metal2 s 386 56200 442 57000 0 FreeSans 224 90 0 0 ccff_tail_0
port 5 nsew signal tristate
flabel metal3 s 50200 25304 51000 25424 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 6 nsew signal input
flabel metal3 s 50200 32104 51000 32224 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 7 nsew signal input
flabel metal3 s 50200 32784 51000 32904 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 8 nsew signal input
flabel metal3 s 50200 33464 51000 33584 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 9 nsew signal input
flabel metal3 s 50200 34144 51000 34264 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 10 nsew signal input
flabel metal3 s 50200 34824 51000 34944 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 11 nsew signal input
flabel metal3 s 50200 35504 51000 35624 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 12 nsew signal input
flabel metal3 s 50200 36184 51000 36304 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 13 nsew signal input
flabel metal3 s 50200 36864 51000 36984 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 14 nsew signal input
flabel metal3 s 50200 37544 51000 37664 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 15 nsew signal input
flabel metal3 s 50200 38224 51000 38344 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 16 nsew signal input
flabel metal3 s 50200 25984 51000 26104 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 17 nsew signal input
flabel metal3 s 50200 38904 51000 39024 0 FreeSans 480 0 0 0 chanx_right_in[20]
port 18 nsew signal input
flabel metal3 s 50200 39584 51000 39704 0 FreeSans 480 0 0 0 chanx_right_in[21]
port 19 nsew signal input
flabel metal3 s 50200 40264 51000 40384 0 FreeSans 480 0 0 0 chanx_right_in[22]
port 20 nsew signal input
flabel metal3 s 50200 40944 51000 41064 0 FreeSans 480 0 0 0 chanx_right_in[23]
port 21 nsew signal input
flabel metal3 s 50200 41624 51000 41744 0 FreeSans 480 0 0 0 chanx_right_in[24]
port 22 nsew signal input
flabel metal3 s 50200 42304 51000 42424 0 FreeSans 480 0 0 0 chanx_right_in[25]
port 23 nsew signal input
flabel metal3 s 50200 42984 51000 43104 0 FreeSans 480 0 0 0 chanx_right_in[26]
port 24 nsew signal input
flabel metal3 s 50200 43664 51000 43784 0 FreeSans 480 0 0 0 chanx_right_in[27]
port 25 nsew signal input
flabel metal3 s 50200 44344 51000 44464 0 FreeSans 480 0 0 0 chanx_right_in[28]
port 26 nsew signal input
flabel metal3 s 50200 45024 51000 45144 0 FreeSans 480 0 0 0 chanx_right_in[29]
port 27 nsew signal input
flabel metal3 s 50200 26664 51000 26784 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 28 nsew signal input
flabel metal3 s 50200 27344 51000 27464 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 29 nsew signal input
flabel metal3 s 50200 28024 51000 28144 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 30 nsew signal input
flabel metal3 s 50200 28704 51000 28824 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 31 nsew signal input
flabel metal3 s 50200 29384 51000 29504 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 32 nsew signal input
flabel metal3 s 50200 30064 51000 30184 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 33 nsew signal input
flabel metal3 s 50200 30744 51000 30864 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 34 nsew signal input
flabel metal3 s 50200 31424 51000 31544 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 35 nsew signal input
flabel metal3 s 50200 4904 51000 5024 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 36 nsew signal tristate
flabel metal3 s 50200 11704 51000 11824 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 37 nsew signal tristate
flabel metal3 s 50200 12384 51000 12504 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 38 nsew signal tristate
flabel metal3 s 50200 13064 51000 13184 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 39 nsew signal tristate
flabel metal3 s 50200 13744 51000 13864 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 40 nsew signal tristate
flabel metal3 s 50200 14424 51000 14544 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 41 nsew signal tristate
flabel metal3 s 50200 15104 51000 15224 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 42 nsew signal tristate
flabel metal3 s 50200 15784 51000 15904 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 43 nsew signal tristate
flabel metal3 s 50200 16464 51000 16584 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 44 nsew signal tristate
flabel metal3 s 50200 17144 51000 17264 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 45 nsew signal tristate
flabel metal3 s 50200 17824 51000 17944 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 46 nsew signal tristate
flabel metal3 s 50200 5584 51000 5704 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 47 nsew signal tristate
flabel metal3 s 50200 18504 51000 18624 0 FreeSans 480 0 0 0 chanx_right_out[20]
port 48 nsew signal tristate
flabel metal3 s 50200 19184 51000 19304 0 FreeSans 480 0 0 0 chanx_right_out[21]
port 49 nsew signal tristate
flabel metal3 s 50200 19864 51000 19984 0 FreeSans 480 0 0 0 chanx_right_out[22]
port 50 nsew signal tristate
flabel metal3 s 50200 20544 51000 20664 0 FreeSans 480 0 0 0 chanx_right_out[23]
port 51 nsew signal tristate
flabel metal3 s 50200 21224 51000 21344 0 FreeSans 480 0 0 0 chanx_right_out[24]
port 52 nsew signal tristate
flabel metal3 s 50200 21904 51000 22024 0 FreeSans 480 0 0 0 chanx_right_out[25]
port 53 nsew signal tristate
flabel metal3 s 50200 22584 51000 22704 0 FreeSans 480 0 0 0 chanx_right_out[26]
port 54 nsew signal tristate
flabel metal3 s 50200 23264 51000 23384 0 FreeSans 480 0 0 0 chanx_right_out[27]
port 55 nsew signal tristate
flabel metal3 s 50200 23944 51000 24064 0 FreeSans 480 0 0 0 chanx_right_out[28]
port 56 nsew signal tristate
flabel metal3 s 50200 24624 51000 24744 0 FreeSans 480 0 0 0 chanx_right_out[29]
port 57 nsew signal tristate
flabel metal3 s 50200 6264 51000 6384 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 58 nsew signal tristate
flabel metal3 s 50200 6944 51000 7064 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 59 nsew signal tristate
flabel metal3 s 50200 7624 51000 7744 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 60 nsew signal tristate
flabel metal3 s 50200 8304 51000 8424 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 61 nsew signal tristate
flabel metal3 s 50200 8984 51000 9104 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 62 nsew signal tristate
flabel metal3 s 50200 9664 51000 9784 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 63 nsew signal tristate
flabel metal3 s 50200 10344 51000 10464 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 64 nsew signal tristate
flabel metal3 s 50200 11024 51000 11144 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 65 nsew signal tristate
flabel metal2 s 754 0 810 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 66 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 67 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 68 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 69 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 70 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 71 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 72 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 73 nsew signal input
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 74 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 75 nsew signal input
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 76 nsew signal input
flabel metal2 s 1490 0 1546 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 77 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_in[20]
port 78 nsew signal input
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_in[21]
port 79 nsew signal input
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_in[22]
port 80 nsew signal input
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_in[23]
port 81 nsew signal input
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_in[24]
port 82 nsew signal input
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_in[25]
port 83 nsew signal input
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 chany_bottom_in[26]
port 84 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 chany_bottom_in[27]
port 85 nsew signal input
flabel metal2 s 21362 0 21418 800 0 FreeSans 224 90 0 0 chany_bottom_in[28]
port 86 nsew signal input
flabel metal2 s 22098 0 22154 800 0 FreeSans 224 90 0 0 chany_bottom_in[29]
port 87 nsew signal input
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 88 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 89 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 90 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 91 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 92 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 93 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 94 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 95 nsew signal input
flabel metal2 s 22834 0 22890 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 96 nsew signal tristate
flabel metal2 s 30194 0 30250 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 97 nsew signal tristate
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 98 nsew signal tristate
flabel metal2 s 31666 0 31722 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 99 nsew signal tristate
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 100 nsew signal tristate
flabel metal2 s 33138 0 33194 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 101 nsew signal tristate
flabel metal2 s 33874 0 33930 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 102 nsew signal tristate
flabel metal2 s 34610 0 34666 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 103 nsew signal tristate
flabel metal2 s 35346 0 35402 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 104 nsew signal tristate
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 105 nsew signal tristate
flabel metal2 s 36818 0 36874 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 106 nsew signal tristate
flabel metal2 s 23570 0 23626 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 107 nsew signal tristate
flabel metal2 s 37554 0 37610 800 0 FreeSans 224 90 0 0 chany_bottom_out[20]
port 108 nsew signal tristate
flabel metal2 s 38290 0 38346 800 0 FreeSans 224 90 0 0 chany_bottom_out[21]
port 109 nsew signal tristate
flabel metal2 s 39026 0 39082 800 0 FreeSans 224 90 0 0 chany_bottom_out[22]
port 110 nsew signal tristate
flabel metal2 s 39762 0 39818 800 0 FreeSans 224 90 0 0 chany_bottom_out[23]
port 111 nsew signal tristate
flabel metal2 s 40498 0 40554 800 0 FreeSans 224 90 0 0 chany_bottom_out[24]
port 112 nsew signal tristate
flabel metal2 s 41234 0 41290 800 0 FreeSans 224 90 0 0 chany_bottom_out[25]
port 113 nsew signal tristate
flabel metal2 s 41970 0 42026 800 0 FreeSans 224 90 0 0 chany_bottom_out[26]
port 114 nsew signal tristate
flabel metal2 s 42706 0 42762 800 0 FreeSans 224 90 0 0 chany_bottom_out[27]
port 115 nsew signal tristate
flabel metal2 s 43442 0 43498 800 0 FreeSans 224 90 0 0 chany_bottom_out[28]
port 116 nsew signal tristate
flabel metal2 s 44178 0 44234 800 0 FreeSans 224 90 0 0 chany_bottom_out[29]
port 117 nsew signal tristate
flabel metal2 s 24306 0 24362 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 118 nsew signal tristate
flabel metal2 s 25042 0 25098 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 119 nsew signal tristate
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 120 nsew signal tristate
flabel metal2 s 26514 0 26570 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 121 nsew signal tristate
flabel metal2 s 27250 0 27306 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 122 nsew signal tristate
flabel metal2 s 27986 0 28042 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 123 nsew signal tristate
flabel metal2 s 28722 0 28778 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 124 nsew signal tristate
flabel metal2 s 29458 0 29514 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 125 nsew signal tristate
flabel metal2 s 23202 56200 23258 57000 0 FreeSans 224 90 0 0 chany_top_in_0[0]
port 126 nsew signal input
flabel metal2 s 30562 56200 30618 57000 0 FreeSans 224 90 0 0 chany_top_in_0[10]
port 127 nsew signal input
flabel metal2 s 31298 56200 31354 57000 0 FreeSans 224 90 0 0 chany_top_in_0[11]
port 128 nsew signal input
flabel metal2 s 32034 56200 32090 57000 0 FreeSans 224 90 0 0 chany_top_in_0[12]
port 129 nsew signal input
flabel metal2 s 32770 56200 32826 57000 0 FreeSans 224 90 0 0 chany_top_in_0[13]
port 130 nsew signal input
flabel metal2 s 33506 56200 33562 57000 0 FreeSans 224 90 0 0 chany_top_in_0[14]
port 131 nsew signal input
flabel metal2 s 34242 56200 34298 57000 0 FreeSans 224 90 0 0 chany_top_in_0[15]
port 132 nsew signal input
flabel metal2 s 34978 56200 35034 57000 0 FreeSans 224 90 0 0 chany_top_in_0[16]
port 133 nsew signal input
flabel metal2 s 35714 56200 35770 57000 0 FreeSans 224 90 0 0 chany_top_in_0[17]
port 134 nsew signal input
flabel metal2 s 36450 56200 36506 57000 0 FreeSans 224 90 0 0 chany_top_in_0[18]
port 135 nsew signal input
flabel metal2 s 37186 56200 37242 57000 0 FreeSans 224 90 0 0 chany_top_in_0[19]
port 136 nsew signal input
flabel metal2 s 23938 56200 23994 57000 0 FreeSans 224 90 0 0 chany_top_in_0[1]
port 137 nsew signal input
flabel metal2 s 37922 56200 37978 57000 0 FreeSans 224 90 0 0 chany_top_in_0[20]
port 138 nsew signal input
flabel metal2 s 38658 56200 38714 57000 0 FreeSans 224 90 0 0 chany_top_in_0[21]
port 139 nsew signal input
flabel metal2 s 39394 56200 39450 57000 0 FreeSans 224 90 0 0 chany_top_in_0[22]
port 140 nsew signal input
flabel metal2 s 40130 56200 40186 57000 0 FreeSans 224 90 0 0 chany_top_in_0[23]
port 141 nsew signal input
flabel metal2 s 40866 56200 40922 57000 0 FreeSans 224 90 0 0 chany_top_in_0[24]
port 142 nsew signal input
flabel metal2 s 41602 56200 41658 57000 0 FreeSans 224 90 0 0 chany_top_in_0[25]
port 143 nsew signal input
flabel metal2 s 42338 56200 42394 57000 0 FreeSans 224 90 0 0 chany_top_in_0[26]
port 144 nsew signal input
flabel metal2 s 43074 56200 43130 57000 0 FreeSans 224 90 0 0 chany_top_in_0[27]
port 145 nsew signal input
flabel metal2 s 43810 56200 43866 57000 0 FreeSans 224 90 0 0 chany_top_in_0[28]
port 146 nsew signal input
flabel metal2 s 44546 56200 44602 57000 0 FreeSans 224 90 0 0 chany_top_in_0[29]
port 147 nsew signal input
flabel metal2 s 24674 56200 24730 57000 0 FreeSans 224 90 0 0 chany_top_in_0[2]
port 148 nsew signal input
flabel metal2 s 25410 56200 25466 57000 0 FreeSans 224 90 0 0 chany_top_in_0[3]
port 149 nsew signal input
flabel metal2 s 26146 56200 26202 57000 0 FreeSans 224 90 0 0 chany_top_in_0[4]
port 150 nsew signal input
flabel metal2 s 26882 56200 26938 57000 0 FreeSans 224 90 0 0 chany_top_in_0[5]
port 151 nsew signal input
flabel metal2 s 27618 56200 27674 57000 0 FreeSans 224 90 0 0 chany_top_in_0[6]
port 152 nsew signal input
flabel metal2 s 28354 56200 28410 57000 0 FreeSans 224 90 0 0 chany_top_in_0[7]
port 153 nsew signal input
flabel metal2 s 29090 56200 29146 57000 0 FreeSans 224 90 0 0 chany_top_in_0[8]
port 154 nsew signal input
flabel metal2 s 29826 56200 29882 57000 0 FreeSans 224 90 0 0 chany_top_in_0[9]
port 155 nsew signal input
flabel metal2 s 1122 56200 1178 57000 0 FreeSans 224 90 0 0 chany_top_out_0[0]
port 156 nsew signal tristate
flabel metal2 s 8482 56200 8538 57000 0 FreeSans 224 90 0 0 chany_top_out_0[10]
port 157 nsew signal tristate
flabel metal2 s 9218 56200 9274 57000 0 FreeSans 224 90 0 0 chany_top_out_0[11]
port 158 nsew signal tristate
flabel metal2 s 9954 56200 10010 57000 0 FreeSans 224 90 0 0 chany_top_out_0[12]
port 159 nsew signal tristate
flabel metal2 s 10690 56200 10746 57000 0 FreeSans 224 90 0 0 chany_top_out_0[13]
port 160 nsew signal tristate
flabel metal2 s 11426 56200 11482 57000 0 FreeSans 224 90 0 0 chany_top_out_0[14]
port 161 nsew signal tristate
flabel metal2 s 12162 56200 12218 57000 0 FreeSans 224 90 0 0 chany_top_out_0[15]
port 162 nsew signal tristate
flabel metal2 s 12898 56200 12954 57000 0 FreeSans 224 90 0 0 chany_top_out_0[16]
port 163 nsew signal tristate
flabel metal2 s 13634 56200 13690 57000 0 FreeSans 224 90 0 0 chany_top_out_0[17]
port 164 nsew signal tristate
flabel metal2 s 14370 56200 14426 57000 0 FreeSans 224 90 0 0 chany_top_out_0[18]
port 165 nsew signal tristate
flabel metal2 s 15106 56200 15162 57000 0 FreeSans 224 90 0 0 chany_top_out_0[19]
port 166 nsew signal tristate
flabel metal2 s 1858 56200 1914 57000 0 FreeSans 224 90 0 0 chany_top_out_0[1]
port 167 nsew signal tristate
flabel metal2 s 15842 56200 15898 57000 0 FreeSans 224 90 0 0 chany_top_out_0[20]
port 168 nsew signal tristate
flabel metal2 s 16578 56200 16634 57000 0 FreeSans 224 90 0 0 chany_top_out_0[21]
port 169 nsew signal tristate
flabel metal2 s 17314 56200 17370 57000 0 FreeSans 224 90 0 0 chany_top_out_0[22]
port 170 nsew signal tristate
flabel metal2 s 18050 56200 18106 57000 0 FreeSans 224 90 0 0 chany_top_out_0[23]
port 171 nsew signal tristate
flabel metal2 s 18786 56200 18842 57000 0 FreeSans 224 90 0 0 chany_top_out_0[24]
port 172 nsew signal tristate
flabel metal2 s 19522 56200 19578 57000 0 FreeSans 224 90 0 0 chany_top_out_0[25]
port 173 nsew signal tristate
flabel metal2 s 20258 56200 20314 57000 0 FreeSans 224 90 0 0 chany_top_out_0[26]
port 174 nsew signal tristate
flabel metal2 s 20994 56200 21050 57000 0 FreeSans 224 90 0 0 chany_top_out_0[27]
port 175 nsew signal tristate
flabel metal2 s 21730 56200 21786 57000 0 FreeSans 224 90 0 0 chany_top_out_0[28]
port 176 nsew signal tristate
flabel metal2 s 22466 56200 22522 57000 0 FreeSans 224 90 0 0 chany_top_out_0[29]
port 177 nsew signal tristate
flabel metal2 s 2594 56200 2650 57000 0 FreeSans 224 90 0 0 chany_top_out_0[2]
port 178 nsew signal tristate
flabel metal2 s 3330 56200 3386 57000 0 FreeSans 224 90 0 0 chany_top_out_0[3]
port 179 nsew signal tristate
flabel metal2 s 4066 56200 4122 57000 0 FreeSans 224 90 0 0 chany_top_out_0[4]
port 180 nsew signal tristate
flabel metal2 s 4802 56200 4858 57000 0 FreeSans 224 90 0 0 chany_top_out_0[5]
port 181 nsew signal tristate
flabel metal2 s 5538 56200 5594 57000 0 FreeSans 224 90 0 0 chany_top_out_0[6]
port 182 nsew signal tristate
flabel metal2 s 6274 56200 6330 57000 0 FreeSans 224 90 0 0 chany_top_out_0[7]
port 183 nsew signal tristate
flabel metal2 s 7010 56200 7066 57000 0 FreeSans 224 90 0 0 chany_top_out_0[8]
port 184 nsew signal tristate
flabel metal2 s 7746 56200 7802 57000 0 FreeSans 224 90 0 0 chany_top_out_0[9]
port 185 nsew signal tristate
flabel metal3 s 0 13336 800 13456 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[0]
port 186 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[1]
port 187 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[2]
port 188 nsew signal tristate
flabel metal3 s 0 20272 800 20392 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_dir[3]
port 189 nsew signal tristate
flabel metal3 s 0 31832 800 31952 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[0]
port 190 nsew signal input
flabel metal3 s 0 34144 800 34264 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[1]
port 191 nsew signal input
flabel metal3 s 0 36456 800 36576 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[2]
port 192 nsew signal input
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_in[3]
port 193 nsew signal input
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[0]
port 194 nsew signal tristate
flabel metal3 s 0 24896 800 25016 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[1]
port 195 nsew signal tristate
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[2]
port 196 nsew signal tristate
flabel metal3 s 0 29520 800 29640 0 FreeSans 480 0 0 0 gfpga_pad_io_soc_out[3]
port 197 nsew signal tristate
flabel metal3 s 0 41080 800 41200 0 FreeSans 480 0 0 0 isol_n
port 198 nsew signal input
flabel metal2 s 44914 0 44970 800 0 FreeSans 224 90 0 0 prog_clk
port 199 nsew signal input
flabel metal2 s 45650 0 45706 800 0 FreeSans 224 90 0 0 prog_reset_bottom_in
port 200 nsew signal input
flabel metal2 s 46386 0 46442 800 0 FreeSans 224 90 0 0 prog_reset_bottom_out
port 201 nsew signal tristate
flabel metal3 s 0 43392 800 43512 0 FreeSans 480 0 0 0 prog_reset_left_in
port 202 nsew signal input
flabel metal3 s 50200 45704 51000 45824 0 FreeSans 480 0 0 0 prog_reset_right_out
port 203 nsew signal tristate
flabel metal2 s 47490 56200 47546 57000 0 FreeSans 224 90 0 0 prog_reset_top_in
port 204 nsew signal input
flabel metal2 s 46754 56200 46810 57000 0 FreeSans 224 90 0 0 prog_reset_top_out
port 205 nsew signal tristate
flabel metal2 s 47122 0 47178 800 0 FreeSans 224 90 0 0 reset_bottom_in
port 206 nsew signal input
flabel metal2 s 47858 0 47914 800 0 FreeSans 224 90 0 0 reset_bottom_out
port 207 nsew signal tristate
flabel metal3 s 50200 46384 51000 46504 0 FreeSans 480 0 0 0 reset_right_in
port 208 nsew signal input
flabel metal2 s 48962 56200 49018 57000 0 FreeSans 224 90 0 0 reset_top_in
port 209 nsew signal input
flabel metal2 s 48226 56200 48282 57000 0 FreeSans 224 90 0 0 reset_top_out
port 210 nsew signal tristate
flabel metal3 s 50200 47064 51000 47184 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
port 211 nsew signal input
flabel metal3 s 50200 47744 51000 47864 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
port 212 nsew signal input
flabel metal3 s 50200 48424 51000 48544 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
port 213 nsew signal input
flabel metal3 s 50200 49104 51000 49224 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
port 214 nsew signal input
flabel metal3 s 50200 49784 51000 49904 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
port 215 nsew signal input
flabel metal3 s 50200 50464 51000 50584 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
port 216 nsew signal input
flabel metal3 s 50200 51144 51000 51264 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
port 217 nsew signal input
flabel metal3 s 50200 51824 51000 51944 0 FreeSans 480 0 0 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
port 218 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_0__pin_inpad_0_
port 219 nsew signal tristate
flabel metal3 s 0 6400 800 6520 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_1__pin_inpad_0_
port 220 nsew signal tristate
flabel metal3 s 0 8712 800 8832 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_2__pin_inpad_0_
port 221 nsew signal tristate
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 right_width_0_height_0_subtile_3__pin_inpad_0_
port 222 nsew signal tristate
flabel metal2 s 48594 0 48650 800 0 FreeSans 224 90 0 0 test_enable_bottom_in
port 223 nsew signal input
flabel metal2 s 49330 0 49386 800 0 FreeSans 224 90 0 0 test_enable_bottom_out
port 224 nsew signal tristate
flabel metal3 s 50200 52504 51000 52624 0 FreeSans 480 0 0 0 test_enable_right_in
port 225 nsew signal input
flabel metal2 s 50434 56200 50490 57000 0 FreeSans 224 90 0 0 test_enable_top_in
port 226 nsew signal input
flabel metal2 s 49698 56200 49754 57000 0 FreeSans 224 90 0 0 test_enable_top_out
port 227 nsew signal tristate
flabel metal3 s 0 45704 800 45824 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
port 228 nsew signal input
flabel metal3 s 0 48016 800 48136 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
port 229 nsew signal input
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
port 230 nsew signal input
flabel metal3 s 0 52640 800 52760 0 FreeSans 480 0 0 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
port 231 nsew signal input
rlabel metal1 25484 54400 25484 54400 0 VGND
rlabel metal1 25484 53856 25484 53856 0 VPWR
rlabel metal1 17986 22576 17986 22576 0 cby_0__1_.cby_0__1_.ccff_tail
rlabel metal1 10028 26418 10028 26418 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_
rlabel metal2 12282 22542 12282 22542 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_
rlabel metal2 10994 20502 10994 20502 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_
rlabel metal2 13478 21692 13478 21692 0 cby_0__1_.cby_0__1_.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_
rlabel metal1 20010 23698 20010 23698 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.ccff_tail
rlabel metal1 17296 8398 17296 8398 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[0\]
rlabel metal2 21390 20978 21390 20978 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[1\]
rlabel metal2 21298 24174 21298 24174 0 cby_0__1_.cby_0__1_.mem_right_ipin_0.mem_out\[2\]
rlabel metal1 21482 19958 21482 19958 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.ccff_tail
rlabel metal1 29348 17102 29348 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[0\]
rlabel metal1 19412 17714 19412 17714 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[1\]
rlabel metal1 23368 19890 23368 19890 0 cby_0__1_.cby_0__1_.mem_right_ipin_1.mem_out\[2\]
rlabel metal1 20700 17714 20700 17714 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.ccff_tail
rlabel metal2 25070 17748 25070 17748 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[0\]
rlabel metal2 21758 18734 21758 18734 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[1\]
rlabel metal1 20056 17102 20056 17102 0 cby_0__1_.cby_0__1_.mem_right_ipin_2.mem_out\[2\]
rlabel metal1 21160 18802 21160 18802 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[0\]
rlabel metal1 20102 21420 20102 21420 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[1\]
rlabel metal1 19918 22610 19918 22610 0 cby_0__1_.cby_0__1_.mem_right_ipin_3.mem_out\[2\]
rlabel metal2 26450 17680 26450 17680 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20240 23834 20240 23834 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 17940 23834 17940 23834 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 26496 17850 26496 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28382 19278 28382 19278 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25714 21658 25714 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22908 19482 22908 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 24426 20026 24426 20026 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 23828 21658 23828 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 20976 21658 20976 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 23322 24480 23322 24480 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 19826 23562 19826 23562 0 cby_0__1_.cby_0__1_.mux_right_ipin_0.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 28198 12954 28198 12954 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 22494 19142 22494 19142 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 18216 19482 18216 19482 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 28014 16558 28014 16558 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 26220 20570 26220 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27186 19822 27186 19822 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20010 17578 20010 17578 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 27186 17374 27186 17374 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24748 18734 24748 18734 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 19044 17782 19044 17782 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 23138 18598 23138 18598 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 21206 19142 21206 19142 0 cby_0__1_.cby_0__1_.mux_right_ipin_1.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 30038 13736 30038 13736 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 19826 17782 19826 17782 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 18676 17850 18676 17850 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 28060 13498 28060 13498 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28014 21862 28014 21862 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 27278 17952 27278 17952 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 21436 20570 21436 20570 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 25484 15130 25484 15130 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 25484 16558 25484 16558 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 19826 19312 19826 19312 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal1 22540 17306 22540 17306 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal2 22034 16694 22034 16694 0 cby_0__1_.cby_0__1_.mux_right_ipin_2.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal1 26542 16218 26542 16218 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 18584 22746 18584 22746 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_10_X
rlabel metal1 15548 21658 15548 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_11_X
rlabel metal1 26128 18394 26128 18394 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 26726 20978 26726 20978 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 23782 21930 23782 21930 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 20102 18938 20102 18938 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 21574 22678 21574 22678 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 23322 22406 23322 22406 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 19642 21658 19642 21658 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_7_X
rlabel metal2 22310 23936 22310 23936 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_8_X
rlabel metal1 19320 22474 19320 22474 0 cby_0__1_.cby_0__1_.mux_right_ipin_3.sky130_fd_sc_hd__mux2_1_9_X
rlabel metal2 12374 24480 12374 24480 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.ccff_tail
rlabel metal1 4600 23086 4600 23086 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_dir
rlabel metal1 6003 28050 6003 28050 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.gfpga_pad_io_soc_out
rlabel metal1 7751 27574 7751 27574 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal1 10902 24344 10902 24344 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.ccff_tail
rlabel metal1 8418 23630 8418 23630 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_dir
rlabel metal2 6302 24548 6302 24548 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.gfpga_pad_io_soc_out
rlabel metal1 7843 26554 7843 26554 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 16468 21658 16468 21658 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.ccff_tail
rlabel metal2 9338 19822 9338 19822 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_dir
rlabel metal2 9706 22066 9706 22066 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.gfpga_pad_io_soc_out
rlabel metal1 8441 24718 8441 24718 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal2 9798 20162 9798 20162 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_dir
rlabel metal2 10258 21794 10258 21794 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.gfpga_pad_io_soc_out
rlabel metal1 9177 23154 9177 23154 0 cby_0__1_.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_0_.SOC_DIR_N
rlabel metal3 1740 55012 1740 55012 0 ccff_head
rlabel metal1 2300 3502 2300 3502 0 ccff_head_0
rlabel metal3 49734 4284 49734 4284 0 ccff_tail
rlabel metal1 1656 55726 1656 55726 0 ccff_tail_0
rlabel metal2 49358 25619 49358 25619 0 chanx_right_in[0]
rlabel metal2 48530 32249 48530 32249 0 chanx_right_in[10]
rlabel via2 49358 32861 49358 32861 0 chanx_right_in[11]
rlabel metal2 49358 33745 49358 33745 0 chanx_right_in[12]
rlabel metal2 49358 34391 49358 34391 0 chanx_right_in[13]
rlabel metal2 49358 34969 49358 34969 0 chanx_right_in[14]
rlabel metal2 49358 35615 49358 35615 0 chanx_right_in[15]
rlabel metal2 49358 36499 49358 36499 0 chanx_right_in[16]
rlabel metal2 48530 37111 48530 37111 0 chanx_right_in[17]
rlabel metal2 49358 37723 49358 37723 0 chanx_right_in[18]
rlabel via2 49358 38301 49358 38301 0 chanx_right_in[19]
rlabel metal2 48530 26197 48530 26197 0 chanx_right_in[1]
rlabel metal2 48530 39185 48530 39185 0 chanx_right_in[20]
rlabel metal2 48530 39797 48530 39797 0 chanx_right_in[21]
rlabel metal2 48530 40409 48530 40409 0 chanx_right_in[22]
rlabel via2 48530 41021 48530 41021 0 chanx_right_in[23]
rlabel metal2 48530 41905 48530 41905 0 chanx_right_in[24]
rlabel metal2 48530 42517 48530 42517 0 chanx_right_in[25]
rlabel metal2 48530 43129 48530 43129 0 chanx_right_in[26]
rlabel via2 48530 43741 48530 43741 0 chanx_right_in[27]
rlabel metal2 48530 44625 48530 44625 0 chanx_right_in[28]
rlabel metal2 49358 44727 49358 44727 0 chanx_right_in[29]
rlabel metal2 48530 26809 48530 26809 0 chanx_right_in[2]
rlabel via2 48530 27421 48530 27421 0 chanx_right_in[3]
rlabel metal2 49358 28305 49358 28305 0 chanx_right_in[4]
rlabel metal2 49358 28951 49358 28951 0 chanx_right_in[5]
rlabel metal2 48530 29529 48530 29529 0 chanx_right_in[6]
rlabel metal2 49358 30175 49358 30175 0 chanx_right_in[7]
rlabel metal2 48530 31025 48530 31025 0 chanx_right_in[8]
rlabel metal1 48300 31790 48300 31790 0 chanx_right_in[9]
rlabel metal3 49734 11764 49734 11764 0 chanx_right_out[10]
rlabel metal2 49174 12597 49174 12597 0 chanx_right_out[11]
rlabel metal3 49734 13124 49734 13124 0 chanx_right_out[12]
rlabel via2 49174 13821 49174 13821 0 chanx_right_out[13]
rlabel metal2 49174 14705 49174 14705 0 chanx_right_out[14]
rlabel metal3 49734 15164 49734 15164 0 chanx_right_out[15]
rlabel metal2 49174 15929 49174 15929 0 chanx_right_out[16]
rlabel via2 49174 16507 49174 16507 0 chanx_right_out[17]
rlabel metal3 49734 17204 49734 17204 0 chanx_right_out[18]
rlabel metal2 49174 18037 49174 18037 0 chanx_right_out[19]
rlabel metal3 49734 5644 49734 5644 0 chanx_right_out[1]
rlabel metal3 49734 18564 49734 18564 0 chanx_right_out[20]
rlabel metal2 49174 19295 49174 19295 0 chanx_right_out[21]
rlabel metal2 49174 20145 49174 20145 0 chanx_right_out[22]
rlabel metal3 49734 20604 49734 20604 0 chanx_right_out[23]
rlabel metal2 49174 21369 49174 21369 0 chanx_right_out[24]
rlabel metal3 49734 21964 49734 21964 0 chanx_right_out[25]
rlabel metal3 49734 22644 49734 22644 0 chanx_right_out[26]
rlabel metal2 49174 23477 49174 23477 0 chanx_right_out[27]
rlabel metal3 49734 24004 49734 24004 0 chanx_right_out[28]
rlabel via2 49174 24701 49174 24701 0 chanx_right_out[29]
rlabel metal3 49734 6324 49734 6324 0 chanx_right_out[2]
rlabel metal2 49174 7157 49174 7157 0 chanx_right_out[3]
rlabel metal3 49734 7684 49734 7684 0 chanx_right_out[4]
rlabel via2 49174 8381 49174 8381 0 chanx_right_out[5]
rlabel metal2 49174 9265 49174 9265 0 chanx_right_out[6]
rlabel metal3 49734 9724 49734 9724 0 chanx_right_out[7]
rlabel metal2 49174 10489 49174 10489 0 chanx_right_out[8]
rlabel metal3 49734 11084 49734 11084 0 chanx_right_out[9]
rlabel metal2 782 1860 782 1860 0 chany_bottom_in[0]
rlabel metal2 8142 823 8142 823 0 chany_bottom_in[10]
rlabel metal2 8878 1554 8878 1554 0 chany_bottom_in[11]
rlabel metal2 9614 1588 9614 1588 0 chany_bottom_in[12]
rlabel metal1 10396 3026 10396 3026 0 chany_bottom_in[13]
rlabel metal2 11086 1554 11086 1554 0 chany_bottom_in[14]
rlabel metal2 11822 1554 11822 1554 0 chany_bottom_in[15]
rlabel metal1 12650 3026 12650 3026 0 chany_bottom_in[16]
rlabel metal2 13294 1554 13294 1554 0 chany_bottom_in[17]
rlabel metal1 14076 3026 14076 3026 0 chany_bottom_in[18]
rlabel metal2 14766 1588 14766 1588 0 chany_bottom_in[19]
rlabel metal2 1518 1894 1518 1894 0 chany_bottom_in[1]
rlabel metal2 15502 1554 15502 1554 0 chany_bottom_in[20]
rlabel metal2 16238 1554 16238 1554 0 chany_bottom_in[21]
rlabel metal2 16974 1554 16974 1554 0 chany_bottom_in[22]
rlabel metal1 17802 3026 17802 3026 0 chany_bottom_in[23]
rlabel metal2 18446 1622 18446 1622 0 chany_bottom_in[24]
rlabel metal1 19228 2958 19228 2958 0 chany_bottom_in[25]
rlabel metal2 19918 1588 19918 1588 0 chany_bottom_in[26]
rlabel metal2 20654 1860 20654 1860 0 chany_bottom_in[27]
rlabel metal2 21390 1622 21390 1622 0 chany_bottom_in[28]
rlabel metal1 22080 2958 22080 2958 0 chany_bottom_in[29]
rlabel metal2 2254 1588 2254 1588 0 chany_bottom_in[2]
rlabel metal2 2990 1554 2990 1554 0 chany_bottom_in[3]
rlabel metal1 3818 3026 3818 3026 0 chany_bottom_in[4]
rlabel metal2 4462 1554 4462 1554 0 chany_bottom_in[5]
rlabel metal1 5290 3026 5290 3026 0 chany_bottom_in[6]
rlabel metal2 5934 1554 5934 1554 0 chany_bottom_in[7]
rlabel metal1 6762 3026 6762 3026 0 chany_bottom_in[8]
rlabel metal2 7406 1588 7406 1588 0 chany_bottom_in[9]
rlabel metal2 22862 1622 22862 1622 0 chany_bottom_out[0]
rlabel metal2 30222 1622 30222 1622 0 chany_bottom_out[10]
rlabel metal2 30958 2166 30958 2166 0 chany_bottom_out[11]
rlabel metal2 31694 1860 31694 1860 0 chany_bottom_out[12]
rlabel metal2 32430 1826 32430 1826 0 chany_bottom_out[13]
rlabel metal2 33166 1520 33166 1520 0 chany_bottom_out[14]
rlabel metal2 33902 2404 33902 2404 0 chany_bottom_out[15]
rlabel metal2 34638 2166 34638 2166 0 chany_bottom_out[16]
rlabel metal2 35374 1622 35374 1622 0 chany_bottom_out[17]
rlabel metal2 36110 2166 36110 2166 0 chany_bottom_out[18]
rlabel metal2 36846 1860 36846 1860 0 chany_bottom_out[19]
rlabel metal1 23690 2958 23690 2958 0 chany_bottom_out[1]
rlabel metal2 37582 1826 37582 1826 0 chany_bottom_out[20]
rlabel metal2 38318 1622 38318 1622 0 chany_bottom_out[21]
rlabel metal2 39054 2404 39054 2404 0 chany_bottom_out[22]
rlabel metal2 39790 2166 39790 2166 0 chany_bottom_out[23]
rlabel metal2 40526 1622 40526 1622 0 chany_bottom_out[24]
rlabel metal2 41262 2166 41262 2166 0 chany_bottom_out[25]
rlabel metal2 41998 1860 41998 1860 0 chany_bottom_out[26]
rlabel metal2 42734 1826 42734 1826 0 chany_bottom_out[27]
rlabel metal2 43470 2404 43470 2404 0 chany_bottom_out[28]
rlabel metal2 44206 2166 44206 2166 0 chany_bottom_out[29]
rlabel metal1 24702 3570 24702 3570 0 chany_bottom_out[2]
rlabel metal1 25346 2958 25346 2958 0 chany_bottom_out[3]
rlabel metal2 25806 1622 25806 1622 0 chany_bottom_out[4]
rlabel metal2 26542 1622 26542 1622 0 chany_bottom_out[5]
rlabel metal1 27554 2958 27554 2958 0 chany_bottom_out[6]
rlabel metal2 28014 823 28014 823 0 chany_bottom_out[7]
rlabel metal1 29210 2958 29210 2958 0 chany_bottom_out[8]
rlabel metal1 29854 3570 29854 3570 0 chany_bottom_out[9]
rlabel metal2 23230 55711 23230 55711 0 chany_top_in_0[0]
rlabel metal1 30636 54162 30636 54162 0 chany_top_in_0[10]
rlabel metal1 31372 54162 31372 54162 0 chany_top_in_0[11]
rlabel metal1 32200 53550 32200 53550 0 chany_top_in_0[12]
rlabel metal1 32890 54230 32890 54230 0 chany_top_in_0[13]
rlabel metal1 33626 54230 33626 54230 0 chany_top_in_0[14]
rlabel metal1 34592 54162 34592 54162 0 chany_top_in_0[15]
rlabel metal1 35144 53550 35144 53550 0 chany_top_in_0[16]
rlabel metal1 35788 54162 35788 54162 0 chany_top_in_0[17]
rlabel metal1 36524 54162 36524 54162 0 chany_top_in_0[18]
rlabel metal1 37398 54230 37398 54230 0 chany_top_in_0[19]
rlabel metal1 24334 53550 24334 53550 0 chany_top_in_0[1]
rlabel metal2 37950 55711 37950 55711 0 chany_top_in_0[20]
rlabel metal1 38732 54162 38732 54162 0 chany_top_in_0[21]
rlabel metal1 39744 54162 39744 54162 0 chany_top_in_0[22]
rlabel metal1 40480 54162 40480 54162 0 chany_top_in_0[23]
rlabel metal1 41308 54162 41308 54162 0 chany_top_in_0[24]
rlabel metal1 41768 53550 41768 53550 0 chany_top_in_0[25]
rlabel metal1 42550 54230 42550 54230 0 chany_top_in_0[26]
rlabel metal1 43424 54162 43424 54162 0 chany_top_in_0[27]
rlabel metal2 44022 56236 44022 56236 0 chany_top_in_0[28]
rlabel metal1 44988 54162 44988 54162 0 chany_top_in_0[29]
rlabel metal1 24748 54162 24748 54162 0 chany_top_in_0[2]
rlabel metal1 25484 54162 25484 54162 0 chany_top_in_0[3]
rlabel metal2 26174 55209 26174 55209 0 chany_top_in_0[4]
rlabel metal1 27048 54162 27048 54162 0 chany_top_in_0[5]
rlabel metal1 27784 54162 27784 54162 0 chany_top_in_0[6]
rlabel metal1 28566 54230 28566 54230 0 chany_top_in_0[7]
rlabel metal1 29532 53550 29532 53550 0 chany_top_in_0[8]
rlabel metal1 29900 54162 29900 54162 0 chany_top_in_0[9]
rlabel metal1 1610 52530 1610 52530 0 chany_top_out_0[0]
rlabel metal1 8464 54230 8464 54230 0 chany_top_out_0[10]
rlabel metal1 9246 52564 9246 52564 0 chany_top_out_0[11]
rlabel metal1 10120 53006 10120 53006 0 chany_top_out_0[12]
rlabel metal1 10810 53618 10810 53618 0 chany_top_out_0[13]
rlabel metal1 11224 54230 11224 54230 0 chany_top_out_0[14]
rlabel metal1 12466 53618 12466 53618 0 chany_top_out_0[15]
rlabel metal2 12926 55711 12926 55711 0 chany_top_out_0[16]
rlabel metal1 13616 54230 13616 54230 0 chany_top_out_0[17]
rlabel metal1 14674 52530 14674 52530 0 chany_top_out_0[18]
rlabel metal1 15272 53006 15272 53006 0 chany_top_out_0[19]
rlabel metal1 2162 53618 2162 53618 0 chany_top_out_0[1]
rlabel metal1 15870 53652 15870 53652 0 chany_top_out_0[20]
rlabel metal2 16606 55226 16606 55226 0 chany_top_out_0[21]
rlabel metal1 17618 53006 17618 53006 0 chany_top_out_0[22]
rlabel metal2 18262 56236 18262 56236 0 chany_top_out_0[23]
rlabel metal1 18768 54230 18768 54230 0 chany_top_out_0[24]
rlabel metal1 19826 53006 19826 53006 0 chany_top_out_0[25]
rlabel metal1 20378 53618 20378 53618 0 chany_top_out_0[26]
rlabel metal2 21022 55226 21022 55226 0 chany_top_out_0[27]
rlabel metal1 22034 53618 22034 53618 0 chany_top_out_0[28]
rlabel metal1 22770 54094 22770 54094 0 chany_top_out_0[29]
rlabel metal1 2898 53006 2898 53006 0 chany_top_out_0[2]
rlabel metal1 3312 54230 3312 54230 0 chany_top_out_0[3]
rlabel metal1 4370 52530 4370 52530 0 chany_top_out_0[4]
rlabel metal2 4830 55711 4830 55711 0 chany_top_out_0[5]
rlabel metal1 5658 53618 5658 53618 0 chany_top_out_0[6]
rlabel metal1 6072 54230 6072 54230 0 chany_top_out_0[7]
rlabel metal1 7314 53618 7314 53618 0 chany_top_out_0[8]
rlabel metal1 8050 53006 8050 53006 0 chany_top_out_0[9]
rlabel metal2 21482 18496 21482 18496 0 clknet_0_prog_clk
rlabel metal1 13662 8534 13662 8534 0 clknet_4_0_0_prog_clk
rlabel via1 38502 21539 38502 21539 0 clknet_4_10_0_prog_clk
rlabel metal1 39284 32334 39284 32334 0 clknet_4_11_0_prog_clk
rlabel metal1 32430 38250 32430 38250 0 clknet_4_12_0_prog_clk
rlabel metal2 24150 41888 24150 41888 0 clknet_4_13_0_prog_clk
rlabel metal1 42366 37298 42366 37298 0 clknet_4_14_0_prog_clk
rlabel metal1 37490 41650 37490 41650 0 clknet_4_15_0_prog_clk
rlabel metal1 17112 22066 17112 22066 0 clknet_4_1_0_prog_clk
rlabel metal1 32338 18156 32338 18156 0 clknet_4_2_0_prog_clk
rlabel metal2 32522 21760 32522 21760 0 clknet_4_3_0_prog_clk
rlabel metal1 21758 28424 21758 28424 0 clknet_4_4_0_prog_clk
rlabel metal2 22034 35360 22034 35360 0 clknet_4_5_0_prog_clk
rlabel metal2 32338 23392 32338 23392 0 clknet_4_6_0_prog_clk
rlabel metal2 24886 26928 24886 26928 0 clknet_4_7_0_prog_clk
rlabel metal1 34546 18122 34546 18122 0 clknet_4_8_0_prog_clk
rlabel metal1 32246 32334 32246 32334 0 clknet_4_9_0_prog_clk
rlabel metal3 1740 13396 1740 13396 0 gfpga_pad_io_soc_dir[0]
rlabel metal3 1004 15708 1004 15708 0 gfpga_pad_io_soc_dir[1]
rlabel metal3 1004 18020 1004 18020 0 gfpga_pad_io_soc_dir[2]
rlabel metal3 1004 20332 1004 20332 0 gfpga_pad_io_soc_dir[3]
rlabel metal3 820 31892 820 31892 0 gfpga_pad_io_soc_in[0]
rlabel metal3 1234 34204 1234 34204 0 gfpga_pad_io_soc_in[1]
rlabel metal3 820 36516 820 36516 0 gfpga_pad_io_soc_in[2]
rlabel metal3 820 38828 820 38828 0 gfpga_pad_io_soc_in[3]
rlabel metal3 1004 22644 1004 22644 0 gfpga_pad_io_soc_out[0]
rlabel metal3 1004 24956 1004 24956 0 gfpga_pad_io_soc_out[1]
rlabel metal3 1004 27268 1004 27268 0 gfpga_pad_io_soc_out[2]
rlabel metal3 1004 29580 1004 29580 0 gfpga_pad_io_soc_out[3]
rlabel metal3 1188 41140 1188 41140 0 isol_n
rlabel metal2 4002 51000 4002 51000 0 net1
rlabel metal2 49174 36414 49174 36414 0 net10
rlabel metal1 46966 53210 46966 53210 0 net100
rlabel metal1 48622 41582 48622 41582 0 net101
rlabel metal1 48668 41786 48668 41786 0 net102
rlabel metal2 48806 50320 48806 50320 0 net103
rlabel metal1 45172 47430 45172 47430 0 net104
rlabel metal1 45034 48518 45034 48518 0 net105
rlabel metal1 33718 17748 33718 17748 0 net106
rlabel metal2 43286 38080 43286 38080 0 net107
rlabel metal1 42918 39372 42918 39372 0 net108
rlabel metal2 31786 14892 31786 14892 0 net109
rlabel metal2 48806 37026 48806 37026 0 net11
rlabel metal2 33994 18445 33994 18445 0 net110
rlabel metal1 43838 51782 43838 51782 0 net111
rlabel metal1 48024 45458 48024 45458 0 net112
rlabel metal1 48530 45322 48530 45322 0 net113
rlabel metal1 47196 48246 47196 48246 0 net114
rlabel metal2 22540 41684 22540 41684 0 net115
rlabel metal2 1886 43656 1886 43656 0 net116
rlabel metal1 1932 50762 1932 50762 0 net117
rlabel metal2 1748 43316 1748 43316 0 net118
rlabel metal1 18492 18938 18492 18938 0 net119
rlabel metal1 42642 37842 42642 37842 0 net12
rlabel metal2 23782 41820 23782 41820 0 net120
rlabel metal2 44758 12444 44758 12444 0 net121
rlabel metal2 46782 12988 46782 12988 0 net122
rlabel metal1 44022 17782 44022 17782 0 net123
rlabel metal1 44666 17578 44666 17578 0 net124
rlabel metal1 45356 17034 45356 17034 0 net125
rlabel metal1 45034 17646 45034 17646 0 net126
rlabel metal1 46138 18666 46138 18666 0 net127
rlabel metal1 45264 19754 45264 19754 0 net128
rlabel metal2 45126 19516 45126 19516 0 net129
rlabel metal2 49174 37808 49174 37808 0 net13
rlabel metal1 47334 18258 47334 18258 0 net130
rlabel metal1 47104 5678 47104 5678 0 net131
rlabel metal1 46230 18734 46230 18734 0 net132
rlabel metal1 46736 19346 46736 19346 0 net133
rlabel metal1 47932 20434 47932 20434 0 net134
rlabel metal1 47472 20910 47472 20910 0 net135
rlabel metal1 47104 21522 47104 21522 0 net136
rlabel metal1 47794 21998 47794 21998 0 net137
rlabel metal1 47840 23086 47840 23086 0 net138
rlabel metal1 47426 23698 47426 23698 0 net139
rlabel metal2 36570 29529 36570 29529 0 net14
rlabel metal1 47932 24174 47932 24174 0 net140
rlabel metal1 47610 24786 47610 24786 0 net141
rlabel metal1 46966 6766 46966 6766 0 net142
rlabel metal1 47886 7378 47886 7378 0 net143
rlabel metal1 47196 7854 47196 7854 0 net144
rlabel metal1 47242 8466 47242 8466 0 net145
rlabel metal1 47426 9554 47426 9554 0 net146
rlabel metal2 45678 10812 45678 10812 0 net147
rlabel metal1 47702 7242 47702 7242 0 net148
rlabel metal2 44298 11594 44298 11594 0 net149
rlabel via2 48806 39491 48806 39491 0 net15
rlabel metal1 23736 15334 23736 15334 0 net150
rlabel metal1 32292 2414 32292 2414 0 net151
rlabel metal1 30866 3502 30866 3502 0 net152
rlabel metal1 32200 3026 32200 3026 0 net153
rlabel metal1 34132 19754 34132 19754 0 net154
rlabel metal1 34362 2414 34362 2414 0 net155
rlabel metal1 33304 9418 33304 9418 0 net156
rlabel metal1 34592 3502 34592 3502 0 net157
rlabel metal1 36386 2414 36386 2414 0 net158
rlabel metal1 36616 18666 36616 18666 0 net159
rlabel metal2 43746 38080 43746 38080 0 net16
rlabel metal1 37858 8330 37858 8330 0 net160
rlabel metal1 25484 16762 25484 16762 0 net161
rlabel metal1 38364 3094 38364 3094 0 net162
rlabel metal1 40066 14348 40066 14348 0 net163
rlabel metal1 38824 4114 38824 4114 0 net164
rlabel metal1 38686 3502 38686 3502 0 net165
rlabel metal1 42044 2414 42044 2414 0 net166
rlabel metal1 40526 12138 40526 12138 0 net167
rlabel metal1 39698 8398 39698 8398 0 net168
rlabel metal1 41492 6698 41492 6698 0 net169
rlabel via2 48806 40579 48806 40579 0 net17
rlabel metal1 38962 6766 38962 6766 0 net170
rlabel metal1 41492 7242 41492 7242 0 net171
rlabel metal1 25300 3502 25300 3502 0 net172
rlabel metal2 25162 6766 25162 6766 0 net173
rlabel metal1 26312 12614 26312 12614 0 net174
rlabel metal1 27692 12682 27692 12682 0 net175
rlabel metal2 29256 13804 29256 13804 0 net176
rlabel metal2 29946 6154 29946 6154 0 net177
rlabel metal2 29210 7582 29210 7582 0 net178
rlabel metal1 29486 13838 29486 13838 0 net179
rlabel metal1 45540 41072 45540 41072 0 net18
rlabel metal1 2760 52462 2760 52462 0 net180
rlabel metal1 12650 43962 12650 43962 0 net181
rlabel metal1 12006 52462 12006 52462 0 net182
rlabel metal1 12098 44506 12098 44506 0 net183
rlabel metal1 12788 45526 12788 45526 0 net184
rlabel metal1 15456 43962 15456 43962 0 net185
rlabel metal1 13570 53550 13570 53550 0 net186
rlabel metal2 16974 48552 16974 48552 0 net187
rlabel metal1 15962 42330 15962 42330 0 net188
rlabel metal2 19182 47940 19182 47940 0 net189
rlabel metal1 47564 42194 47564 42194 0 net19
rlabel metal1 15134 53074 15134 53074 0 net190
rlabel metal1 2162 53516 2162 53516 0 net191
rlabel metal2 20470 48688 20470 48688 0 net192
rlabel metal2 20378 44479 20378 44479 0 net193
rlabel metal1 17618 53108 17618 53108 0 net194
rlabel metal1 18078 53550 18078 53550 0 net195
rlabel metal2 17710 52326 17710 52326 0 net196
rlabel metal1 21298 43894 21298 43894 0 net197
rlabel metal1 20194 53516 20194 53516 0 net198
rlabel metal1 20332 54162 20332 54162 0 net199
rlabel metal1 3588 3706 3588 3706 0 net2
rlabel metal1 40526 42568 40526 42568 0 net20
rlabel metal1 23782 51578 23782 51578 0 net200
rlabel metal1 23184 52122 23184 52122 0 net201
rlabel metal1 2898 53108 2898 53108 0 net202
rlabel metal1 2254 54128 2254 54128 0 net203
rlabel metal1 6808 52462 6808 52462 0 net204
rlabel metal1 5865 53074 5865 53074 0 net205
rlabel metal1 6187 53550 6187 53550 0 net206
rlabel metal1 4830 54230 4830 54230 0 net207
rlabel metal1 10580 43418 10580 43418 0 net208
rlabel metal1 8878 53074 8878 53074 0 net209
rlabel metal2 41446 39202 41446 39202 0 net21
rlabel metal1 3726 13906 3726 13906 0 net210
rlabel metal1 3772 18598 3772 18598 0 net211
rlabel metal1 2346 18258 2346 18258 0 net212
rlabel metal1 2300 20434 2300 20434 0 net213
rlabel metal1 2668 23086 2668 23086 0 net214
rlabel metal1 2990 25262 2990 25262 0 net215
rlabel metal1 3358 27438 3358 27438 0 net216
rlabel metal2 4922 28900 4922 28900 0 net217
rlabel metal2 47794 3162 47794 3162 0 net218
rlabel metal2 48622 45764 48622 45764 0 net219
rlabel metal1 48806 43724 48806 43724 0 net22
rlabel metal2 46138 53380 46138 53380 0 net220
rlabel metal1 47886 3060 47886 3060 0 net221
rlabel metal1 47932 54162 47932 54162 0 net222
rlabel metal1 47840 3502 47840 3502 0 net223
rlabel metal1 48254 53074 48254 53074 0 net224
rlabel metal1 30590 20502 30590 20502 0 net225
rlabel metal1 29026 27438 29026 27438 0 net226
rlabel metal1 42918 31450 42918 31450 0 net227
rlabel metal1 39422 23086 39422 23086 0 net228
rlabel metal1 32108 36142 32108 36142 0 net229
rlabel metal1 42067 44846 42067 44846 0 net23
rlabel metal1 31970 22610 31970 22610 0 net230
rlabel metal1 38870 28526 38870 28526 0 net231
rlabel metal1 31234 33490 31234 33490 0 net232
rlabel metal1 32614 34170 32614 34170 0 net233
rlabel metal1 32246 35666 32246 35666 0 net234
rlabel metal1 29670 37230 29670 37230 0 net235
rlabel metal2 27370 36550 27370 36550 0 net236
rlabel metal1 41906 34578 41906 34578 0 net237
rlabel metal1 28750 32334 28750 32334 0 net238
rlabel metal1 26220 29614 26220 29614 0 net239
rlabel metal1 43286 37978 43286 37978 0 net24
rlabel metal1 26542 25874 26542 25874 0 net240
rlabel metal2 25806 25296 25806 25296 0 net241
rlabel metal2 24978 23290 24978 23290 0 net242
rlabel metal1 25438 23732 25438 23732 0 net243
rlabel metal1 24794 25874 24794 25874 0 net244
rlabel metal2 23138 27268 23138 27268 0 net245
rlabel metal1 13938 11118 13938 11118 0 net246
rlabel metal2 30222 14586 30222 14586 0 net247
rlabel metal1 34914 32878 34914 32878 0 net248
rlabel metal2 32246 14790 32246 14790 0 net249
rlabel metal1 32890 25942 32890 25942 0 net25
rlabel metal2 33442 15674 33442 15674 0 net250
rlabel metal1 35604 17170 35604 17170 0 net251
rlabel metal1 37996 16422 37996 16422 0 net252
rlabel metal1 33856 16082 33856 16082 0 net253
rlabel metal1 38088 14382 38088 14382 0 net254
rlabel metal1 36800 12954 36800 12954 0 net255
rlabel metal1 37766 15130 37766 15130 0 net256
rlabel metal1 40618 36074 40618 36074 0 net257
rlabel metal2 38870 39236 38870 39236 0 net258
rlabel metal2 22862 36346 22862 36346 0 net259
rlabel metal1 35052 25806 35052 25806 0 net26
rlabel metal2 21850 31246 21850 31246 0 net260
rlabel metal1 24334 31450 24334 31450 0 net261
rlabel metal2 31326 37434 31326 37434 0 net262
rlabel metal1 23920 30226 23920 30226 0 net263
rlabel metal1 18216 32402 18216 32402 0 net264
rlabel metal2 22494 37434 22494 37434 0 net265
rlabel metal1 26496 35054 26496 35054 0 net266
rlabel metal1 24242 37230 24242 37230 0 net267
rlabel metal2 29118 33796 29118 33796 0 net268
rlabel metal1 21942 31314 21942 31314 0 net269
rlabel metal1 39284 33558 39284 33558 0 net27
rlabel via2 49358 4981 49358 4981 0 net270
rlabel metal1 24518 25262 24518 25262 0 net271
rlabel metal1 25484 22610 25484 22610 0 net272
rlabel metal2 23322 17476 23322 17476 0 net273
rlabel metal2 22678 25466 22678 25466 0 net274
rlabel metal1 29210 21658 29210 21658 0 net275
rlabel metal2 29118 24786 29118 24786 0 net276
rlabel metal2 36938 25432 36938 25432 0 net277
rlabel metal1 40342 24786 40342 24786 0 net278
rlabel metal1 36432 28526 36432 28526 0 net279
rlabel metal1 39100 34986 39100 34986 0 net28
rlabel metal1 37490 34034 37490 34034 0 net29
rlabel metal1 37766 24174 37766 24174 0 net3
rlabel metal2 43516 32164 43516 32164 0 net30
rlabel metal1 34638 37094 34638 37094 0 net31
rlabel metal2 41538 32164 41538 32164 0 net32
rlabel metal1 2346 3128 2346 3128 0 net33
rlabel metal2 21942 40052 21942 40052 0 net34
rlabel metal2 13478 43418 13478 43418 0 net35
rlabel metal2 10074 3706 10074 3706 0 net36
rlabel metal1 12558 3162 12558 3162 0 net37
rlabel metal2 14950 41276 14950 41276 0 net38
rlabel metal2 21022 43520 21022 43520 0 net39
rlabel metal2 48806 32742 48806 32742 0 net4
rlabel metal2 12926 3230 12926 3230 0 net40
rlabel metal1 18446 43690 18446 43690 0 net41
rlabel metal1 17342 42194 17342 42194 0 net42
rlabel metal1 16652 2618 16652 2618 0 net43
rlabel metal1 1794 2924 1794 2924 0 net44
rlabel metal2 17342 2108 17342 2108 0 net45
rlabel metal1 20424 43690 20424 43690 0 net46
rlabel metal2 17434 2074 17434 2074 0 net47
rlabel metal1 18308 3026 18308 3026 0 net48
rlabel metal1 33718 17646 33718 17646 0 net49
rlabel metal2 49174 32504 49174 32504 0 net5
rlabel metal1 19550 2924 19550 2924 0 net50
rlabel metal1 22494 43690 22494 43690 0 net51
rlabel metal1 20930 3094 20930 3094 0 net52
rlabel metal1 25691 2346 25691 2346 0 net53
rlabel metal1 33672 17170 33672 17170 0 net54
rlabel metal2 2438 2074 2438 2074 0 net55
rlabel metal1 7958 42160 7958 42160 0 net56
rlabel metal1 17710 2856 17710 2856 0 net57
rlabel metal2 21160 6900 21160 6900 0 net58
rlabel metal2 5750 2975 5750 2975 0 net59
rlabel metal1 48898 33830 48898 33830 0 net6
rlabel metal2 10718 35700 10718 35700 0 net60
rlabel metal2 20010 5031 20010 5031 0 net61
rlabel metal2 21574 37808 21574 37808 0 net62
rlabel metal1 25392 53686 25392 53686 0 net63
rlabel metal1 30820 53958 30820 53958 0 net64
rlabel metal1 28934 43860 28934 43860 0 net65
rlabel metal1 33028 45526 33028 45526 0 net66
rlabel via2 41814 36227 41814 36227 0 net67
rlabel metal1 33948 19822 33948 19822 0 net68
rlabel metal1 33856 44778 33856 44778 0 net69
rlabel metal1 49174 34476 49174 34476 0 net7
rlabel metal1 35236 53414 35236 53414 0 net70
rlabel metal1 36294 53958 36294 53958 0 net71
rlabel metal2 36754 48824 36754 48824 0 net72
rlabel metal1 36662 18598 36662 18598 0 net73
rlabel metal1 24932 53482 24932 53482 0 net74
rlabel metal1 37352 53414 37352 53414 0 net75
rlabel metal2 36938 18258 36938 18258 0 net76
rlabel metal1 36386 20774 36386 20774 0 net77
rlabel metal1 41446 42194 41446 42194 0 net78
rlabel metal1 39652 43758 39652 43758 0 net79
rlabel metal2 43654 34782 43654 34782 0 net8
rlabel metal1 39974 44506 39974 44506 0 net80
rlabel metal3 38755 12308 38755 12308 0 net81
rlabel metal1 40986 54026 40986 54026 0 net82
rlabel metal1 42366 42670 42366 42670 0 net83
rlabel metal2 41630 43935 41630 43935 0 net84
rlabel metal3 25047 53924 25047 53924 0 net85
rlabel metal1 25576 13294 25576 13294 0 net86
rlabel metal1 28198 43690 28198 43690 0 net87
rlabel metal1 27416 53958 27416 53958 0 net88
rlabel metal1 28336 53958 28336 53958 0 net89
rlabel metal2 41998 34238 41998 34238 0 net9
rlabel metal1 29302 54026 29302 54026 0 net90
rlabel metal1 31234 45458 31234 45458 0 net91
rlabel metal1 30084 53958 30084 53958 0 net92
rlabel metal2 7682 26047 7682 26047 0 net93
rlabel metal2 7866 30838 7866 30838 0 net94
rlabel metal1 4600 36550 4600 36550 0 net95
rlabel metal1 4508 38726 4508 38726 0 net96
rlabel metal2 10626 24718 10626 24718 0 net97
rlabel metal1 38555 18666 38555 18666 0 net98
rlabel metal2 2070 43520 2070 43520 0 net99
rlabel metal2 44942 2115 44942 2115 0 prog_clk
rlabel metal2 45678 1554 45678 1554 0 prog_reset_bottom_in
rlabel metal2 46414 1792 46414 1792 0 prog_reset_bottom_out
rlabel metal3 820 43452 820 43452 0 prog_reset_left_in
rlabel metal3 49734 45764 49734 45764 0 prog_reset_right_out
rlabel metal1 47380 54162 47380 54162 0 prog_reset_top_in
rlabel metal1 47058 53618 47058 53618 0 prog_reset_top_out
rlabel metal2 47150 1894 47150 1894 0 reset_bottom_in
rlabel metal2 47886 1860 47886 1860 0 reset_bottom_out
rlabel metal2 49358 46495 49358 46495 0 reset_right_in
rlabel metal1 49128 53550 49128 53550 0 reset_top_in
rlabel metal2 48300 54604 48300 54604 0 reset_top_out
rlabel metal2 49082 47379 49082 47379 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_
rlabel metal2 49082 48263 49082 48263 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_
rlabel metal1 49174 49198 49174 49198 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_
rlabel metal1 49128 49810 49128 49810 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_
rlabel metal2 49082 50065 49082 50065 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_
rlabel metal2 48990 50711 48990 50711 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_
rlabel metal2 49082 51289 49082 51289 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_
rlabel metal2 49082 51935 49082 51935 0 right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_
rlabel metal3 2062 4148 2062 4148 0 right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 2062 6460 2062 6460 0 right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 2016 8772 2016 8772 0 right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 2016 11084 2016 11084 0 right_width_0_height_0_subtile_3__pin_inpad_0_
rlabel metal1 36800 16422 36800 16422 0 sb_0__1_.mem_bottom_track_1.ccff_head
rlabel metal2 31786 21216 31786 21216 0 sb_0__1_.mem_bottom_track_1.ccff_tail
rlabel metal1 33764 19890 33764 19890 0 sb_0__1_.mem_bottom_track_1.mem_out\[0\]
rlabel metal2 31878 24310 31878 24310 0 sb_0__1_.mem_bottom_track_1.mem_out\[1\]
rlabel metal2 34270 23698 34270 23698 0 sb_0__1_.mem_bottom_track_11.ccff_head
rlabel metal1 33258 26554 33258 26554 0 sb_0__1_.mem_bottom_track_11.ccff_tail
rlabel metal2 38962 31654 38962 31654 0 sb_0__1_.mem_bottom_track_11.mem_out\[0\]
rlabel metal2 32430 26044 32430 26044 0 sb_0__1_.mem_bottom_track_11.mem_out\[1\]
rlabel metal2 39514 25874 39514 25874 0 sb_0__1_.mem_bottom_track_13.ccff_tail
rlabel metal1 37490 32742 37490 32742 0 sb_0__1_.mem_bottom_track_13.mem_out\[0\]
rlabel metal1 38640 27574 38640 27574 0 sb_0__1_.mem_bottom_track_13.mem_out\[1\]
rlabel metal2 40434 26690 40434 26690 0 sb_0__1_.mem_bottom_track_21.ccff_tail
rlabel metal1 37766 26418 37766 26418 0 sb_0__1_.mem_bottom_track_21.mem_out\[0\]
rlabel metal2 40710 27846 40710 27846 0 sb_0__1_.mem_bottom_track_21.mem_out\[1\]
rlabel metal1 35466 29274 35466 29274 0 sb_0__1_.mem_bottom_track_29.ccff_tail
rlabel metal1 40802 34442 40802 34442 0 sb_0__1_.mem_bottom_track_29.mem_out\[0\]
rlabel metal1 36110 31858 36110 31858 0 sb_0__1_.mem_bottom_track_29.mem_out\[1\]
rlabel metal1 33672 20366 33672 20366 0 sb_0__1_.mem_bottom_track_3.ccff_tail
rlabel metal1 33856 26894 33856 26894 0 sb_0__1_.mem_bottom_track_3.mem_out\[0\]
rlabel metal1 32522 21454 32522 21454 0 sb_0__1_.mem_bottom_track_3.mem_out\[1\]
rlabel metal1 31510 27914 31510 27914 0 sb_0__1_.mem_bottom_track_37.ccff_tail
rlabel metal1 35604 32266 35604 32266 0 sb_0__1_.mem_bottom_track_37.mem_out\[0\]
rlabel metal1 34638 32266 34638 32266 0 sb_0__1_.mem_bottom_track_37.mem_out\[1\]
rlabel metal1 40618 32198 40618 32198 0 sb_0__1_.mem_bottom_track_45.ccff_tail
rlabel metal2 41906 34816 41906 34816 0 sb_0__1_.mem_bottom_track_45.mem_out\[0\]
rlabel metal1 42136 33286 42136 33286 0 sb_0__1_.mem_bottom_track_45.mem_out\[1\]
rlabel metal1 38134 20978 38134 20978 0 sb_0__1_.mem_bottom_track_5.ccff_tail
rlabel metal1 37214 22066 37214 22066 0 sb_0__1_.mem_bottom_track_5.mem_out\[0\]
rlabel metal1 39652 23494 39652 23494 0 sb_0__1_.mem_bottom_track_5.mem_out\[1\]
rlabel metal1 21659 41786 21659 41786 0 sb_0__1_.mem_bottom_track_53.mem_out\[0\]
rlabel metal1 35604 28594 35604 28594 0 sb_0__1_.mem_bottom_track_7.mem_out\[0\]
rlabel metal1 35236 23630 35236 23630 0 sb_0__1_.mem_bottom_track_7.mem_out\[1\]
rlabel metal1 33948 35258 33948 35258 0 sb_0__1_.mem_right_track_0.ccff_head
rlabel metal1 42458 31858 42458 31858 0 sb_0__1_.mem_right_track_0.ccff_tail
rlabel metal1 38778 31280 38778 31280 0 sb_0__1_.mem_right_track_0.mem_out\[0\]
rlabel metal1 40388 30022 40388 30022 0 sb_0__1_.mem_right_track_0.mem_out\[1\]
rlabel metal1 39468 42126 39468 42126 0 sb_0__1_.mem_right_track_10.ccff_head
rlabel metal1 37030 41514 37030 41514 0 sb_0__1_.mem_right_track_10.ccff_tail
rlabel metal1 38134 43826 38134 43826 0 sb_0__1_.mem_right_track_10.mem_out\[0\]
rlabel metal1 35328 38250 35328 38250 0 sb_0__1_.mem_right_track_10.mem_out\[1\]
rlabel metal1 35512 41446 35512 41446 0 sb_0__1_.mem_right_track_12.ccff_tail
rlabel metal1 36432 42738 36432 42738 0 sb_0__1_.mem_right_track_12.mem_out\[0\]
rlabel metal1 37122 42534 37122 42534 0 sb_0__1_.mem_right_track_12.mem_out\[1\]
rlabel metal1 35052 40902 35052 40902 0 sb_0__1_.mem_right_track_14.ccff_tail
rlabel metal2 35558 43350 35558 43350 0 sb_0__1_.mem_right_track_14.mem_out\[0\]
rlabel metal1 33166 41174 33166 41174 0 sb_0__1_.mem_right_track_14.mem_out\[1\]
rlabel metal1 33626 41446 33626 41446 0 sb_0__1_.mem_right_track_16.ccff_tail
rlabel metal1 33120 43214 33120 43214 0 sb_0__1_.mem_right_track_16.mem_out\[0\]
rlabel metal1 31464 41514 31464 41514 0 sb_0__1_.mem_right_track_16.mem_out\[1\]
rlabel metal1 31832 41990 31832 41990 0 sb_0__1_.mem_right_track_18.ccff_tail
rlabel metal1 32246 43826 32246 43826 0 sb_0__1_.mem_right_track_18.mem_out\[0\]
rlabel metal1 30314 42296 30314 42296 0 sb_0__1_.mem_right_track_18.mem_out\[1\]
rlabel metal1 43148 37094 43148 37094 0 sb_0__1_.mem_right_track_2.ccff_tail
rlabel metal1 42872 42126 42872 42126 0 sb_0__1_.mem_right_track_2.mem_out\[0\]
rlabel metal1 43286 36210 43286 36210 0 sb_0__1_.mem_right_track_2.mem_out\[1\]
rlabel metal1 29992 34510 29992 34510 0 sb_0__1_.mem_right_track_20.ccff_tail
rlabel via1 29026 43843 29026 43843 0 sb_0__1_.mem_right_track_20.mem_out\[0\]
rlabel metal1 32223 37298 32223 37298 0 sb_0__1_.mem_right_track_20.mem_out\[1\]
rlabel metal2 28842 29920 28842 29920 0 sb_0__1_.mem_right_track_22.ccff_tail
rlabel metal1 28152 35258 28152 35258 0 sb_0__1_.mem_right_track_22.mem_out\[0\]
rlabel metal1 30498 33388 30498 33388 0 sb_0__1_.mem_right_track_22.mem_out\[1\]
rlabel metal1 29026 26894 29026 26894 0 sb_0__1_.mem_right_track_24.ccff_tail
rlabel metal1 27968 28118 27968 28118 0 sb_0__1_.mem_right_track_24.mem_out\[0\]
rlabel metal1 30038 25670 30038 25670 0 sb_0__1_.mem_right_track_26.ccff_tail
rlabel metal1 32131 29682 32131 29682 0 sb_0__1_.mem_right_track_26.mem_out\[0\]
rlabel metal1 28244 22542 28244 22542 0 sb_0__1_.mem_right_track_28.ccff_tail
rlabel metal2 31142 25772 31142 25772 0 sb_0__1_.mem_right_track_28.mem_out\[0\]
rlabel metal1 30314 24276 30314 24276 0 sb_0__1_.mem_right_track_30.ccff_tail
rlabel metal1 27600 24242 27600 24242 0 sb_0__1_.mem_right_track_30.mem_out\[0\]
rlabel metal1 26956 27302 26956 27302 0 sb_0__1_.mem_right_track_32.ccff_tail
rlabel metal1 28888 25466 28888 25466 0 sb_0__1_.mem_right_track_32.mem_out\[0\]
rlabel metal1 24288 27846 24288 27846 0 sb_0__1_.mem_right_track_34.ccff_tail
rlabel metal1 26910 28186 26910 28186 0 sb_0__1_.mem_right_track_34.mem_out\[0\]
rlabel metal1 21160 14926 21160 14926 0 sb_0__1_.mem_right_track_36.ccff_tail
rlabel metal1 23736 26486 23736 26486 0 sb_0__1_.mem_right_track_36.mem_out\[0\]
rlabel metal1 16698 11186 16698 11186 0 sb_0__1_.mem_right_track_36.mem_out\[1\]
rlabel metal1 28060 14586 28060 14586 0 sb_0__1_.mem_right_track_38.ccff_tail
rlabel metal2 26174 15164 26174 15164 0 sb_0__1_.mem_right_track_38.mem_out\[0\]
rlabel metal2 39974 36244 39974 36244 0 sb_0__1_.mem_right_track_4.ccff_tail
rlabel metal1 43102 36720 43102 36720 0 sb_0__1_.mem_right_track_4.mem_out\[0\]
rlabel metal1 40480 37298 40480 37298 0 sb_0__1_.mem_right_track_4.mem_out\[1\]
rlabel metal2 32890 15402 32890 15402 0 sb_0__1_.mem_right_track_40.ccff_tail
rlabel metal1 29164 16014 29164 16014 0 sb_0__1_.mem_right_track_40.mem_out\[0\]
rlabel metal1 32706 17102 32706 17102 0 sb_0__1_.mem_right_track_44.ccff_tail
rlabel metal2 30314 16218 30314 16218 0 sb_0__1_.mem_right_track_44.mem_out\[0\]
rlabel metal1 35052 18190 35052 18190 0 sb_0__1_.mem_right_track_46.ccff_tail
rlabel metal2 32614 18564 32614 18564 0 sb_0__1_.mem_right_track_46.mem_out\[0\]
rlabel metal1 37260 17850 37260 17850 0 sb_0__1_.mem_right_track_48.ccff_tail
rlabel metal2 36110 17816 36110 17816 0 sb_0__1_.mem_right_track_48.mem_out\[0\]
rlabel metal1 38318 18190 38318 18190 0 sb_0__1_.mem_right_track_50.ccff_tail
rlabel metal1 37674 19278 37674 19278 0 sb_0__1_.mem_right_track_50.mem_out\[0\]
rlabel metal2 37720 14450 37720 14450 0 sb_0__1_.mem_right_track_52.ccff_tail
rlabel metal2 37122 17170 37122 17170 0 sb_0__1_.mem_right_track_52.mem_out\[0\]
rlabel metal1 36478 12818 36478 12818 0 sb_0__1_.mem_right_track_54.ccff_tail
rlabel metal2 33994 13668 33994 13668 0 sb_0__1_.mem_right_track_54.mem_out\[0\]
rlabel metal1 35098 16626 35098 16626 0 sb_0__1_.mem_right_track_56.mem_out\[0\]
rlabel metal1 43056 38522 43056 38522 0 sb_0__1_.mem_right_track_6.ccff_tail
rlabel metal1 40572 43214 40572 43214 0 sb_0__1_.mem_right_track_6.mem_out\[0\]
rlabel metal1 41768 38250 41768 38250 0 sb_0__1_.mem_right_track_6.mem_out\[1\]
rlabel metal2 39330 42851 39330 42851 0 sb_0__1_.mem_right_track_8.mem_out\[0\]
rlabel metal1 39698 40562 39698 40562 0 sb_0__1_.mem_right_track_8.mem_out\[1\]
rlabel metal2 27370 43044 27370 43044 0 sb_0__1_.mem_top_track_0.ccff_tail
rlabel metal2 22172 41548 22172 41548 0 sb_0__1_.mem_top_track_0.mem_out\[0\]
rlabel metal2 25898 42466 25898 42466 0 sb_0__1_.mem_top_track_0.mem_out\[1\]
rlabel metal1 24932 37638 24932 37638 0 sb_0__1_.mem_top_track_10.ccff_head
rlabel metal1 23828 35802 23828 35802 0 sb_0__1_.mem_top_track_10.ccff_tail
rlabel metal2 36202 35649 36202 35649 0 sb_0__1_.mem_top_track_10.mem_out\[0\]
rlabel metal1 23736 35190 23736 35190 0 sb_0__1_.mem_top_track_10.mem_out\[1\]
rlabel metal1 25484 32538 25484 32538 0 sb_0__1_.mem_top_track_12.ccff_tail
rlabel metal2 35834 32853 35834 32853 0 sb_0__1_.mem_top_track_12.mem_out\[0\]
rlabel metal1 26680 31450 26680 31450 0 sb_0__1_.mem_top_track_12.mem_out\[1\]
rlabel metal1 30038 41004 30038 41004 0 sb_0__1_.mem_top_track_2.ccff_tail
rlabel metal1 29670 41990 29670 41990 0 sb_0__1_.mem_top_track_2.mem_out\[0\]
rlabel metal1 32568 39474 32568 39474 0 sb_0__1_.mem_top_track_2.mem_out\[1\]
rlabel metal2 23966 33014 23966 33014 0 sb_0__1_.mem_top_track_20.ccff_tail
rlabel metal1 27830 31892 27830 31892 0 sb_0__1_.mem_top_track_20.mem_out\[0\]
rlabel metal2 29026 32759 29026 32759 0 sb_0__1_.mem_top_track_20.mem_out\[1\]
rlabel metal1 20746 36686 20746 36686 0 sb_0__1_.mem_top_track_28.ccff_tail
rlabel metal2 28658 34034 28658 34034 0 sb_0__1_.mem_top_track_28.mem_out\[0\]
rlabel metal1 18860 35598 18860 35598 0 sb_0__1_.mem_top_track_28.mem_out\[1\]
rlabel metal2 25070 40596 25070 40596 0 sb_0__1_.mem_top_track_36.ccff_tail
rlabel metal1 26680 39474 26680 39474 0 sb_0__1_.mem_top_track_36.mem_out\[0\]
rlabel metal2 23598 38624 23598 38624 0 sb_0__1_.mem_top_track_36.mem_out\[1\]
rlabel metal1 27646 37774 27646 37774 0 sb_0__1_.mem_top_track_4.ccff_tail
rlabel metal1 32982 38828 32982 38828 0 sb_0__1_.mem_top_track_4.mem_out\[0\]
rlabel metal1 32338 36652 32338 36652 0 sb_0__1_.mem_top_track_4.mem_out\[1\]
rlabel metal1 32154 39916 32154 39916 0 sb_0__1_.mem_top_track_44.ccff_tail
rlabel metal2 32890 37638 32890 37638 0 sb_0__1_.mem_top_track_44.mem_out\[0\]
rlabel metal2 43194 38080 43194 38080 0 sb_0__1_.mem_top_track_52.mem_out\[0\]
rlabel metal1 32430 35122 32430 35122 0 sb_0__1_.mem_top_track_52.mem_out\[1\]
rlabel metal1 25024 35734 25024 35734 0 sb_0__1_.mem_top_track_6.mem_out\[0\]
rlabel metal1 27370 38386 27370 38386 0 sb_0__1_.mem_top_track_6.mem_out\[1\]
rlabel metal1 29946 17510 29946 17510 0 sb_0__1_.mux_bottom_track_1.out
rlabel metal1 32200 25262 32200 25262 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33442 25194 33442 25194 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 25622 21726 25622 21726 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 31050 20774 31050 20774 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 30682 21114 30682 21114 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 30176 17578 30176 17578 0 sb_0__1_.mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 31786 10302 31786 10302 0 sb_0__1_.mux_bottom_track_11.out
rlabel metal1 33488 28594 33488 28594 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36018 33082 36018 33082 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31878 26010 31878 26010 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29578 25126 29578 25126 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 32890 25483 32890 25483 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 30958 25296 30958 25296 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 32476 17170 32476 17170 0 sb_0__1_.mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 35466 9622 35466 9622 0 sb_0__1_.mux_bottom_track_13.out
rlabel metal2 37398 29308 37398 29308 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40296 32742 40296 32742 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36524 25330 36524 25330 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 37582 24786 37582 24786 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37214 24922 37214 24922 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36248 24582 36248 24582 0 sb_0__1_.mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 37858 12206 37858 12206 0 sb_0__1_.mux_bottom_track_21.out
rlabel metal1 40526 28628 40526 28628 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41308 32742 41308 32742 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 40526 25942 40526 25942 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40434 24242 40434 24242 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 40250 24174 40250 24174 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 39468 16082 39468 16082 0 sb_0__1_.mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 32062 20774 32062 20774 0 sb_0__1_.mux_bottom_track_29.out
rlabel metal1 34960 31858 34960 31858 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37996 31722 37996 31722 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37812 28186 37812 28186 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35328 31926 35328 31926 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 35374 27370 35374 27370 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33718 20910 33718 20910 0 sb_0__1_.mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 35006 6698 35006 6698 0 sb_0__1_.mux_bottom_track_3.out
rlabel metal2 33994 26044 33994 26044 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33902 25330 33902 25330 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32844 20570 32844 20570 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32269 20502 32269 20502 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 32476 20230 32476 20230 0 sb_0__1_.mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 28474 21386 28474 21386 0 sb_0__1_.mux_bottom_track_37.out
rlabel metal1 35420 32470 35420 32470 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35834 32538 35834 32538 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33442 32198 33442 32198 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28612 27574 28612 27574 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 29486 21114 29486 21114 0 sb_0__1_.mux_bottom_track_37.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 33764 19958 33764 19958 0 sb_0__1_.mux_bottom_track_45.out
rlabel metal1 42090 33830 42090 33830 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40802 33830 40802 33830 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 39698 30090 39698 30090 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 36294 19822 36294 19822 0 sb_0__1_.mux_bottom_track_45.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 37260 6766 37260 6766 0 sb_0__1_.mux_bottom_track_5.out
rlabel metal1 39468 25874 39468 25874 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39698 26010 39698 26010 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38042 23018 38042 23018 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38318 20808 38318 20808 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 38272 20910 38272 20910 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 36570 20842 36570 20842 0 sb_0__1_.mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 23828 17306 23828 17306 0 sb_0__1_.mux_bottom_track_53.out
rlabel metal1 30406 36720 30406 36720 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 27462 36516 27462 36516 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25714 36550 25714 36550 0 sb_0__1_.mux_bottom_track_53.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32384 17068 32384 17068 0 sb_0__1_.mux_bottom_track_7.out
rlabel metal1 35236 25194 35236 25194 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36018 25126 36018 25126 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 34454 23766 34454 23766 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32706 23188 32706 23188 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 34684 22678 34684 22678 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 34316 22746 34316 22746 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 33028 22406 33028 22406 0 sb_0__1_.mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 45632 26350 45632 26350 0 sb_0__1_.mux_right_track_0.out
rlabel metal1 40296 30770 40296 30770 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40434 30906 40434 30906 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 41262 29920 41262 29920 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 39928 28730 39928 28730 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 44022 28220 44022 28220 0 sb_0__1_.mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 41354 30600 41354 30600 0 sb_0__1_.mux_right_track_10.out
rlabel metal1 37628 39066 37628 39066 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37674 37978 37674 37978 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36984 35054 36984 35054 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36386 34510 36386 34510 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 41538 31178 41538 31178 0 sb_0__1_.mux_right_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 44804 25942 44804 25942 0 sb_0__1_.mux_right_track_12.out
rlabel metal1 36432 39066 36432 39066 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 36616 36210 36616 36210 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33396 34714 33396 34714 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 41906 30702 41906 30702 0 sb_0__1_.mux_right_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 42826 31144 42826 31144 0 sb_0__1_.mux_right_track_14.out
rlabel metal1 35190 39066 35190 39066 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35282 36210 35282 36210 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 32752 35802 32752 35802 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35972 36006 35972 36006 0 sb_0__1_.mux_right_track_14.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 41400 31994 41400 31994 0 sb_0__1_.mux_right_track_16.out
rlabel metal1 33810 40562 33810 40562 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 33948 37978 33948 37978 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33902 37774 33902 37774 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 34362 34816 34362 34816 0 sb_0__1_.mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 39698 31212 39698 31212 0 sb_0__1_.mux_right_track_18.out
rlabel metal1 32522 45254 32522 45254 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 33350 39406 33350 39406 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 29670 37145 29670 37145 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 36432 32436 36432 32436 0 sb_0__1_.mux_right_track_18.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 48024 28050 48024 28050 0 sb_0__1_.mux_right_track_2.out
rlabel metal1 43286 36142 43286 36142 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 42918 35734 42918 35734 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 38686 33592 38686 33592 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42688 36006 42688 36006 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 42412 34714 42412 34714 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 43976 34510 43976 34510 0 sb_0__1_.mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 38410 24990 38410 24990 0 sb_0__1_.mux_right_track_20.out
rlabel metal1 30268 43962 30268 43962 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 31372 32946 31372 32946 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 31326 32640 31326 32640 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 32476 29546 32476 29546 0 sb_0__1_.mux_right_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 43838 21760 43838 21760 0 sb_0__1_.mux_right_track_22.out
rlabel metal1 29992 33422 29992 33422 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 30176 29682 30176 29682 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 27738 29546 27738 29546 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 33810 27574 33810 27574 0 sb_0__1_.mux_right_track_22.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 42688 19822 42688 19822 0 sb_0__1_.mux_right_track_24.out
rlabel metal1 30912 26418 30912 26418 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29762 26282 29762 26282 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 33994 22984 33994 22984 0 sb_0__1_.mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42780 18734 42780 18734 0 sb_0__1_.mux_right_track_26.out
rlabel metal2 31786 27370 31786 27370 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27232 24582 27232 24582 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36938 21896 36938 21896 0 sb_0__1_.mux_right_track_26.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 44482 17544 44482 17544 0 sb_0__1_.mux_right_track_28.out
rlabel metal1 30314 22746 30314 22746 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27324 22746 27324 22746 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35742 20434 35742 20434 0 sb_0__1_.mux_right_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 43746 19142 43746 19142 0 sb_0__1_.mux_right_track_30.out
rlabel metal2 30222 25772 30222 25772 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 29210 24038 29210 24038 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 36846 20944 36846 20944 0 sb_0__1_.mux_right_track_30.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 37122 19550 37122 19550 0 sb_0__1_.mux_right_track_32.out
rlabel metal1 28934 25262 28934 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 28520 25262 28520 25262 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 32246 25024 32246 25024 0 sb_0__1_.mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38594 21352 38594 21352 0 sb_0__1_.mux_right_track_34.out
rlabel metal1 27600 25874 27600 25874 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 25852 26010 25852 26010 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 35374 21284 35374 21284 0 sb_0__1_.mux_right_track_34.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 38226 13872 38226 13872 0 sb_0__1_.mux_right_track_36.out
rlabel metal1 21482 19720 21482 19720 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 20148 15130 20148 15130 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 15456 11322 15456 11322 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20470 14688 20470 14688 0 sb_0__1_.mux_right_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 43746 13464 43746 13464 0 sb_0__1_.mux_right_track_38.out
rlabel metal1 30130 14246 30130 14246 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 36938 14076 36938 14076 0 sb_0__1_.mux_right_track_38.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 46276 26962 46276 26962 0 sb_0__1_.mux_right_track_4.out
rlabel metal1 40158 42534 40158 42534 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39514 37162 39514 37162 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 39514 35904 39514 35904 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 35466 33014 35466 33014 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 42550 34510 42550 34510 0 sb_0__1_.mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 44482 12240 44482 12240 0 sb_0__1_.mux_right_track_40.out
rlabel metal2 29670 15266 29670 15266 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 38318 14076 38318 14076 0 sb_0__1_.mux_right_track_40.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 43792 11730 43792 11730 0 sb_0__1_.mux_right_track_44.out
rlabel metal1 33626 15470 33626 15470 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 39146 14926 39146 14926 0 sb_0__1_.mux_right_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 45494 11698 45494 11698 0 sb_0__1_.mux_right_track_46.out
rlabel metal1 34040 17306 34040 17306 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 40250 15708 40250 15708 0 sb_0__1_.mux_right_track_46.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44390 12444 44390 12444 0 sb_0__1_.mux_right_track_48.out
rlabel metal1 37904 16558 37904 16558 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37490 16456 37490 16456 0 sb_0__1_.mux_right_track_48.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 44206 13294 44206 13294 0 sb_0__1_.mux_right_track_50.out
rlabel metal1 37858 18394 37858 18394 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37628 18258 37628 18258 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 39652 18054 39652 18054 0 sb_0__1_.mux_right_track_50.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 44206 10540 44206 10540 0 sb_0__1_.mux_right_track_52.out
rlabel metal1 33626 16456 33626 16456 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 41492 11730 41492 11730 0 sb_0__1_.mux_right_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 42734 9486 42734 9486 0 sb_0__1_.mux_right_track_54.out
rlabel metal2 34362 13634 34362 13634 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40388 10642 40388 10642 0 sb_0__1_.mux_right_track_54.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 43378 10506 43378 10506 0 sb_0__1_.mux_right_track_56.out
rlabel metal1 37398 15062 37398 15062 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 41262 13498 41262 13498 0 sb_0__1_.mux_right_track_56.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 46276 27030 46276 27030 0 sb_0__1_.mux_right_track_6.out
rlabel metal1 40572 43078 40572 43078 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 40618 38522 40618 38522 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 37743 34170 37743 34170 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 42780 36890 42780 36890 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 40710 36346 40710 36346 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 43378 36550 43378 36550 0 sb_0__1_.mux_right_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 45034 32742 45034 32742 0 sb_0__1_.mux_right_track_8.out
rlabel metal1 39008 40562 39008 40562 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 39238 39066 39238 39066 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 35190 35530 35190 35530 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 40802 37910 40802 37910 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 41262 38352 41262 38352 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 43838 35292 43838 35292 0 sb_0__1_.mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 24242 47770 24242 47770 0 sb_0__1_.mux_top_track_0.out
rlabel metal1 24173 41446 24173 41446 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 34040 41514 34040 41514 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 31050 34476 31050 34476 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 24380 36346 24380 36346 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26680 41786 26680 41786 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 25944 41412 25944 41412 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 25392 43418 25392 43418 0 sb_0__1_.mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21252 50218 21252 50218 0 sb_0__1_.mux_top_track_10.out
rlabel metal2 25990 38352 25990 38352 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35374 35802 35374 35802 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 24978 33490 24978 33490 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21482 32198 21482 32198 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 25530 37808 25530 37808 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 23690 35904 23690 35904 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 22908 43758 22908 43758 0 sb_0__1_.mux_top_track_10.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal1 21252 49130 21252 49130 0 sb_0__1_.mux_top_track_12.out
rlabel via2 28934 32827 28934 32827 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 35834 30906 35834 30906 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22862 30260 22862 30260 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 28152 33082 28152 33082 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24242 33898 24242 33898 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 22402 41797 22402 41797 0 sb_0__1_.mux_top_track_12.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 26726 48756 26726 48756 0 sb_0__1_.mux_top_track_2.out
rlabel metal2 33626 39168 33626 39168 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38134 34918 38134 34918 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 29302 34952 29302 34952 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 32614 40358 32614 40358 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 30912 37094 30912 37094 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 27324 45934 27324 45934 0 sb_0__1_.mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19320 49198 19320 49198 0 sb_0__1_.mux_top_track_20.out
rlabel metal2 30222 33932 30222 33932 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 32798 32776 32798 32776 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 23138 28730 23138 28730 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 23782 33422 23782 33422 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 23552 33830 23552 33830 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 20838 38182 20838 38182 0 sb_0__1_.mux_top_track_20.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal2 16882 46614 16882 46614 0 sb_0__1_.mux_top_track_28.out
rlabel metal1 25668 35054 25668 35054 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal2 28474 33456 28474 33456 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20884 36754 20884 36754 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 18538 36754 18538 36754 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 19458 40052 19458 40052 0 sb_0__1_.mux_top_track_28.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal2 15962 48722 15962 48722 0 sb_0__1_.mux_top_track_36.out
rlabel metal1 28750 38386 28750 38386 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 27554 38454 27554 38454 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal2 22126 38896 22126 38896 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 20102 45866 20102 45866 0 sb_0__1_.mux_top_track_36.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 24610 45050 24610 45050 0 sb_0__1_.mux_top_track_4.out
rlabel metal1 32614 36890 32614 36890 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 38962 33286 38962 33286 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 25576 34918 25576 34918 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 29854 37944 29854 37944 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 26450 38794 26450 38794 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 26220 44846 26220 44846 0 sb_0__1_.mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 19550 45832 19550 45832 0 sb_0__1_.mux_top_track_44.out
rlabel metal1 33442 37128 33442 37128 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 23368 37094 23368 37094 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 20884 45934 20884 45934 0 sb_0__1_.mux_top_track_44.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 20930 46648 20930 46648 0 sb_0__1_.mux_top_track_52.out
rlabel metal1 42044 37638 42044 37638 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37398 34952 37398 34952 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 28888 33626 28888 33626 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal2 21758 39678 21758 39678 0 sb_0__1_.mux_top_track_52.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal1 22862 45050 22862 45050 0 sb_0__1_.mux_top_track_6.out
rlabel metal1 27278 38182 27278 38182 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_0_X
rlabel metal1 37398 36346 37398 36346 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_1_X
rlabel metal1 29440 30022 29440 30022 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_2_X
rlabel metal1 25392 34578 25392 34578 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_3_X
rlabel metal2 27094 38760 27094 38760 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_4_X
rlabel metal1 25162 34714 25162 34714 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_5_X
rlabel metal1 23828 44846 23828 44846 0 sb_0__1_.mux_top_track_6.sky130_fd_sc_hd__mux2_1_6_X
rlabel metal2 48622 2438 48622 2438 0 test_enable_bottom_in
rlabel metal2 49358 2098 49358 2098 0 test_enable_bottom_out
rlabel metal2 49358 52513 49358 52513 0 test_enable_right_in
rlabel metal1 48668 55726 48668 55726 0 test_enable_top_in
rlabel metal1 49450 53142 49450 53142 0 test_enable_top_out
rlabel metal3 820 45764 820 45764 0 top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_
rlabel metal3 820 48076 820 48076 0 top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_
rlabel metal3 820 50388 820 50388 0 top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_
rlabel metal3 820 52700 820 52700 0 top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_
<< properties >>
string FIXED_BBOX 0 0 51000 57000
<< end >>
