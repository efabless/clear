magic
tech sky130A
magscale 1 2
timestamp 1656574955
<< viali >>
rect 2053 20553 2087 20587
rect 17049 20553 17083 20587
rect 18889 20553 18923 20587
rect 20177 20553 20211 20587
rect 15577 20485 15611 20519
rect 1685 20417 1719 20451
rect 2237 20417 2271 20451
rect 2697 20417 2731 20451
rect 2973 20417 3007 20451
rect 4169 20417 4203 20451
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 16865 20417 16899 20451
rect 17785 20417 17819 20451
rect 18705 20417 18739 20451
rect 19533 20417 19567 20451
rect 19993 20417 20027 20451
rect 20545 20417 20579 20451
rect 21097 20417 21131 20451
rect 3801 20349 3835 20383
rect 4537 20349 4571 20383
rect 7849 20349 7883 20383
rect 17877 20349 17911 20383
rect 17969 20349 18003 20383
rect 2513 20281 2547 20315
rect 6009 20281 6043 20315
rect 15945 20281 15979 20315
rect 1501 20213 1535 20247
rect 3157 20213 3191 20247
rect 12449 20213 12483 20247
rect 16221 20213 16255 20247
rect 17417 20213 17451 20247
rect 19717 20213 19751 20247
rect 20729 20213 20763 20247
rect 21281 20213 21315 20247
rect 2053 20009 2087 20043
rect 12725 20009 12759 20043
rect 15301 20009 15335 20043
rect 20177 20009 20211 20043
rect 9965 19941 9999 19975
rect 13737 19941 13771 19975
rect 20729 19941 20763 19975
rect 7665 19873 7699 19907
rect 10517 19873 10551 19907
rect 11805 19873 11839 19907
rect 11897 19873 11931 19907
rect 14749 19873 14783 19907
rect 16681 19873 16715 19907
rect 17325 19873 17359 19907
rect 18705 19873 18739 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2689 19805 2723 19839
rect 3249 19805 3283 19839
rect 7849 19805 7883 19839
rect 12541 19805 12575 19839
rect 13001 19805 13035 19839
rect 13553 19805 13587 19839
rect 15117 19805 15151 19839
rect 19257 19805 19291 19839
rect 19993 19805 20027 19839
rect 20545 19805 20579 19839
rect 21097 19805 21131 19839
rect 4537 19737 4571 19771
rect 10333 19737 10367 19771
rect 14473 19737 14507 19771
rect 1501 19669 1535 19703
rect 2513 19669 2547 19703
rect 3065 19669 3099 19703
rect 3893 19669 3927 19703
rect 4261 19669 4295 19703
rect 4905 19669 4939 19703
rect 7757 19669 7791 19703
rect 8217 19669 8251 19703
rect 10425 19669 10459 19703
rect 11069 19669 11103 19703
rect 11345 19669 11379 19703
rect 11713 19669 11747 19703
rect 13185 19669 13219 19703
rect 14105 19669 14139 19703
rect 14565 19669 14599 19703
rect 15853 19669 15887 19703
rect 16129 19669 16163 19703
rect 16497 19669 16531 19703
rect 16589 19669 16623 19703
rect 17509 19669 17543 19703
rect 17601 19669 17635 19703
rect 17969 19669 18003 19703
rect 18245 19669 18279 19703
rect 19441 19669 19475 19703
rect 21281 19669 21315 19703
rect 2973 19465 3007 19499
rect 4169 19465 4203 19499
rect 4721 19465 4755 19499
rect 5181 19465 5215 19499
rect 7573 19465 7607 19499
rect 7941 19465 7975 19499
rect 10425 19465 10459 19499
rect 11805 19465 11839 19499
rect 14381 19465 14415 19499
rect 14841 19465 14875 19499
rect 17417 19465 17451 19499
rect 17785 19465 17819 19499
rect 18889 19465 18923 19499
rect 19349 19465 19383 19499
rect 19809 19465 19843 19499
rect 20729 19465 20763 19499
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 2697 19329 2731 19363
rect 3157 19329 3191 19363
rect 5089 19329 5123 19363
rect 9413 19329 9447 19363
rect 10057 19329 10091 19363
rect 14473 19329 14507 19363
rect 18705 19329 18739 19363
rect 19165 19329 19199 19363
rect 19625 19329 19659 19363
rect 20085 19329 20119 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 3893 19261 3927 19295
rect 5273 19261 5307 19295
rect 8033 19261 8067 19295
rect 8217 19261 8251 19295
rect 9873 19261 9907 19295
rect 9965 19261 9999 19295
rect 10701 19261 10735 19295
rect 12357 19261 12391 19295
rect 14289 19261 14323 19295
rect 16773 19261 16807 19295
rect 17877 19261 17911 19295
rect 18061 19261 18095 19295
rect 2053 19193 2087 19227
rect 2513 19193 2547 19227
rect 1501 19125 1535 19159
rect 3525 19125 3559 19159
rect 5733 19125 5767 19159
rect 6469 19125 6503 19159
rect 12817 19125 12851 19159
rect 15485 19125 15519 19159
rect 17049 19125 17083 19159
rect 20269 19125 20303 19159
rect 21281 19125 21315 19159
rect 2421 18921 2455 18955
rect 3341 18921 3375 18955
rect 5273 18921 5307 18955
rect 11069 18921 11103 18955
rect 14565 18921 14599 18955
rect 16589 18921 16623 18955
rect 17693 18921 17727 18955
rect 18797 18921 18831 18955
rect 19993 18853 20027 18887
rect 4353 18785 4387 18819
rect 5917 18785 5951 18819
rect 6837 18785 6871 18819
rect 11897 18785 11931 18819
rect 11989 18785 12023 18819
rect 12633 18785 12667 18819
rect 15117 18785 15151 18819
rect 16129 18785 16163 18819
rect 17233 18785 17267 18819
rect 18429 18785 18463 18819
rect 19349 18785 19383 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 3065 18717 3099 18751
rect 5733 18717 5767 18751
rect 8953 18717 8987 18751
rect 11805 18717 11839 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 5641 18649 5675 18683
rect 6285 18649 6319 18683
rect 14933 18649 14967 18683
rect 17049 18649 17083 18683
rect 19533 18649 19567 18683
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 2881 18581 2915 18615
rect 3801 18581 3835 18615
rect 4169 18581 4203 18615
rect 4261 18581 4295 18615
rect 4813 18581 4847 18615
rect 7205 18581 7239 18615
rect 9505 18581 9539 18615
rect 11437 18581 11471 18615
rect 12725 18581 12759 18615
rect 12817 18581 12851 18615
rect 13185 18581 13219 18615
rect 15025 18581 15059 18615
rect 15577 18581 15611 18615
rect 15945 18581 15979 18615
rect 16037 18581 16071 18615
rect 16957 18581 16991 18615
rect 17969 18581 18003 18615
rect 19625 18581 19659 18615
rect 20269 18581 20303 18615
rect 20821 18581 20855 18615
rect 21281 18581 21315 18615
rect 1961 18377 1995 18411
rect 3617 18377 3651 18411
rect 4261 18377 4295 18411
rect 5273 18377 5307 18411
rect 7573 18377 7607 18411
rect 7941 18377 7975 18411
rect 9321 18377 9355 18411
rect 10149 18377 10183 18411
rect 12357 18377 12391 18411
rect 14105 18377 14139 18411
rect 15209 18377 15243 18411
rect 15301 18377 15335 18411
rect 15669 18377 15703 18411
rect 19165 18377 19199 18411
rect 5641 18309 5675 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2605 18241 2639 18275
rect 3249 18241 3283 18275
rect 5733 18241 5767 18275
rect 8309 18241 8343 18275
rect 8401 18241 8435 18275
rect 9965 18241 9999 18275
rect 11161 18241 11195 18275
rect 11989 18241 12023 18275
rect 12633 18241 12667 18275
rect 13645 18241 13679 18275
rect 18153 18241 18187 18275
rect 20085 18241 20119 18275
rect 20545 18241 20579 18275
rect 21097 18241 21131 18275
rect 2973 18173 3007 18207
rect 3157 18173 3191 18207
rect 3985 18173 4019 18207
rect 4169 18173 4203 18207
rect 5825 18173 5859 18207
rect 7021 18173 7055 18207
rect 8493 18173 8527 18207
rect 9413 18173 9447 18207
rect 9505 18173 9539 18207
rect 11805 18173 11839 18207
rect 11897 18173 11931 18207
rect 15117 18173 15151 18207
rect 17417 18173 17451 18207
rect 17969 18173 18003 18207
rect 18061 18173 18095 18207
rect 19257 18173 19291 18207
rect 19349 18173 19383 18207
rect 4997 18105 5031 18139
rect 13829 18105 13863 18139
rect 20269 18105 20303 18139
rect 1501 18037 1535 18071
rect 2421 18037 2455 18071
rect 4629 18037 4663 18071
rect 6469 18037 6503 18071
rect 8953 18037 8987 18071
rect 13185 18037 13219 18071
rect 16221 18037 16255 18071
rect 16773 18037 16807 18071
rect 17141 18037 17175 18071
rect 18521 18037 18555 18071
rect 18797 18037 18831 18071
rect 20729 18037 20763 18071
rect 21281 18037 21315 18071
rect 2513 17833 2547 17867
rect 3433 17833 3467 17867
rect 5641 17833 5675 17867
rect 9597 17833 9631 17867
rect 16129 17833 16163 17867
rect 19257 17833 19291 17867
rect 21281 17833 21315 17867
rect 7481 17765 7515 17799
rect 17601 17765 17635 17799
rect 3801 17697 3835 17731
rect 4721 17697 4755 17731
rect 6285 17697 6319 17731
rect 6929 17697 6963 17731
rect 7941 17697 7975 17731
rect 10241 17697 10275 17731
rect 12173 17697 12207 17731
rect 15577 17697 15611 17731
rect 18153 17697 18187 17731
rect 19901 17697 19935 17731
rect 20821 17697 20855 17731
rect 1685 17629 1719 17663
rect 2237 17629 2271 17663
rect 2697 17629 2731 17663
rect 2973 17629 3007 17663
rect 11989 17629 12023 17663
rect 16405 17629 16439 17663
rect 16865 17629 16899 17663
rect 17969 17629 18003 17663
rect 20729 17629 20763 17663
rect 4905 17561 4939 17595
rect 8125 17561 8159 17595
rect 8953 17561 8987 17595
rect 11897 17561 11931 17595
rect 12541 17561 12575 17595
rect 17325 17561 17359 17595
rect 19625 17561 19659 17595
rect 1501 17493 1535 17527
rect 2053 17493 2087 17527
rect 4261 17493 4295 17527
rect 4997 17493 5031 17527
rect 5365 17493 5399 17527
rect 6009 17493 6043 17527
rect 6101 17493 6135 17527
rect 7021 17493 7055 17527
rect 7113 17493 7147 17527
rect 8033 17493 8067 17527
rect 8493 17493 8527 17527
rect 9965 17493 9999 17527
rect 10057 17493 10091 17527
rect 10701 17493 10735 17527
rect 11161 17493 11195 17527
rect 11529 17493 11563 17527
rect 13093 17493 13127 17527
rect 15117 17493 15151 17527
rect 15669 17493 15703 17527
rect 15761 17493 15795 17527
rect 16589 17493 16623 17527
rect 18061 17493 18095 17527
rect 18613 17493 18647 17527
rect 19717 17493 19751 17527
rect 20269 17493 20303 17527
rect 20637 17493 20671 17527
rect 2881 17289 2915 17323
rect 3985 17289 4019 17323
rect 4445 17289 4479 17323
rect 5181 17289 5215 17323
rect 6929 17289 6963 17323
rect 8309 17289 8343 17323
rect 8401 17289 8435 17323
rect 9045 17289 9079 17323
rect 9505 17289 9539 17323
rect 10701 17289 10735 17323
rect 14749 17289 14783 17323
rect 19073 17289 19107 17323
rect 20821 17289 20855 17323
rect 4077 17221 4111 17255
rect 5089 17221 5123 17255
rect 13645 17221 13679 17255
rect 14289 17221 14323 17255
rect 20729 17221 20763 17255
rect 1685 17153 1719 17187
rect 1961 17153 1995 17187
rect 2605 17153 2639 17187
rect 3065 17153 3099 17187
rect 3433 17153 3467 17187
rect 9413 17153 9447 17187
rect 10149 17153 10183 17187
rect 10793 17153 10827 17187
rect 11989 17153 12023 17187
rect 12633 17153 12667 17187
rect 14381 17153 14415 17187
rect 15025 17153 15059 17187
rect 16681 17153 16715 17187
rect 17141 17153 17175 17187
rect 18889 17153 18923 17187
rect 19349 17153 19383 17187
rect 19809 17153 19843 17187
rect 3801 17085 3835 17119
rect 5365 17085 5399 17119
rect 6745 17085 6779 17119
rect 6837 17085 6871 17119
rect 8217 17085 8251 17119
rect 9597 17085 9631 17119
rect 10517 17085 10551 17119
rect 11805 17085 11839 17119
rect 11897 17085 11931 17119
rect 14197 17085 14231 17119
rect 21005 17085 21039 17119
rect 2145 17017 2179 17051
rect 4721 17017 4755 17051
rect 16865 17017 16899 17051
rect 19533 17017 19567 17051
rect 1501 16949 1535 16983
rect 2421 16949 2455 16983
rect 5825 16949 5859 16983
rect 7297 16949 7331 16983
rect 7665 16949 7699 16983
rect 8769 16949 8803 16983
rect 11161 16949 11195 16983
rect 12357 16949 12391 16983
rect 17509 16949 17543 16983
rect 18613 16949 18647 16983
rect 19993 16949 20027 16983
rect 20361 16949 20395 16983
rect 16221 16745 16255 16779
rect 19533 16745 19567 16779
rect 6009 16677 6043 16711
rect 9505 16677 9539 16711
rect 3985 16609 4019 16643
rect 4077 16609 4111 16643
rect 5641 16609 5675 16643
rect 6377 16609 6411 16643
rect 9137 16609 9171 16643
rect 10057 16609 10091 16643
rect 11069 16609 11103 16643
rect 12817 16609 12851 16643
rect 12909 16609 12943 16643
rect 15853 16609 15887 16643
rect 16865 16609 16899 16643
rect 17785 16609 17819 16643
rect 18889 16609 18923 16643
rect 20453 16609 20487 16643
rect 20545 16609 20579 16643
rect 1685 16541 1719 16575
rect 2145 16541 2179 16575
rect 2881 16541 2915 16575
rect 3341 16541 3375 16575
rect 8493 16541 8527 16575
rect 10241 16541 10275 16575
rect 13001 16541 13035 16575
rect 16681 16541 16715 16575
rect 17693 16541 17727 16575
rect 18337 16541 18371 16575
rect 19717 16541 19751 16575
rect 21097 16541 21131 16575
rect 4169 16473 4203 16507
rect 7389 16473 7423 16507
rect 17601 16473 17635 16507
rect 1501 16405 1535 16439
rect 1961 16405 1995 16439
rect 2697 16405 2731 16439
rect 3157 16405 3191 16439
rect 4537 16405 4571 16439
rect 4905 16405 4939 16439
rect 5273 16405 5307 16439
rect 6745 16405 6779 16439
rect 7849 16405 7883 16439
rect 8125 16405 8159 16439
rect 10149 16405 10183 16439
rect 10609 16405 10643 16439
rect 11161 16405 11195 16439
rect 11253 16405 11287 16439
rect 11621 16405 11655 16439
rect 11989 16405 12023 16439
rect 13369 16405 13403 16439
rect 16589 16405 16623 16439
rect 17233 16405 17267 16439
rect 18521 16405 18555 16439
rect 19993 16405 20027 16439
rect 20361 16405 20395 16439
rect 21281 16405 21315 16439
rect 2513 16201 2547 16235
rect 3341 16201 3375 16235
rect 5089 16201 5123 16235
rect 6561 16201 6595 16235
rect 7573 16201 7607 16235
rect 7941 16201 7975 16235
rect 14565 16201 14599 16235
rect 16681 16201 16715 16235
rect 17693 16201 17727 16235
rect 18337 16201 18371 16235
rect 18797 16201 18831 16235
rect 20177 16201 20211 16235
rect 3065 16133 3099 16167
rect 6929 16133 6963 16167
rect 14105 16133 14139 16167
rect 1685 16065 1719 16099
rect 2237 16065 2271 16099
rect 2697 16065 2731 16099
rect 4445 16065 4479 16099
rect 5457 16065 5491 16099
rect 10261 16065 10295 16099
rect 14197 16065 14231 16099
rect 17601 16065 17635 16099
rect 18705 16065 18739 16099
rect 19349 16065 19383 16099
rect 19993 16065 20027 16099
rect 20545 16065 20579 16099
rect 21097 16065 21131 16099
rect 4537 15997 4571 16031
rect 4721 15997 4755 16031
rect 5549 15997 5583 16031
rect 5641 15997 5675 16031
rect 7021 15997 7055 16031
rect 7205 15997 7239 16031
rect 8033 15997 8067 16031
rect 8125 15997 8159 16031
rect 10517 15997 10551 16031
rect 14013 15997 14047 16031
rect 17509 15997 17543 16031
rect 18889 15997 18923 16031
rect 2053 15929 2087 15963
rect 3709 15929 3743 15963
rect 11621 15929 11655 15963
rect 18061 15929 18095 15963
rect 20729 15929 20763 15963
rect 1501 15861 1535 15895
rect 4077 15861 4111 15895
rect 8585 15861 8619 15895
rect 9137 15861 9171 15895
rect 10793 15861 10827 15895
rect 13461 15861 13495 15895
rect 14933 15861 14967 15895
rect 21281 15861 21315 15895
rect 4445 15657 4479 15691
rect 8217 15657 8251 15691
rect 10609 15657 10643 15691
rect 12357 15657 12391 15691
rect 13645 15657 13679 15691
rect 16957 15657 16991 15691
rect 18521 15657 18555 15691
rect 19809 15657 19843 15691
rect 6929 15589 6963 15623
rect 11989 15589 12023 15623
rect 4905 15521 4939 15555
rect 5089 15521 5123 15555
rect 6377 15521 6411 15555
rect 6469 15521 6503 15555
rect 7665 15521 7699 15555
rect 11713 15521 11747 15555
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 2605 15453 2639 15487
rect 7757 15453 7791 15487
rect 8493 15453 8527 15487
rect 9229 15453 9263 15487
rect 10885 15453 10919 15487
rect 16589 15453 16623 15487
rect 17233 15453 17267 15487
rect 17693 15453 17727 15487
rect 18797 15453 18831 15487
rect 19625 15453 19659 15487
rect 20085 15453 20119 15487
rect 20545 15453 20579 15487
rect 21097 15453 21131 15487
rect 4813 15385 4847 15419
rect 5457 15385 5491 15419
rect 9496 15385 9530 15419
rect 16322 15385 16356 15419
rect 18153 15385 18187 15419
rect 1501 15317 1535 15351
rect 1961 15317 1995 15351
rect 2421 15317 2455 15351
rect 2881 15317 2915 15351
rect 3341 15317 3375 15351
rect 3985 15317 4019 15351
rect 6561 15317 6595 15351
rect 7849 15317 7883 15351
rect 11345 15317 11379 15351
rect 15209 15317 15243 15351
rect 19349 15317 19383 15351
rect 20269 15317 20303 15351
rect 20729 15317 20763 15351
rect 21281 15317 21315 15351
rect 2513 15113 2547 15147
rect 4353 15113 4387 15147
rect 6653 15113 6687 15147
rect 7021 15113 7055 15147
rect 7665 15113 7699 15147
rect 11529 15113 11563 15147
rect 16681 15113 16715 15147
rect 7757 15045 7791 15079
rect 8309 15045 8343 15079
rect 8769 15045 8803 15079
rect 18337 15045 18371 15079
rect 18889 15045 18923 15079
rect 1685 14977 1719 15011
rect 1961 14977 1995 15011
rect 2697 14977 2731 15011
rect 3157 14977 3191 15011
rect 4997 14977 5031 15011
rect 5089 14977 5123 15011
rect 9689 14977 9723 15011
rect 9956 14977 9990 15011
rect 12265 14977 12299 15011
rect 13461 14977 13495 15011
rect 13728 14977 13762 15011
rect 17794 14977 17828 15011
rect 18061 14977 18095 15011
rect 19441 14977 19475 15011
rect 19901 14977 19935 15011
rect 20157 14977 20191 15011
rect 5273 14909 5307 14943
rect 7941 14909 7975 14943
rect 9045 14909 9079 14943
rect 2973 14841 3007 14875
rect 3801 14841 3835 14875
rect 14841 14841 14875 14875
rect 1501 14773 1535 14807
rect 2145 14773 2179 14807
rect 3525 14773 3559 14807
rect 4629 14773 4663 14807
rect 6009 14773 6043 14807
rect 7297 14773 7331 14807
rect 11069 14773 11103 14807
rect 11989 14773 12023 14807
rect 12725 14773 12759 14807
rect 13001 14773 13035 14807
rect 15117 14773 15151 14807
rect 15577 14773 15611 14807
rect 16037 14773 16071 14807
rect 19625 14773 19659 14807
rect 21281 14773 21315 14807
rect 5089 14569 5123 14603
rect 6653 14569 6687 14603
rect 7941 14569 7975 14603
rect 14105 14569 14139 14603
rect 17141 14569 17175 14603
rect 19257 14569 19291 14603
rect 3801 14501 3835 14535
rect 11621 14501 11655 14535
rect 4353 14433 4387 14467
rect 5733 14433 5767 14467
rect 7021 14433 7055 14467
rect 7205 14433 7239 14467
rect 10241 14433 10275 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 2789 14365 2823 14399
rect 4261 14365 4295 14399
rect 5457 14365 5491 14399
rect 7297 14365 7331 14399
rect 10508 14365 10542 14399
rect 13277 14365 13311 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 18797 14365 18831 14399
rect 20637 14365 20671 14399
rect 21097 14365 21131 14399
rect 4169 14297 4203 14331
rect 8953 14297 8987 14331
rect 9413 14297 9447 14331
rect 13010 14297 13044 14331
rect 15218 14297 15252 14331
rect 16006 14297 16040 14331
rect 18530 14297 18564 14331
rect 20392 14297 20426 14331
rect 1501 14229 1535 14263
rect 2145 14229 2179 14263
rect 2605 14229 2639 14263
rect 3065 14229 3099 14263
rect 5549 14229 5583 14263
rect 6193 14229 6227 14263
rect 7665 14229 7699 14263
rect 8309 14229 8343 14263
rect 9689 14229 9723 14263
rect 11897 14229 11931 14263
rect 13645 14229 13679 14263
rect 17417 14229 17451 14263
rect 21281 14229 21315 14263
rect 2881 14025 2915 14059
rect 3157 14025 3191 14059
rect 3985 14025 4019 14059
rect 4445 14025 4479 14059
rect 5089 14025 5123 14059
rect 6837 14025 6871 14059
rect 8033 14025 8067 14059
rect 8493 14025 8527 14059
rect 10885 14025 10919 14059
rect 11713 14025 11747 14059
rect 15945 14025 15979 14059
rect 18981 14025 19015 14059
rect 19625 14025 19659 14059
rect 2145 13957 2179 13991
rect 4353 13957 4387 13991
rect 8861 13957 8895 13991
rect 9496 13957 9530 13991
rect 17868 13957 17902 13991
rect 2053 13889 2087 13923
rect 2697 13889 2731 13923
rect 3341 13889 3375 13923
rect 5549 13889 5583 13923
rect 9229 13889 9263 13923
rect 12173 13889 12207 13923
rect 13165 13889 13199 13923
rect 14565 13889 14599 13923
rect 14821 13889 14855 13923
rect 19441 13889 19475 13923
rect 21014 13889 21048 13923
rect 21281 13889 21315 13923
rect 2237 13821 2271 13855
rect 4629 13821 4663 13855
rect 5825 13821 5859 13855
rect 6929 13821 6963 13855
rect 7113 13821 7147 13855
rect 12909 13821 12943 13855
rect 16957 13821 16991 13855
rect 17325 13821 17359 13855
rect 17601 13821 17635 13855
rect 7757 13753 7791 13787
rect 10609 13753 10643 13787
rect 14289 13753 14323 13787
rect 19901 13753 19935 13787
rect 1685 13685 1719 13719
rect 3617 13685 3651 13719
rect 6469 13685 6503 13719
rect 12449 13685 12483 13719
rect 16221 13685 16255 13719
rect 2421 13481 2455 13515
rect 3433 13481 3467 13515
rect 6469 13481 6503 13515
rect 9045 13481 9079 13515
rect 10793 13481 10827 13515
rect 11069 13481 11103 13515
rect 12541 13481 12575 13515
rect 17417 13481 17451 13515
rect 18061 13481 18095 13515
rect 21281 13481 21315 13515
rect 3801 13413 3835 13447
rect 6193 13413 6227 13447
rect 8493 13413 8527 13447
rect 1869 13345 1903 13379
rect 4445 13345 4479 13379
rect 5641 13345 5675 13379
rect 7113 13345 7147 13379
rect 8125 13345 8159 13379
rect 9413 13345 9447 13379
rect 13369 13345 13403 13379
rect 15761 13345 15795 13379
rect 2053 13277 2087 13311
rect 2697 13277 2731 13311
rect 3249 13277 3283 13311
rect 5825 13277 5859 13311
rect 6929 13277 6963 13311
rect 7941 13277 7975 13311
rect 16037 13277 16071 13311
rect 17785 13277 17819 13311
rect 18889 13277 18923 13311
rect 20729 13277 20763 13311
rect 21097 13277 21131 13311
rect 5181 13209 5215 13243
rect 5733 13209 5767 13243
rect 9669 13209 9703 13243
rect 11529 13209 11563 13243
rect 12173 13209 12207 13243
rect 16304 13209 16338 13243
rect 18429 13209 18463 13243
rect 20484 13209 20518 13243
rect 1961 13141 1995 13175
rect 2881 13141 2915 13175
rect 4169 13141 4203 13175
rect 4261 13141 4295 13175
rect 6837 13141 6871 13175
rect 7481 13141 7515 13175
rect 7849 13141 7883 13175
rect 11805 13141 11839 13175
rect 13001 13141 13035 13175
rect 13737 13141 13771 13175
rect 14381 13141 14415 13175
rect 14933 13141 14967 13175
rect 15301 13141 15335 13175
rect 19349 13141 19383 13175
rect 2697 12937 2731 12971
rect 5273 12937 5307 12971
rect 5733 12937 5767 12971
rect 7021 12937 7055 12971
rect 7665 12937 7699 12971
rect 8677 12937 8711 12971
rect 9229 12937 9263 12971
rect 10885 12937 10919 12971
rect 11529 12937 11563 12971
rect 16221 12937 16255 12971
rect 17233 12937 17267 12971
rect 20177 12937 20211 12971
rect 10342 12869 10376 12903
rect 11897 12869 11931 12903
rect 15218 12869 15252 12903
rect 1961 12801 1995 12835
rect 2513 12801 2547 12835
rect 3709 12801 3743 12835
rect 5641 12801 5675 12835
rect 10609 12801 10643 12835
rect 13481 12801 13515 12835
rect 18133 12801 18167 12835
rect 19717 12801 19751 12835
rect 19993 12801 20027 12835
rect 20821 12801 20855 12835
rect 2237 12733 2271 12767
rect 2973 12733 3007 12767
rect 3525 12733 3559 12767
rect 3617 12733 3651 12767
rect 4353 12733 4387 12767
rect 5917 12733 5951 12767
rect 7757 12733 7791 12767
rect 7849 12733 7883 12767
rect 13737 12733 13771 12767
rect 15485 12733 15519 12767
rect 16865 12733 16899 12767
rect 17877 12733 17911 12767
rect 20545 12733 20579 12767
rect 7297 12665 7331 12699
rect 12357 12665 12391 12699
rect 19533 12665 19567 12699
rect 4077 12597 4111 12631
rect 4813 12597 4847 12631
rect 6377 12597 6411 12631
rect 8309 12597 8343 12631
rect 14105 12597 14139 12631
rect 15761 12597 15795 12631
rect 17601 12597 17635 12631
rect 19257 12597 19291 12631
rect 3893 12393 3927 12427
rect 6101 12393 6135 12427
rect 6929 12393 6963 12427
rect 8493 12393 8527 12427
rect 9229 12393 9263 12427
rect 12265 12393 12299 12427
rect 14933 12393 14967 12427
rect 19717 12393 19751 12427
rect 20545 12393 20579 12427
rect 5273 12325 5307 12359
rect 12909 12325 12943 12359
rect 1961 12257 1995 12291
rect 3065 12257 3099 12291
rect 4445 12257 4479 12291
rect 7389 12257 7423 12291
rect 7573 12257 7607 12291
rect 17693 12257 17727 12291
rect 19993 12257 20027 12291
rect 21097 12257 21131 12291
rect 2237 12189 2271 12223
rect 2973 12189 3007 12223
rect 6469 12189 6503 12223
rect 8125 12189 8159 12223
rect 10609 12189 10643 12223
rect 10885 12189 10919 12223
rect 13369 12189 13403 12223
rect 15669 12189 15703 12223
rect 19533 12189 19567 12223
rect 5641 12121 5675 12155
rect 10342 12121 10376 12155
rect 11130 12121 11164 12155
rect 12633 12121 12667 12155
rect 14105 12121 14139 12155
rect 15936 12121 15970 12155
rect 18061 12121 18095 12155
rect 18429 12121 18463 12155
rect 18797 12121 18831 12155
rect 20177 12121 20211 12155
rect 20913 12121 20947 12155
rect 2513 12053 2547 12087
rect 2881 12053 2915 12087
rect 4261 12053 4295 12087
rect 4353 12053 4387 12087
rect 4997 12053 5031 12087
rect 7297 12053 7331 12087
rect 13645 12053 13679 12087
rect 14473 12053 14507 12087
rect 15393 12053 15427 12087
rect 17049 12053 17083 12087
rect 17325 12053 17359 12087
rect 21005 12053 21039 12087
rect 3525 11849 3559 11883
rect 4261 11849 4295 11883
rect 5273 11849 5307 11883
rect 7297 11849 7331 11883
rect 9505 11849 9539 11883
rect 13185 11849 13219 11883
rect 13553 11849 13587 11883
rect 15761 11849 15795 11883
rect 16957 11849 16991 11883
rect 19717 11849 19751 11883
rect 20085 11849 20119 11883
rect 20821 11849 20855 11883
rect 21281 11849 21315 11883
rect 3157 11781 3191 11815
rect 4169 11781 4203 11815
rect 7205 11781 7239 11815
rect 10618 11781 10652 11815
rect 12050 11781 12084 11815
rect 1961 11713 1995 11747
rect 5641 11713 5675 11747
rect 5733 11713 5767 11747
rect 14105 11713 14139 11747
rect 14372 11713 14406 11747
rect 16313 11713 16347 11747
rect 18236 11713 18270 11747
rect 20177 11713 20211 11747
rect 20913 11713 20947 11747
rect 2237 11645 2271 11679
rect 2973 11645 3007 11679
rect 3065 11645 3099 11679
rect 4445 11645 4479 11679
rect 4905 11645 4939 11679
rect 5825 11645 5859 11679
rect 6653 11645 6687 11679
rect 7113 11645 7147 11679
rect 10885 11645 10919 11679
rect 11805 11645 11839 11679
rect 17969 11645 18003 11679
rect 20729 11645 20763 11679
rect 3801 11577 3835 11611
rect 7665 11577 7699 11611
rect 8769 11577 8803 11611
rect 17233 11577 17267 11611
rect 19349 11577 19383 11611
rect 7941 11509 7975 11543
rect 8309 11509 8343 11543
rect 9137 11509 9171 11543
rect 15485 11509 15519 11543
rect 17601 11509 17635 11543
rect 1685 11305 1719 11339
rect 3985 11305 4019 11339
rect 9229 11305 9263 11339
rect 11713 11305 11747 11339
rect 13093 11305 13127 11339
rect 14105 11305 14139 11339
rect 14841 11305 14875 11339
rect 15301 11305 15335 11339
rect 2973 11237 3007 11271
rect 5365 11237 5399 11271
rect 14565 11237 14599 11271
rect 16957 11237 16991 11271
rect 18705 11237 18739 11271
rect 19441 11237 19475 11271
rect 2237 11169 2271 11203
rect 4813 11169 4847 11203
rect 6101 11169 6135 11203
rect 6193 11169 6227 11203
rect 7297 11169 7331 11203
rect 8493 11169 8527 11203
rect 12541 11169 12575 11203
rect 15577 11169 15611 11203
rect 2053 11101 2087 11135
rect 2789 11101 2823 11135
rect 3801 11101 3835 11135
rect 4997 11101 5031 11135
rect 6009 11101 6043 11135
rect 7021 11101 7055 11135
rect 8217 11101 8251 11135
rect 10342 11101 10376 11135
rect 10609 11101 10643 11135
rect 12081 11101 12115 11135
rect 15833 11101 15867 11135
rect 17325 11101 17359 11135
rect 17581 11101 17615 11135
rect 20821 11101 20855 11135
rect 21281 11101 21315 11135
rect 2145 11033 2179 11067
rect 4353 11033 4387 11067
rect 4905 11033 4939 11067
rect 7113 11033 7147 11067
rect 20576 11033 20610 11067
rect 21097 11033 21131 11067
rect 3249 10965 3283 10999
rect 5641 10965 5675 10999
rect 6653 10965 6687 10999
rect 7849 10965 7883 10999
rect 8309 10965 8343 10999
rect 11069 10965 11103 10999
rect 11345 10965 11379 10999
rect 13369 10965 13403 10999
rect 2513 10761 2547 10795
rect 3893 10761 3927 10795
rect 4537 10761 4571 10795
rect 4997 10761 5031 10795
rect 6837 10761 6871 10795
rect 7481 10761 7515 10795
rect 7941 10761 7975 10795
rect 9229 10761 9263 10795
rect 11529 10761 11563 10795
rect 14933 10761 14967 10795
rect 15485 10761 15519 10795
rect 15853 10761 15887 10795
rect 16221 10761 16255 10795
rect 17141 10761 17175 10795
rect 17509 10761 17543 10795
rect 19257 10761 19291 10795
rect 20913 10761 20947 10795
rect 21189 10761 21223 10795
rect 8769 10693 8803 10727
rect 18122 10693 18156 10727
rect 19800 10693 19834 10727
rect 1961 10625 1995 10659
rect 2237 10625 2271 10659
rect 2881 10625 2915 10659
rect 5457 10625 5491 10659
rect 7849 10625 7883 10659
rect 10353 10625 10387 10659
rect 12642 10625 12676 10659
rect 12909 10625 12943 10659
rect 13277 10625 13311 10659
rect 13533 10625 13567 10659
rect 17877 10625 17911 10659
rect 21373 10625 21407 10659
rect 2973 10557 3007 10591
rect 3065 10557 3099 10591
rect 3985 10557 4019 10591
rect 4077 10557 4111 10591
rect 6653 10557 6687 10591
rect 6745 10557 6779 10591
rect 8125 10557 8159 10591
rect 10609 10557 10643 10591
rect 19533 10557 19567 10591
rect 14657 10489 14691 10523
rect 3525 10421 3559 10455
rect 5273 10421 5307 10455
rect 5825 10421 5859 10455
rect 7205 10421 7239 10455
rect 10977 10421 11011 10455
rect 16865 10421 16899 10455
rect 6561 10217 6595 10251
rect 7297 10217 7331 10251
rect 14657 10217 14691 10251
rect 17693 10217 17727 10251
rect 19533 10217 19567 10251
rect 8309 10149 8343 10183
rect 10793 10149 10827 10183
rect 15669 10149 15703 10183
rect 1961 10081 1995 10115
rect 3157 10081 3191 10115
rect 3801 10081 3835 10115
rect 5089 10081 5123 10115
rect 7941 10081 7975 10115
rect 11621 10081 11655 10115
rect 20085 10081 20119 10115
rect 20545 10081 20579 10115
rect 20821 10081 20855 10115
rect 2237 10013 2271 10047
rect 9413 10013 9447 10047
rect 12173 10013 12207 10047
rect 14197 10013 14231 10047
rect 15393 10013 15427 10047
rect 16037 10013 16071 10047
rect 16293 10013 16327 10047
rect 18429 10013 18463 10047
rect 18705 10013 18739 10047
rect 19901 10013 19935 10047
rect 4905 9945 4939 9979
rect 7665 9945 7699 9979
rect 7757 9945 7791 9979
rect 9658 9945 9692 9979
rect 12418 9945 12452 9979
rect 15025 9945 15059 9979
rect 2513 9877 2547 9911
rect 2881 9877 2915 9911
rect 2973 9877 3007 9911
rect 4445 9877 4479 9911
rect 4813 9877 4847 9911
rect 5549 9877 5583 9911
rect 6193 9877 6227 9911
rect 6929 9877 6963 9911
rect 9045 9877 9079 9911
rect 11253 9877 11287 9911
rect 13553 9877 13587 9911
rect 17417 9877 17451 9911
rect 18245 9877 18279 9911
rect 18889 9877 18923 9911
rect 19993 9877 20027 9911
rect 2421 9673 2455 9707
rect 7297 9673 7331 9707
rect 8125 9673 8159 9707
rect 4353 9605 4387 9639
rect 7389 9605 7423 9639
rect 9260 9605 9294 9639
rect 10026 9605 10060 9639
rect 13062 9605 13096 9639
rect 15678 9605 15712 9639
rect 2053 9537 2087 9571
rect 3249 9537 3283 9571
rect 4445 9537 4479 9571
rect 5549 9537 5583 9571
rect 6377 9537 6411 9571
rect 12817 9537 12851 9571
rect 15945 9537 15979 9571
rect 16221 9537 16255 9571
rect 19082 9537 19116 9571
rect 20177 9537 20211 9571
rect 20821 9537 20855 9571
rect 1869 9469 1903 9503
rect 1961 9469 1995 9503
rect 3065 9469 3099 9503
rect 3157 9469 3191 9503
rect 4261 9469 4295 9503
rect 5273 9469 5307 9503
rect 5457 9469 5491 9503
rect 7573 9469 7607 9503
rect 9505 9469 9539 9503
rect 9781 9469 9815 9503
rect 12541 9469 12575 9503
rect 16957 9469 16991 9503
rect 19349 9469 19383 9503
rect 19717 9469 19751 9503
rect 20545 9469 20579 9503
rect 4813 9401 4847 9435
rect 11161 9401 11195 9435
rect 14197 9401 14231 9435
rect 14565 9401 14599 9435
rect 3617 9333 3651 9367
rect 5917 9333 5951 9367
rect 6929 9333 6963 9367
rect 11529 9333 11563 9367
rect 11989 9333 12023 9367
rect 17325 9333 17359 9367
rect 17969 9333 18003 9367
rect 20085 9333 20119 9367
rect 2605 9129 2639 9163
rect 3985 9129 4019 9163
rect 10793 9129 10827 9163
rect 13737 9129 13771 9163
rect 17417 9129 17451 9163
rect 20453 9129 20487 9163
rect 3341 9061 3375 9095
rect 1961 8993 1995 9027
rect 4353 8993 4387 9027
rect 5457 8993 5491 9027
rect 5549 8993 5583 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 8217 8993 8251 9027
rect 11989 8993 12023 9027
rect 14197 8993 14231 9027
rect 14565 8993 14599 9027
rect 15761 8993 15795 9027
rect 19625 8993 19659 9027
rect 19717 8993 19751 9027
rect 20913 8993 20947 9027
rect 21005 8993 21039 9027
rect 2237 8925 2271 8959
rect 3157 8925 3191 8959
rect 3801 8925 3835 8959
rect 4629 8925 4663 8959
rect 6653 8925 6687 8959
rect 7941 8925 7975 8959
rect 9413 8925 9447 8959
rect 12357 8925 12391 8959
rect 15301 8925 15335 8959
rect 16017 8925 16051 8959
rect 18797 8925 18831 8959
rect 2697 8857 2731 8891
rect 5641 8857 5675 8891
rect 9658 8857 9692 8891
rect 12602 8857 12636 8891
rect 15025 8857 15059 8891
rect 18530 8857 18564 8891
rect 20821 8857 20855 8891
rect 4537 8789 4571 8823
rect 4997 8789 5031 8823
rect 6009 8789 6043 8823
rect 6285 8789 6319 8823
rect 7573 8789 7607 8823
rect 8033 8789 8067 8823
rect 8953 8789 8987 8823
rect 11069 8789 11103 8823
rect 11713 8789 11747 8823
rect 15485 8789 15519 8823
rect 17141 8789 17175 8823
rect 19809 8789 19843 8823
rect 20177 8789 20211 8823
rect 2513 8585 2547 8619
rect 2973 8585 3007 8619
rect 4537 8585 4571 8619
rect 4905 8585 4939 8619
rect 8033 8585 8067 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 12725 8585 12759 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 15853 8585 15887 8619
rect 17417 8585 17451 8619
rect 19809 8585 19843 8619
rect 10793 8517 10827 8551
rect 11989 8517 12023 8551
rect 13093 8517 13127 8551
rect 20922 8517 20956 8551
rect 1961 8449 1995 8483
rect 2881 8449 2915 8483
rect 8769 8449 8803 8483
rect 10057 8449 10091 8483
rect 15218 8449 15252 8483
rect 15485 8449 15519 8483
rect 17233 8449 17267 8483
rect 17693 8449 17727 8483
rect 18409 8449 18443 8483
rect 21189 8449 21223 8483
rect 2237 8381 2271 8415
rect 3065 8381 3099 8415
rect 3525 8381 3559 8415
rect 4997 8381 5031 8415
rect 5181 8381 5215 8415
rect 6009 8381 6043 8415
rect 7941 8381 7975 8415
rect 18153 8381 18187 8415
rect 4169 8313 4203 8347
rect 5641 8313 5675 8347
rect 6469 8313 6503 8347
rect 6837 8313 6871 8347
rect 7481 8313 7515 8347
rect 9137 8313 9171 8347
rect 9689 8313 9723 8347
rect 10517 8313 10551 8347
rect 11529 8313 11563 8347
rect 12265 8313 12299 8347
rect 14105 8313 14139 8347
rect 16129 8313 16163 8347
rect 17877 8313 17911 8347
rect 16957 8245 16991 8279
rect 19533 8245 19567 8279
rect 2237 8041 2271 8075
rect 4997 8041 5031 8075
rect 8953 8041 8987 8075
rect 10609 8041 10643 8075
rect 15025 8041 15059 8075
rect 15853 8041 15887 8075
rect 16589 8041 16623 8075
rect 18705 8041 18739 8075
rect 4721 7973 4755 8007
rect 7665 7973 7699 8007
rect 13001 7973 13035 8007
rect 19993 7973 20027 8007
rect 1685 7905 1719 7939
rect 2697 7905 2731 7939
rect 5549 7905 5583 7939
rect 5733 7905 5767 7939
rect 7113 7905 7147 7939
rect 7297 7905 7331 7939
rect 8309 7905 8343 7939
rect 20453 7905 20487 7939
rect 20545 7905 20579 7939
rect 1777 7837 1811 7871
rect 2881 7837 2915 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 10066 7837 10100 7871
rect 10333 7837 10367 7871
rect 11989 7837 12023 7871
rect 12265 7837 12299 7871
rect 13645 7837 13679 7871
rect 17969 7837 18003 7871
rect 21281 7837 21315 7871
rect 2789 7769 2823 7803
rect 8033 7769 8067 7803
rect 11722 7769 11756 7803
rect 13369 7769 13403 7803
rect 17724 7769 17758 7803
rect 18797 7769 18831 7803
rect 19625 7769 19659 7803
rect 20361 7769 20395 7803
rect 21097 7769 21131 7803
rect 1869 7701 1903 7735
rect 3249 7701 3283 7735
rect 3801 7701 3835 7735
rect 5825 7701 5859 7735
rect 6193 7701 6227 7735
rect 6653 7701 6687 7735
rect 7021 7701 7055 7735
rect 8125 7701 8159 7735
rect 14289 7701 14323 7735
rect 14657 7701 14691 7735
rect 15485 7701 15519 7735
rect 16221 7701 16255 7735
rect 18337 7701 18371 7735
rect 19533 7701 19567 7735
rect 1593 7497 1627 7531
rect 2329 7497 2363 7531
rect 3341 7497 3375 7531
rect 3985 7497 4019 7531
rect 4353 7497 4387 7531
rect 6009 7497 6043 7531
rect 15393 7497 15427 7531
rect 16313 7497 16347 7531
rect 18061 7497 18095 7531
rect 19257 7497 19291 7531
rect 19625 7497 19659 7531
rect 5641 7429 5675 7463
rect 7389 7429 7423 7463
rect 13185 7429 13219 7463
rect 16948 7429 16982 7463
rect 19165 7429 19199 7463
rect 19901 7429 19935 7463
rect 20085 7429 20119 7463
rect 1501 7361 1535 7395
rect 3433 7361 3467 7395
rect 7941 7361 7975 7395
rect 8493 7361 8527 7395
rect 10526 7361 10560 7395
rect 12642 7361 12676 7395
rect 12909 7361 12943 7395
rect 13645 7361 13679 7395
rect 13912 7361 13946 7395
rect 16129 7361 16163 7395
rect 16681 7361 16715 7395
rect 20545 7361 20579 7395
rect 2053 7293 2087 7327
rect 2237 7293 2271 7327
rect 3617 7293 3651 7327
rect 4445 7293 4479 7327
rect 4629 7293 4663 7327
rect 5365 7293 5399 7327
rect 5549 7293 5583 7327
rect 10793 7293 10827 7327
rect 18337 7293 18371 7327
rect 18981 7293 19015 7327
rect 20821 7293 20855 7327
rect 8861 7225 8895 7259
rect 2697 7157 2731 7191
rect 2973 7157 3007 7191
rect 6377 7157 6411 7191
rect 7021 7157 7055 7191
rect 8125 7157 8159 7191
rect 9413 7157 9447 7191
rect 11069 7157 11103 7191
rect 11529 7157 11563 7191
rect 15025 7157 15059 7191
rect 15761 7157 15795 7191
rect 2145 6953 2179 6987
rect 2421 6953 2455 6987
rect 7481 6953 7515 6987
rect 8493 6953 8527 6987
rect 9229 6953 9263 6987
rect 18889 6953 18923 6987
rect 12081 6885 12115 6919
rect 3065 6817 3099 6851
rect 4813 6817 4847 6851
rect 5825 6817 5859 6851
rect 6653 6817 6687 6851
rect 8125 6817 8159 6851
rect 13461 6817 13495 6851
rect 14105 6817 14139 6851
rect 14565 6817 14599 6851
rect 17601 6817 17635 6851
rect 18245 6817 18279 6851
rect 19625 6817 19659 6851
rect 19809 6817 19843 6851
rect 20821 6817 20855 6851
rect 1501 6749 1535 6783
rect 1961 6749 1995 6783
rect 2789 6749 2823 6783
rect 4629 6749 4663 6783
rect 5641 6749 5675 6783
rect 10342 6749 10376 6783
rect 10609 6749 10643 6783
rect 13194 6749 13228 6783
rect 14832 6749 14866 6783
rect 16681 6749 16715 6783
rect 17325 6749 17359 6783
rect 20545 6749 20579 6783
rect 1685 6681 1719 6715
rect 6745 6681 6779 6715
rect 7941 6681 7975 6715
rect 11805 6681 11839 6715
rect 17417 6681 17451 6715
rect 19901 6681 19935 6715
rect 2881 6613 2915 6647
rect 3893 6613 3927 6647
rect 4169 6613 4203 6647
rect 4537 6613 4571 6647
rect 5181 6613 5215 6647
rect 5549 6613 5583 6647
rect 6837 6613 6871 6647
rect 7205 6613 7239 6647
rect 7849 6613 7883 6647
rect 10977 6613 11011 6647
rect 11253 6613 11287 6647
rect 15945 6613 15979 6647
rect 16497 6613 16531 6647
rect 16957 6613 16991 6647
rect 18429 6613 18463 6647
rect 18521 6613 18555 6647
rect 20269 6613 20303 6647
rect 2605 6409 2639 6443
rect 3065 6409 3099 6443
rect 4353 6409 4387 6443
rect 13461 6409 13495 6443
rect 13737 6409 13771 6443
rect 15117 6409 15151 6443
rect 16313 6409 16347 6443
rect 16957 6409 16991 6443
rect 17417 6409 17451 6443
rect 20637 6409 20671 6443
rect 21097 6409 21131 6443
rect 1869 6341 1903 6375
rect 5641 6341 5675 6375
rect 8585 6341 8619 6375
rect 17049 6341 17083 6375
rect 18337 6341 18371 6375
rect 20094 6341 20128 6375
rect 1961 6273 1995 6307
rect 2973 6273 3007 6307
rect 3709 6273 3743 6307
rect 4169 6273 4203 6307
rect 4629 6273 4663 6307
rect 5733 6273 5767 6307
rect 6561 6273 6595 6307
rect 7573 6273 7607 6307
rect 9873 6273 9907 6307
rect 12348 6273 12382 6307
rect 14657 6273 14691 6307
rect 15301 6273 15335 6307
rect 15945 6273 15979 6307
rect 21005 6273 21039 6307
rect 1777 6205 1811 6239
rect 3249 6205 3283 6239
rect 5825 6205 5859 6239
rect 7389 6205 7423 6239
rect 7481 6205 7515 6239
rect 8309 6205 8343 6239
rect 8493 6205 8527 6239
rect 12081 6205 12115 6239
rect 15669 6205 15703 6239
rect 15853 6205 15887 6239
rect 16865 6205 16899 6239
rect 18153 6205 18187 6239
rect 18245 6205 18279 6239
rect 20361 6205 20395 6239
rect 21189 6205 21223 6239
rect 2329 6137 2363 6171
rect 3893 6137 3927 6171
rect 4813 6137 4847 6171
rect 6377 6137 6411 6171
rect 7941 6137 7975 6171
rect 8953 6137 8987 6171
rect 18705 6137 18739 6171
rect 5273 6069 5307 6103
rect 6929 6069 6963 6103
rect 9229 6069 9263 6103
rect 10241 6069 10275 6103
rect 10517 6069 10551 6103
rect 10977 6069 11011 6103
rect 11529 6069 11563 6103
rect 14381 6069 14415 6103
rect 14841 6069 14875 6103
rect 18981 6069 19015 6103
rect 3801 5865 3835 5899
rect 4261 5865 4295 5899
rect 4721 5865 4755 5899
rect 5825 5865 5859 5899
rect 16129 5865 16163 5899
rect 17969 5865 18003 5899
rect 6837 5797 6871 5831
rect 7941 5797 7975 5831
rect 9229 5797 9263 5831
rect 9597 5797 9631 5831
rect 19349 5797 19383 5831
rect 21097 5797 21131 5831
rect 1869 5729 1903 5763
rect 1961 5729 1995 5763
rect 3341 5729 3375 5763
rect 6469 5729 6503 5763
rect 12173 5729 12207 5763
rect 3985 5661 4019 5695
rect 4445 5661 4479 5695
rect 4905 5661 4939 5695
rect 7021 5661 7055 5695
rect 8401 5661 8435 5695
rect 10977 5661 11011 5695
rect 11253 5661 11287 5695
rect 13277 5661 13311 5695
rect 13737 5661 13771 5695
rect 15577 5661 15611 5695
rect 17509 5661 17543 5695
rect 17785 5661 17819 5695
rect 18245 5661 18279 5695
rect 18881 5661 18915 5695
rect 20729 5661 20763 5695
rect 3065 5593 3099 5627
rect 6193 5593 6227 5627
rect 7573 5593 7607 5627
rect 10710 5593 10744 5627
rect 15310 5593 15344 5627
rect 17242 5593 17276 5627
rect 20462 5593 20496 5627
rect 21281 5593 21315 5627
rect 2053 5525 2087 5559
rect 2421 5525 2455 5559
rect 2697 5525 2731 5559
rect 3157 5525 3191 5559
rect 5365 5525 5399 5559
rect 6285 5525 6319 5559
rect 8217 5525 8251 5559
rect 11621 5525 11655 5559
rect 12725 5525 12759 5559
rect 13553 5525 13587 5559
rect 14197 5525 14231 5559
rect 18429 5525 18463 5559
rect 18705 5525 18739 5559
rect 3249 5321 3283 5355
rect 4261 5321 4295 5355
rect 4353 5321 4387 5355
rect 5365 5321 5399 5355
rect 6377 5321 6411 5355
rect 7573 5321 7607 5355
rect 8309 5321 8343 5355
rect 11529 5321 11563 5355
rect 11897 5321 11931 5355
rect 16865 5321 16899 5355
rect 19993 5321 20027 5355
rect 20361 5321 20395 5355
rect 20637 5321 20671 5355
rect 21097 5321 21131 5355
rect 1501 5253 1535 5287
rect 2605 5253 2639 5287
rect 13584 5253 13618 5287
rect 21005 5253 21039 5287
rect 5457 5185 5491 5219
rect 6561 5185 6595 5219
rect 7113 5185 7147 5219
rect 7757 5185 7791 5219
rect 8125 5185 8159 5219
rect 8585 5185 8619 5219
rect 9413 5185 9447 5219
rect 9669 5185 9703 5219
rect 14381 5185 14415 5219
rect 14841 5185 14875 5219
rect 15485 5185 15519 5219
rect 15761 5185 15795 5219
rect 16681 5185 16715 5219
rect 17141 5185 17175 5219
rect 17601 5185 17635 5219
rect 18337 5185 18371 5219
rect 18889 5185 18923 5219
rect 2329 5117 2363 5151
rect 2513 5117 2547 5151
rect 4169 5117 4203 5151
rect 5641 5117 5675 5151
rect 13829 5117 13863 5151
rect 19717 5117 19751 5151
rect 19901 5117 19935 5151
rect 21189 5117 21223 5151
rect 8769 5049 8803 5083
rect 12449 5049 12483 5083
rect 15301 5049 15335 5083
rect 18521 5049 18555 5083
rect 1593 4981 1627 5015
rect 2973 4981 3007 5015
rect 4721 4981 4755 5015
rect 4997 4981 5031 5015
rect 7297 4981 7331 5015
rect 9137 4981 9171 5015
rect 10793 4981 10827 5015
rect 11161 4981 11195 5015
rect 14565 4981 14599 5015
rect 15025 4981 15059 5015
rect 15945 4981 15979 5015
rect 16313 4981 16347 5015
rect 17325 4981 17359 5015
rect 17785 4981 17819 5015
rect 19073 4981 19107 5015
rect 3249 4777 3283 4811
rect 3985 4777 4019 4811
rect 6377 4777 6411 4811
rect 7573 4777 7607 4811
rect 9965 4777 9999 4811
rect 10425 4777 10459 4811
rect 14841 4777 14875 4811
rect 15117 4777 15151 4811
rect 7297 4709 7331 4743
rect 9689 4709 9723 4743
rect 19441 4709 19475 4743
rect 21097 4709 21131 4743
rect 1961 4641 1995 4675
rect 2697 4641 2731 4675
rect 4629 4641 4663 4675
rect 4813 4641 4847 4675
rect 5825 4641 5859 4675
rect 5917 4641 5951 4675
rect 9137 4641 9171 4675
rect 11805 4641 11839 4675
rect 2237 4573 2271 4607
rect 2881 4573 2915 4607
rect 3801 4573 3835 4607
rect 4905 4573 4939 4607
rect 6837 4573 6871 4607
rect 7113 4573 7147 4607
rect 7757 4573 7791 4607
rect 8401 4573 8435 4607
rect 11549 4573 11583 4607
rect 13645 4573 13679 4607
rect 14381 4573 14415 4607
rect 14657 4573 14691 4607
rect 16497 4573 16531 4607
rect 18245 4573 18279 4607
rect 18521 4573 18555 4607
rect 20821 4573 20855 4607
rect 21281 4573 21315 4607
rect 2789 4505 2823 4539
rect 6009 4505 6043 4539
rect 9321 4505 9355 4539
rect 13378 4505 13412 4539
rect 16230 4505 16264 4539
rect 18000 4505 18034 4539
rect 20576 4505 20610 4539
rect 5273 4437 5307 4471
rect 6653 4437 6687 4471
rect 8217 4437 8251 4471
rect 9229 4437 9263 4471
rect 12265 4437 12299 4471
rect 14197 4437 14231 4471
rect 16865 4437 16899 4471
rect 18705 4437 18739 4471
rect 1593 4233 1627 4267
rect 3801 4233 3835 4267
rect 6009 4233 6043 4267
rect 7849 4233 7883 4267
rect 17509 4233 17543 4267
rect 3249 4165 3283 4199
rect 3893 4165 3927 4199
rect 8953 4165 8987 4199
rect 10894 4165 10928 4199
rect 11713 4165 11747 4199
rect 20729 4165 20763 4199
rect 1409 4097 1443 4131
rect 2513 4097 2547 4131
rect 4537 4097 4571 4131
rect 4905 4097 4939 4131
rect 5365 4097 5399 4131
rect 5825 4097 5859 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 7665 4097 7699 4131
rect 8309 4097 8343 4131
rect 11529 4097 11563 4131
rect 12265 4097 12299 4131
rect 12817 4097 12851 4131
rect 13277 4097 13311 4131
rect 13737 4097 13771 4131
rect 15310 4097 15344 4131
rect 15577 4097 15611 4131
rect 15853 4097 15887 4131
rect 16681 4097 16715 4131
rect 17601 4097 17635 4131
rect 18153 4097 18187 4131
rect 19645 4097 19679 4131
rect 19901 4097 19935 4131
rect 20821 4097 20855 4131
rect 2329 4029 2363 4063
rect 2421 4029 2455 4063
rect 3709 4029 3743 4063
rect 8677 4029 8711 4063
rect 8861 4029 8895 4063
rect 11161 4029 11195 4063
rect 17785 4029 17819 4063
rect 20913 4029 20947 4063
rect 2881 3961 2915 3995
rect 5089 3961 5123 3995
rect 6561 3961 6595 3995
rect 9321 3961 9355 3995
rect 9781 3961 9815 3995
rect 13921 3961 13955 3995
rect 14197 3961 14231 3995
rect 16865 3961 16899 3995
rect 18521 3961 18555 3995
rect 4261 3893 4295 3927
rect 5549 3893 5583 3927
rect 7205 3893 7239 3927
rect 8125 3893 8159 3927
rect 12081 3893 12115 3927
rect 13001 3893 13035 3927
rect 13461 3893 13495 3927
rect 16037 3893 16071 3927
rect 17141 3893 17175 3927
rect 20361 3893 20395 3927
rect 2605 3689 2639 3723
rect 2973 3689 3007 3723
rect 4905 3689 4939 3723
rect 8125 3689 8159 3723
rect 13737 3689 13771 3723
rect 14381 3689 14415 3723
rect 15577 3689 15611 3723
rect 17877 3689 17911 3723
rect 19625 3689 19659 3723
rect 20637 3689 20671 3723
rect 3893 3621 3927 3655
rect 10701 3621 10735 3655
rect 12541 3621 12575 3655
rect 16773 3621 16807 3655
rect 19349 3621 19383 3655
rect 2053 3553 2087 3587
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 5457 3553 5491 3587
rect 6101 3553 6135 3587
rect 9413 3553 9447 3587
rect 9505 3553 9539 3587
rect 12081 3553 12115 3587
rect 15025 3553 15059 3587
rect 17233 3553 17267 3587
rect 17417 3553 17451 3587
rect 18797 3553 18831 3587
rect 20269 3553 20303 3587
rect 21189 3553 21223 3587
rect 2145 3485 2179 3519
rect 3249 3485 3283 3519
rect 4261 3485 4295 3519
rect 6377 3485 6411 3519
rect 7021 3485 7055 3519
rect 7481 3485 7515 3519
rect 7941 3485 7975 3519
rect 8585 3485 8619 3519
rect 10149 3485 10183 3519
rect 12357 3485 12391 3519
rect 13001 3485 13035 3519
rect 13553 3485 13587 3519
rect 14749 3485 14783 3519
rect 15393 3485 15427 3519
rect 16037 3485 16071 3519
rect 16589 3485 16623 3519
rect 17509 3485 17543 3519
rect 21005 3485 21039 3519
rect 21097 3485 21131 3519
rect 1593 3417 1627 3451
rect 2237 3417 2271 3451
rect 11836 3417 11870 3451
rect 14841 3417 14875 3451
rect 18521 3417 18555 3451
rect 18613 3417 18647 3451
rect 20085 3417 20119 3451
rect 3433 3349 3467 3383
rect 5273 3349 5307 3383
rect 5365 3349 5399 3383
rect 6285 3349 6319 3383
rect 6745 3349 6779 3383
rect 7205 3349 7239 3383
rect 7665 3349 7699 3383
rect 8401 3349 8435 3383
rect 8953 3349 8987 3383
rect 9321 3349 9355 3383
rect 10333 3349 10367 3383
rect 12817 3349 12851 3383
rect 16221 3349 16255 3383
rect 18153 3349 18187 3383
rect 19993 3349 20027 3383
rect 2789 3145 2823 3179
rect 3249 3145 3283 3179
rect 3801 3145 3835 3179
rect 4261 3145 4295 3179
rect 13553 3145 13587 3179
rect 13921 3145 13955 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 17693 3145 17727 3179
rect 6837 3077 6871 3111
rect 10894 3077 10928 3111
rect 18061 3077 18095 3111
rect 18153 3077 18187 3111
rect 1961 3009 1995 3043
rect 2605 3009 2639 3043
rect 3065 3009 3099 3043
rect 3893 3009 3927 3043
rect 5365 3009 5399 3043
rect 5825 3009 5859 3043
rect 6745 3009 6779 3043
rect 7389 3009 7423 3043
rect 7849 3009 7883 3043
rect 8493 2993 8527 3027
rect 8953 3009 8987 3043
rect 9229 3009 9263 3043
rect 11161 3009 11195 3043
rect 12642 3009 12676 3043
rect 12909 3009 12943 3043
rect 14197 3009 14231 3043
rect 14749 3009 14783 3043
rect 15301 3009 15335 3043
rect 15853 3009 15887 3043
rect 19073 3009 19107 3043
rect 20177 3009 20211 3043
rect 2237 2941 2271 2975
rect 3617 2941 3651 2975
rect 5089 2941 5123 2975
rect 7021 2941 7055 2975
rect 13277 2941 13311 2975
rect 13461 2941 13495 2975
rect 17141 2941 17175 2975
rect 17325 2941 17359 2975
rect 18245 2941 18279 2975
rect 19165 2941 19199 2975
rect 19349 2941 19383 2975
rect 20361 2941 20395 2975
rect 6009 2873 6043 2907
rect 11529 2873 11563 2907
rect 16037 2873 16071 2907
rect 18705 2873 18739 2907
rect 6377 2805 6411 2839
rect 7573 2805 7607 2839
rect 8033 2805 8067 2839
rect 8309 2805 8343 2839
rect 8769 2805 8803 2839
rect 9413 2805 9447 2839
rect 9781 2805 9815 2839
rect 14381 2805 14415 2839
rect 14933 2805 14967 2839
rect 15485 2805 15519 2839
rect 21281 2805 21315 2839
rect 1869 2601 1903 2635
rect 9045 2601 9079 2635
rect 13645 2601 13679 2635
rect 15945 2601 15979 2635
rect 20545 2601 20579 2635
rect 2421 2533 2455 2567
rect 2973 2533 3007 2567
rect 6837 2533 6871 2567
rect 9781 2533 9815 2567
rect 15393 2533 15427 2567
rect 16865 2533 16899 2567
rect 4629 2465 4663 2499
rect 5457 2465 5491 2499
rect 7941 2465 7975 2499
rect 11989 2465 12023 2499
rect 13093 2465 13127 2499
rect 13185 2465 13219 2499
rect 1685 2397 1719 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 4353 2397 4387 2431
rect 5733 2397 5767 2431
rect 6653 2397 6687 2431
rect 7665 2397 7699 2431
rect 8585 2397 8619 2431
rect 9505 2397 9539 2431
rect 10333 2397 10367 2431
rect 10609 2397 10643 2431
rect 13277 2397 13311 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 19257 2397 19291 2431
rect 19809 2397 19843 2431
rect 20361 2397 20395 2431
rect 20913 2397 20947 2431
rect 2237 2329 2271 2363
rect 9965 2329 9999 2363
rect 3433 2261 3467 2295
rect 8401 2261 8435 2295
rect 9321 2261 9355 2295
rect 11621 2261 11655 2295
rect 12173 2261 12207 2295
rect 12265 2261 12299 2295
rect 12633 2261 12667 2295
rect 14289 2261 14323 2295
rect 14841 2261 14875 2295
rect 17417 2261 17451 2295
rect 17969 2261 18003 2295
rect 18521 2261 18555 2295
rect 19441 2261 19475 2295
rect 19993 2261 20027 2295
rect 21097 2261 21131 2295
<< metal1 >>
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 1104 20624 22056 20646
rect 2038 20584 2044 20596
rect 1999 20556 2044 20584
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 17037 20587 17095 20593
rect 17037 20553 17049 20587
rect 17083 20584 17095 20587
rect 17218 20584 17224 20596
rect 17083 20556 17224 20584
rect 17083 20553 17095 20556
rect 17037 20547 17095 20553
rect 17218 20544 17224 20556
rect 17276 20544 17282 20596
rect 18877 20587 18935 20593
rect 18877 20553 18889 20587
rect 18923 20553 18935 20587
rect 20162 20584 20168 20596
rect 20123 20556 20168 20584
rect 18877 20547 18935 20553
rect 15565 20519 15623 20525
rect 15565 20485 15577 20519
rect 15611 20516 15623 20519
rect 18892 20516 18920 20547
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 21174 20516 21180 20528
rect 15611 20488 18736 20516
rect 18892 20488 21180 20516
rect 15611 20485 15623 20488
rect 15565 20479 15623 20485
rect 18708 20460 18736 20488
rect 21174 20476 21180 20488
rect 21232 20476 21238 20528
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 2130 20448 2136 20460
rect 1719 20420 2136 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 2130 20408 2136 20420
rect 2188 20408 2194 20460
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20448 2283 20451
rect 2685 20451 2743 20457
rect 2271 20420 2544 20448
rect 2271 20417 2283 20420
rect 2225 20411 2283 20417
rect 2516 20321 2544 20420
rect 2685 20417 2697 20451
rect 2731 20417 2743 20451
rect 2958 20448 2964 20460
rect 2919 20420 2964 20448
rect 2685 20411 2743 20417
rect 2700 20380 2728 20411
rect 2958 20408 2964 20420
rect 3016 20448 3022 20460
rect 4157 20451 4215 20457
rect 4157 20448 4169 20451
rect 3016 20420 4169 20448
rect 3016 20408 3022 20420
rect 4157 20417 4169 20420
rect 4203 20417 4215 20451
rect 4157 20411 4215 20417
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5859 20420 6377 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 16850 20448 16856 20460
rect 16811 20420 16856 20448
rect 6365 20411 6423 20417
rect 16850 20408 16856 20420
rect 16908 20408 16914 20460
rect 17770 20448 17776 20460
rect 17731 20420 17776 20448
rect 17770 20408 17776 20420
rect 17828 20408 17834 20460
rect 18690 20448 18696 20460
rect 18651 20420 18696 20448
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 19518 20448 19524 20460
rect 19479 20420 19524 20448
rect 19518 20408 19524 20420
rect 19576 20408 19582 20460
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20417 20039 20451
rect 20530 20448 20536 20460
rect 20491 20420 20536 20448
rect 19981 20411 20039 20417
rect 3789 20383 3847 20389
rect 3789 20380 3801 20383
rect 2700 20352 3801 20380
rect 3789 20349 3801 20352
rect 3835 20380 3847 20383
rect 4062 20380 4068 20392
rect 3835 20352 4068 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 4062 20340 4068 20352
rect 4120 20340 4126 20392
rect 4522 20380 4528 20392
rect 4483 20352 4528 20380
rect 4522 20340 4528 20352
rect 4580 20340 4586 20392
rect 7834 20380 7840 20392
rect 7795 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 17865 20383 17923 20389
rect 17865 20380 17877 20383
rect 15856 20352 17877 20380
rect 2501 20315 2559 20321
rect 2501 20281 2513 20315
rect 2547 20281 2559 20315
rect 2501 20275 2559 20281
rect 5997 20315 6055 20321
rect 5997 20281 6009 20315
rect 6043 20312 6055 20315
rect 14642 20312 14648 20324
rect 6043 20284 14648 20312
rect 6043 20281 6055 20284
rect 5997 20275 6055 20281
rect 14642 20272 14648 20284
rect 14700 20272 14706 20324
rect 1486 20244 1492 20256
rect 1447 20216 1492 20244
rect 1486 20204 1492 20216
rect 1544 20204 1550 20256
rect 3142 20244 3148 20256
rect 3103 20216 3148 20244
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 12437 20247 12495 20253
rect 12437 20213 12449 20247
rect 12483 20244 12495 20247
rect 12526 20244 12532 20256
rect 12483 20216 12532 20244
rect 12483 20213 12495 20216
rect 12437 20207 12495 20213
rect 12526 20204 12532 20216
rect 12584 20204 12590 20256
rect 12986 20204 12992 20256
rect 13044 20244 13050 20256
rect 15856 20244 15884 20352
rect 17865 20349 17877 20352
rect 17911 20349 17923 20383
rect 17865 20343 17923 20349
rect 17957 20383 18015 20389
rect 17957 20349 17969 20383
rect 18003 20349 18015 20383
rect 17957 20343 18015 20349
rect 15933 20315 15991 20321
rect 15933 20281 15945 20315
rect 15979 20312 15991 20315
rect 16390 20312 16396 20324
rect 15979 20284 16396 20312
rect 15979 20281 15991 20284
rect 15933 20275 15991 20281
rect 16390 20272 16396 20284
rect 16448 20312 16454 20324
rect 17972 20312 18000 20343
rect 19996 20312 20024 20411
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 16448 20284 18000 20312
rect 18156 20284 20024 20312
rect 16448 20272 16454 20284
rect 16209 20247 16267 20253
rect 16209 20244 16221 20247
rect 13044 20216 16221 20244
rect 13044 20204 13050 20216
rect 16209 20213 16221 20216
rect 16255 20213 16267 20247
rect 16209 20207 16267 20213
rect 16482 20204 16488 20256
rect 16540 20244 16546 20256
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 16540 20216 17417 20244
rect 16540 20204 16546 20216
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17405 20207 17463 20213
rect 17678 20204 17684 20256
rect 17736 20244 17742 20256
rect 18156 20244 18184 20284
rect 17736 20216 18184 20244
rect 19705 20247 19763 20253
rect 17736 20204 17742 20216
rect 19705 20213 19717 20247
rect 19751 20244 19763 20247
rect 20438 20244 20444 20256
rect 19751 20216 20444 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 20438 20204 20444 20216
rect 20496 20204 20502 20256
rect 20714 20244 20720 20256
rect 20675 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21266 20244 21272 20256
rect 21227 20216 21272 20244
rect 21266 20204 21272 20216
rect 21324 20204 21330 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1946 20000 1952 20052
rect 2004 20040 2010 20052
rect 2041 20043 2099 20049
rect 2041 20040 2053 20043
rect 2004 20012 2053 20040
rect 2004 20000 2010 20012
rect 2041 20009 2053 20012
rect 2087 20009 2099 20043
rect 2041 20003 2099 20009
rect 12713 20043 12771 20049
rect 12713 20009 12725 20043
rect 12759 20040 12771 20043
rect 15289 20043 15347 20049
rect 12759 20012 15148 20040
rect 12759 20009 12771 20012
rect 12713 20003 12771 20009
rect 9953 19975 10011 19981
rect 9953 19941 9965 19975
rect 9999 19972 10011 19975
rect 12894 19972 12900 19984
rect 9999 19944 12900 19972
rect 9999 19941 10011 19944
rect 9953 19935 10011 19941
rect 12894 19932 12900 19944
rect 12952 19932 12958 19984
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 15010 19972 15016 19984
rect 13771 19944 15016 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 15010 19932 15016 19944
rect 15068 19932 15074 19984
rect 7653 19907 7711 19913
rect 7653 19873 7665 19907
rect 7699 19904 7711 19907
rect 8478 19904 8484 19916
rect 7699 19876 8484 19904
rect 7699 19873 7711 19876
rect 7653 19867 7711 19873
rect 8478 19864 8484 19876
rect 8536 19864 8542 19916
rect 10502 19904 10508 19916
rect 10463 19876 10508 19904
rect 10502 19864 10508 19876
rect 10560 19864 10566 19916
rect 11238 19864 11244 19916
rect 11296 19904 11302 19916
rect 11790 19904 11796 19916
rect 11296 19876 11796 19904
rect 11296 19864 11302 19876
rect 11790 19864 11796 19876
rect 11848 19864 11854 19916
rect 11885 19907 11943 19913
rect 11885 19873 11897 19907
rect 11931 19873 11943 19907
rect 14734 19904 14740 19916
rect 14695 19876 14740 19904
rect 11885 19867 11943 19873
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 1673 19799 1731 19805
rect 1688 19768 1716 19799
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2677 19839 2735 19845
rect 2677 19805 2689 19839
rect 2723 19805 2735 19839
rect 2677 19799 2735 19805
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 4706 19836 4712 19848
rect 3283 19808 4712 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 2700 19768 2728 19799
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 9858 19796 9864 19848
rect 9916 19836 9922 19848
rect 11900 19836 11928 19867
rect 14734 19864 14740 19876
rect 14792 19864 14798 19916
rect 15120 19904 15148 20012
rect 15289 20009 15301 20043
rect 15335 20040 15347 20043
rect 19518 20040 19524 20052
rect 15335 20012 19524 20040
rect 15335 20009 15347 20012
rect 15289 20003 15347 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 20165 20043 20223 20049
rect 20165 20009 20177 20043
rect 20211 20040 20223 20043
rect 21082 20040 21088 20052
rect 20211 20012 21088 20040
rect 20211 20009 20223 20012
rect 20165 20003 20223 20009
rect 21082 20000 21088 20012
rect 21140 20000 21146 20052
rect 15194 19932 15200 19984
rect 15252 19972 15258 19984
rect 16206 19972 16212 19984
rect 15252 19944 16212 19972
rect 15252 19932 15258 19944
rect 16206 19932 16212 19944
rect 16264 19932 16270 19984
rect 20530 19972 20536 19984
rect 16316 19944 20536 19972
rect 16316 19904 16344 19944
rect 20530 19932 20536 19944
rect 20588 19932 20594 19984
rect 20622 19932 20628 19984
rect 20680 19972 20686 19984
rect 20717 19975 20775 19981
rect 20717 19972 20729 19975
rect 20680 19944 20729 19972
rect 20680 19932 20686 19944
rect 20717 19941 20729 19944
rect 20763 19941 20775 19975
rect 20717 19935 20775 19941
rect 16669 19907 16727 19913
rect 16669 19904 16681 19907
rect 15120 19876 16344 19904
rect 16546 19876 16681 19904
rect 12526 19836 12532 19848
rect 9916 19808 11928 19836
rect 12487 19808 12532 19836
rect 9916 19796 9922 19808
rect 12526 19796 12532 19808
rect 12584 19796 12590 19848
rect 12986 19836 12992 19848
rect 12947 19808 12992 19836
rect 12986 19796 12992 19808
rect 13044 19796 13050 19848
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19836 13599 19839
rect 13587 19808 14136 19836
rect 13587 19805 13599 19808
rect 13541 19799 13599 19805
rect 4522 19768 4528 19780
rect 1688 19740 2544 19768
rect 2700 19740 3096 19768
rect 4483 19740 4528 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2516 19709 2544 19740
rect 3068 19709 3096 19740
rect 4522 19728 4528 19740
rect 4580 19728 4586 19780
rect 10321 19771 10379 19777
rect 10321 19737 10333 19771
rect 10367 19768 10379 19771
rect 10367 19740 11376 19768
rect 10367 19737 10379 19740
rect 10321 19731 10379 19737
rect 2501 19703 2559 19709
rect 2501 19669 2513 19703
rect 2547 19669 2559 19703
rect 2501 19663 2559 19669
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19669 3111 19703
rect 3878 19700 3884 19712
rect 3839 19672 3884 19700
rect 3053 19663 3111 19669
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 4246 19700 4252 19712
rect 4207 19672 4252 19700
rect 4246 19660 4252 19672
rect 4304 19660 4310 19712
rect 4890 19700 4896 19712
rect 4851 19672 4896 19700
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 5442 19660 5448 19712
rect 5500 19700 5506 19712
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 5500 19672 7757 19700
rect 5500 19660 5506 19672
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 7745 19663 7803 19669
rect 7926 19660 7932 19712
rect 7984 19700 7990 19712
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7984 19672 8217 19700
rect 7984 19660 7990 19672
rect 8205 19669 8217 19672
rect 8251 19669 8263 19703
rect 8205 19663 8263 19669
rect 10410 19660 10416 19712
rect 10468 19700 10474 19712
rect 11057 19703 11115 19709
rect 10468 19672 10513 19700
rect 10468 19660 10474 19672
rect 11057 19669 11069 19703
rect 11103 19700 11115 19703
rect 11238 19700 11244 19712
rect 11103 19672 11244 19700
rect 11103 19669 11115 19672
rect 11057 19663 11115 19669
rect 11238 19660 11244 19672
rect 11296 19660 11302 19712
rect 11348 19709 11376 19740
rect 11333 19703 11391 19709
rect 11333 19669 11345 19703
rect 11379 19669 11391 19703
rect 11698 19700 11704 19712
rect 11659 19672 11704 19700
rect 11333 19663 11391 19669
rect 11698 19660 11704 19672
rect 11756 19660 11762 19712
rect 13170 19700 13176 19712
rect 13131 19672 13176 19700
rect 13170 19660 13176 19672
rect 13228 19660 13234 19712
rect 14108 19709 14136 19808
rect 14826 19796 14832 19848
rect 14884 19836 14890 19848
rect 15105 19839 15163 19845
rect 15105 19836 15117 19839
rect 14884 19808 15117 19836
rect 14884 19796 14890 19808
rect 15105 19805 15117 19808
rect 15151 19805 15163 19839
rect 15105 19799 15163 19805
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16546 19836 16574 19876
rect 16669 19873 16681 19876
rect 16715 19873 16727 19907
rect 17310 19904 17316 19916
rect 17271 19876 17316 19904
rect 16669 19867 16727 19873
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 17770 19864 17776 19916
rect 17828 19904 17834 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 17828 19876 18705 19904
rect 17828 19864 17834 19876
rect 18693 19873 18705 19876
rect 18739 19873 18751 19907
rect 18693 19867 18751 19873
rect 18874 19864 18880 19916
rect 18932 19904 18938 19916
rect 18932 19876 21128 19904
rect 18932 19864 18938 19876
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 15988 19808 16574 19836
rect 17972 19808 19257 19836
rect 15988 19796 15994 19808
rect 14461 19771 14519 19777
rect 14461 19737 14473 19771
rect 14507 19768 14519 19771
rect 14507 19740 16160 19768
rect 14507 19737 14519 19740
rect 14461 19731 14519 19737
rect 14093 19703 14151 19709
rect 14093 19669 14105 19703
rect 14139 19669 14151 19703
rect 14550 19700 14556 19712
rect 14511 19672 14556 19700
rect 14093 19663 14151 19669
rect 14550 19660 14556 19672
rect 14608 19660 14614 19712
rect 15841 19703 15899 19709
rect 15841 19669 15853 19703
rect 15887 19700 15899 19703
rect 15930 19700 15936 19712
rect 15887 19672 15936 19700
rect 15887 19669 15899 19672
rect 15841 19663 15899 19669
rect 15930 19660 15936 19672
rect 15988 19660 15994 19712
rect 16132 19709 16160 19740
rect 16206 19728 16212 19780
rect 16264 19768 16270 19780
rect 17862 19768 17868 19780
rect 16264 19740 17868 19768
rect 16264 19728 16270 19740
rect 17862 19728 17868 19740
rect 17920 19728 17926 19780
rect 16117 19703 16175 19709
rect 16117 19669 16129 19703
rect 16163 19669 16175 19703
rect 16482 19700 16488 19712
rect 16443 19672 16488 19700
rect 16117 19663 16175 19669
rect 16482 19660 16488 19672
rect 16540 19660 16546 19712
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19700 16635 19703
rect 16942 19700 16948 19712
rect 16623 19672 16948 19700
rect 16623 19669 16635 19672
rect 16577 19663 16635 19669
rect 16942 19660 16948 19672
rect 17000 19660 17006 19712
rect 17494 19700 17500 19712
rect 17455 19672 17500 19700
rect 17494 19660 17500 19672
rect 17552 19660 17558 19712
rect 17586 19660 17592 19712
rect 17644 19700 17650 19712
rect 17972 19709 18000 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19245 19799 19303 19805
rect 19444 19808 19993 19836
rect 17957 19703 18015 19709
rect 17644 19672 17689 19700
rect 17644 19660 17650 19672
rect 17957 19669 17969 19703
rect 18003 19669 18015 19703
rect 18230 19700 18236 19712
rect 18191 19672 18236 19700
rect 17957 19663 18015 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 19444 19709 19472 19808
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 20530 19836 20536 19848
rect 20491 19808 20536 19836
rect 19981 19799 20039 19805
rect 20530 19796 20536 19808
rect 20588 19796 20594 19848
rect 21100 19845 21128 19876
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 19429 19703 19487 19709
rect 19429 19669 19441 19703
rect 19475 19669 19487 19703
rect 19429 19663 19487 19669
rect 21269 19703 21327 19709
rect 21269 19669 21281 19703
rect 21315 19700 21327 19703
rect 21358 19700 21364 19712
rect 21315 19672 21364 19700
rect 21315 19669 21327 19672
rect 21269 19663 21327 19669
rect 21358 19660 21364 19672
rect 21416 19660 21422 19712
rect 1104 19610 22056 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2222 19456 2228 19508
rect 2280 19496 2286 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2280 19468 2973 19496
rect 2280 19456 2286 19468
rect 2961 19465 2973 19468
rect 3007 19465 3019 19499
rect 2961 19459 3019 19465
rect 3694 19456 3700 19508
rect 3752 19496 3758 19508
rect 4157 19499 4215 19505
rect 4157 19496 4169 19499
rect 3752 19468 4169 19496
rect 3752 19456 3758 19468
rect 4157 19465 4169 19468
rect 4203 19465 4215 19499
rect 4706 19496 4712 19508
rect 4667 19468 4712 19496
rect 4157 19459 4215 19465
rect 2130 19388 2136 19440
rect 2188 19428 2194 19440
rect 2188 19400 2544 19428
rect 2188 19388 2194 19400
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 1946 19360 1952 19372
rect 1719 19332 1952 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 2222 19360 2228 19372
rect 2183 19332 2228 19360
rect 2222 19320 2228 19332
rect 2280 19320 2286 19372
rect 1210 19184 1216 19236
rect 1268 19224 1274 19236
rect 2038 19224 2044 19236
rect 1268 19196 1624 19224
rect 1999 19196 2044 19224
rect 1268 19184 1274 19196
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1596 19156 1624 19196
rect 2038 19184 2044 19196
rect 2096 19184 2102 19236
rect 2516 19233 2544 19400
rect 2682 19360 2688 19372
rect 2643 19332 2688 19360
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 3145 19363 3203 19369
rect 3145 19329 3157 19363
rect 3191 19360 3203 19363
rect 3510 19360 3516 19372
rect 3191 19332 3516 19360
rect 3191 19329 3203 19332
rect 3145 19323 3203 19329
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 4172 19360 4200 19459
rect 4706 19456 4712 19468
rect 4764 19456 4770 19508
rect 5166 19496 5172 19508
rect 5127 19468 5172 19496
rect 5166 19456 5172 19468
rect 5224 19456 5230 19508
rect 7558 19496 7564 19508
rect 7519 19468 7564 19496
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 7926 19496 7932 19508
rect 7887 19468 7932 19496
rect 7926 19456 7932 19468
rect 7984 19456 7990 19508
rect 10410 19496 10416 19508
rect 10371 19468 10416 19496
rect 10410 19456 10416 19468
rect 10468 19456 10474 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 11793 19499 11851 19505
rect 11793 19496 11805 19499
rect 11756 19468 11805 19496
rect 11756 19456 11762 19468
rect 11793 19465 11805 19468
rect 11839 19465 11851 19499
rect 14366 19496 14372 19508
rect 14327 19468 14372 19496
rect 11793 19459 11851 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14826 19496 14832 19508
rect 14787 19468 14832 19496
rect 14826 19456 14832 19468
rect 14884 19456 14890 19508
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 17586 19496 17592 19508
rect 17451 19468 17592 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 17773 19499 17831 19505
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 18230 19496 18236 19508
rect 17819 19468 18236 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 18230 19456 18236 19468
rect 18288 19456 18294 19508
rect 18877 19499 18935 19505
rect 18877 19465 18889 19499
rect 18923 19465 18935 19499
rect 18877 19459 18935 19465
rect 19337 19499 19395 19505
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 19702 19496 19708 19508
rect 19383 19468 19708 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 5258 19388 5264 19440
rect 5316 19388 5322 19440
rect 13170 19388 13176 19440
rect 13228 19428 13234 19440
rect 17678 19428 17684 19440
rect 13228 19400 17684 19428
rect 13228 19388 13234 19400
rect 17678 19388 17684 19400
rect 17736 19388 17742 19440
rect 17862 19388 17868 19440
rect 17920 19428 17926 19440
rect 18892 19428 18920 19459
rect 19702 19456 19708 19468
rect 19760 19456 19766 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 20530 19496 20536 19508
rect 19843 19468 20536 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 20530 19456 20536 19468
rect 20588 19456 20594 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 20717 19499 20775 19505
rect 20717 19496 20729 19499
rect 20680 19468 20729 19496
rect 20680 19456 20686 19468
rect 20717 19465 20729 19468
rect 20763 19465 20775 19499
rect 20717 19459 20775 19465
rect 17920 19400 18828 19428
rect 18892 19400 20576 19428
rect 17920 19388 17926 19400
rect 5074 19360 5080 19372
rect 4172 19332 4292 19360
rect 5035 19332 5080 19360
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19292 3939 19295
rect 4154 19292 4160 19304
rect 3927 19264 4160 19292
rect 3927 19261 3939 19264
rect 3881 19255 3939 19261
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4264 19292 4292 19332
rect 5074 19320 5080 19332
rect 5132 19320 5138 19372
rect 4982 19292 4988 19304
rect 4264 19264 4988 19292
rect 4982 19252 4988 19264
rect 5040 19252 5046 19304
rect 5276 19301 5304 19388
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 9401 19363 9459 19369
rect 9401 19360 9413 19363
rect 8628 19332 9413 19360
rect 8628 19320 8634 19332
rect 9401 19329 9413 19332
rect 9447 19360 9459 19363
rect 10045 19363 10103 19369
rect 10045 19360 10057 19363
rect 9447 19332 10057 19360
rect 9447 19329 9459 19332
rect 9401 19323 9459 19329
rect 10045 19329 10057 19332
rect 10091 19329 10103 19363
rect 14458 19360 14464 19372
rect 14419 19332 14464 19360
rect 10045 19323 10103 19329
rect 14458 19320 14464 19332
rect 14516 19320 14522 19372
rect 18064 19360 18184 19364
rect 18690 19360 18696 19372
rect 17788 19336 18184 19360
rect 17788 19332 18092 19336
rect 5261 19295 5319 19301
rect 5261 19261 5273 19295
rect 5307 19261 5319 19295
rect 5261 19255 5319 19261
rect 5350 19252 5356 19304
rect 5408 19292 5414 19304
rect 8018 19292 8024 19304
rect 5408 19264 6776 19292
rect 7979 19264 8024 19292
rect 5408 19252 5414 19264
rect 2501 19227 2559 19233
rect 2501 19193 2513 19227
rect 2547 19193 2559 19227
rect 6362 19224 6368 19236
rect 2501 19187 2559 19193
rect 2746 19196 6368 19224
rect 2746 19156 2774 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 6748 19224 6776 19264
rect 8018 19252 8024 19264
rect 8076 19252 8082 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19292 8263 19295
rect 9490 19292 9496 19304
rect 8251 19264 9496 19292
rect 8251 19261 8263 19264
rect 8205 19255 8263 19261
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 9858 19292 9864 19304
rect 9819 19264 9864 19292
rect 9858 19252 9864 19264
rect 9916 19252 9922 19304
rect 9953 19295 10011 19301
rect 9953 19261 9965 19295
rect 9999 19292 10011 19295
rect 10689 19295 10747 19301
rect 10689 19292 10701 19295
rect 9999 19264 10701 19292
rect 9999 19261 10011 19264
rect 9953 19255 10011 19261
rect 10689 19261 10701 19264
rect 10735 19261 10747 19295
rect 12342 19292 12348 19304
rect 12303 19264 12348 19292
rect 10689 19255 10747 19261
rect 9968 19224 9996 19255
rect 12342 19252 12348 19264
rect 12400 19252 12406 19304
rect 14277 19295 14335 19301
rect 14277 19261 14289 19295
rect 14323 19292 14335 19295
rect 15470 19292 15476 19304
rect 14323 19264 15476 19292
rect 14323 19261 14335 19264
rect 14277 19255 14335 19261
rect 15470 19252 15476 19264
rect 15528 19252 15534 19304
rect 16761 19295 16819 19301
rect 16761 19261 16773 19295
rect 16807 19292 16819 19295
rect 17788 19292 17816 19332
rect 16807 19264 17816 19292
rect 16807 19261 16819 19264
rect 16761 19255 16819 19261
rect 17862 19252 17868 19304
rect 17920 19292 17926 19304
rect 18049 19295 18107 19301
rect 17920 19264 17965 19292
rect 17920 19252 17926 19264
rect 18049 19261 18061 19295
rect 18095 19261 18107 19295
rect 18156 19292 18184 19336
rect 18651 19332 18696 19360
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18800 19360 18828 19400
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 18800 19332 19165 19360
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 20070 19360 20076 19372
rect 19613 19323 19671 19329
rect 19720 19332 20076 19360
rect 18230 19292 18236 19304
rect 18156 19264 18236 19292
rect 18049 19255 18107 19261
rect 6748 19196 9996 19224
rect 15838 19184 15844 19236
rect 15896 19224 15902 19236
rect 16390 19224 16396 19236
rect 15896 19196 16396 19224
rect 15896 19184 15902 19196
rect 16390 19184 16396 19196
rect 16448 19224 16454 19236
rect 17218 19224 17224 19236
rect 16448 19196 17224 19224
rect 16448 19184 16454 19196
rect 17218 19184 17224 19196
rect 17276 19184 17282 19236
rect 17770 19184 17776 19236
rect 17828 19224 17834 19236
rect 18064 19224 18092 19255
rect 18230 19252 18236 19264
rect 18288 19292 18294 19304
rect 19628 19292 19656 19323
rect 18288 19264 19656 19292
rect 18288 19252 18294 19264
rect 19720 19224 19748 19332
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20548 19369 20576 19400
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20956 19332 21097 19360
rect 20956 19320 20962 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 17828 19196 18092 19224
rect 19536 19196 19748 19224
rect 17828 19184 17834 19196
rect 3510 19156 3516 19168
rect 1596 19128 2774 19156
rect 3423 19128 3516 19156
rect 3510 19116 3516 19128
rect 3568 19156 3574 19168
rect 4062 19156 4068 19168
rect 3568 19128 4068 19156
rect 3568 19116 3574 19128
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 4154 19116 4160 19168
rect 4212 19156 4218 19168
rect 4706 19156 4712 19168
rect 4212 19128 4712 19156
rect 4212 19116 4218 19128
rect 4706 19116 4712 19128
rect 4764 19156 4770 19168
rect 5350 19156 5356 19168
rect 4764 19128 5356 19156
rect 4764 19116 4770 19128
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 5718 19156 5724 19168
rect 5679 19128 5724 19156
rect 5718 19116 5724 19128
rect 5776 19116 5782 19168
rect 6457 19159 6515 19165
rect 6457 19125 6469 19159
rect 6503 19156 6515 19159
rect 6546 19156 6552 19168
rect 6503 19128 6552 19156
rect 6503 19125 6515 19128
rect 6457 19119 6515 19125
rect 6546 19116 6552 19128
rect 6604 19116 6610 19168
rect 11882 19116 11888 19168
rect 11940 19156 11946 19168
rect 12805 19159 12863 19165
rect 12805 19156 12817 19159
rect 11940 19128 12817 19156
rect 11940 19116 11946 19128
rect 12805 19125 12817 19128
rect 12851 19156 12863 19159
rect 12986 19156 12992 19168
rect 12851 19128 12992 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 13078 19116 13084 19168
rect 13136 19156 13142 19168
rect 15473 19159 15531 19165
rect 15473 19156 15485 19159
rect 13136 19128 15485 19156
rect 13136 19116 13142 19128
rect 15473 19125 15485 19128
rect 15519 19156 15531 19159
rect 15654 19156 15660 19168
rect 15519 19128 15660 19156
rect 15519 19125 15531 19128
rect 15473 19119 15531 19125
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 17034 19156 17040 19168
rect 16995 19128 17040 19156
rect 17034 19116 17040 19128
rect 17092 19156 17098 19168
rect 17862 19156 17868 19168
rect 17092 19128 17868 19156
rect 17092 19116 17098 19128
rect 17862 19116 17868 19128
rect 17920 19156 17926 19168
rect 19536 19156 19564 19196
rect 20254 19156 20260 19168
rect 17920 19128 19564 19156
rect 20215 19128 20260 19156
rect 17920 19116 17926 19128
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 21266 19156 21272 19168
rect 21227 19128 21272 19156
rect 21266 19116 21272 19128
rect 21324 19116 21330 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 2222 18912 2228 18964
rect 2280 18952 2286 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 2280 18924 2421 18952
rect 2280 18912 2286 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 2498 18912 2504 18964
rect 2556 18952 2562 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 2556 18924 3341 18952
rect 2556 18912 2562 18924
rect 3329 18921 3341 18924
rect 3375 18952 3387 18955
rect 3375 18924 4936 18952
rect 3375 18921 3387 18924
rect 3329 18915 3387 18921
rect 4154 18816 4160 18828
rect 2746 18788 4160 18816
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 2038 18748 2044 18760
rect 1719 18720 2044 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 2038 18708 2044 18720
rect 2096 18708 2102 18760
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18748 2651 18751
rect 2746 18748 2774 18788
rect 4154 18776 4160 18788
rect 4212 18776 4218 18828
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18785 4399 18819
rect 4908 18816 4936 18924
rect 5074 18912 5080 18964
rect 5132 18952 5138 18964
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 5132 18924 5273 18952
rect 5132 18912 5138 18924
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 7190 18952 7196 18964
rect 5261 18915 5319 18921
rect 5736 18924 7196 18952
rect 5736 18816 5764 18924
rect 7190 18912 7196 18924
rect 7248 18912 7254 18964
rect 11057 18955 11115 18961
rect 11057 18952 11069 18955
rect 9508 18924 11069 18952
rect 5994 18884 6000 18896
rect 4908 18788 5764 18816
rect 5828 18856 6000 18884
rect 4341 18779 4399 18785
rect 2639 18720 2774 18748
rect 3053 18751 3111 18757
rect 2639 18717 2651 18720
rect 2593 18711 2651 18717
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3099 18720 3832 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 2148 18680 2176 18711
rect 2148 18652 2774 18680
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1728 18584 1961 18612
rect 1728 18572 1734 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 2746 18612 2774 18652
rect 3804 18621 3832 18720
rect 4356 18680 4384 18779
rect 5721 18751 5779 18757
rect 5721 18717 5733 18751
rect 5767 18748 5779 18751
rect 5828 18748 5856 18856
rect 5994 18844 6000 18856
rect 6052 18844 6058 18896
rect 6362 18844 6368 18896
rect 6420 18884 6426 18896
rect 9508 18884 9536 18924
rect 11057 18921 11069 18924
rect 11103 18952 11115 18955
rect 11882 18952 11888 18964
rect 11103 18924 11888 18952
rect 11103 18921 11115 18924
rect 11057 18915 11115 18921
rect 11882 18912 11888 18924
rect 11940 18912 11946 18964
rect 14458 18912 14464 18964
rect 14516 18952 14522 18964
rect 14553 18955 14611 18961
rect 14553 18952 14565 18955
rect 14516 18924 14565 18952
rect 14516 18912 14522 18924
rect 14553 18921 14565 18924
rect 14599 18921 14611 18955
rect 14553 18915 14611 18921
rect 14642 18912 14648 18964
rect 14700 18952 14706 18964
rect 16298 18952 16304 18964
rect 14700 18924 16304 18952
rect 14700 18912 14706 18924
rect 16298 18912 16304 18924
rect 16356 18912 16362 18964
rect 16577 18955 16635 18961
rect 16577 18921 16589 18955
rect 16623 18952 16635 18955
rect 16942 18952 16948 18964
rect 16623 18924 16948 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 17681 18955 17739 18961
rect 17681 18921 17693 18955
rect 17727 18952 17739 18955
rect 17954 18952 17960 18964
rect 17727 18924 17960 18952
rect 17727 18921 17739 18924
rect 17681 18915 17739 18921
rect 17954 18912 17960 18924
rect 18012 18952 18018 18964
rect 18138 18952 18144 18964
rect 18012 18924 18144 18952
rect 18012 18912 18018 18924
rect 18138 18912 18144 18924
rect 18196 18952 18202 18964
rect 18690 18952 18696 18964
rect 18196 18924 18696 18952
rect 18196 18912 18202 18924
rect 18690 18912 18696 18924
rect 18748 18952 18754 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18748 18924 18797 18952
rect 18748 18912 18754 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 6420 18856 9536 18884
rect 6420 18844 6426 18856
rect 5905 18819 5963 18825
rect 5905 18785 5917 18819
rect 5951 18816 5963 18819
rect 6546 18816 6552 18828
rect 5951 18788 6552 18816
rect 5951 18785 5963 18788
rect 5905 18779 5963 18785
rect 6546 18776 6552 18788
rect 6604 18776 6610 18828
rect 6822 18816 6828 18828
rect 6735 18788 6828 18816
rect 6822 18776 6828 18788
rect 6880 18816 6886 18828
rect 10042 18816 10048 18828
rect 6880 18788 10048 18816
rect 6880 18776 6886 18788
rect 10042 18776 10048 18788
rect 10100 18776 10106 18828
rect 11900 18825 11928 18912
rect 12066 18844 12072 18896
rect 12124 18884 12130 18896
rect 18874 18884 18880 18896
rect 12124 18856 18880 18884
rect 12124 18844 12130 18856
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 19981 18887 20039 18893
rect 19981 18853 19993 18887
rect 20027 18884 20039 18887
rect 20806 18884 20812 18896
rect 20027 18856 20812 18884
rect 20027 18853 20039 18856
rect 19981 18847 20039 18853
rect 20806 18844 20812 18856
rect 20864 18844 20870 18896
rect 11885 18819 11943 18825
rect 11885 18785 11897 18819
rect 11931 18785 11943 18819
rect 11885 18779 11943 18785
rect 11974 18776 11980 18828
rect 12032 18816 12038 18828
rect 12621 18819 12679 18825
rect 12032 18788 12077 18816
rect 12032 18776 12038 18788
rect 12621 18785 12633 18819
rect 12667 18785 12679 18819
rect 12621 18779 12679 18785
rect 5767 18720 5856 18748
rect 5767 18717 5779 18720
rect 5721 18711 5779 18717
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8941 18751 8999 18757
rect 8941 18748 8953 18751
rect 8168 18720 8953 18748
rect 8168 18708 8174 18720
rect 8941 18717 8953 18720
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 11793 18751 11851 18757
rect 11793 18717 11805 18751
rect 11839 18748 11851 18751
rect 12342 18748 12348 18760
rect 11839 18720 12348 18748
rect 11839 18717 11851 18720
rect 11793 18711 11851 18717
rect 12342 18708 12348 18720
rect 12400 18708 12406 18760
rect 12636 18748 12664 18779
rect 14366 18776 14372 18828
rect 14424 18816 14430 18828
rect 15105 18819 15163 18825
rect 15105 18816 15117 18819
rect 14424 18788 15117 18816
rect 14424 18776 14430 18788
rect 15105 18785 15117 18788
rect 15151 18785 15163 18819
rect 16114 18816 16120 18828
rect 16075 18788 16120 18816
rect 15105 18779 15163 18785
rect 16114 18776 16120 18788
rect 16172 18776 16178 18828
rect 17218 18816 17224 18828
rect 16224 18788 17080 18816
rect 17131 18788 17224 18816
rect 16224 18748 16252 18788
rect 12636 18720 16252 18748
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 16942 18748 16948 18760
rect 16356 18720 16948 18748
rect 16356 18708 16362 18720
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17052 18748 17080 18788
rect 17218 18776 17224 18788
rect 17276 18816 17282 18828
rect 18417 18819 18475 18825
rect 18417 18816 18429 18819
rect 17276 18788 18429 18816
rect 17276 18776 17282 18788
rect 18417 18785 18429 18788
rect 18463 18785 18475 18819
rect 18417 18779 18475 18785
rect 18690 18776 18696 18828
rect 18748 18816 18754 18828
rect 19337 18819 19395 18825
rect 19337 18816 19349 18819
rect 18748 18788 19349 18816
rect 18748 18776 18754 18788
rect 19337 18785 19349 18788
rect 19383 18785 19395 18819
rect 19337 18779 19395 18785
rect 20254 18776 20260 18828
rect 20312 18816 20318 18828
rect 20312 18788 21128 18816
rect 20312 18776 20318 18788
rect 18708 18748 18736 18776
rect 17052 18720 18736 18748
rect 19978 18708 19984 18760
rect 20036 18748 20042 18760
rect 21100 18757 21128 18788
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20036 18720 20637 18748
rect 20036 18708 20042 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 5629 18683 5687 18689
rect 4356 18652 4936 18680
rect 2869 18615 2927 18621
rect 2869 18612 2881 18615
rect 2746 18584 2881 18612
rect 1949 18575 2007 18581
rect 2869 18581 2881 18584
rect 2915 18581 2927 18615
rect 2869 18575 2927 18581
rect 3789 18615 3847 18621
rect 3789 18581 3801 18615
rect 3835 18581 3847 18615
rect 3789 18575 3847 18581
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3936 18584 4169 18612
rect 3936 18572 3942 18584
rect 4157 18581 4169 18584
rect 4203 18581 4215 18615
rect 4157 18575 4215 18581
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4522 18612 4528 18624
rect 4295 18584 4528 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4522 18572 4528 18584
rect 4580 18572 4586 18624
rect 4798 18612 4804 18624
rect 4759 18584 4804 18612
rect 4798 18572 4804 18584
rect 4856 18572 4862 18624
rect 4908 18612 4936 18652
rect 5629 18649 5641 18683
rect 5675 18680 5687 18683
rect 6273 18683 6331 18689
rect 6273 18680 6285 18683
rect 5675 18652 6285 18680
rect 5675 18649 5687 18652
rect 5629 18643 5687 18649
rect 6273 18649 6285 18652
rect 6319 18649 6331 18683
rect 6273 18643 6331 18649
rect 6380 18652 7788 18680
rect 6380 18612 6408 18652
rect 4908 18584 6408 18612
rect 7193 18615 7251 18621
rect 7193 18581 7205 18615
rect 7239 18612 7251 18615
rect 7650 18612 7656 18624
rect 7239 18584 7656 18612
rect 7239 18581 7251 18584
rect 7193 18575 7251 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 7760 18612 7788 18652
rect 8294 18640 8300 18692
rect 8352 18680 8358 18692
rect 14642 18680 14648 18692
rect 8352 18652 14648 18680
rect 8352 18640 8358 18652
rect 14642 18640 14648 18652
rect 14700 18640 14706 18692
rect 14921 18683 14979 18689
rect 14921 18649 14933 18683
rect 14967 18680 14979 18683
rect 15746 18680 15752 18692
rect 14967 18652 15752 18680
rect 14967 18649 14979 18652
rect 14921 18643 14979 18649
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 16206 18640 16212 18692
rect 16264 18680 16270 18692
rect 17037 18683 17095 18689
rect 17037 18680 17049 18683
rect 16264 18652 17049 18680
rect 16264 18640 16270 18652
rect 17037 18649 17049 18652
rect 17083 18649 17095 18683
rect 17037 18643 17095 18649
rect 17218 18640 17224 18692
rect 17276 18680 17282 18692
rect 19426 18680 19432 18692
rect 17276 18652 19432 18680
rect 17276 18640 17282 18652
rect 19426 18640 19432 18652
rect 19484 18640 19490 18692
rect 19521 18683 19579 18689
rect 19521 18649 19533 18683
rect 19567 18680 19579 18683
rect 19567 18652 20668 18680
rect 19567 18649 19579 18652
rect 19521 18643 19579 18649
rect 20640 18624 20668 18652
rect 9214 18612 9220 18624
rect 7760 18584 9220 18612
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 9493 18615 9551 18621
rect 9493 18581 9505 18615
rect 9539 18612 9551 18615
rect 9766 18612 9772 18624
rect 9539 18584 9772 18612
rect 9539 18581 9551 18584
rect 9493 18575 9551 18581
rect 9766 18572 9772 18584
rect 9824 18572 9830 18624
rect 11425 18615 11483 18621
rect 11425 18581 11437 18615
rect 11471 18612 11483 18615
rect 11698 18612 11704 18624
rect 11471 18584 11704 18612
rect 11471 18581 11483 18584
rect 11425 18575 11483 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12710 18612 12716 18624
rect 12671 18584 12716 18612
rect 12710 18572 12716 18584
rect 12768 18572 12774 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13170 18612 13176 18624
rect 12860 18584 12905 18612
rect 13131 18584 13176 18612
rect 12860 18572 12866 18584
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 15068 18584 15113 18612
rect 15068 18572 15074 18584
rect 15194 18572 15200 18624
rect 15252 18612 15258 18624
rect 15565 18615 15623 18621
rect 15565 18612 15577 18615
rect 15252 18584 15577 18612
rect 15252 18572 15258 18584
rect 15565 18581 15577 18584
rect 15611 18581 15623 18615
rect 15565 18575 15623 18581
rect 15654 18572 15660 18624
rect 15712 18612 15718 18624
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 15712 18584 15945 18612
rect 15712 18572 15718 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 15933 18575 15991 18581
rect 16022 18572 16028 18624
rect 16080 18612 16086 18624
rect 16942 18612 16948 18624
rect 16080 18584 16125 18612
rect 16903 18584 16948 18612
rect 16080 18572 16086 18584
rect 16942 18572 16948 18584
rect 17000 18572 17006 18624
rect 17954 18612 17960 18624
rect 17915 18584 17960 18612
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 19610 18572 19616 18624
rect 19668 18612 19674 18624
rect 20254 18612 20260 18624
rect 19668 18584 19713 18612
rect 20215 18584 20260 18612
rect 19668 18572 19674 18584
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 20622 18572 20628 18624
rect 20680 18572 20686 18624
rect 20809 18615 20867 18621
rect 20809 18581 20821 18615
rect 20855 18612 20867 18615
rect 21082 18612 21088 18624
rect 20855 18584 21088 18612
rect 20855 18581 20867 18584
rect 20809 18575 20867 18581
rect 21082 18572 21088 18584
rect 21140 18572 21146 18624
rect 21269 18615 21327 18621
rect 21269 18581 21281 18615
rect 21315 18612 21327 18615
rect 21358 18612 21364 18624
rect 21315 18584 21364 18612
rect 21315 18581 21327 18584
rect 21269 18575 21327 18581
rect 21358 18572 21364 18584
rect 21416 18572 21422 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 1104 18448 22056 18470
rect 1946 18408 1952 18420
rect 1907 18380 1952 18408
rect 1946 18368 1952 18380
rect 2004 18368 2010 18420
rect 3605 18411 3663 18417
rect 3605 18377 3617 18411
rect 3651 18408 3663 18411
rect 4249 18411 4307 18417
rect 4249 18408 4261 18411
rect 3651 18380 4261 18408
rect 3651 18377 3663 18380
rect 3605 18371 3663 18377
rect 4249 18377 4261 18380
rect 4295 18377 4307 18411
rect 5258 18408 5264 18420
rect 5219 18380 5264 18408
rect 4249 18371 4307 18377
rect 5258 18368 5264 18380
rect 5316 18368 5322 18420
rect 5442 18368 5448 18420
rect 5500 18408 5506 18420
rect 7561 18411 7619 18417
rect 7561 18408 7573 18411
rect 5500 18380 7573 18408
rect 5500 18368 5506 18380
rect 7561 18377 7573 18380
rect 7607 18377 7619 18411
rect 7561 18371 7619 18377
rect 7929 18411 7987 18417
rect 7929 18377 7941 18411
rect 7975 18408 7987 18411
rect 8018 18408 8024 18420
rect 7975 18380 8024 18408
rect 7975 18377 7987 18380
rect 7929 18371 7987 18377
rect 1026 18300 1032 18352
rect 1084 18340 1090 18352
rect 4798 18340 4804 18352
rect 1084 18312 4804 18340
rect 1084 18300 1090 18312
rect 4798 18300 4804 18312
rect 4856 18300 4862 18352
rect 5629 18343 5687 18349
rect 5629 18309 5641 18343
rect 5675 18340 5687 18343
rect 5675 18312 7144 18340
rect 5675 18309 5687 18312
rect 5629 18303 5687 18309
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 2133 18275 2191 18281
rect 2133 18241 2145 18275
rect 2179 18272 2191 18275
rect 2498 18272 2504 18284
rect 2179 18244 2504 18272
rect 2179 18241 2191 18244
rect 2133 18235 2191 18241
rect 2498 18232 2504 18244
rect 2556 18232 2562 18284
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 3050 18272 3056 18284
rect 2639 18244 3056 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 3234 18272 3240 18284
rect 3195 18244 3240 18272
rect 3234 18232 3240 18244
rect 3292 18232 3298 18284
rect 4062 18232 4068 18284
rect 4120 18272 4126 18284
rect 5644 18272 5672 18303
rect 4120 18244 5672 18272
rect 5721 18275 5779 18281
rect 4120 18232 4126 18244
rect 5721 18241 5733 18275
rect 5767 18272 5779 18275
rect 6822 18272 6828 18284
rect 5767 18244 6828 18272
rect 5767 18241 5779 18244
rect 5721 18235 5779 18241
rect 2866 18164 2872 18216
rect 2924 18204 2930 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2924 18176 2973 18204
rect 2924 18164 2930 18176
rect 2961 18173 2973 18176
rect 3007 18173 3019 18207
rect 2961 18167 3019 18173
rect 3145 18207 3203 18213
rect 3145 18173 3157 18207
rect 3191 18173 3203 18207
rect 3970 18204 3976 18216
rect 3931 18176 3976 18204
rect 3145 18167 3203 18173
rect 1578 18096 1584 18148
rect 1636 18136 1642 18148
rect 3160 18136 3188 18167
rect 3970 18164 3976 18176
rect 4028 18164 4034 18216
rect 4154 18204 4160 18216
rect 4115 18176 4160 18204
rect 4154 18164 4160 18176
rect 4212 18164 4218 18216
rect 5736 18204 5764 18235
rect 6822 18232 6828 18244
rect 6880 18232 6886 18284
rect 4264 18176 5764 18204
rect 5813 18207 5871 18213
rect 3418 18136 3424 18148
rect 1636 18108 2544 18136
rect 3160 18108 3424 18136
rect 1636 18096 1642 18108
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2130 18028 2136 18080
rect 2188 18068 2194 18080
rect 2409 18071 2467 18077
rect 2409 18068 2421 18071
rect 2188 18040 2421 18068
rect 2188 18028 2194 18040
rect 2409 18037 2421 18040
rect 2455 18037 2467 18071
rect 2516 18068 2544 18108
rect 3418 18096 3424 18108
rect 3476 18096 3482 18148
rect 4062 18096 4068 18148
rect 4120 18136 4126 18148
rect 4264 18136 4292 18176
rect 5813 18173 5825 18207
rect 5859 18173 5871 18207
rect 7006 18204 7012 18216
rect 6967 18176 7012 18204
rect 5813 18167 5871 18173
rect 4985 18139 5043 18145
rect 4120 18108 4292 18136
rect 4448 18108 4936 18136
rect 4120 18096 4126 18108
rect 4448 18068 4476 18108
rect 4614 18068 4620 18080
rect 2516 18040 4476 18068
rect 4575 18040 4620 18068
rect 2409 18031 2467 18037
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 4908 18068 4936 18108
rect 4985 18105 4997 18139
rect 5031 18136 5043 18139
rect 5828 18136 5856 18167
rect 7006 18164 7012 18176
rect 7064 18164 7070 18216
rect 7116 18204 7144 18312
rect 7576 18272 7604 18371
rect 8018 18368 8024 18380
rect 8076 18368 8082 18420
rect 8110 18368 8116 18420
rect 8168 18408 8174 18420
rect 9306 18408 9312 18420
rect 8168 18380 9312 18408
rect 8168 18368 8174 18380
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 10137 18411 10195 18417
rect 10137 18377 10149 18411
rect 10183 18408 10195 18411
rect 12066 18408 12072 18420
rect 10183 18380 12072 18408
rect 10183 18377 10195 18380
rect 10137 18371 10195 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 12345 18411 12403 18417
rect 12345 18377 12357 18411
rect 12391 18408 12403 18411
rect 12802 18408 12808 18420
rect 12391 18380 12808 18408
rect 12391 18377 12403 18380
rect 12345 18371 12403 18377
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 14093 18411 14151 18417
rect 14093 18408 14105 18411
rect 13688 18380 14105 18408
rect 13688 18368 13694 18380
rect 14093 18377 14105 18380
rect 14139 18377 14151 18411
rect 15194 18408 15200 18420
rect 15155 18380 15200 18408
rect 14093 18371 14151 18377
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15654 18408 15660 18420
rect 15344 18380 15389 18408
rect 15615 18380 15660 18408
rect 15344 18368 15350 18380
rect 15654 18368 15660 18380
rect 15712 18368 15718 18420
rect 16850 18368 16856 18420
rect 16908 18408 16914 18420
rect 17678 18408 17684 18420
rect 16908 18380 17684 18408
rect 16908 18368 16914 18380
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 17862 18368 17868 18420
rect 17920 18408 17926 18420
rect 19153 18411 19211 18417
rect 19153 18408 19165 18411
rect 17920 18380 19165 18408
rect 17920 18368 17926 18380
rect 19153 18377 19165 18380
rect 19199 18377 19211 18411
rect 19153 18371 19211 18377
rect 7650 18300 7656 18352
rect 7708 18340 7714 18352
rect 7708 18312 12756 18340
rect 7708 18300 7714 18312
rect 8294 18272 8300 18284
rect 7576 18244 8300 18272
rect 8294 18232 8300 18244
rect 8352 18232 8358 18284
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8662 18272 8668 18284
rect 8435 18244 8668 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9232 18244 9904 18272
rect 7650 18204 7656 18216
rect 7116 18176 7656 18204
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 8478 18204 8484 18216
rect 8439 18176 8484 18204
rect 8478 18164 8484 18176
rect 8536 18204 8542 18216
rect 9232 18204 9260 18244
rect 9398 18204 9404 18216
rect 8536 18176 9260 18204
rect 9359 18176 9404 18204
rect 8536 18164 8542 18176
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9493 18207 9551 18213
rect 9493 18173 9505 18207
rect 9539 18173 9551 18207
rect 9876 18204 9904 18244
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 11149 18275 11207 18281
rect 10008 18244 10053 18272
rect 10008 18232 10014 18244
rect 11149 18241 11161 18275
rect 11195 18272 11207 18275
rect 11977 18275 12035 18281
rect 11195 18244 11928 18272
rect 11195 18241 11207 18244
rect 11149 18235 11207 18241
rect 11900 18216 11928 18244
rect 11977 18241 11989 18275
rect 12023 18272 12035 18275
rect 12621 18275 12679 18281
rect 12621 18272 12633 18275
rect 12023 18244 12633 18272
rect 12023 18241 12035 18244
rect 11977 18235 12035 18241
rect 12621 18241 12633 18244
rect 12667 18241 12679 18275
rect 12621 18235 12679 18241
rect 10962 18204 10968 18216
rect 9876 18176 10968 18204
rect 9493 18167 9551 18173
rect 5994 18136 6000 18148
rect 5031 18108 6000 18136
rect 5031 18105 5043 18108
rect 4985 18099 5043 18105
rect 5994 18096 6000 18108
rect 6052 18096 6058 18148
rect 8110 18136 8116 18148
rect 6196 18108 8116 18136
rect 6196 18068 6224 18108
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 8202 18096 8208 18148
rect 8260 18136 8266 18148
rect 9508 18136 9536 18167
rect 10962 18164 10968 18176
rect 11020 18164 11026 18216
rect 11793 18207 11851 18213
rect 11793 18173 11805 18207
rect 11839 18173 11851 18207
rect 11793 18167 11851 18173
rect 8260 18108 9536 18136
rect 8260 18096 8266 18108
rect 10778 18096 10784 18148
rect 10836 18136 10842 18148
rect 11808 18136 11836 18167
rect 11882 18164 11888 18216
rect 11940 18204 11946 18216
rect 12526 18204 12532 18216
rect 11940 18176 12532 18204
rect 11940 18164 11946 18176
rect 12526 18164 12532 18176
rect 12584 18164 12590 18216
rect 12728 18204 12756 18312
rect 13170 18300 13176 18352
rect 13228 18340 13234 18352
rect 17218 18340 17224 18352
rect 13228 18312 17224 18340
rect 13228 18300 13234 18312
rect 17218 18300 17224 18312
rect 17276 18300 17282 18352
rect 17402 18300 17408 18352
rect 17460 18300 17466 18352
rect 18598 18340 18604 18352
rect 17972 18312 18604 18340
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13630 18272 13636 18284
rect 13044 18244 13636 18272
rect 13044 18232 13050 18244
rect 13630 18232 13636 18244
rect 13688 18232 13694 18284
rect 16850 18272 16856 18284
rect 13740 18244 16856 18272
rect 13740 18204 13768 18244
rect 16850 18232 16856 18244
rect 16908 18232 16914 18284
rect 17420 18272 17448 18300
rect 16960 18244 17448 18272
rect 12728 18176 13768 18204
rect 15105 18207 15163 18213
rect 15105 18173 15117 18207
rect 15151 18173 15163 18207
rect 16960 18204 16988 18244
rect 15105 18167 15163 18173
rect 15764 18176 16988 18204
rect 13817 18139 13875 18145
rect 10836 18108 13216 18136
rect 10836 18096 10842 18108
rect 4908 18040 6224 18068
rect 6270 18028 6276 18080
rect 6328 18068 6334 18080
rect 6457 18071 6515 18077
rect 6457 18068 6469 18071
rect 6328 18040 6469 18068
rect 6328 18028 6334 18040
rect 6457 18037 6469 18040
rect 6503 18068 6515 18071
rect 6546 18068 6552 18080
rect 6503 18040 6552 18068
rect 6503 18037 6515 18040
rect 6457 18031 6515 18037
rect 6546 18028 6552 18040
rect 6604 18028 6610 18080
rect 8294 18028 8300 18080
rect 8352 18068 8358 18080
rect 8941 18071 8999 18077
rect 8941 18068 8953 18071
rect 8352 18040 8953 18068
rect 8352 18028 8358 18040
rect 8941 18037 8953 18040
rect 8987 18037 8999 18071
rect 8941 18031 8999 18037
rect 9306 18028 9312 18080
rect 9364 18068 9370 18080
rect 12986 18068 12992 18080
rect 9364 18040 12992 18068
rect 9364 18028 9370 18040
rect 12986 18028 12992 18040
rect 13044 18028 13050 18080
rect 13188 18077 13216 18108
rect 13817 18105 13829 18139
rect 13863 18136 13875 18139
rect 15120 18136 15148 18167
rect 15764 18136 15792 18176
rect 17034 18164 17040 18216
rect 17092 18204 17098 18216
rect 17405 18207 17463 18213
rect 17405 18204 17417 18207
rect 17092 18176 17417 18204
rect 17092 18164 17098 18176
rect 17405 18173 17417 18176
rect 17451 18204 17463 18207
rect 17586 18204 17592 18216
rect 17451 18176 17592 18204
rect 17451 18173 17463 18176
rect 17405 18167 17463 18173
rect 17586 18164 17592 18176
rect 17644 18164 17650 18216
rect 17972 18213 18000 18312
rect 18598 18300 18604 18312
rect 18656 18300 18662 18352
rect 18138 18272 18144 18284
rect 18099 18244 18144 18272
rect 18138 18232 18144 18244
rect 18196 18232 18202 18284
rect 20073 18275 20131 18281
rect 20073 18272 20085 18275
rect 18524 18244 20085 18272
rect 17957 18207 18015 18213
rect 17957 18173 17969 18207
rect 18003 18173 18015 18207
rect 17957 18167 18015 18173
rect 18046 18164 18052 18216
rect 18104 18204 18110 18216
rect 18524 18204 18552 18244
rect 20073 18241 20085 18244
rect 20119 18272 20131 18275
rect 20254 18272 20260 18284
rect 20119 18244 20260 18272
rect 20119 18241 20131 18244
rect 20073 18235 20131 18241
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 20438 18232 20444 18284
rect 20496 18272 20502 18284
rect 20533 18275 20591 18281
rect 20533 18272 20545 18275
rect 20496 18244 20545 18272
rect 20496 18232 20502 18244
rect 20533 18241 20545 18244
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 18104 18176 18552 18204
rect 18104 18164 18110 18176
rect 19058 18164 19064 18216
rect 19116 18204 19122 18216
rect 19245 18207 19303 18213
rect 19245 18204 19257 18207
rect 19116 18176 19257 18204
rect 19116 18164 19122 18176
rect 19245 18173 19257 18176
rect 19291 18173 19303 18207
rect 19245 18167 19303 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18173 19395 18207
rect 21100 18204 21128 18235
rect 19337 18167 19395 18173
rect 19444 18176 21128 18204
rect 13863 18108 15056 18136
rect 15120 18108 15792 18136
rect 15856 18108 18920 18136
rect 13863 18105 13875 18108
rect 13817 18099 13875 18105
rect 13173 18071 13231 18077
rect 13173 18037 13185 18071
rect 13219 18068 13231 18071
rect 13354 18068 13360 18080
rect 13219 18040 13360 18068
rect 13219 18037 13231 18040
rect 13173 18031 13231 18037
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 15028 18068 15056 18108
rect 15856 18068 15884 18108
rect 16206 18068 16212 18080
rect 15028 18040 15884 18068
rect 16167 18040 16212 18068
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16761 18071 16819 18077
rect 16761 18037 16773 18071
rect 16807 18068 16819 18071
rect 16942 18068 16948 18080
rect 16807 18040 16948 18068
rect 16807 18037 16819 18040
rect 16761 18031 16819 18037
rect 16942 18028 16948 18040
rect 17000 18028 17006 18080
rect 17126 18068 17132 18080
rect 17087 18040 17132 18068
rect 17126 18028 17132 18040
rect 17184 18068 17190 18080
rect 18046 18068 18052 18080
rect 17184 18040 18052 18068
rect 17184 18028 17190 18040
rect 18046 18028 18052 18040
rect 18104 18028 18110 18080
rect 18506 18068 18512 18080
rect 18467 18040 18512 18068
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 18782 18068 18788 18080
rect 18743 18040 18788 18068
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18892 18068 18920 18108
rect 18966 18096 18972 18148
rect 19024 18136 19030 18148
rect 19352 18136 19380 18167
rect 19024 18108 19380 18136
rect 19024 18096 19030 18108
rect 19444 18068 19472 18176
rect 20257 18139 20315 18145
rect 20257 18105 20269 18139
rect 20303 18136 20315 18139
rect 20990 18136 20996 18148
rect 20303 18108 20996 18136
rect 20303 18105 20315 18108
rect 20257 18099 20315 18105
rect 20990 18096 20996 18108
rect 21048 18096 21054 18148
rect 20714 18068 20720 18080
rect 18892 18040 19472 18068
rect 20675 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21266 18068 21272 18080
rect 21227 18040 21272 18068
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 2501 17867 2559 17873
rect 2501 17864 2513 17867
rect 2096 17836 2513 17864
rect 2096 17824 2102 17836
rect 2501 17833 2513 17836
rect 2547 17833 2559 17867
rect 2501 17827 2559 17833
rect 3050 17824 3056 17876
rect 3108 17864 3114 17876
rect 3421 17867 3479 17873
rect 3421 17864 3433 17867
rect 3108 17836 3433 17864
rect 3108 17824 3114 17836
rect 3421 17833 3433 17836
rect 3467 17864 3479 17867
rect 4062 17864 4068 17876
rect 3467 17836 4068 17864
rect 3467 17833 3479 17836
rect 3421 17827 3479 17833
rect 4062 17824 4068 17836
rect 4120 17824 4126 17876
rect 5166 17824 5172 17876
rect 5224 17864 5230 17876
rect 5629 17867 5687 17873
rect 5629 17864 5641 17867
rect 5224 17836 5641 17864
rect 5224 17824 5230 17836
rect 5629 17833 5641 17836
rect 5675 17833 5687 17867
rect 5629 17827 5687 17833
rect 6270 17824 6276 17876
rect 6328 17864 6334 17876
rect 6328 17836 7604 17864
rect 6328 17824 6334 17836
rect 7466 17796 7472 17808
rect 2976 17768 7328 17796
rect 7427 17768 7472 17796
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 2130 17660 2136 17672
rect 1719 17632 2136 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2222 17620 2228 17672
rect 2280 17660 2286 17672
rect 2976 17669 3004 17768
rect 3234 17688 3240 17740
rect 3292 17728 3298 17740
rect 3789 17731 3847 17737
rect 3789 17728 3801 17731
rect 3292 17700 3801 17728
rect 3292 17688 3298 17700
rect 3789 17697 3801 17700
rect 3835 17697 3847 17731
rect 3789 17691 3847 17697
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 4709 17731 4767 17737
rect 4709 17728 4721 17731
rect 4028 17700 4721 17728
rect 4028 17688 4034 17700
rect 4709 17697 4721 17700
rect 4755 17728 4767 17731
rect 5442 17728 5448 17740
rect 4755 17700 5448 17728
rect 4755 17697 4767 17700
rect 4709 17691 4767 17697
rect 5442 17688 5448 17700
rect 5500 17688 5506 17740
rect 6270 17728 6276 17740
rect 6231 17700 6276 17728
rect 6270 17688 6276 17700
rect 6328 17688 6334 17740
rect 6822 17688 6828 17740
rect 6880 17728 6886 17740
rect 6917 17731 6975 17737
rect 6917 17728 6929 17731
rect 6880 17700 6929 17728
rect 6880 17688 6886 17700
rect 6917 17697 6929 17700
rect 6963 17697 6975 17731
rect 7300 17728 7328 17768
rect 7466 17756 7472 17768
rect 7524 17756 7530 17808
rect 7576 17796 7604 17836
rect 9398 17824 9404 17876
rect 9456 17864 9462 17876
rect 9585 17867 9643 17873
rect 9585 17864 9597 17867
rect 9456 17836 9597 17864
rect 9456 17824 9462 17836
rect 9585 17833 9597 17836
rect 9631 17833 9643 17867
rect 9585 17827 9643 17833
rect 9674 17824 9680 17876
rect 9732 17864 9738 17876
rect 13078 17864 13084 17876
rect 9732 17836 13084 17864
rect 9732 17824 9738 17836
rect 13078 17824 13084 17836
rect 13136 17824 13142 17876
rect 16117 17867 16175 17873
rect 16117 17833 16129 17867
rect 16163 17864 16175 17867
rect 17862 17864 17868 17876
rect 16163 17836 17868 17864
rect 16163 17833 16175 17836
rect 16117 17827 16175 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 19116 17836 19257 17864
rect 19116 17824 19122 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 20070 17824 20076 17876
rect 20128 17864 20134 17876
rect 21269 17867 21327 17873
rect 21269 17864 21281 17867
rect 20128 17836 21281 17864
rect 20128 17824 20134 17836
rect 21269 17833 21281 17836
rect 21315 17833 21327 17867
rect 21269 17827 21327 17833
rect 10870 17796 10876 17808
rect 7576 17768 10876 17796
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 15746 17756 15752 17808
rect 15804 17796 15810 17808
rect 17589 17799 17647 17805
rect 17589 17796 17601 17799
rect 15804 17768 17601 17796
rect 15804 17756 15810 17768
rect 17589 17765 17601 17768
rect 17635 17765 17647 17799
rect 20898 17796 20904 17808
rect 17589 17759 17647 17765
rect 17788 17768 20904 17796
rect 7650 17728 7656 17740
rect 7300 17700 7656 17728
rect 6917 17691 6975 17697
rect 2685 17663 2743 17669
rect 2280 17632 2325 17660
rect 2280 17620 2286 17632
rect 2685 17629 2697 17663
rect 2731 17660 2743 17663
rect 2961 17663 3019 17669
rect 2961 17660 2973 17663
rect 2731 17632 2973 17660
rect 2731 17629 2743 17632
rect 2685 17623 2743 17629
rect 2961 17629 2973 17632
rect 3007 17629 3019 17663
rect 2961 17623 3019 17629
rect 4798 17620 4804 17672
rect 4856 17660 4862 17672
rect 6932 17660 6960 17691
rect 7650 17688 7656 17700
rect 7708 17688 7714 17740
rect 7929 17731 7987 17737
rect 7929 17697 7941 17731
rect 7975 17728 7987 17731
rect 8202 17728 8208 17740
rect 7975 17700 8208 17728
rect 7975 17697 7987 17700
rect 7929 17691 7987 17697
rect 8202 17688 8208 17700
rect 8260 17688 8266 17740
rect 10226 17728 10232 17740
rect 10187 17700 10232 17728
rect 10226 17688 10232 17700
rect 10284 17688 10290 17740
rect 12161 17731 12219 17737
rect 12161 17697 12173 17731
rect 12207 17728 12219 17731
rect 15562 17728 15568 17740
rect 12207 17700 13124 17728
rect 15523 17700 15568 17728
rect 12207 17697 12219 17700
rect 12161 17691 12219 17697
rect 7374 17660 7380 17672
rect 4856 17632 6868 17660
rect 6932 17632 7380 17660
rect 4856 17620 4862 17632
rect 4893 17595 4951 17601
rect 4893 17561 4905 17595
rect 4939 17592 4951 17595
rect 6730 17592 6736 17604
rect 4939 17564 6736 17592
rect 4939 17561 4951 17564
rect 4893 17555 4951 17561
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 6840 17592 6868 17632
rect 7374 17620 7380 17632
rect 7432 17620 7438 17672
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 9950 17660 9956 17672
rect 7800 17632 9956 17660
rect 7800 17620 7806 17632
rect 9950 17620 9956 17632
rect 10008 17660 10014 17672
rect 11977 17663 12035 17669
rect 11977 17660 11989 17663
rect 10008 17632 11989 17660
rect 10008 17620 10014 17632
rect 11977 17629 11989 17632
rect 12023 17629 12035 17663
rect 11977 17623 12035 17629
rect 8113 17595 8171 17601
rect 6840 17564 8064 17592
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2038 17524 2044 17536
rect 1999 17496 2044 17524
rect 2038 17484 2044 17496
rect 2096 17484 2102 17536
rect 4246 17524 4252 17536
rect 4207 17496 4252 17524
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5040 17496 5085 17524
rect 5040 17484 5046 17496
rect 5166 17484 5172 17536
rect 5224 17524 5230 17536
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 5224 17496 5365 17524
rect 5224 17484 5230 17496
rect 5353 17493 5365 17496
rect 5399 17493 5411 17527
rect 5353 17487 5411 17493
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5960 17496 6009 17524
rect 5960 17484 5966 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6089 17527 6147 17533
rect 6089 17493 6101 17527
rect 6135 17524 6147 17527
rect 6546 17524 6552 17536
rect 6135 17496 6552 17524
rect 6135 17493 6147 17496
rect 6089 17487 6147 17493
rect 6546 17484 6552 17496
rect 6604 17484 6610 17536
rect 6914 17484 6920 17536
rect 6972 17524 6978 17536
rect 7009 17527 7067 17533
rect 7009 17524 7021 17527
rect 6972 17496 7021 17524
rect 6972 17484 6978 17496
rect 7009 17493 7021 17496
rect 7055 17493 7067 17527
rect 7009 17487 7067 17493
rect 7098 17484 7104 17536
rect 7156 17524 7162 17536
rect 8036 17533 8064 17564
rect 8113 17561 8125 17595
rect 8159 17592 8171 17595
rect 8941 17595 8999 17601
rect 8941 17592 8953 17595
rect 8159 17564 8953 17592
rect 8159 17561 8171 17564
rect 8113 17555 8171 17561
rect 8941 17561 8953 17564
rect 8987 17561 8999 17595
rect 8941 17555 8999 17561
rect 9030 17552 9036 17604
rect 9088 17592 9094 17604
rect 11885 17595 11943 17601
rect 9088 17564 11652 17592
rect 9088 17552 9094 17564
rect 8021 17527 8079 17533
rect 7156 17496 7201 17524
rect 7156 17484 7162 17496
rect 8021 17493 8033 17527
rect 8067 17493 8079 17527
rect 8478 17524 8484 17536
rect 8439 17496 8484 17524
rect 8021 17487 8079 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 9766 17484 9772 17536
rect 9824 17524 9830 17536
rect 9953 17527 10011 17533
rect 9953 17524 9965 17527
rect 9824 17496 9965 17524
rect 9824 17484 9830 17496
rect 9953 17493 9965 17496
rect 9999 17493 10011 17527
rect 9953 17487 10011 17493
rect 10042 17484 10048 17536
rect 10100 17524 10106 17536
rect 10686 17524 10692 17536
rect 10100 17496 10692 17524
rect 10100 17484 10106 17496
rect 10686 17484 10692 17496
rect 10744 17484 10750 17536
rect 11146 17524 11152 17536
rect 11107 17496 11152 17524
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11514 17524 11520 17536
rect 11475 17496 11520 17524
rect 11514 17484 11520 17496
rect 11572 17484 11578 17536
rect 11624 17524 11652 17564
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 12529 17595 12587 17601
rect 12529 17592 12541 17595
rect 11931 17564 12541 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 12529 17561 12541 17564
rect 12575 17561 12587 17595
rect 12529 17555 12587 17561
rect 12066 17524 12072 17536
rect 11624 17496 12072 17524
rect 12066 17484 12072 17496
rect 12124 17484 12130 17536
rect 13096 17533 13124 17700
rect 15562 17688 15568 17700
rect 15620 17688 15626 17740
rect 16390 17660 16396 17672
rect 16351 17632 16396 17660
rect 16390 17620 16396 17632
rect 16448 17660 16454 17672
rect 16853 17663 16911 17669
rect 16853 17660 16865 17663
rect 16448 17632 16865 17660
rect 16448 17620 16454 17632
rect 16853 17629 16865 17632
rect 16899 17629 16911 17663
rect 17788 17660 17816 17768
rect 20898 17756 20904 17768
rect 20956 17756 20962 17808
rect 17862 17688 17868 17740
rect 17920 17728 17926 17740
rect 18141 17731 18199 17737
rect 18141 17728 18153 17731
rect 17920 17700 18153 17728
rect 17920 17688 17926 17700
rect 18141 17697 18153 17700
rect 18187 17697 18199 17731
rect 19886 17728 19892 17740
rect 19847 17700 19892 17728
rect 18141 17691 18199 17697
rect 19886 17688 19892 17700
rect 19944 17688 19950 17740
rect 20809 17731 20867 17737
rect 20809 17728 20821 17731
rect 19996 17700 20821 17728
rect 17954 17660 17960 17672
rect 16853 17623 16911 17629
rect 17236 17632 17816 17660
rect 17915 17632 17960 17660
rect 13081 17527 13139 17533
rect 13081 17493 13093 17527
rect 13127 17524 13139 17527
rect 13446 17524 13452 17536
rect 13127 17496 13452 17524
rect 13127 17493 13139 17496
rect 13081 17487 13139 17493
rect 13446 17484 13452 17496
rect 13504 17484 13510 17536
rect 15102 17524 15108 17536
rect 15063 17496 15108 17524
rect 15102 17484 15108 17496
rect 15160 17524 15166 17536
rect 15657 17527 15715 17533
rect 15657 17524 15669 17527
rect 15160 17496 15669 17524
rect 15160 17484 15166 17496
rect 15657 17493 15669 17496
rect 15703 17493 15715 17527
rect 15657 17487 15715 17493
rect 15746 17484 15752 17536
rect 15804 17524 15810 17536
rect 16577 17527 16635 17533
rect 15804 17496 15849 17524
rect 15804 17484 15810 17496
rect 16577 17493 16589 17527
rect 16623 17524 16635 17527
rect 17236 17524 17264 17632
rect 17954 17620 17960 17632
rect 18012 17620 18018 17672
rect 18046 17620 18052 17672
rect 18104 17660 18110 17672
rect 19996 17660 20024 17700
rect 20809 17697 20821 17700
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 18104 17632 20024 17660
rect 18104 17620 18110 17632
rect 20254 17620 20260 17672
rect 20312 17660 20318 17672
rect 20717 17663 20775 17669
rect 20717 17660 20729 17663
rect 20312 17632 20729 17660
rect 20312 17620 20318 17632
rect 20717 17629 20729 17632
rect 20763 17629 20775 17663
rect 20717 17623 20775 17629
rect 20898 17620 20904 17672
rect 20956 17660 20962 17672
rect 21174 17660 21180 17672
rect 20956 17632 21180 17660
rect 20956 17620 20962 17632
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 17313 17595 17371 17601
rect 17313 17561 17325 17595
rect 17359 17592 17371 17595
rect 18230 17592 18236 17604
rect 17359 17564 18236 17592
rect 17359 17561 17371 17564
rect 17313 17555 17371 17561
rect 16623 17496 17264 17524
rect 16623 17493 16635 17496
rect 16577 17487 16635 17493
rect 17586 17484 17592 17536
rect 17644 17524 17650 17536
rect 17862 17524 17868 17536
rect 17644 17496 17868 17524
rect 17644 17484 17650 17496
rect 17862 17484 17868 17496
rect 17920 17484 17926 17536
rect 18064 17533 18092 17564
rect 18230 17552 18236 17564
rect 18288 17552 18294 17604
rect 19613 17595 19671 17601
rect 19613 17561 19625 17595
rect 19659 17592 19671 17595
rect 20070 17592 20076 17604
rect 19659 17564 20076 17592
rect 19659 17561 19671 17564
rect 19613 17555 19671 17561
rect 20070 17552 20076 17564
rect 20128 17552 20134 17604
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18598 17524 18604 17536
rect 18095 17496 18129 17524
rect 18559 17496 18604 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18598 17484 18604 17496
rect 18656 17484 18662 17536
rect 19702 17524 19708 17536
rect 19663 17496 19708 17524
rect 19702 17484 19708 17496
rect 19760 17484 19766 17536
rect 20257 17527 20315 17533
rect 20257 17493 20269 17527
rect 20303 17524 20315 17527
rect 20438 17524 20444 17536
rect 20303 17496 20444 17524
rect 20303 17493 20315 17496
rect 20257 17487 20315 17493
rect 20438 17484 20444 17496
rect 20496 17484 20502 17536
rect 20622 17524 20628 17536
rect 20583 17496 20628 17524
rect 20622 17484 20628 17496
rect 20680 17484 20686 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2869 17323 2927 17329
rect 2869 17320 2881 17323
rect 2280 17292 2881 17320
rect 2280 17280 2286 17292
rect 2869 17289 2881 17292
rect 2915 17289 2927 17323
rect 2869 17283 2927 17289
rect 3142 17280 3148 17332
rect 3200 17320 3206 17332
rect 3970 17320 3976 17332
rect 3200 17292 3976 17320
rect 3200 17280 3206 17292
rect 3970 17280 3976 17292
rect 4028 17280 4034 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 4212 17292 4445 17320
rect 4212 17280 4218 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 5166 17320 5172 17332
rect 5127 17292 5172 17320
rect 4433 17283 4491 17289
rect 5166 17280 5172 17292
rect 5224 17280 5230 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7006 17320 7012 17332
rect 6963 17292 7012 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8389 17323 8447 17329
rect 8389 17289 8401 17323
rect 8435 17320 8447 17323
rect 8478 17320 8484 17332
rect 8435 17292 8484 17320
rect 8435 17289 8447 17292
rect 8389 17283 8447 17289
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8720 17292 9045 17320
rect 8720 17280 8726 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 9398 17280 9404 17332
rect 9456 17320 9462 17332
rect 9493 17323 9551 17329
rect 9493 17320 9505 17323
rect 9456 17292 9505 17320
rect 9456 17280 9462 17292
rect 9493 17289 9505 17292
rect 9539 17289 9551 17323
rect 10686 17320 10692 17332
rect 10647 17292 10692 17320
rect 9493 17283 9551 17289
rect 10686 17280 10692 17292
rect 10744 17320 10750 17332
rect 11146 17320 11152 17332
rect 10744 17292 11152 17320
rect 10744 17280 10750 17292
rect 11146 17280 11152 17292
rect 11204 17280 11210 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 15286 17320 15292 17332
rect 14783 17292 15292 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 17862 17320 17868 17332
rect 15620 17292 17868 17320
rect 15620 17280 15626 17292
rect 17862 17280 17868 17292
rect 17920 17280 17926 17332
rect 19061 17323 19119 17329
rect 19061 17289 19073 17323
rect 19107 17320 19119 17323
rect 19978 17320 19984 17332
rect 19107 17292 19984 17320
rect 19107 17289 19119 17292
rect 19061 17283 19119 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20806 17320 20812 17332
rect 20767 17292 20812 17320
rect 20806 17280 20812 17292
rect 20864 17280 20870 17332
rect 2958 17212 2964 17264
rect 3016 17252 3022 17264
rect 4065 17255 4123 17261
rect 4065 17252 4077 17255
rect 3016 17224 4077 17252
rect 3016 17212 3022 17224
rect 4065 17221 4077 17224
rect 4111 17221 4123 17255
rect 4065 17215 4123 17221
rect 4614 17212 4620 17264
rect 4672 17252 4678 17264
rect 5077 17255 5135 17261
rect 5077 17252 5089 17255
rect 4672 17224 5089 17252
rect 4672 17212 4678 17224
rect 5077 17221 5089 17224
rect 5123 17221 5135 17255
rect 5077 17215 5135 17221
rect 8754 17212 8760 17264
rect 8812 17252 8818 17264
rect 13633 17255 13691 17261
rect 13633 17252 13645 17255
rect 8812 17224 13645 17252
rect 8812 17212 8818 17224
rect 13633 17221 13645 17224
rect 13679 17252 13691 17255
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 13679 17224 14289 17252
rect 13679 17221 13691 17224
rect 13633 17215 13691 17221
rect 14277 17221 14289 17224
rect 14323 17252 14335 17255
rect 18230 17252 18236 17264
rect 14323 17224 18236 17252
rect 14323 17221 14335 17224
rect 14277 17215 14335 17221
rect 18230 17212 18236 17224
rect 18288 17212 18294 17264
rect 19610 17212 19616 17264
rect 19668 17252 19674 17264
rect 20717 17255 20775 17261
rect 20717 17252 20729 17255
rect 19668 17224 20729 17252
rect 19668 17212 19674 17224
rect 20717 17221 20729 17224
rect 20763 17221 20775 17255
rect 20717 17215 20775 17221
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17184 2007 17187
rect 2314 17184 2320 17196
rect 1995 17156 2320 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 2314 17144 2320 17156
rect 2372 17144 2378 17196
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17153 2651 17187
rect 2593 17147 2651 17153
rect 3053 17187 3111 17193
rect 3053 17153 3065 17187
rect 3099 17184 3111 17187
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 3099 17156 3433 17184
rect 3099 17153 3111 17156
rect 3053 17147 3111 17153
rect 3421 17153 3433 17156
rect 3467 17184 3479 17187
rect 7006 17184 7012 17196
rect 3467 17156 7012 17184
rect 3467 17153 3479 17156
rect 3421 17147 3479 17153
rect 2133 17051 2191 17057
rect 2133 17017 2145 17051
rect 2179 17048 2191 17051
rect 2608 17048 2636 17147
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 9122 17144 9128 17196
rect 9180 17184 9186 17196
rect 9401 17187 9459 17193
rect 9401 17184 9413 17187
rect 9180 17156 9413 17184
rect 9180 17144 9186 17156
rect 9401 17153 9413 17156
rect 9447 17184 9459 17187
rect 9674 17184 9680 17196
rect 9447 17156 9680 17184
rect 9447 17153 9459 17156
rect 9401 17147 9459 17153
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10137 17187 10195 17193
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10781 17187 10839 17193
rect 10781 17184 10793 17187
rect 10183 17156 10793 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10781 17153 10793 17156
rect 10827 17184 10839 17187
rect 11054 17184 11060 17196
rect 10827 17156 11060 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12023 17156 12633 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 14369 17187 14427 17193
rect 14369 17153 14381 17187
rect 14415 17184 14427 17187
rect 15013 17187 15071 17193
rect 15013 17184 15025 17187
rect 14415 17156 15025 17184
rect 14415 17153 14427 17156
rect 14369 17147 14427 17153
rect 15013 17153 15025 17156
rect 15059 17153 15071 17187
rect 15013 17147 15071 17153
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16942 17184 16948 17196
rect 16715 17156 16948 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16942 17144 16948 17156
rect 17000 17184 17006 17196
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 17000 17156 17141 17184
rect 17000 17144 17006 17156
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 18874 17184 18880 17196
rect 18835 17156 18880 17184
rect 17129 17147 17187 17153
rect 18874 17144 18880 17156
rect 18932 17144 18938 17196
rect 19337 17187 19395 17193
rect 19337 17153 19349 17187
rect 19383 17184 19395 17187
rect 19518 17184 19524 17196
rect 19383 17156 19524 17184
rect 19383 17153 19395 17156
rect 19337 17147 19395 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3789 17119 3847 17125
rect 3789 17116 3801 17119
rect 2924 17088 3801 17116
rect 2924 17076 2930 17088
rect 3789 17085 3801 17088
rect 3835 17116 3847 17119
rect 4062 17116 4068 17128
rect 3835 17088 4068 17116
rect 3835 17085 3847 17088
rect 3789 17079 3847 17085
rect 4062 17076 4068 17088
rect 4120 17076 4126 17128
rect 5353 17119 5411 17125
rect 5353 17085 5365 17119
rect 5399 17116 5411 17119
rect 6086 17116 6092 17128
rect 5399 17088 6092 17116
rect 5399 17085 5411 17088
rect 5353 17079 5411 17085
rect 6086 17076 6092 17088
rect 6144 17076 6150 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17085 6791 17119
rect 6733 17079 6791 17085
rect 6825 17119 6883 17125
rect 6825 17085 6837 17119
rect 6871 17116 6883 17119
rect 7098 17116 7104 17128
rect 6871 17088 7104 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 4709 17051 4767 17057
rect 4709 17048 4721 17051
rect 2179 17020 2544 17048
rect 2608 17020 4721 17048
rect 2179 17017 2191 17020
rect 2133 17011 2191 17017
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2406 16980 2412 16992
rect 2367 16952 2412 16980
rect 2406 16940 2412 16952
rect 2464 16940 2470 16992
rect 2516 16980 2544 17020
rect 4709 17017 4721 17020
rect 4755 17017 4767 17051
rect 6748 17048 6776 17079
rect 7098 17076 7104 17088
rect 7156 17116 7162 17128
rect 7742 17116 7748 17128
rect 7156 17088 7748 17116
rect 7156 17076 7162 17088
rect 7742 17076 7748 17088
rect 7800 17076 7806 17128
rect 8205 17119 8263 17125
rect 8205 17085 8217 17119
rect 8251 17116 8263 17119
rect 8294 17116 8300 17128
rect 8251 17088 8300 17116
rect 8251 17085 8263 17088
rect 8205 17079 8263 17085
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9582 17076 9588 17128
rect 9640 17116 9646 17128
rect 9640 17088 9685 17116
rect 9640 17076 9646 17088
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10505 17119 10563 17125
rect 10505 17116 10517 17119
rect 10468 17088 10517 17116
rect 10468 17076 10474 17088
rect 10505 17085 10517 17088
rect 10551 17085 10563 17119
rect 11790 17116 11796 17128
rect 11751 17088 11796 17116
rect 10505 17079 10563 17085
rect 11790 17076 11796 17088
rect 11848 17076 11854 17128
rect 11882 17076 11888 17128
rect 11940 17116 11946 17128
rect 12526 17116 12532 17128
rect 11940 17088 12532 17116
rect 11940 17076 11946 17088
rect 12526 17076 12532 17088
rect 12584 17076 12590 17128
rect 14185 17119 14243 17125
rect 14185 17085 14197 17119
rect 14231 17116 14243 17119
rect 15194 17116 15200 17128
rect 14231 17088 15200 17116
rect 14231 17085 14243 17088
rect 14185 17079 14243 17085
rect 15194 17076 15200 17088
rect 15252 17116 15258 17128
rect 16114 17116 16120 17128
rect 15252 17088 16120 17116
rect 15252 17076 15258 17088
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 19812 17116 19840 17147
rect 16868 17088 19840 17116
rect 20993 17119 21051 17125
rect 7834 17048 7840 17060
rect 6748 17020 7840 17048
rect 4709 17011 4767 17017
rect 7834 17008 7840 17020
rect 7892 17008 7898 17060
rect 8496 17020 8892 17048
rect 3050 16980 3056 16992
rect 2516 16952 3056 16980
rect 3050 16940 3056 16952
rect 3108 16940 3114 16992
rect 5810 16980 5816 16992
rect 5771 16952 5816 16980
rect 5810 16940 5816 16952
rect 5868 16940 5874 16992
rect 7282 16980 7288 16992
rect 7243 16952 7288 16980
rect 7282 16940 7288 16952
rect 7340 16940 7346 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 7653 16983 7711 16989
rect 7653 16980 7665 16983
rect 7432 16952 7665 16980
rect 7432 16940 7438 16952
rect 7653 16949 7665 16952
rect 7699 16980 7711 16983
rect 8496 16980 8524 17020
rect 7699 16952 8524 16980
rect 7699 16949 7711 16952
rect 7653 16943 7711 16949
rect 8570 16940 8576 16992
rect 8628 16980 8634 16992
rect 8757 16983 8815 16989
rect 8757 16980 8769 16983
rect 8628 16952 8769 16980
rect 8628 16940 8634 16952
rect 8757 16949 8769 16952
rect 8803 16949 8815 16983
rect 8864 16980 8892 17020
rect 8938 17008 8944 17060
rect 8996 17048 9002 17060
rect 10134 17048 10140 17060
rect 8996 17020 10140 17048
rect 8996 17008 9002 17020
rect 10134 17008 10140 17020
rect 10192 17008 10198 17060
rect 16868 17057 16896 17088
rect 20993 17085 21005 17119
rect 21039 17116 21051 17119
rect 21174 17116 21180 17128
rect 21039 17088 21180 17116
rect 21039 17085 21051 17088
rect 20993 17079 21051 17085
rect 21174 17076 21180 17088
rect 21232 17076 21238 17128
rect 16853 17051 16911 17057
rect 16853 17017 16865 17051
rect 16899 17017 16911 17051
rect 16853 17011 16911 17017
rect 19521 17051 19579 17057
rect 19521 17017 19533 17051
rect 19567 17048 19579 17051
rect 20898 17048 20904 17060
rect 19567 17020 20904 17048
rect 19567 17017 19579 17020
rect 19521 17011 19579 17017
rect 20898 17008 20904 17020
rect 20956 17008 20962 17060
rect 10778 16980 10784 16992
rect 8864 16952 10784 16980
rect 8757 16943 8815 16949
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 12345 16983 12403 16989
rect 12345 16949 12357 16983
rect 12391 16980 12403 16983
rect 12986 16980 12992 16992
rect 12391 16952 12992 16980
rect 12391 16949 12403 16952
rect 12345 16943 12403 16949
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 17494 16980 17500 16992
rect 17455 16952 17500 16980
rect 17494 16940 17500 16952
rect 17552 16940 17558 16992
rect 18598 16980 18604 16992
rect 18559 16952 18604 16980
rect 18598 16940 18604 16952
rect 18656 16940 18662 16992
rect 19981 16983 20039 16989
rect 19981 16949 19993 16983
rect 20027 16980 20039 16983
rect 20162 16980 20168 16992
rect 20027 16952 20168 16980
rect 20027 16949 20039 16952
rect 19981 16943 20039 16949
rect 20162 16940 20168 16952
rect 20220 16940 20226 16992
rect 20346 16980 20352 16992
rect 20307 16952 20352 16980
rect 20346 16940 20352 16952
rect 20404 16940 20410 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2130 16736 2136 16788
rect 2188 16776 2194 16788
rect 8478 16776 8484 16788
rect 2188 16748 8484 16776
rect 2188 16736 2194 16748
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 9950 16776 9956 16788
rect 8588 16748 9956 16776
rect 4338 16708 4344 16720
rect 3988 16680 4344 16708
rect 3988 16649 4016 16680
rect 4338 16668 4344 16680
rect 4396 16668 4402 16720
rect 4430 16668 4436 16720
rect 4488 16708 4494 16720
rect 5997 16711 6055 16717
rect 5997 16708 6009 16711
rect 4488 16680 6009 16708
rect 4488 16668 4494 16680
rect 5997 16677 6009 16680
rect 6043 16677 6055 16711
rect 5997 16671 6055 16677
rect 6086 16668 6092 16720
rect 6144 16708 6150 16720
rect 8588 16708 8616 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 11974 16776 11980 16788
rect 10060 16748 11980 16776
rect 6144 16680 8616 16708
rect 6144 16668 6150 16680
rect 8662 16668 8668 16720
rect 8720 16708 8726 16720
rect 9493 16711 9551 16717
rect 9493 16708 9505 16711
rect 8720 16680 9505 16708
rect 8720 16668 8726 16680
rect 9493 16677 9505 16680
rect 9539 16677 9551 16711
rect 9493 16671 9551 16677
rect 3973 16643 4031 16649
rect 3973 16609 3985 16643
rect 4019 16609 4031 16643
rect 3973 16603 4031 16609
rect 4065 16643 4123 16649
rect 4065 16609 4077 16643
rect 4111 16640 4123 16643
rect 5258 16640 5264 16652
rect 4111 16612 5264 16640
rect 4111 16609 4123 16612
rect 4065 16603 4123 16609
rect 5258 16600 5264 16612
rect 5316 16600 5322 16652
rect 5626 16640 5632 16652
rect 5587 16612 5632 16640
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 5718 16600 5724 16652
rect 5776 16640 5782 16652
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 5776 16612 6377 16640
rect 5776 16600 5782 16612
rect 6365 16609 6377 16612
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 7374 16600 7380 16652
rect 7432 16640 7438 16652
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 7432 16612 9137 16640
rect 7432 16600 7438 16612
rect 9125 16609 9137 16612
rect 9171 16640 9183 16643
rect 9398 16640 9404 16652
rect 9171 16612 9404 16640
rect 9171 16609 9183 16612
rect 9125 16603 9183 16609
rect 9398 16600 9404 16612
rect 9456 16600 9462 16652
rect 9508 16640 9536 16671
rect 10060 16649 10088 16748
rect 11974 16736 11980 16748
rect 12032 16776 12038 16788
rect 15562 16776 15568 16788
rect 12032 16748 15568 16776
rect 12032 16736 12038 16748
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 15746 16736 15752 16788
rect 15804 16776 15810 16788
rect 16209 16779 16267 16785
rect 16209 16776 16221 16779
rect 15804 16748 16221 16776
rect 15804 16736 15810 16748
rect 16209 16745 16221 16748
rect 16255 16745 16267 16779
rect 19518 16776 19524 16788
rect 19479 16748 19524 16776
rect 16209 16739 16267 16745
rect 19518 16736 19524 16748
rect 19576 16736 19582 16788
rect 11146 16668 11152 16720
rect 11204 16708 11210 16720
rect 17494 16708 17500 16720
rect 11204 16680 12940 16708
rect 11204 16668 11210 16680
rect 10045 16643 10103 16649
rect 9508 16612 9628 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16541 1731 16575
rect 1673 16535 1731 16541
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16572 2191 16575
rect 2406 16572 2412 16584
rect 2179 16544 2412 16572
rect 2179 16541 2191 16544
rect 2133 16535 2191 16541
rect 1688 16504 1716 16535
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2866 16572 2872 16584
rect 2827 16544 2872 16572
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3050 16532 3056 16584
rect 3108 16572 3114 16584
rect 3329 16575 3387 16581
rect 3329 16572 3341 16575
rect 3108 16544 3341 16572
rect 3108 16532 3114 16544
rect 3329 16541 3341 16544
rect 3375 16541 3387 16575
rect 3329 16535 3387 16541
rect 6638 16532 6644 16584
rect 6696 16572 6702 16584
rect 8481 16575 8539 16581
rect 8481 16572 8493 16575
rect 6696 16544 8493 16572
rect 6696 16532 6702 16544
rect 8481 16541 8493 16544
rect 8527 16572 8539 16575
rect 9030 16572 9036 16584
rect 8527 16544 9036 16572
rect 8527 16541 8539 16544
rect 8481 16535 8539 16541
rect 9030 16532 9036 16544
rect 9088 16532 9094 16584
rect 9600 16572 9628 16612
rect 10045 16609 10057 16643
rect 10091 16609 10103 16643
rect 10045 16603 10103 16609
rect 11057 16643 11115 16649
rect 11057 16609 11069 16643
rect 11103 16640 11115 16643
rect 11698 16640 11704 16652
rect 11103 16612 11704 16640
rect 11103 16609 11115 16612
rect 11057 16603 11115 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 12802 16640 12808 16652
rect 12763 16612 12808 16640
rect 12802 16600 12808 16612
rect 12860 16600 12866 16652
rect 12912 16649 12940 16680
rect 16868 16680 17500 16708
rect 12897 16643 12955 16649
rect 12897 16609 12909 16643
rect 12943 16609 12955 16643
rect 12897 16603 12955 16609
rect 15102 16600 15108 16652
rect 15160 16640 15166 16652
rect 15841 16643 15899 16649
rect 15841 16640 15853 16643
rect 15160 16612 15853 16640
rect 15160 16600 15166 16612
rect 15841 16609 15853 16612
rect 15887 16640 15899 16643
rect 16390 16640 16396 16652
rect 15887 16612 16396 16640
rect 15887 16609 15899 16612
rect 15841 16603 15899 16609
rect 16390 16600 16396 16612
rect 16448 16640 16454 16652
rect 16868 16649 16896 16680
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 17678 16668 17684 16720
rect 17736 16708 17742 16720
rect 21450 16708 21456 16720
rect 17736 16680 17908 16708
rect 17736 16668 17742 16680
rect 16853 16643 16911 16649
rect 16448 16612 16620 16640
rect 16448 16600 16454 16612
rect 10229 16575 10287 16581
rect 10229 16572 10241 16575
rect 9600 16544 10241 16572
rect 10229 16541 10241 16544
rect 10275 16541 10287 16575
rect 10229 16535 10287 16541
rect 10686 16532 10692 16584
rect 10744 16572 10750 16584
rect 12158 16572 12164 16584
rect 10744 16544 12164 16572
rect 10744 16532 10750 16544
rect 12158 16532 12164 16544
rect 12216 16532 12222 16584
rect 12986 16572 12992 16584
rect 12947 16544 12992 16572
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 16592 16572 16620 16612
rect 16853 16609 16865 16643
rect 16899 16609 16911 16643
rect 16853 16603 16911 16609
rect 16942 16600 16948 16652
rect 17000 16640 17006 16652
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 17000 16612 17785 16640
rect 17000 16600 17006 16612
rect 17773 16609 17785 16612
rect 17819 16609 17831 16643
rect 17880 16640 17908 16680
rect 19720 16680 21456 16708
rect 18877 16643 18935 16649
rect 18877 16640 18889 16643
rect 17880 16612 18889 16640
rect 17773 16603 17831 16609
rect 18877 16609 18889 16612
rect 18923 16640 18935 16643
rect 19720 16640 19748 16680
rect 21450 16668 21456 16680
rect 21508 16668 21514 16720
rect 20438 16640 20444 16652
rect 18923 16612 19748 16640
rect 20399 16612 20444 16640
rect 18923 16609 18935 16612
rect 18877 16603 18935 16609
rect 20438 16600 20444 16612
rect 20496 16600 20502 16652
rect 20530 16600 20536 16652
rect 20588 16640 20594 16652
rect 20588 16612 20633 16640
rect 20588 16600 20594 16612
rect 16669 16575 16727 16581
rect 16669 16572 16681 16575
rect 16592 16544 16681 16572
rect 16669 16541 16681 16544
rect 16715 16541 16727 16575
rect 17678 16572 17684 16584
rect 17639 16544 17684 16572
rect 16669 16535 16727 16541
rect 17678 16532 17684 16544
rect 17736 16532 17742 16584
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16572 18383 16575
rect 18782 16572 18788 16584
rect 18371 16544 18788 16572
rect 18371 16541 18383 16544
rect 18325 16535 18383 16541
rect 18782 16532 18788 16544
rect 18840 16532 18846 16584
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16572 19763 16575
rect 20346 16572 20352 16584
rect 19751 16544 20352 16572
rect 19751 16541 19763 16544
rect 19705 16535 19763 16541
rect 20346 16532 20352 16544
rect 20404 16532 20410 16584
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 21048 16544 21097 16572
rect 21048 16532 21054 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 4154 16504 4160 16516
rect 1688 16476 3188 16504
rect 4115 16476 4160 16504
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 1949 16439 2007 16445
rect 1949 16405 1961 16439
rect 1995 16436 2007 16439
rect 2038 16436 2044 16448
rect 1995 16408 2044 16436
rect 1995 16405 2007 16408
rect 1949 16399 2007 16405
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 2222 16396 2228 16448
rect 2280 16436 2286 16448
rect 3160 16445 3188 16476
rect 4154 16464 4160 16476
rect 4212 16464 4218 16516
rect 6454 16464 6460 16516
rect 6512 16504 6518 16516
rect 7377 16507 7435 16513
rect 7377 16504 7389 16507
rect 6512 16476 7389 16504
rect 6512 16464 6518 16476
rect 7377 16473 7389 16476
rect 7423 16473 7435 16507
rect 15286 16504 15292 16516
rect 7377 16467 7435 16473
rect 11624 16476 15292 16504
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 2280 16408 2697 16436
rect 2280 16396 2286 16408
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16405 3203 16439
rect 4522 16436 4528 16448
rect 4483 16408 4528 16436
rect 3145 16399 3203 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 4890 16436 4896 16448
rect 4851 16408 4896 16436
rect 4890 16396 4896 16408
rect 4948 16396 4954 16448
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5261 16439 5319 16445
rect 5261 16436 5273 16439
rect 5132 16408 5273 16436
rect 5132 16396 5138 16408
rect 5261 16405 5273 16408
rect 5307 16405 5319 16439
rect 5261 16399 5319 16405
rect 6638 16396 6644 16448
rect 6696 16436 6702 16448
rect 6733 16439 6791 16445
rect 6733 16436 6745 16439
rect 6696 16408 6745 16436
rect 6696 16396 6702 16408
rect 6733 16405 6745 16408
rect 6779 16405 6791 16439
rect 6733 16399 6791 16405
rect 7837 16439 7895 16445
rect 7837 16405 7849 16439
rect 7883 16436 7895 16439
rect 7926 16436 7932 16448
rect 7883 16408 7932 16436
rect 7883 16405 7895 16408
rect 7837 16399 7895 16405
rect 7926 16396 7932 16408
rect 7984 16396 7990 16448
rect 8110 16436 8116 16448
rect 8071 16408 8116 16436
rect 8110 16396 8116 16408
rect 8168 16396 8174 16448
rect 8662 16396 8668 16448
rect 8720 16436 8726 16448
rect 10137 16439 10195 16445
rect 10137 16436 10149 16439
rect 8720 16408 10149 16436
rect 8720 16396 8726 16408
rect 10137 16405 10149 16408
rect 10183 16436 10195 16439
rect 10410 16436 10416 16448
rect 10183 16408 10416 16436
rect 10183 16405 10195 16408
rect 10137 16399 10195 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 10597 16439 10655 16445
rect 10597 16405 10609 16439
rect 10643 16436 10655 16439
rect 11149 16439 11207 16445
rect 11149 16436 11161 16439
rect 10643 16408 11161 16436
rect 10643 16405 10655 16408
rect 10597 16399 10655 16405
rect 11149 16405 11161 16408
rect 11195 16405 11207 16439
rect 11149 16399 11207 16405
rect 11241 16439 11299 16445
rect 11241 16405 11253 16439
rect 11287 16436 11299 16439
rect 11514 16436 11520 16448
rect 11287 16408 11520 16436
rect 11287 16405 11299 16408
rect 11241 16399 11299 16405
rect 11514 16396 11520 16408
rect 11572 16396 11578 16448
rect 11624 16445 11652 16476
rect 15286 16464 15292 16476
rect 15344 16464 15350 16516
rect 16022 16464 16028 16516
rect 16080 16504 16086 16516
rect 17589 16507 17647 16513
rect 16080 16476 17264 16504
rect 16080 16464 16086 16476
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16405 11667 16439
rect 11609 16399 11667 16405
rect 11977 16439 12035 16445
rect 11977 16405 11989 16439
rect 12023 16436 12035 16439
rect 12526 16436 12532 16448
rect 12023 16408 12532 16436
rect 12023 16405 12035 16408
rect 11977 16399 12035 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13357 16439 13415 16445
rect 13357 16405 13369 16439
rect 13403 16436 13415 16439
rect 13446 16436 13452 16448
rect 13403 16408 13452 16436
rect 13403 16405 13415 16408
rect 13357 16399 13415 16405
rect 13446 16396 13452 16408
rect 13504 16396 13510 16448
rect 16390 16396 16396 16448
rect 16448 16436 16454 16448
rect 17236 16445 17264 16476
rect 17589 16473 17601 16507
rect 17635 16504 17647 16507
rect 17635 16476 20116 16504
rect 17635 16473 17647 16476
rect 17589 16467 17647 16473
rect 20088 16448 20116 16476
rect 16577 16439 16635 16445
rect 16577 16436 16589 16439
rect 16448 16408 16589 16436
rect 16448 16396 16454 16408
rect 16577 16405 16589 16408
rect 16623 16405 16635 16439
rect 16577 16399 16635 16405
rect 17221 16439 17279 16445
rect 17221 16405 17233 16439
rect 17267 16405 17279 16439
rect 17221 16399 17279 16405
rect 18509 16439 18567 16445
rect 18509 16405 18521 16439
rect 18555 16436 18567 16439
rect 18690 16436 18696 16448
rect 18555 16408 18696 16436
rect 18555 16405 18567 16408
rect 18509 16399 18567 16405
rect 18690 16396 18696 16408
rect 18748 16396 18754 16448
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 19981 16439 20039 16445
rect 19981 16436 19993 16439
rect 18932 16408 19993 16436
rect 18932 16396 18938 16408
rect 19981 16405 19993 16408
rect 20027 16405 20039 16439
rect 19981 16399 20039 16405
rect 20070 16396 20076 16448
rect 20128 16396 20134 16448
rect 20346 16436 20352 16448
rect 20307 16408 20352 16436
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1670 16192 1676 16244
rect 1728 16232 1734 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 1728 16204 2513 16232
rect 1728 16192 1734 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 2501 16195 2559 16201
rect 2866 16192 2872 16244
rect 2924 16232 2930 16244
rect 3329 16235 3387 16241
rect 3329 16232 3341 16235
rect 2924 16204 3341 16232
rect 2924 16192 2930 16204
rect 3329 16201 3341 16204
rect 3375 16232 3387 16235
rect 4706 16232 4712 16244
rect 3375 16204 4712 16232
rect 3375 16201 3387 16204
rect 3329 16195 3387 16201
rect 4706 16192 4712 16204
rect 4764 16192 4770 16244
rect 4982 16192 4988 16244
rect 5040 16232 5046 16244
rect 5077 16235 5135 16241
rect 5077 16232 5089 16235
rect 5040 16204 5089 16232
rect 5040 16192 5046 16204
rect 5077 16201 5089 16204
rect 5123 16201 5135 16235
rect 6546 16232 6552 16244
rect 6507 16204 6552 16232
rect 5077 16195 5135 16201
rect 6546 16192 6552 16204
rect 6604 16192 6610 16244
rect 6730 16192 6736 16244
rect 6788 16232 6794 16244
rect 7561 16235 7619 16241
rect 7561 16232 7573 16235
rect 6788 16204 7573 16232
rect 6788 16192 6794 16204
rect 7561 16201 7573 16204
rect 7607 16201 7619 16235
rect 7926 16232 7932 16244
rect 7887 16204 7932 16232
rect 7561 16195 7619 16201
rect 7926 16192 7932 16204
rect 7984 16192 7990 16244
rect 8478 16192 8484 16244
rect 8536 16232 8542 16244
rect 10686 16232 10692 16244
rect 8536 16204 10692 16232
rect 8536 16192 8542 16204
rect 10686 16192 10692 16204
rect 10744 16192 10750 16244
rect 14553 16235 14611 16241
rect 14553 16201 14565 16235
rect 14599 16232 14611 16235
rect 15010 16232 15016 16244
rect 14599 16204 15016 16232
rect 14599 16201 14611 16204
rect 14553 16195 14611 16201
rect 15010 16192 15016 16204
rect 15068 16192 15074 16244
rect 16390 16192 16396 16244
rect 16448 16232 16454 16244
rect 16669 16235 16727 16241
rect 16669 16232 16681 16235
rect 16448 16204 16681 16232
rect 16448 16192 16454 16204
rect 16669 16201 16681 16204
rect 16715 16201 16727 16235
rect 16669 16195 16727 16201
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17586 16232 17592 16244
rect 17368 16204 17592 16232
rect 17368 16192 17374 16204
rect 17586 16192 17592 16204
rect 17644 16192 17650 16244
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 18325 16235 18383 16241
rect 18325 16232 18337 16235
rect 17727 16204 18337 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18325 16201 18337 16204
rect 18371 16201 18383 16235
rect 18325 16195 18383 16201
rect 18506 16192 18512 16244
rect 18564 16232 18570 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18564 16204 18797 16232
rect 18564 16192 18570 16204
rect 18785 16201 18797 16204
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 20714 16232 20720 16244
rect 20211 16204 20720 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 3053 16167 3111 16173
rect 3053 16133 3065 16167
rect 3099 16164 3111 16167
rect 6917 16167 6975 16173
rect 3099 16136 6868 16164
rect 3099 16133 3111 16136
rect 3053 16127 3111 16133
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2222 16096 2228 16108
rect 2183 16068 2228 16096
rect 2222 16056 2228 16068
rect 2280 16056 2286 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 3068 16096 3096 16127
rect 4430 16096 4436 16108
rect 2731 16068 3096 16096
rect 4391 16068 4436 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 4430 16056 4436 16068
rect 4488 16056 4494 16108
rect 5442 16096 5448 16108
rect 5403 16068 5448 16096
rect 5442 16056 5448 16068
rect 5500 16056 5506 16108
rect 6840 16096 6868 16136
rect 6917 16133 6929 16167
rect 6963 16164 6975 16167
rect 7742 16164 7748 16176
rect 6963 16136 7748 16164
rect 6963 16133 6975 16136
rect 6917 16127 6975 16133
rect 7742 16124 7748 16136
rect 7800 16124 7806 16176
rect 10134 16124 10140 16176
rect 10192 16124 10198 16176
rect 10410 16124 10416 16176
rect 10468 16164 10474 16176
rect 14093 16167 14151 16173
rect 14093 16164 14105 16167
rect 10468 16136 11376 16164
rect 10468 16124 10474 16136
rect 7374 16096 7380 16108
rect 6840 16068 7380 16096
rect 7374 16056 7380 16068
rect 7432 16056 7438 16108
rect 7466 16056 7472 16108
rect 7524 16096 7530 16108
rect 9674 16096 9680 16108
rect 7524 16068 9680 16096
rect 7524 16056 7530 16068
rect 4062 15988 4068 16040
rect 4120 15988 4126 16040
rect 4522 16028 4528 16040
rect 4483 16000 4528 16028
rect 4522 15988 4528 16000
rect 4580 15988 4586 16040
rect 4709 16031 4767 16037
rect 4709 15997 4721 16031
rect 4755 16028 4767 16031
rect 4890 16028 4896 16040
rect 4755 16000 4896 16028
rect 4755 15997 4767 16000
rect 4709 15991 4767 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 5350 15988 5356 16040
rect 5408 16028 5414 16040
rect 5537 16031 5595 16037
rect 5537 16028 5549 16031
rect 5408 16000 5549 16028
rect 5408 15988 5414 16000
rect 5537 15997 5549 16000
rect 5583 15997 5595 16031
rect 5537 15991 5595 15997
rect 5629 16031 5687 16037
rect 5629 15997 5641 16031
rect 5675 15997 5687 16031
rect 7006 16028 7012 16040
rect 6967 16000 7012 16028
rect 5629 15991 5687 15997
rect 1394 15920 1400 15972
rect 1452 15960 1458 15972
rect 2041 15963 2099 15969
rect 2041 15960 2053 15963
rect 1452 15932 2053 15960
rect 1452 15920 1458 15932
rect 2041 15929 2053 15932
rect 2087 15929 2099 15963
rect 2041 15923 2099 15929
rect 2774 15920 2780 15972
rect 2832 15960 2838 15972
rect 3697 15963 3755 15969
rect 3697 15960 3709 15963
rect 2832 15932 3709 15960
rect 2832 15920 2838 15932
rect 3697 15929 3709 15932
rect 3743 15929 3755 15963
rect 4080 15960 4108 15988
rect 5644 15960 5672 15991
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7193 16031 7251 16037
rect 7193 15997 7205 16031
rect 7239 16028 7251 16031
rect 7558 16028 7564 16040
rect 7239 16000 7564 16028
rect 7239 15997 7251 16000
rect 7193 15991 7251 15997
rect 7558 15988 7564 16000
rect 7616 16028 7622 16040
rect 8018 16028 8024 16040
rect 7616 16000 7709 16028
rect 7979 16000 8024 16028
rect 7616 15988 7622 16000
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 8128 16037 8156 16068
rect 9674 16056 9680 16068
rect 9732 16056 9738 16108
rect 10152 16096 10180 16124
rect 10249 16099 10307 16105
rect 10249 16096 10261 16099
rect 10152 16068 10261 16096
rect 10249 16065 10261 16068
rect 10295 16096 10307 16099
rect 11238 16096 11244 16108
rect 10295 16068 11244 16096
rect 10295 16065 10307 16068
rect 10249 16059 10307 16065
rect 11238 16056 11244 16068
rect 11296 16056 11302 16108
rect 8113 16031 8171 16037
rect 8113 15997 8125 16031
rect 8159 15997 8171 16031
rect 8113 15991 8171 15997
rect 10505 16031 10563 16037
rect 10505 15997 10517 16031
rect 10551 16028 10563 16031
rect 11348 16028 11376 16136
rect 13280 16136 14105 16164
rect 10551 16000 10824 16028
rect 11348 16000 11652 16028
rect 10551 15997 10563 16000
rect 10505 15991 10563 15997
rect 6730 15960 6736 15972
rect 4080 15932 6736 15960
rect 3697 15923 3755 15929
rect 6730 15920 6736 15932
rect 6788 15920 6794 15972
rect 7576 15960 7604 15988
rect 7576 15932 9444 15960
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 4062 15892 4068 15904
rect 4023 15864 4068 15892
rect 4062 15852 4068 15864
rect 4120 15852 4126 15904
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 6914 15892 6920 15904
rect 4212 15864 6920 15892
rect 4212 15852 4218 15864
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7006 15852 7012 15904
rect 7064 15892 7070 15904
rect 7742 15892 7748 15904
rect 7064 15864 7748 15892
rect 7064 15852 7070 15864
rect 7742 15852 7748 15864
rect 7800 15892 7806 15904
rect 8110 15892 8116 15904
rect 7800 15864 8116 15892
rect 7800 15852 7806 15864
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 8573 15895 8631 15901
rect 8573 15892 8585 15895
rect 8536 15864 8585 15892
rect 8536 15852 8542 15864
rect 8573 15861 8585 15864
rect 8619 15861 8631 15895
rect 9122 15892 9128 15904
rect 9083 15864 9128 15892
rect 8573 15855 8631 15861
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 9416 15892 9444 15932
rect 10796 15904 10824 16000
rect 11624 15969 11652 16000
rect 11609 15963 11667 15969
rect 11609 15929 11621 15963
rect 11655 15960 11667 15963
rect 13170 15960 13176 15972
rect 11655 15932 13176 15960
rect 11655 15929 11667 15932
rect 11609 15923 11667 15929
rect 13170 15920 13176 15932
rect 13228 15920 13234 15972
rect 10594 15892 10600 15904
rect 9416 15864 10600 15892
rect 10594 15852 10600 15864
rect 10652 15852 10658 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 10870 15852 10876 15904
rect 10928 15892 10934 15904
rect 12066 15892 12072 15904
rect 10928 15864 12072 15892
rect 10928 15852 10934 15864
rect 12066 15852 12072 15864
rect 12124 15852 12130 15904
rect 12618 15852 12624 15904
rect 12676 15892 12682 15904
rect 13280 15892 13308 16136
rect 14093 16133 14105 16136
rect 14139 16133 14151 16167
rect 17034 16164 17040 16176
rect 14093 16127 14151 16133
rect 15396 16136 17040 16164
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13688 16068 14197 16096
rect 13688 16056 13694 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 15396 16040 15424 16136
rect 17034 16124 17040 16136
rect 17092 16124 17098 16176
rect 17310 16056 17316 16108
rect 17368 16096 17374 16108
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 17368 16068 17601 16096
rect 17368 16056 17374 16068
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 17589 16059 17647 16065
rect 18046 16056 18052 16108
rect 18104 16056 18110 16108
rect 18693 16099 18751 16105
rect 18693 16065 18705 16099
rect 18739 16096 18751 16099
rect 19337 16099 19395 16105
rect 19337 16096 19349 16099
rect 18739 16068 19349 16096
rect 18739 16065 18751 16068
rect 18693 16059 18751 16065
rect 19337 16065 19349 16068
rect 19383 16065 19395 16099
rect 19978 16096 19984 16108
rect 19939 16068 19984 16096
rect 19337 16059 19395 16065
rect 19978 16056 19984 16068
rect 20036 16056 20042 16108
rect 20530 16096 20536 16108
rect 20491 16068 20536 16096
rect 20530 16056 20536 16068
rect 20588 16056 20594 16108
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20956 16068 21097 16096
rect 20956 16056 20962 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 15378 16028 15384 16040
rect 14047 16000 15384 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 15378 15988 15384 16000
rect 15436 15988 15442 16040
rect 17497 16031 17555 16037
rect 17497 15997 17509 16031
rect 17543 16028 17555 16031
rect 18064 16028 18092 16056
rect 18874 16028 18880 16040
rect 17543 16000 18092 16028
rect 18835 16000 18880 16028
rect 17543 15997 17555 16000
rect 17497 15991 17555 15997
rect 18874 15988 18880 16000
rect 18932 15988 18938 16040
rect 13354 15920 13360 15972
rect 13412 15960 13418 15972
rect 17678 15960 17684 15972
rect 13412 15932 17684 15960
rect 13412 15920 13418 15932
rect 17678 15920 17684 15932
rect 17736 15920 17742 15972
rect 18049 15963 18107 15969
rect 18049 15929 18061 15963
rect 18095 15960 18107 15963
rect 20346 15960 20352 15972
rect 18095 15932 20352 15960
rect 18095 15929 18107 15932
rect 18049 15923 18107 15929
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 20714 15960 20720 15972
rect 20675 15932 20720 15960
rect 20714 15920 20720 15932
rect 20772 15920 20778 15972
rect 13449 15895 13507 15901
rect 13449 15892 13461 15895
rect 12676 15864 13461 15892
rect 12676 15852 12682 15864
rect 13449 15861 13461 15864
rect 13495 15861 13507 15895
rect 13449 15855 13507 15861
rect 14921 15895 14979 15901
rect 14921 15861 14933 15895
rect 14967 15892 14979 15895
rect 15378 15892 15384 15904
rect 14967 15864 15384 15892
rect 14967 15861 14979 15864
rect 14921 15855 14979 15861
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 4430 15688 4436 15700
rect 4391 15660 4436 15688
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4706 15648 4712 15700
rect 4764 15688 4770 15700
rect 4764 15660 7604 15688
rect 4764 15648 4770 15660
rect 842 15580 848 15632
rect 900 15620 906 15632
rect 5442 15620 5448 15632
rect 900 15592 5448 15620
rect 900 15580 906 15592
rect 5442 15580 5448 15592
rect 5500 15620 5506 15632
rect 6917 15623 6975 15629
rect 5500 15592 6500 15620
rect 5500 15580 5506 15592
rect 3418 15512 3424 15564
rect 3476 15552 3482 15564
rect 4893 15555 4951 15561
rect 4893 15552 4905 15555
rect 3476 15524 4905 15552
rect 3476 15512 3482 15524
rect 4893 15521 4905 15524
rect 4939 15521 4951 15555
rect 5074 15552 5080 15564
rect 5035 15524 5080 15552
rect 4893 15515 4951 15521
rect 5074 15512 5080 15524
rect 5132 15512 5138 15564
rect 6472 15561 6500 15592
rect 6917 15589 6929 15623
rect 6963 15589 6975 15623
rect 6917 15583 6975 15589
rect 6365 15555 6423 15561
rect 6365 15521 6377 15555
rect 6411 15521 6423 15555
rect 6365 15515 6423 15521
rect 6457 15555 6515 15561
rect 6457 15521 6469 15555
rect 6503 15521 6515 15555
rect 6457 15515 6515 15521
rect 1394 15444 1400 15496
rect 1452 15484 1458 15496
rect 1673 15487 1731 15493
rect 1673 15484 1685 15487
rect 1452 15456 1685 15484
rect 1452 15444 1458 15456
rect 1673 15453 1685 15456
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 2133 15487 2191 15493
rect 2133 15453 2145 15487
rect 2179 15484 2191 15487
rect 2590 15484 2596 15496
rect 2179 15456 2452 15484
rect 2551 15456 2596 15484
rect 2179 15453 2191 15456
rect 2133 15447 2191 15453
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 1946 15348 1952 15360
rect 1907 15320 1952 15348
rect 1946 15308 1952 15320
rect 2004 15308 2010 15360
rect 2424 15357 2452 15456
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 5166 15444 5172 15496
rect 5224 15484 5230 15496
rect 6380 15484 6408 15515
rect 6822 15484 6828 15496
rect 5224 15456 6316 15484
rect 6380 15456 6828 15484
rect 5224 15444 5230 15456
rect 4801 15419 4859 15425
rect 4801 15385 4813 15419
rect 4847 15416 4859 15419
rect 5445 15419 5503 15425
rect 5445 15416 5457 15419
rect 4847 15388 5457 15416
rect 4847 15385 4859 15388
rect 4801 15379 4859 15385
rect 5445 15385 5457 15388
rect 5491 15385 5503 15419
rect 6288 15416 6316 15456
rect 6822 15444 6828 15456
rect 6880 15444 6886 15496
rect 6932 15416 6960 15583
rect 7006 15444 7012 15496
rect 7064 15484 7070 15496
rect 7466 15484 7472 15496
rect 7064 15456 7472 15484
rect 7064 15444 7070 15456
rect 7466 15444 7472 15456
rect 7524 15444 7530 15496
rect 7576 15484 7604 15660
rect 8018 15648 8024 15700
rect 8076 15688 8082 15700
rect 8205 15691 8263 15697
rect 8205 15688 8217 15691
rect 8076 15660 8217 15688
rect 8076 15648 8082 15660
rect 8205 15657 8217 15660
rect 8251 15657 8263 15691
rect 8205 15651 8263 15657
rect 9122 15648 9128 15700
rect 9180 15648 9186 15700
rect 10226 15648 10232 15700
rect 10284 15688 10290 15700
rect 10597 15691 10655 15697
rect 10597 15688 10609 15691
rect 10284 15660 10609 15688
rect 10284 15648 10290 15660
rect 10597 15657 10609 15660
rect 10643 15657 10655 15691
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 10597 15651 10655 15657
rect 10704 15660 12357 15688
rect 8110 15580 8116 15632
rect 8168 15620 8174 15632
rect 9140 15620 9168 15648
rect 8168 15592 9168 15620
rect 8168 15580 8174 15592
rect 10410 15580 10416 15632
rect 10468 15620 10474 15632
rect 10704 15620 10732 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 13630 15688 13636 15700
rect 13591 15660 13636 15688
rect 12345 15651 12403 15657
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 16945 15691 17003 15697
rect 16945 15688 16957 15691
rect 13740 15660 16957 15688
rect 11974 15620 11980 15632
rect 10468 15592 10732 15620
rect 11935 15592 11980 15620
rect 10468 15580 10474 15592
rect 11974 15580 11980 15592
rect 12032 15580 12038 15632
rect 12066 15580 12072 15632
rect 12124 15620 12130 15632
rect 13740 15620 13768 15660
rect 16945 15657 16957 15660
rect 16991 15688 17003 15691
rect 17218 15688 17224 15700
rect 16991 15660 17224 15688
rect 16991 15657 17003 15660
rect 16945 15651 17003 15657
rect 17218 15648 17224 15660
rect 17276 15648 17282 15700
rect 17678 15648 17684 15700
rect 17736 15688 17742 15700
rect 18509 15691 18567 15697
rect 18509 15688 18521 15691
rect 17736 15660 18521 15688
rect 17736 15648 17742 15660
rect 18509 15657 18521 15660
rect 18555 15688 18567 15691
rect 19702 15688 19708 15700
rect 18555 15660 19708 15688
rect 18555 15657 18567 15660
rect 18509 15651 18567 15657
rect 19702 15648 19708 15660
rect 19760 15648 19766 15700
rect 19797 15691 19855 15697
rect 19797 15657 19809 15691
rect 19843 15688 19855 15691
rect 20530 15688 20536 15700
rect 19843 15660 20536 15688
rect 19843 15657 19855 15660
rect 19797 15651 19855 15657
rect 20530 15648 20536 15660
rect 20588 15648 20594 15700
rect 12124 15592 13768 15620
rect 12124 15580 12130 15592
rect 7653 15555 7711 15561
rect 7653 15521 7665 15555
rect 7699 15552 7711 15555
rect 9122 15552 9128 15564
rect 7699 15524 9128 15552
rect 7699 15521 7711 15524
rect 7653 15515 7711 15521
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15552 11759 15555
rect 12434 15552 12440 15564
rect 11747 15524 12440 15552
rect 11747 15521 11759 15524
rect 11701 15515 11759 15521
rect 12434 15512 12440 15524
rect 12492 15512 12498 15564
rect 7745 15487 7803 15493
rect 7745 15484 7757 15487
rect 7576 15456 7757 15484
rect 7745 15453 7757 15456
rect 7791 15484 7803 15487
rect 8481 15487 8539 15493
rect 8481 15484 8493 15487
rect 7791 15456 8493 15484
rect 7791 15453 7803 15456
rect 7745 15447 7803 15453
rect 8481 15453 8493 15456
rect 8527 15453 8539 15487
rect 9214 15484 9220 15496
rect 9175 15456 9220 15484
rect 8481 15447 8539 15453
rect 9214 15444 9220 15456
rect 9272 15484 9278 15496
rect 10778 15484 10784 15496
rect 9272 15456 10784 15484
rect 9272 15444 9278 15456
rect 10778 15444 10784 15456
rect 10836 15484 10842 15496
rect 10873 15487 10931 15493
rect 10873 15484 10885 15487
rect 10836 15456 10885 15484
rect 10836 15444 10842 15456
rect 10873 15453 10885 15456
rect 10919 15453 10931 15487
rect 12710 15484 12716 15496
rect 10873 15447 10931 15453
rect 10980 15456 12716 15484
rect 9490 15425 9496 15428
rect 6288 15388 6868 15416
rect 6932 15388 9444 15416
rect 5445 15379 5503 15385
rect 2409 15351 2467 15357
rect 2409 15317 2421 15351
rect 2455 15317 2467 15351
rect 2409 15311 2467 15317
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 2869 15351 2927 15357
rect 2869 15348 2881 15351
rect 2740 15320 2881 15348
rect 2740 15308 2746 15320
rect 2869 15317 2881 15320
rect 2915 15317 2927 15351
rect 2869 15311 2927 15317
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 3108 15320 3341 15348
rect 3108 15308 3114 15320
rect 3329 15317 3341 15320
rect 3375 15317 3387 15351
rect 3329 15311 3387 15317
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 3973 15351 4031 15357
rect 3973 15348 3985 15351
rect 3844 15320 3985 15348
rect 3844 15308 3850 15320
rect 3973 15317 3985 15320
rect 4019 15317 4031 15351
rect 6546 15348 6552 15360
rect 6507 15320 6552 15348
rect 3973 15311 4031 15317
rect 6546 15308 6552 15320
rect 6604 15308 6610 15360
rect 6840 15348 6868 15388
rect 7837 15351 7895 15357
rect 7837 15348 7849 15351
rect 6840 15320 7849 15348
rect 7837 15317 7849 15320
rect 7883 15348 7895 15351
rect 8478 15348 8484 15360
rect 7883 15320 8484 15348
rect 7883 15317 7895 15320
rect 7837 15311 7895 15317
rect 8478 15308 8484 15320
rect 8536 15308 8542 15360
rect 9416 15348 9444 15388
rect 9484 15379 9496 15425
rect 9548 15416 9554 15428
rect 10686 15416 10692 15428
rect 9548 15388 10692 15416
rect 9490 15376 9496 15379
rect 9548 15376 9554 15388
rect 10686 15376 10692 15388
rect 10744 15376 10750 15428
rect 10980 15348 11008 15456
rect 12710 15444 12716 15456
rect 12768 15444 12774 15496
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13044 15456 16436 15484
rect 13044 15444 13050 15456
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 13814 15416 13820 15428
rect 11296 15388 13820 15416
rect 11296 15376 11302 15388
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 16310 15419 16368 15425
rect 16310 15385 16322 15419
rect 16356 15385 16368 15419
rect 16408 15416 16436 15456
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16632 15456 17233 15484
rect 16632 15444 16638 15456
rect 17221 15453 17233 15456
rect 17267 15484 17279 15487
rect 17678 15484 17684 15496
rect 17267 15456 17684 15484
rect 17267 15453 17279 15456
rect 17221 15447 17279 15453
rect 17678 15444 17684 15456
rect 17736 15484 17742 15496
rect 18785 15487 18843 15493
rect 18785 15484 18797 15487
rect 17736 15456 18797 15484
rect 17736 15444 17742 15456
rect 18785 15453 18797 15456
rect 18831 15453 18843 15487
rect 18785 15447 18843 15453
rect 19518 15444 19524 15496
rect 19576 15484 19582 15496
rect 19613 15487 19671 15493
rect 19613 15484 19625 15487
rect 19576 15456 19625 15484
rect 19576 15444 19582 15456
rect 19613 15453 19625 15456
rect 19659 15453 19671 15487
rect 19613 15447 19671 15453
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20533 15487 20591 15493
rect 20533 15484 20545 15487
rect 20073 15447 20131 15453
rect 20272 15456 20545 15484
rect 18141 15419 18199 15425
rect 18141 15416 18153 15419
rect 16408 15388 18153 15416
rect 16310 15379 16368 15385
rect 18141 15385 18153 15388
rect 18187 15416 18199 15419
rect 20088 15416 20116 15447
rect 18187 15388 20116 15416
rect 18187 15385 18199 15388
rect 18141 15379 18199 15385
rect 9416 15320 11008 15348
rect 11333 15351 11391 15357
rect 11333 15317 11345 15351
rect 11379 15348 11391 15351
rect 11882 15348 11888 15360
rect 11379 15320 11888 15348
rect 11379 15317 11391 15320
rect 11333 15311 11391 15317
rect 11882 15308 11888 15320
rect 11940 15308 11946 15360
rect 15194 15348 15200 15360
rect 15107 15320 15200 15348
rect 15194 15308 15200 15320
rect 15252 15348 15258 15360
rect 16114 15348 16120 15360
rect 15252 15320 16120 15348
rect 15252 15308 15258 15320
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16316 15348 16344 15379
rect 16758 15348 16764 15360
rect 16316 15320 16764 15348
rect 16758 15308 16764 15320
rect 16816 15308 16822 15360
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 19518 15348 19524 15360
rect 19383 15320 19524 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 20272 15357 20300 15456
rect 20533 15453 20545 15456
rect 20579 15453 20591 15487
rect 20533 15447 20591 15453
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 20346 15376 20352 15428
rect 20404 15416 20410 15428
rect 21100 15416 21128 15447
rect 20404 15388 21128 15416
rect 20404 15376 20410 15388
rect 20257 15351 20315 15357
rect 20257 15317 20269 15351
rect 20303 15317 20315 15351
rect 20257 15311 20315 15317
rect 20717 15351 20775 15357
rect 20717 15317 20729 15351
rect 20763 15348 20775 15351
rect 20806 15348 20812 15360
rect 20763 15320 20812 15348
rect 20763 15317 20775 15320
rect 20717 15311 20775 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 2501 15147 2559 15153
rect 2501 15113 2513 15147
rect 2547 15113 2559 15147
rect 2501 15107 2559 15113
rect 2516 15076 2544 15107
rect 4246 15104 4252 15156
rect 4304 15144 4310 15156
rect 4341 15147 4399 15153
rect 4341 15144 4353 15147
rect 4304 15116 4353 15144
rect 4304 15104 4310 15116
rect 4341 15113 4353 15116
rect 4387 15144 4399 15147
rect 5534 15144 5540 15156
rect 4387 15116 5540 15144
rect 4387 15113 4399 15116
rect 4341 15107 4399 15113
rect 5534 15104 5540 15116
rect 5592 15104 5598 15156
rect 5902 15104 5908 15156
rect 5960 15104 5966 15156
rect 6641 15147 6699 15153
rect 6641 15113 6653 15147
rect 6687 15144 6699 15147
rect 6822 15144 6828 15156
rect 6687 15116 6828 15144
rect 6687 15113 6699 15116
rect 6641 15107 6699 15113
rect 6822 15104 6828 15116
rect 6880 15104 6886 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7009 15147 7067 15153
rect 7009 15144 7021 15147
rect 6972 15116 7021 15144
rect 6972 15104 6978 15116
rect 7009 15113 7021 15116
rect 7055 15144 7067 15147
rect 7653 15147 7711 15153
rect 7653 15144 7665 15147
rect 7055 15116 7665 15144
rect 7055 15113 7067 15116
rect 7009 15107 7067 15113
rect 7653 15113 7665 15116
rect 7699 15144 7711 15147
rect 9674 15144 9680 15156
rect 7699 15116 9680 15144
rect 7699 15113 7711 15116
rect 7653 15107 7711 15113
rect 9674 15104 9680 15116
rect 9732 15104 9738 15156
rect 9876 15116 10088 15144
rect 1688 15048 2544 15076
rect 5920 15076 5948 15104
rect 5920 15048 7052 15076
rect 1688 15017 1716 15048
rect 7024 15020 7052 15048
rect 7190 15036 7196 15088
rect 7248 15076 7254 15088
rect 7745 15079 7803 15085
rect 7745 15076 7757 15079
rect 7248 15048 7757 15076
rect 7248 15036 7254 15048
rect 7745 15045 7757 15048
rect 7791 15076 7803 15079
rect 7926 15076 7932 15088
rect 7791 15048 7932 15076
rect 7791 15045 7803 15048
rect 7745 15039 7803 15045
rect 7926 15036 7932 15048
rect 7984 15076 7990 15088
rect 8297 15079 8355 15085
rect 8297 15076 8309 15079
rect 7984 15048 8309 15076
rect 7984 15036 7990 15048
rect 8297 15045 8309 15048
rect 8343 15045 8355 15079
rect 8297 15039 8355 15045
rect 8662 15036 8668 15088
rect 8720 15036 8726 15088
rect 8757 15079 8815 15085
rect 8757 15045 8769 15079
rect 8803 15076 8815 15079
rect 9876 15076 9904 15116
rect 8803 15048 9904 15076
rect 10060 15076 10088 15116
rect 10778 15104 10784 15156
rect 10836 15144 10842 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 10836 15116 11529 15144
rect 10836 15104 10842 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 12802 15104 12808 15156
rect 12860 15144 12866 15156
rect 13722 15144 13728 15156
rect 12860 15116 13728 15144
rect 12860 15104 12866 15116
rect 13722 15104 13728 15116
rect 13780 15104 13786 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15144 16727 15147
rect 16942 15144 16948 15156
rect 16715 15116 16948 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 19702 15104 19708 15156
rect 19760 15144 19766 15156
rect 20530 15144 20536 15156
rect 19760 15116 20536 15144
rect 19760 15104 19766 15116
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 11238 15076 11244 15088
rect 10060 15048 11244 15076
rect 8803 15045 8815 15048
rect 8757 15039 8815 15045
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 18325 15079 18383 15085
rect 18325 15076 18337 15079
rect 17736 15048 18337 15076
rect 17736 15036 17742 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 1949 15011 2007 15017
rect 1949 14977 1961 15011
rect 1995 15008 2007 15011
rect 2038 15008 2044 15020
rect 1995 14980 2044 15008
rect 1995 14977 2007 14980
rect 1949 14971 2007 14977
rect 2038 14968 2044 14980
rect 2096 14968 2102 15020
rect 2682 15008 2688 15020
rect 2643 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 14968 2746 15020
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 4982 15008 4988 15020
rect 3191 14980 3280 15008
rect 4943 14980 4988 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 2961 14875 3019 14881
rect 2961 14872 2973 14875
rect 1728 14844 2973 14872
rect 1728 14832 1734 14844
rect 2961 14841 2973 14844
rect 3007 14841 3019 14875
rect 2961 14835 3019 14841
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2130 14804 2136 14816
rect 2091 14776 2136 14804
rect 2130 14764 2136 14776
rect 2188 14764 2194 14816
rect 3252 14804 3280 14980
rect 4982 14968 4988 14980
rect 5040 14968 5046 15020
rect 5077 15011 5135 15017
rect 5077 14977 5089 15011
rect 5123 15008 5135 15011
rect 5902 15008 5908 15020
rect 5123 14980 5908 15008
rect 5123 14977 5135 14980
rect 5077 14971 5135 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 8680 15008 8708 15036
rect 7064 14980 8708 15008
rect 7064 14968 7070 14980
rect 9214 14968 9220 15020
rect 9272 15008 9278 15020
rect 9674 15008 9680 15020
rect 9272 14980 9680 15008
rect 9272 14968 9278 14980
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 9766 14968 9772 15020
rect 9824 15008 9830 15020
rect 9944 15011 10002 15017
rect 9944 15008 9956 15011
rect 9824 14980 9956 15008
rect 9824 14968 9830 14980
rect 9944 14977 9956 14980
rect 9990 14977 10002 15011
rect 9944 14971 10002 14977
rect 10318 14968 10324 15020
rect 10376 15008 10382 15020
rect 12253 15011 12311 15017
rect 12253 15008 12265 15011
rect 10376 14980 12265 15008
rect 10376 14968 10382 14980
rect 12253 14977 12265 14980
rect 12299 14977 12311 15011
rect 12253 14971 12311 14977
rect 13449 15011 13507 15017
rect 13449 14977 13461 15011
rect 13495 14977 13507 15011
rect 13449 14971 13507 14977
rect 13716 15011 13774 15017
rect 13716 14977 13728 15011
rect 13762 15008 13774 15011
rect 15930 15008 15936 15020
rect 13762 14980 15936 15008
rect 13762 14977 13774 14980
rect 13716 14971 13774 14977
rect 4890 14900 4896 14952
rect 4948 14940 4954 14952
rect 5261 14943 5319 14949
rect 5261 14940 5273 14943
rect 4948 14912 5273 14940
rect 4948 14900 4954 14912
rect 5261 14909 5273 14912
rect 5307 14940 5319 14943
rect 5350 14940 5356 14952
rect 5307 14912 5356 14940
rect 5307 14909 5319 14912
rect 5261 14903 5319 14909
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 7834 14900 7840 14952
rect 7892 14940 7898 14952
rect 7929 14943 7987 14949
rect 7929 14940 7941 14943
rect 7892 14912 7941 14940
rect 7892 14900 7898 14912
rect 7929 14909 7941 14912
rect 7975 14940 7987 14943
rect 7975 14912 8432 14940
rect 7975 14909 7987 14912
rect 7929 14903 7987 14909
rect 3326 14832 3332 14884
rect 3384 14872 3390 14884
rect 3789 14875 3847 14881
rect 3789 14872 3801 14875
rect 3384 14844 3801 14872
rect 3384 14832 3390 14844
rect 3789 14841 3801 14844
rect 3835 14841 3847 14875
rect 3789 14835 3847 14841
rect 3988 14844 4936 14872
rect 3513 14807 3571 14813
rect 3513 14804 3525 14807
rect 3252 14776 3525 14804
rect 3513 14773 3525 14776
rect 3559 14804 3571 14807
rect 3988 14804 4016 14844
rect 4908 14816 4936 14844
rect 3559 14776 4016 14804
rect 3559 14773 3571 14776
rect 3513 14767 3571 14773
rect 4430 14764 4436 14816
rect 4488 14804 4494 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4488 14776 4629 14804
rect 4488 14764 4494 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 4890 14764 4896 14816
rect 4948 14764 4954 14816
rect 5997 14807 6055 14813
rect 5997 14773 6009 14807
rect 6043 14804 6055 14807
rect 6546 14804 6552 14816
rect 6043 14776 6552 14804
rect 6043 14773 6055 14776
rect 5997 14767 6055 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 7285 14807 7343 14813
rect 7285 14804 7297 14807
rect 7248 14776 7297 14804
rect 7248 14764 7254 14776
rect 7285 14773 7297 14776
rect 7331 14773 7343 14807
rect 8404 14804 8432 14912
rect 8662 14900 8668 14952
rect 8720 14940 8726 14952
rect 9033 14943 9091 14949
rect 9033 14940 9045 14943
rect 8720 14912 9045 14940
rect 8720 14900 8726 14912
rect 9033 14909 9045 14912
rect 9079 14909 9091 14943
rect 9033 14903 9091 14909
rect 11606 14900 11612 14952
rect 11664 14940 11670 14952
rect 12986 14940 12992 14952
rect 11664 14912 12992 14940
rect 11664 14900 11670 14912
rect 12986 14900 12992 14912
rect 13044 14900 13050 14952
rect 10778 14832 10784 14884
rect 10836 14872 10842 14884
rect 13464 14872 13492 14971
rect 15930 14968 15936 14980
rect 15988 14968 15994 15020
rect 17218 14968 17224 15020
rect 17276 15008 17282 15020
rect 18064 15017 18092 15048
rect 18325 15045 18337 15048
rect 18371 15076 18383 15079
rect 18877 15079 18935 15085
rect 18877 15076 18889 15079
rect 18371 15048 18889 15076
rect 18371 15045 18383 15048
rect 18325 15039 18383 15045
rect 18877 15045 18889 15048
rect 18923 15045 18935 15079
rect 20714 15076 20720 15088
rect 18877 15039 18935 15045
rect 19904 15048 20720 15076
rect 17782 15011 17840 15017
rect 17782 15008 17794 15011
rect 17276 14980 17794 15008
rect 17276 14968 17282 14980
rect 17782 14977 17794 14980
rect 17828 14977 17840 15011
rect 17782 14971 17840 14977
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18690 14968 18696 15020
rect 18748 15008 18754 15020
rect 19904 15017 19932 15048
rect 20714 15036 20720 15048
rect 20772 15036 20778 15088
rect 19429 15011 19487 15017
rect 19429 15008 19441 15011
rect 18748 14980 19441 15008
rect 18748 14968 18754 14980
rect 19429 14977 19441 14980
rect 19475 14977 19487 15011
rect 19429 14971 19487 14977
rect 19889 15011 19947 15017
rect 19889 14977 19901 15011
rect 19935 14977 19947 15011
rect 20145 15011 20203 15017
rect 20145 15008 20157 15011
rect 19889 14971 19947 14977
rect 19996 14980 20157 15008
rect 10836 14844 13492 14872
rect 14476 14912 16574 14940
rect 10836 14832 10842 14844
rect 10042 14804 10048 14816
rect 8404 14776 10048 14804
rect 7285 14767 7343 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11422 14804 11428 14816
rect 11103 14776 11428 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 11974 14804 11980 14816
rect 11935 14776 11980 14804
rect 11974 14764 11980 14776
rect 12032 14764 12038 14816
rect 12710 14804 12716 14816
rect 12671 14776 12716 14804
rect 12710 14764 12716 14776
rect 12768 14764 12774 14816
rect 12986 14804 12992 14816
rect 12947 14776 12992 14804
rect 12986 14764 12992 14776
rect 13044 14764 13050 14816
rect 13078 14764 13084 14816
rect 13136 14804 13142 14816
rect 14476 14804 14504 14912
rect 14734 14832 14740 14884
rect 14792 14872 14798 14884
rect 14829 14875 14887 14881
rect 14829 14872 14841 14875
rect 14792 14844 14841 14872
rect 14792 14832 14798 14844
rect 14829 14841 14841 14844
rect 14875 14872 14887 14875
rect 15010 14872 15016 14884
rect 14875 14844 15016 14872
rect 14875 14841 14887 14844
rect 14829 14835 14887 14841
rect 15010 14832 15016 14844
rect 15068 14832 15074 14884
rect 16390 14872 16396 14884
rect 15580 14844 16396 14872
rect 13136 14776 14504 14804
rect 13136 14764 13142 14776
rect 14918 14764 14924 14816
rect 14976 14804 14982 14816
rect 15580 14813 15608 14844
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 15105 14807 15163 14813
rect 15105 14804 15117 14807
rect 14976 14776 15117 14804
rect 14976 14764 14982 14776
rect 15105 14773 15117 14776
rect 15151 14804 15163 14807
rect 15565 14807 15623 14813
rect 15565 14804 15577 14807
rect 15151 14776 15577 14804
rect 15151 14773 15163 14776
rect 15105 14767 15163 14773
rect 15565 14773 15577 14776
rect 15611 14773 15623 14807
rect 16022 14804 16028 14816
rect 15983 14776 16028 14804
rect 15565 14767 15623 14773
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 16546 14804 16574 14912
rect 19794 14900 19800 14952
rect 19852 14940 19858 14952
rect 19996 14940 20024 14980
rect 20145 14977 20157 14980
rect 20191 14977 20203 15011
rect 20145 14971 20203 14977
rect 19852 14912 20024 14940
rect 19852 14900 19858 14912
rect 18690 14804 18696 14816
rect 16546 14776 18696 14804
rect 18690 14764 18696 14776
rect 18748 14764 18754 14816
rect 19613 14807 19671 14813
rect 19613 14773 19625 14807
rect 19659 14804 19671 14807
rect 19886 14804 19892 14816
rect 19659 14776 19892 14804
rect 19659 14773 19671 14776
rect 19613 14767 19671 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20990 14764 20996 14816
rect 21048 14804 21054 14816
rect 21174 14804 21180 14816
rect 21048 14776 21180 14804
rect 21048 14764 21054 14776
rect 21174 14764 21180 14776
rect 21232 14804 21238 14816
rect 21269 14807 21327 14813
rect 21269 14804 21281 14807
rect 21232 14776 21281 14804
rect 21232 14764 21238 14776
rect 21269 14773 21281 14776
rect 21315 14773 21327 14807
rect 21269 14767 21327 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 4982 14560 4988 14612
rect 5040 14600 5046 14612
rect 5077 14603 5135 14609
rect 5077 14600 5089 14603
rect 5040 14572 5089 14600
rect 5040 14560 5046 14572
rect 5077 14569 5089 14572
rect 5123 14569 5135 14603
rect 6638 14600 6644 14612
rect 6599 14572 6644 14600
rect 5077 14563 5135 14569
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7929 14603 7987 14609
rect 7929 14600 7941 14603
rect 6748 14572 7941 14600
rect 14 14492 20 14544
rect 72 14532 78 14544
rect 1670 14532 1676 14544
rect 72 14504 1676 14532
rect 72 14492 78 14504
rect 1670 14492 1676 14504
rect 1728 14492 1734 14544
rect 3234 14492 3240 14544
rect 3292 14532 3298 14544
rect 3789 14535 3847 14541
rect 3789 14532 3801 14535
rect 3292 14504 3801 14532
rect 3292 14492 3298 14504
rect 3789 14501 3801 14504
rect 3835 14501 3847 14535
rect 3789 14495 3847 14501
rect 3970 14492 3976 14544
rect 4028 14532 4034 14544
rect 4028 14504 4108 14532
rect 4028 14492 4034 14504
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1673 14359 1731 14365
rect 1688 14328 1716 14359
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2777 14399 2835 14405
rect 2777 14365 2789 14399
rect 2823 14396 2835 14399
rect 3970 14396 3976 14408
rect 2823 14368 3976 14396
rect 2823 14365 2835 14368
rect 2777 14359 2835 14365
rect 3970 14356 3976 14368
rect 4028 14356 4034 14408
rect 3142 14328 3148 14340
rect 1688 14300 3148 14328
rect 3142 14288 3148 14300
rect 3200 14288 3206 14340
rect 4080 14328 4108 14504
rect 5166 14492 5172 14544
rect 5224 14532 5230 14544
rect 6748 14532 6776 14572
rect 7929 14569 7941 14572
rect 7975 14569 7987 14603
rect 7929 14563 7987 14569
rect 8386 14560 8392 14612
rect 8444 14600 8450 14612
rect 8846 14600 8852 14612
rect 8444 14572 8852 14600
rect 8444 14560 8450 14572
rect 8846 14560 8852 14572
rect 8904 14600 8910 14612
rect 11514 14600 11520 14612
rect 8904 14572 11520 14600
rect 8904 14560 8910 14572
rect 11514 14560 11520 14572
rect 11572 14560 11578 14612
rect 11698 14560 11704 14612
rect 11756 14600 11762 14612
rect 11756 14572 13768 14600
rect 11756 14560 11762 14572
rect 9306 14532 9312 14544
rect 5224 14504 6776 14532
rect 7024 14504 9312 14532
rect 5224 14492 5230 14504
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4341 14467 4399 14473
rect 4341 14464 4353 14467
rect 4212 14436 4353 14464
rect 4212 14424 4218 14436
rect 4341 14433 4353 14436
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 5074 14424 5080 14476
rect 5132 14464 5138 14476
rect 5721 14467 5779 14473
rect 5721 14464 5733 14467
rect 5132 14436 5733 14464
rect 5132 14424 5138 14436
rect 5721 14433 5733 14436
rect 5767 14464 5779 14467
rect 6638 14464 6644 14476
rect 5767 14436 6644 14464
rect 5767 14433 5779 14436
rect 5721 14427 5779 14433
rect 6638 14424 6644 14436
rect 6696 14424 6702 14476
rect 7024 14473 7052 14504
rect 9306 14492 9312 14504
rect 9364 14492 9370 14544
rect 11609 14535 11667 14541
rect 11609 14501 11621 14535
rect 11655 14532 11667 14535
rect 11790 14532 11796 14544
rect 11655 14504 11796 14532
rect 11655 14501 11667 14504
rect 11609 14495 11667 14501
rect 11790 14492 11796 14504
rect 11848 14532 11854 14544
rect 12250 14532 12256 14544
rect 11848 14504 12256 14532
rect 11848 14492 11854 14504
rect 12250 14492 12256 14504
rect 12308 14492 12314 14544
rect 13740 14532 13768 14572
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13872 14572 14105 14600
rect 13872 14560 13878 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 16390 14600 16396 14612
rect 14093 14563 14151 14569
rect 14568 14572 16396 14600
rect 14568 14532 14596 14572
rect 16390 14560 16396 14572
rect 16448 14600 16454 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 16448 14572 17141 14600
rect 16448 14560 16454 14572
rect 17129 14569 17141 14572
rect 17175 14569 17187 14603
rect 17129 14563 17187 14569
rect 19245 14603 19303 14609
rect 19245 14569 19257 14603
rect 19291 14600 19303 14603
rect 19702 14600 19708 14612
rect 19291 14572 19708 14600
rect 19291 14569 19303 14572
rect 19245 14563 19303 14569
rect 19702 14560 19708 14572
rect 19760 14560 19766 14612
rect 13740 14504 14596 14532
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14433 7067 14467
rect 7190 14464 7196 14476
rect 7151 14436 7196 14464
rect 7009 14427 7067 14433
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 9674 14424 9680 14476
rect 9732 14464 9738 14476
rect 10226 14464 10232 14476
rect 9732 14436 10232 14464
rect 9732 14424 9738 14436
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 14458 14464 14464 14476
rect 13197 14436 14464 14464
rect 4246 14396 4252 14408
rect 4207 14368 4252 14396
rect 4246 14356 4252 14368
rect 4304 14356 4310 14408
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5534 14396 5540 14408
rect 5491 14368 5540 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 7282 14396 7288 14408
rect 7243 14368 7288 14396
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 10502 14405 10508 14408
rect 10496 14396 10508 14405
rect 7392 14368 10180 14396
rect 10463 14368 10508 14396
rect 4157 14331 4215 14337
rect 4157 14328 4169 14331
rect 4080 14300 4169 14328
rect 4157 14297 4169 14300
rect 4203 14328 4215 14331
rect 4203 14300 4384 14328
rect 4203 14297 4215 14300
rect 4157 14291 4215 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2130 14260 2136 14272
rect 2091 14232 2136 14260
rect 2130 14220 2136 14232
rect 2188 14220 2194 14272
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 2593 14263 2651 14269
rect 2593 14260 2605 14263
rect 2556 14232 2605 14260
rect 2556 14220 2562 14232
rect 2593 14229 2605 14232
rect 2639 14229 2651 14263
rect 2593 14223 2651 14229
rect 3053 14263 3111 14269
rect 3053 14229 3065 14263
rect 3099 14260 3111 14263
rect 3418 14260 3424 14272
rect 3099 14232 3424 14260
rect 3099 14229 3111 14232
rect 3053 14223 3111 14229
rect 3418 14220 3424 14232
rect 3476 14220 3482 14272
rect 4356 14260 4384 14300
rect 5074 14288 5080 14340
rect 5132 14328 5138 14340
rect 7392 14328 7420 14368
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 5132 14300 7420 14328
rect 7484 14300 8953 14328
rect 5132 14288 5138 14300
rect 5537 14263 5595 14269
rect 5537 14260 5549 14263
rect 4356 14232 5549 14260
rect 5537 14229 5549 14232
rect 5583 14229 5595 14263
rect 5537 14223 5595 14229
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14260 6239 14263
rect 6638 14260 6644 14272
rect 6227 14232 6644 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6638 14220 6644 14232
rect 6696 14220 6702 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7484 14260 7512 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 9401 14331 9459 14337
rect 9401 14297 9413 14331
rect 9447 14328 9459 14331
rect 10042 14328 10048 14340
rect 9447 14300 10048 14328
rect 9447 14297 9459 14300
rect 9401 14291 9459 14297
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10152 14328 10180 14368
rect 10496 14359 10508 14368
rect 10502 14356 10508 14359
rect 10560 14356 10566 14408
rect 13197 14396 13225 14436
rect 14458 14424 14464 14436
rect 14516 14424 14522 14476
rect 10612 14368 13225 14396
rect 13265 14399 13323 14405
rect 10612 14328 10640 14368
rect 13265 14365 13277 14399
rect 13311 14396 13323 14399
rect 14918 14396 14924 14408
rect 13311 14368 14924 14396
rect 13311 14365 13323 14368
rect 13265 14359 13323 14365
rect 10152 14300 10640 14328
rect 10962 14288 10968 14340
rect 11020 14328 11026 14340
rect 12998 14331 13056 14337
rect 12998 14328 13010 14331
rect 11020 14300 13010 14328
rect 11020 14288 11026 14300
rect 12998 14297 13010 14300
rect 13044 14297 13056 14331
rect 12998 14291 13056 14297
rect 7650 14260 7656 14272
rect 6788 14232 7512 14260
rect 7611 14232 7656 14260
rect 6788 14220 6794 14232
rect 7650 14220 7656 14232
rect 7708 14220 7714 14272
rect 8294 14260 8300 14272
rect 8255 14232 8300 14260
rect 8294 14220 8300 14232
rect 8352 14220 8358 14272
rect 9674 14260 9680 14272
rect 9635 14232 9680 14260
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 10686 14220 10692 14272
rect 10744 14260 10750 14272
rect 11885 14263 11943 14269
rect 11885 14260 11897 14263
rect 10744 14232 11897 14260
rect 10744 14220 10750 14232
rect 11885 14229 11897 14232
rect 11931 14229 11943 14263
rect 11885 14223 11943 14229
rect 12066 14220 12072 14272
rect 12124 14260 12130 14272
rect 13078 14260 13084 14272
rect 12124 14232 13084 14260
rect 12124 14220 12130 14232
rect 13078 14220 13084 14232
rect 13136 14220 13142 14272
rect 13648 14269 13676 14368
rect 14918 14356 14924 14368
rect 14976 14396 14982 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 14976 14368 15485 14396
rect 14976 14356 14982 14368
rect 15473 14365 15485 14368
rect 15519 14396 15531 14399
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15519 14368 15761 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15749 14359 15807 14365
rect 18785 14399 18843 14405
rect 18785 14365 18797 14399
rect 18831 14396 18843 14399
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 18831 14368 20637 14396
rect 18831 14365 18843 14368
rect 18785 14359 18843 14365
rect 20625 14365 20637 14368
rect 20671 14396 20683 14399
rect 20714 14396 20720 14408
rect 20671 14368 20720 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 20714 14356 20720 14368
rect 20772 14356 20778 14408
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 15102 14288 15108 14340
rect 15160 14328 15166 14340
rect 15206 14331 15264 14337
rect 15206 14328 15218 14331
rect 15160 14300 15218 14328
rect 15160 14288 15166 14300
rect 15206 14297 15218 14300
rect 15252 14297 15264 14331
rect 15206 14291 15264 14297
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 15930 14328 15936 14340
rect 15620 14300 15936 14328
rect 15620 14288 15626 14300
rect 15930 14288 15936 14300
rect 15988 14337 15994 14340
rect 15988 14331 16052 14337
rect 15988 14297 16006 14331
rect 16040 14297 16052 14331
rect 15988 14291 16052 14297
rect 15988 14288 15994 14291
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 18518 14331 18576 14337
rect 18518 14328 18530 14331
rect 16172 14300 18530 14328
rect 16172 14288 16178 14300
rect 18518 14297 18530 14300
rect 18564 14297 18576 14331
rect 18518 14291 18576 14297
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 20380 14331 20438 14337
rect 20380 14328 20392 14331
rect 19484 14300 20392 14328
rect 19484 14288 19490 14300
rect 20380 14297 20392 14300
rect 20426 14328 20438 14331
rect 20530 14328 20536 14340
rect 20426 14300 20536 14328
rect 20426 14297 20438 14300
rect 20380 14291 20438 14297
rect 20530 14288 20536 14300
rect 20588 14288 20594 14340
rect 13633 14263 13691 14269
rect 13633 14229 13645 14263
rect 13679 14260 13691 14263
rect 13814 14260 13820 14272
rect 13679 14232 13820 14260
rect 13679 14229 13691 14232
rect 13633 14223 13691 14229
rect 13814 14220 13820 14232
rect 13872 14220 13878 14272
rect 17402 14260 17408 14272
rect 17363 14232 17408 14260
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 2869 14059 2927 14065
rect 2869 14025 2881 14059
rect 2915 14025 2927 14059
rect 3142 14056 3148 14068
rect 3103 14028 3148 14056
rect 2869 14019 2927 14025
rect 2133 13991 2191 13997
rect 2133 13957 2145 13991
rect 2179 13988 2191 13991
rect 2314 13988 2320 14000
rect 2179 13960 2320 13988
rect 2179 13957 2191 13960
rect 2133 13951 2191 13957
rect 2314 13948 2320 13960
rect 2372 13948 2378 14000
rect 2041 13923 2099 13929
rect 2041 13889 2053 13923
rect 2087 13920 2099 13923
rect 2406 13920 2412 13932
rect 2087 13892 2412 13920
rect 2087 13889 2099 13892
rect 2041 13883 2099 13889
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 2682 13920 2688 13932
rect 2643 13892 2688 13920
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 2884 13920 2912 14019
rect 3142 14016 3148 14028
rect 3200 14016 3206 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4430 14056 4436 14068
rect 4391 14028 4436 14056
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 5074 14056 5080 14068
rect 5035 14028 5080 14056
rect 5074 14016 5080 14028
rect 5132 14016 5138 14068
rect 6825 14059 6883 14065
rect 6825 14025 6837 14059
rect 6871 14056 6883 14059
rect 7006 14056 7012 14068
rect 6871 14028 7012 14056
rect 6871 14025 6883 14028
rect 6825 14019 6883 14025
rect 7006 14016 7012 14028
rect 7064 14056 7070 14068
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 7064 14028 8033 14056
rect 7064 14016 7070 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 8481 14059 8539 14065
rect 8481 14025 8493 14059
rect 8527 14056 8539 14059
rect 8527 14028 10180 14056
rect 8527 14025 8539 14028
rect 8481 14019 8539 14025
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 4341 13991 4399 13997
rect 4341 13988 4353 13991
rect 4120 13960 4353 13988
rect 4120 13948 4126 13960
rect 4341 13957 4353 13960
rect 4387 13957 4399 13991
rect 8496 13988 8524 14019
rect 8846 13988 8852 14000
rect 4341 13951 4399 13957
rect 7300 13960 8524 13988
rect 8807 13960 8852 13988
rect 7300 13944 7328 13960
rect 8846 13948 8852 13960
rect 8904 13948 8910 14000
rect 9484 13991 9542 13997
rect 9484 13957 9496 13991
rect 9530 13988 9542 13991
rect 9582 13988 9588 14000
rect 9530 13960 9588 13988
rect 9530 13957 9542 13960
rect 9484 13951 9542 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 10152 13988 10180 14028
rect 10226 14016 10232 14068
rect 10284 14056 10290 14068
rect 10870 14056 10876 14068
rect 10284 14028 10876 14056
rect 10284 14016 10290 14028
rect 10870 14016 10876 14028
rect 10928 14056 10934 14068
rect 11701 14059 11759 14065
rect 11701 14056 11713 14059
rect 10928 14028 11713 14056
rect 10928 14016 10934 14028
rect 11701 14025 11713 14028
rect 11747 14025 11759 14059
rect 11701 14019 11759 14025
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 15746 14056 15752 14068
rect 14516 14028 15752 14056
rect 14516 14016 14522 14028
rect 15746 14016 15752 14028
rect 15804 14016 15810 14068
rect 15930 14056 15936 14068
rect 15891 14028 15936 14056
rect 15930 14016 15936 14028
rect 15988 14016 15994 14068
rect 18966 14056 18972 14068
rect 18927 14028 18972 14056
rect 18966 14016 18972 14028
rect 19024 14016 19030 14068
rect 19613 14059 19671 14065
rect 19613 14025 19625 14059
rect 19659 14056 19671 14059
rect 20346 14056 20352 14068
rect 19659 14028 20352 14056
rect 19659 14025 19671 14028
rect 19613 14019 19671 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 11882 13988 11888 14000
rect 10152 13960 11888 13988
rect 11882 13948 11888 13960
rect 11940 13948 11946 14000
rect 13814 13948 13820 14000
rect 13872 13988 13878 14000
rect 17862 13997 17868 14000
rect 17856 13988 17868 13997
rect 13872 13960 16068 13988
rect 17775 13960 17868 13988
rect 13872 13948 13878 13960
rect 3329 13923 3387 13929
rect 3329 13920 3341 13923
rect 2884 13892 3341 13920
rect 3329 13889 3341 13892
rect 3375 13889 3387 13923
rect 3329 13883 3387 13889
rect 5350 13880 5356 13932
rect 5408 13920 5414 13932
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 5408 13892 5549 13920
rect 5408 13880 5414 13892
rect 5537 13889 5549 13892
rect 5583 13920 5595 13923
rect 5583 13892 6868 13920
rect 5583 13889 5595 13892
rect 5537 13883 5595 13889
rect 2130 13812 2136 13864
rect 2188 13852 2194 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2188 13824 2237 13852
rect 2188 13812 2194 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 2225 13815 2283 13821
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13852 4675 13855
rect 5074 13852 5080 13864
rect 4663 13824 5080 13852
rect 4663 13821 4675 13824
rect 4617 13815 4675 13821
rect 5074 13812 5080 13824
rect 5132 13812 5138 13864
rect 5810 13852 5816 13864
rect 5771 13824 5816 13852
rect 5810 13812 5816 13824
rect 5868 13812 5874 13864
rect 6546 13812 6552 13864
rect 6604 13852 6610 13864
rect 6730 13852 6736 13864
rect 6604 13824 6736 13852
rect 6604 13812 6610 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 5442 13744 5448 13796
rect 5500 13784 5506 13796
rect 6638 13784 6644 13796
rect 5500 13756 6644 13784
rect 5500 13744 5506 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 1670 13716 1676 13728
rect 1631 13688 1676 13716
rect 1670 13676 1676 13688
rect 1728 13676 1734 13728
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 3605 13719 3663 13725
rect 3605 13716 3617 13719
rect 3200 13688 3617 13716
rect 3200 13676 3206 13688
rect 3605 13685 3617 13688
rect 3651 13685 3663 13719
rect 3605 13679 3663 13685
rect 5718 13676 5724 13728
rect 5776 13716 5782 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 5776 13688 6469 13716
rect 5776 13676 5782 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6840 13716 6868 13892
rect 7116 13916 7328 13944
rect 9214 13920 9220 13932
rect 7116 13861 7144 13916
rect 9175 13892 9220 13920
rect 9214 13880 9220 13892
rect 9272 13880 9278 13932
rect 10778 13920 10784 13932
rect 9324 13892 10784 13920
rect 6917 13855 6975 13861
rect 6917 13821 6929 13855
rect 6963 13852 6975 13855
rect 7101 13855 7159 13861
rect 6963 13824 7052 13852
rect 6963 13821 6975 13824
rect 6917 13815 6975 13821
rect 7024 13784 7052 13824
rect 7101 13821 7113 13855
rect 7147 13821 7159 13855
rect 7101 13815 7159 13821
rect 7466 13812 7472 13864
rect 7524 13852 7530 13864
rect 9324 13852 9352 13892
rect 10778 13880 10784 13892
rect 10836 13880 10842 13932
rect 12161 13923 12219 13929
rect 12161 13889 12173 13923
rect 12207 13920 12219 13923
rect 12250 13920 12256 13932
rect 12207 13892 12256 13920
rect 12207 13889 12219 13892
rect 12161 13883 12219 13889
rect 12250 13880 12256 13892
rect 12308 13880 12314 13932
rect 12342 13880 12348 13932
rect 12400 13920 12406 13932
rect 13153 13923 13211 13929
rect 13153 13920 13165 13923
rect 12400 13892 13165 13920
rect 12400 13880 12406 13892
rect 13153 13889 13165 13892
rect 13199 13889 13211 13923
rect 13153 13883 13211 13889
rect 13722 13880 13728 13932
rect 13780 13920 13786 13932
rect 14568 13929 14596 13960
rect 14553 13923 14611 13929
rect 13780 13892 14320 13920
rect 13780 13880 13786 13892
rect 10962 13852 10968 13864
rect 7524 13824 9352 13852
rect 10612 13824 10968 13852
rect 7524 13812 7530 13824
rect 7374 13784 7380 13796
rect 7024 13756 7380 13784
rect 7374 13744 7380 13756
rect 7432 13784 7438 13796
rect 10612 13793 10640 13824
rect 10962 13812 10968 13824
rect 11020 13812 11026 13864
rect 12897 13855 12955 13861
rect 12897 13852 12909 13855
rect 12406 13824 12909 13852
rect 7745 13787 7803 13793
rect 7745 13784 7757 13787
rect 7432 13756 7757 13784
rect 7432 13744 7438 13756
rect 7745 13753 7757 13756
rect 7791 13784 7803 13787
rect 10597 13787 10655 13793
rect 7791 13756 8248 13784
rect 7791 13753 7803 13756
rect 7745 13747 7803 13753
rect 7466 13716 7472 13728
rect 6840 13688 7472 13716
rect 6457 13679 6515 13685
rect 7466 13676 7472 13688
rect 7524 13676 7530 13728
rect 8220 13716 8248 13756
rect 10597 13753 10609 13787
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 10870 13744 10876 13796
rect 10928 13784 10934 13796
rect 12406 13784 12434 13824
rect 12897 13821 12909 13824
rect 12943 13821 12955 13855
rect 12897 13815 12955 13821
rect 14292 13852 14320 13892
rect 14553 13889 14565 13923
rect 14599 13889 14611 13923
rect 14809 13923 14867 13929
rect 14809 13920 14821 13923
rect 14553 13883 14611 13889
rect 14660 13892 14821 13920
rect 14660 13852 14688 13892
rect 14809 13889 14821 13892
rect 14855 13889 14867 13923
rect 14809 13883 14867 13889
rect 14292 13824 14688 13852
rect 14292 13793 14320 13824
rect 10928 13756 12434 13784
rect 14277 13787 14335 13793
rect 10928 13744 10934 13756
rect 14277 13753 14289 13787
rect 14323 13753 14335 13787
rect 14277 13747 14335 13753
rect 16040 13728 16068 13960
rect 17856 13951 17868 13960
rect 17920 13988 17926 14000
rect 19978 13988 19984 14000
rect 17920 13960 19984 13988
rect 17862 13948 17868 13951
rect 17920 13948 17926 13960
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13889 19487 13923
rect 19429 13883 19487 13889
rect 16945 13855 17003 13861
rect 16945 13821 16957 13855
rect 16991 13852 17003 13855
rect 17313 13855 17371 13861
rect 17313 13852 17325 13855
rect 16991 13824 17325 13852
rect 16991 13821 17003 13824
rect 16945 13815 17003 13821
rect 17313 13821 17325 13824
rect 17359 13852 17371 13855
rect 17586 13852 17592 13864
rect 17359 13824 17592 13852
rect 17359 13821 17371 13824
rect 17313 13815 17371 13821
rect 12066 13716 12072 13728
rect 8220 13688 12072 13716
rect 12066 13676 12072 13688
rect 12124 13676 12130 13728
rect 12434 13716 12440 13728
rect 12395 13688 12440 13716
rect 12434 13676 12440 13688
rect 12492 13676 12498 13728
rect 16022 13676 16028 13728
rect 16080 13716 16086 13728
rect 16209 13719 16267 13725
rect 16209 13716 16221 13719
rect 16080 13688 16221 13716
rect 16080 13676 16086 13688
rect 16209 13685 16221 13688
rect 16255 13716 16267 13719
rect 16960 13716 16988 13815
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 19444 13852 19472 13883
rect 19260 13824 19472 13852
rect 19260 13784 19288 13824
rect 19904 13793 19932 13960
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20714 13948 20720 14000
rect 20772 13988 20778 14000
rect 20772 13960 21312 13988
rect 20772 13948 20778 13960
rect 21284 13929 21312 13960
rect 21002 13923 21060 13929
rect 21002 13920 21014 13923
rect 19996 13892 21014 13920
rect 19996 13864 20024 13892
rect 21002 13889 21014 13892
rect 21048 13889 21060 13923
rect 21002 13883 21060 13889
rect 21269 13923 21327 13929
rect 21269 13889 21281 13923
rect 21315 13889 21327 13923
rect 21269 13883 21327 13889
rect 19978 13812 19984 13864
rect 20036 13812 20042 13864
rect 18524 13756 19288 13784
rect 19889 13787 19947 13793
rect 18524 13728 18552 13756
rect 19889 13753 19901 13787
rect 19935 13753 19947 13787
rect 19889 13747 19947 13753
rect 16255 13688 16988 13716
rect 16255 13685 16267 13688
rect 16209 13679 16267 13685
rect 18506 13676 18512 13728
rect 18564 13676 18570 13728
rect 20162 13676 20168 13728
rect 20220 13716 20226 13728
rect 20346 13716 20352 13728
rect 20220 13688 20352 13716
rect 20220 13676 20226 13688
rect 20346 13676 20352 13688
rect 20404 13676 20410 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2409 13515 2467 13521
rect 2409 13481 2421 13515
rect 2455 13512 2467 13515
rect 2590 13512 2596 13524
rect 2455 13484 2596 13512
rect 2455 13481 2467 13484
rect 2409 13475 2467 13481
rect 2590 13472 2596 13484
rect 2648 13472 2654 13524
rect 3421 13515 3479 13521
rect 3421 13481 3433 13515
rect 3467 13512 3479 13515
rect 4798 13512 4804 13524
rect 3467 13484 4804 13512
rect 3467 13481 3479 13484
rect 3421 13475 3479 13481
rect 4798 13472 4804 13484
rect 4856 13472 4862 13524
rect 5902 13472 5908 13524
rect 5960 13512 5966 13524
rect 6457 13515 6515 13521
rect 6457 13512 6469 13515
rect 5960 13484 6469 13512
rect 5960 13472 5966 13484
rect 6457 13481 6469 13484
rect 6503 13481 6515 13515
rect 6457 13475 6515 13481
rect 6638 13472 6644 13524
rect 6696 13512 6702 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 6696 13484 9045 13512
rect 6696 13472 6702 13484
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 2280 13416 3801 13444
rect 2280 13404 2286 13416
rect 3789 13413 3801 13416
rect 3835 13413 3847 13447
rect 3789 13407 3847 13413
rect 6181 13447 6239 13453
rect 6181 13413 6193 13447
rect 6227 13444 6239 13447
rect 7006 13444 7012 13456
rect 6227 13416 7012 13444
rect 6227 13413 6239 13416
rect 6181 13407 6239 13413
rect 7006 13404 7012 13416
rect 7064 13404 7070 13456
rect 1854 13376 1860 13388
rect 1815 13348 1860 13376
rect 1854 13336 1860 13348
rect 1912 13336 1918 13388
rect 4430 13376 4436 13388
rect 4391 13348 4436 13376
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 7116 13385 7144 13484
rect 9033 13481 9045 13484
rect 9079 13512 9091 13515
rect 9079 13484 10364 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 7742 13404 7748 13456
rect 7800 13444 7806 13456
rect 8481 13447 8539 13453
rect 8481 13444 8493 13447
rect 7800 13416 8493 13444
rect 7800 13404 7806 13416
rect 8481 13413 8493 13416
rect 8527 13413 8539 13447
rect 10336 13444 10364 13484
rect 10502 13472 10508 13524
rect 10560 13512 10566 13524
rect 10781 13515 10839 13521
rect 10781 13512 10793 13515
rect 10560 13484 10793 13512
rect 10560 13472 10566 13484
rect 10781 13481 10793 13484
rect 10827 13481 10839 13515
rect 10781 13475 10839 13481
rect 10870 13472 10876 13524
rect 10928 13512 10934 13524
rect 11057 13515 11115 13521
rect 11057 13512 11069 13515
rect 10928 13484 11069 13512
rect 10928 13472 10934 13484
rect 11057 13481 11069 13484
rect 11103 13481 11115 13515
rect 11057 13475 11115 13481
rect 11882 13472 11888 13524
rect 11940 13512 11946 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 11940 13484 12541 13512
rect 11940 13472 11946 13484
rect 12529 13481 12541 13484
rect 12575 13512 12587 13515
rect 12802 13512 12808 13524
rect 12575 13484 12808 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13170 13472 13176 13524
rect 13228 13512 13234 13524
rect 16942 13512 16948 13524
rect 13228 13484 16948 13512
rect 13228 13472 13234 13484
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17034 13472 17040 13524
rect 17092 13512 17098 13524
rect 17405 13515 17463 13521
rect 17405 13512 17417 13515
rect 17092 13484 17417 13512
rect 17092 13472 17098 13484
rect 17405 13481 17417 13484
rect 17451 13481 17463 13515
rect 17405 13475 17463 13481
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 18049 13515 18107 13521
rect 18049 13512 18061 13515
rect 17552 13484 18061 13512
rect 17552 13472 17558 13484
rect 18049 13481 18061 13484
rect 18095 13512 18107 13515
rect 19978 13512 19984 13524
rect 18095 13484 19984 13512
rect 18095 13481 18107 13484
rect 18049 13475 18107 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 15194 13444 15200 13456
rect 10336 13416 15200 13444
rect 8481 13407 8539 13413
rect 15194 13404 15200 13416
rect 15252 13404 15258 13456
rect 5629 13379 5687 13385
rect 5629 13345 5641 13379
rect 5675 13376 5687 13379
rect 7101 13379 7159 13385
rect 5675 13348 7052 13376
rect 5675 13345 5687 13348
rect 5629 13339 5687 13345
rect 1670 13268 1676 13320
rect 1728 13308 1734 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 1728 13280 2053 13308
rect 1728 13268 1734 13280
rect 2041 13277 2053 13280
rect 2087 13277 2099 13311
rect 2682 13308 2688 13320
rect 2643 13280 2688 13308
rect 2041 13271 2099 13277
rect 2682 13268 2688 13280
rect 2740 13268 2746 13320
rect 3142 13268 3148 13320
rect 3200 13308 3206 13320
rect 3237 13311 3295 13317
rect 3237 13308 3249 13311
rect 3200 13280 3249 13308
rect 3200 13268 3206 13280
rect 3237 13277 3249 13280
rect 3283 13277 3295 13311
rect 5810 13308 5816 13320
rect 5771 13280 5816 13308
rect 3237 13271 3295 13277
rect 5810 13268 5816 13280
rect 5868 13268 5874 13320
rect 6822 13268 6828 13320
rect 6880 13308 6886 13320
rect 6917 13311 6975 13317
rect 6917 13308 6929 13311
rect 6880 13280 6929 13308
rect 6880 13268 6886 13280
rect 6917 13277 6929 13280
rect 6963 13277 6975 13311
rect 7024 13308 7052 13348
rect 7101 13345 7113 13379
rect 7147 13345 7159 13379
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7101 13339 7159 13345
rect 7668 13348 8125 13376
rect 7668 13308 7696 13348
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 7024 13280 7696 13308
rect 6917 13271 6975 13277
rect 7742 13268 7748 13320
rect 7800 13308 7806 13320
rect 7929 13311 7987 13317
rect 7929 13308 7941 13311
rect 7800 13280 7941 13308
rect 7800 13268 7806 13280
rect 7929 13277 7941 13280
rect 7975 13308 7987 13311
rect 8018 13308 8024 13320
rect 7975 13280 8024 13308
rect 7975 13277 7987 13280
rect 7929 13271 7987 13277
rect 8018 13268 8024 13280
rect 8076 13268 8082 13320
rect 8128 13308 8156 13339
rect 9214 13336 9220 13388
rect 9272 13376 9278 13388
rect 9401 13379 9459 13385
rect 9401 13376 9413 13379
rect 9272 13348 9413 13376
rect 9272 13336 9278 13348
rect 9401 13345 9413 13348
rect 9447 13345 9459 13379
rect 9401 13339 9459 13345
rect 13357 13379 13415 13385
rect 13357 13345 13369 13379
rect 13403 13376 13415 13379
rect 15654 13376 15660 13388
rect 13403 13348 15660 13376
rect 13403 13345 13415 13348
rect 13357 13339 13415 13345
rect 15654 13336 15660 13348
rect 15712 13336 15718 13388
rect 15749 13379 15807 13385
rect 15749 13345 15761 13379
rect 15795 13376 15807 13379
rect 15795 13348 16160 13376
rect 15795 13345 15807 13348
rect 15749 13339 15807 13345
rect 16022 13308 16028 13320
rect 8128 13280 9976 13308
rect 5169 13243 5227 13249
rect 5169 13240 5181 13243
rect 1688 13212 5181 13240
rect 1688 13184 1716 13212
rect 5169 13209 5181 13212
rect 5215 13240 5227 13243
rect 5721 13243 5779 13249
rect 5721 13240 5733 13243
rect 5215 13212 5733 13240
rect 5215 13209 5227 13212
rect 5169 13203 5227 13209
rect 5721 13209 5733 13212
rect 5767 13240 5779 13243
rect 8754 13240 8760 13252
rect 5767 13212 8760 13240
rect 5767 13209 5779 13212
rect 5721 13203 5779 13209
rect 8754 13200 8760 13212
rect 8812 13200 8818 13252
rect 9657 13243 9715 13249
rect 9657 13209 9669 13243
rect 9703 13209 9715 13243
rect 9948 13240 9976 13280
rect 12176 13280 12434 13308
rect 10226 13240 10232 13252
rect 9948 13212 10232 13240
rect 9657 13203 9715 13209
rect 1670 13132 1676 13184
rect 1728 13132 1734 13184
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 2866 13172 2872 13184
rect 2827 13144 2872 13172
rect 2866 13132 2872 13144
rect 2924 13132 2930 13184
rect 4154 13172 4160 13184
rect 4115 13144 4160 13172
rect 4154 13132 4160 13144
rect 4212 13132 4218 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4304 13144 4349 13172
rect 4304 13132 4310 13144
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 6730 13172 6736 13184
rect 5868 13144 6736 13172
rect 5868 13132 5874 13144
rect 6730 13132 6736 13144
rect 6788 13132 6794 13184
rect 6825 13175 6883 13181
rect 6825 13141 6837 13175
rect 6871 13172 6883 13175
rect 7006 13172 7012 13184
rect 6871 13144 7012 13172
rect 6871 13141 6883 13144
rect 6825 13135 6883 13141
rect 7006 13132 7012 13144
rect 7064 13132 7070 13184
rect 7466 13172 7472 13184
rect 7427 13144 7472 13172
rect 7466 13132 7472 13144
rect 7524 13132 7530 13184
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 7837 13175 7895 13181
rect 7837 13172 7849 13175
rect 7800 13144 7849 13172
rect 7800 13132 7806 13144
rect 7837 13141 7849 13144
rect 7883 13141 7895 13175
rect 9683 13172 9711 13203
rect 10226 13200 10232 13212
rect 10284 13200 10290 13252
rect 12176 13249 12204 13280
rect 12406 13252 12434 13280
rect 15304 13280 16028 13308
rect 11517 13243 11575 13249
rect 11517 13209 11529 13243
rect 11563 13240 11575 13243
rect 12161 13243 12219 13249
rect 12161 13240 12173 13243
rect 11563 13212 12173 13240
rect 11563 13209 11575 13212
rect 11517 13203 11575 13209
rect 12161 13209 12173 13212
rect 12207 13209 12219 13243
rect 12406 13240 12440 13252
rect 12347 13212 12440 13240
rect 12161 13203 12219 13209
rect 12434 13200 12440 13212
rect 12492 13240 12498 13252
rect 13078 13240 13084 13252
rect 12492 13212 13084 13240
rect 12492 13200 12498 13212
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 9766 13172 9772 13184
rect 9683 13144 9772 13172
rect 7837 13135 7895 13141
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11606 13172 11612 13184
rect 11020 13144 11612 13172
rect 11020 13132 11026 13144
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11790 13172 11796 13184
rect 11751 13144 11796 13172
rect 11790 13132 11796 13144
rect 11848 13132 11854 13184
rect 12986 13172 12992 13184
rect 12947 13144 12992 13172
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 13722 13172 13728 13184
rect 13683 13144 13728 13172
rect 13722 13132 13728 13144
rect 13780 13172 13786 13184
rect 15304 13181 15332 13280
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16132 13308 16160 13348
rect 16132 13280 17540 13308
rect 16292 13243 16350 13249
rect 16292 13209 16304 13243
rect 16338 13240 16350 13243
rect 16390 13240 16396 13252
rect 16338 13212 16396 13240
rect 16338 13209 16350 13212
rect 16292 13203 16350 13209
rect 16390 13200 16396 13212
rect 16448 13200 16454 13252
rect 14369 13175 14427 13181
rect 14369 13172 14381 13175
rect 13780 13144 14381 13172
rect 13780 13132 13786 13144
rect 14369 13141 14381 13144
rect 14415 13172 14427 13175
rect 14921 13175 14979 13181
rect 14921 13172 14933 13175
rect 14415 13144 14933 13172
rect 14415 13141 14427 13144
rect 14369 13135 14427 13141
rect 14921 13141 14933 13144
rect 14967 13172 14979 13175
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 14967 13144 15301 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 17512 13172 17540 13280
rect 17586 13268 17592 13320
rect 17644 13308 17650 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17644 13280 17785 13308
rect 17644 13268 17650 13280
rect 17773 13277 17785 13280
rect 17819 13308 17831 13311
rect 18877 13311 18935 13317
rect 18877 13308 18889 13311
rect 17819 13280 18889 13308
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 18877 13277 18889 13280
rect 18923 13308 18935 13311
rect 20714 13308 20720 13320
rect 18923 13280 20720 13308
rect 18923 13277 18935 13280
rect 18877 13271 18935 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 21085 13311 21143 13317
rect 21085 13277 21097 13311
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 18414 13240 18420 13252
rect 18375 13212 18420 13240
rect 18414 13200 18420 13212
rect 18472 13200 18478 13252
rect 20472 13243 20530 13249
rect 20472 13209 20484 13243
rect 20518 13240 20530 13243
rect 20990 13240 20996 13252
rect 20518 13212 20996 13240
rect 20518 13209 20530 13212
rect 20472 13203 20530 13209
rect 20990 13200 20996 13212
rect 21048 13200 21054 13252
rect 18322 13172 18328 13184
rect 17512 13144 18328 13172
rect 15289 13135 15347 13141
rect 18322 13132 18328 13144
rect 18380 13132 18386 13184
rect 19334 13172 19340 13184
rect 19295 13144 19340 13172
rect 19334 13132 19340 13144
rect 19392 13132 19398 13184
rect 19702 13132 19708 13184
rect 19760 13172 19766 13184
rect 21100 13172 21128 13271
rect 19760 13144 21128 13172
rect 19760 13132 19766 13144
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 2682 12968 2688 12980
rect 2643 12940 2688 12968
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 4246 12928 4252 12980
rect 4304 12968 4310 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4304 12940 5273 12968
rect 4304 12928 4310 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5261 12931 5319 12937
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7009 12971 7067 12977
rect 7009 12937 7021 12971
rect 7055 12968 7067 12971
rect 7190 12968 7196 12980
rect 7055 12940 7196 12968
rect 7055 12937 7067 12940
rect 7009 12931 7067 12937
rect 7190 12928 7196 12940
rect 7248 12968 7254 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7248 12940 7665 12968
rect 7248 12928 7254 12940
rect 7653 12937 7665 12940
rect 7699 12968 7711 12971
rect 8478 12968 8484 12980
rect 7699 12940 8484 12968
rect 7699 12937 7711 12940
rect 7653 12931 7711 12937
rect 8478 12928 8484 12940
rect 8536 12968 8542 12980
rect 8665 12971 8723 12977
rect 8665 12968 8677 12971
rect 8536 12940 8677 12968
rect 8536 12928 8542 12940
rect 8665 12937 8677 12940
rect 8711 12937 8723 12971
rect 9217 12971 9275 12977
rect 9217 12968 9229 12971
rect 8665 12931 8723 12937
rect 8772 12940 9229 12968
rect 4062 12900 4068 12912
rect 3620 12872 4068 12900
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2038 12832 2044 12844
rect 1995 12804 2044 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2038 12792 2044 12804
rect 2096 12792 2102 12844
rect 2498 12832 2504 12844
rect 2459 12804 2504 12832
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3620 12832 3648 12872
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 8202 12860 8208 12912
rect 8260 12900 8266 12912
rect 8772 12900 8800 12940
rect 9217 12937 9229 12940
rect 9263 12968 9275 12971
rect 10870 12968 10876 12980
rect 9263 12940 10548 12968
rect 10831 12940 10876 12968
rect 9263 12937 9275 12940
rect 9217 12931 9275 12937
rect 8260 12872 8800 12900
rect 8260 12860 8266 12872
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 10226 12900 10232 12912
rect 9916 12872 10232 12900
rect 9916 12860 9922 12872
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10318 12860 10324 12912
rect 10376 12909 10382 12912
rect 10376 12900 10388 12909
rect 10376 12872 10421 12900
rect 10376 12863 10388 12872
rect 10376 12860 10382 12863
rect 3528 12804 3648 12832
rect 3697 12835 3755 12841
rect 2222 12764 2228 12776
rect 2183 12736 2228 12764
rect 2222 12724 2228 12736
rect 2280 12764 2286 12776
rect 3528 12773 3556 12804
rect 3697 12801 3709 12835
rect 3743 12832 3755 12835
rect 4614 12832 4620 12844
rect 3743 12804 4620 12832
rect 3743 12801 3755 12804
rect 3697 12795 3755 12801
rect 4614 12792 4620 12804
rect 4672 12792 4678 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12832 5687 12835
rect 6638 12832 6644 12844
rect 5675 12804 6644 12832
rect 5675 12801 5687 12804
rect 5629 12795 5687 12801
rect 6638 12792 6644 12804
rect 6696 12792 6702 12844
rect 8478 12792 8484 12844
rect 8536 12832 8542 12844
rect 9490 12832 9496 12844
rect 8536 12804 9496 12832
rect 8536 12792 8542 12804
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 2961 12767 3019 12773
rect 2961 12764 2973 12767
rect 2280 12736 2973 12764
rect 2280 12724 2286 12736
rect 2961 12733 2973 12736
rect 3007 12733 3019 12767
rect 2961 12727 3019 12733
rect 3513 12767 3571 12773
rect 3513 12733 3525 12767
rect 3559 12733 3571 12767
rect 3513 12727 3571 12733
rect 3605 12767 3663 12773
rect 3605 12733 3617 12767
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3620 12696 3648 12727
rect 3970 12724 3976 12776
rect 4028 12764 4034 12776
rect 4341 12767 4399 12773
rect 4341 12764 4353 12767
rect 4028 12736 4353 12764
rect 4028 12724 4034 12736
rect 4341 12733 4353 12736
rect 4387 12733 4399 12767
rect 5902 12764 5908 12776
rect 5863 12736 5908 12764
rect 4341 12727 4399 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 6546 12724 6552 12776
rect 6604 12764 6610 12776
rect 7742 12764 7748 12776
rect 6604 12736 7420 12764
rect 7703 12736 7748 12764
rect 6604 12724 6610 12736
rect 3620 12668 4844 12696
rect 4816 12640 4844 12668
rect 5994 12656 6000 12708
rect 6052 12696 6058 12708
rect 7285 12699 7343 12705
rect 7285 12696 7297 12699
rect 6052 12668 7297 12696
rect 6052 12656 6058 12668
rect 7285 12665 7297 12668
rect 7331 12665 7343 12699
rect 7392 12696 7420 12736
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7837 12767 7895 12773
rect 7837 12733 7849 12767
rect 7883 12733 7895 12767
rect 10520 12764 10548 12940
rect 10870 12928 10876 12940
rect 10928 12968 10934 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 10928 12940 11529 12968
rect 10928 12928 10934 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 15102 12968 15108 12980
rect 11517 12931 11575 12937
rect 13096 12940 15108 12968
rect 10597 12835 10655 12841
rect 10597 12801 10609 12835
rect 10643 12832 10655 12835
rect 10888 12832 10916 12928
rect 11054 12860 11060 12912
rect 11112 12900 11118 12912
rect 11698 12900 11704 12912
rect 11112 12872 11704 12900
rect 11112 12860 11118 12872
rect 11698 12860 11704 12872
rect 11756 12900 11762 12912
rect 11885 12903 11943 12909
rect 11885 12900 11897 12903
rect 11756 12872 11897 12900
rect 11756 12860 11762 12872
rect 11885 12869 11897 12872
rect 11931 12869 11943 12903
rect 13096 12900 13124 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 16206 12968 16212 12980
rect 16167 12940 16212 12968
rect 16206 12928 16212 12940
rect 16264 12928 16270 12980
rect 17221 12971 17279 12977
rect 17221 12937 17233 12971
rect 17267 12968 17279 12971
rect 20165 12971 20223 12977
rect 17267 12940 20024 12968
rect 17267 12937 17279 12940
rect 17221 12931 17279 12937
rect 11885 12863 11943 12869
rect 11992 12872 13124 12900
rect 10643 12804 10916 12832
rect 10643 12801 10655 12804
rect 10597 12795 10655 12801
rect 11992 12764 12020 12872
rect 13170 12860 13176 12912
rect 13228 12900 13234 12912
rect 15206 12903 15264 12909
rect 15206 12900 15218 12903
rect 13228 12872 15218 12900
rect 13228 12860 13234 12872
rect 15206 12869 15218 12872
rect 15252 12869 15264 12903
rect 15838 12900 15844 12912
rect 15206 12863 15264 12869
rect 15304 12872 15844 12900
rect 13469 12835 13527 12841
rect 13469 12801 13481 12835
rect 13515 12832 13527 12835
rect 14458 12832 14464 12844
rect 13515 12804 14464 12832
rect 13515 12801 13527 12804
rect 13469 12795 13527 12801
rect 14458 12792 14464 12804
rect 14516 12792 14522 12844
rect 14918 12792 14924 12844
rect 14976 12832 14982 12844
rect 15304 12832 15332 12872
rect 15838 12860 15844 12872
rect 15896 12900 15902 12912
rect 19334 12900 19340 12912
rect 15896 12872 19340 12900
rect 15896 12860 15902 12872
rect 19334 12860 19340 12872
rect 19392 12860 19398 12912
rect 19996 12900 20024 12940
rect 20165 12937 20177 12971
rect 20211 12968 20223 12971
rect 20530 12968 20536 12980
rect 20211 12940 20536 12968
rect 20211 12937 20223 12940
rect 20165 12931 20223 12937
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 19996 12872 20576 12900
rect 14976 12804 15332 12832
rect 14976 12792 14982 12804
rect 15654 12792 15660 12844
rect 15712 12832 15718 12844
rect 16390 12832 16396 12844
rect 15712 12804 16396 12832
rect 15712 12792 15718 12804
rect 16390 12792 16396 12804
rect 16448 12792 16454 12844
rect 17494 12792 17500 12844
rect 17552 12832 17558 12844
rect 18121 12835 18179 12841
rect 18121 12832 18133 12835
rect 17552 12804 18133 12832
rect 17552 12792 17558 12804
rect 18121 12801 18133 12804
rect 18167 12832 18179 12835
rect 18874 12832 18880 12844
rect 18167 12804 18880 12832
rect 18167 12801 18179 12804
rect 18121 12795 18179 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 19705 12835 19763 12841
rect 19705 12801 19717 12835
rect 19751 12832 19763 12835
rect 19794 12832 19800 12844
rect 19751 12804 19800 12832
rect 19751 12801 19763 12804
rect 19705 12795 19763 12801
rect 19794 12792 19800 12804
rect 19852 12792 19858 12844
rect 19886 12792 19892 12844
rect 19944 12832 19950 12844
rect 19981 12835 20039 12841
rect 19981 12832 19993 12835
rect 19944 12804 19993 12832
rect 19944 12792 19950 12804
rect 19981 12801 19993 12804
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20548 12776 20576 12872
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21450 12832 21456 12844
rect 20855 12804 21456 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21450 12792 21456 12804
rect 21508 12792 21514 12844
rect 13722 12764 13728 12776
rect 10520 12736 12020 12764
rect 13683 12736 13728 12764
rect 7837 12727 7895 12733
rect 7852 12696 7880 12727
rect 13722 12724 13728 12736
rect 13780 12724 13786 12776
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 16853 12767 16911 12773
rect 16853 12764 16865 12767
rect 15519 12736 16865 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 7392 12668 7880 12696
rect 7285 12659 7343 12665
rect 10594 12656 10600 12708
rect 10652 12696 10658 12708
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 10652 12668 12357 12696
rect 10652 12656 10658 12668
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 12345 12659 12403 12665
rect 13740 12668 14228 12696
rect 4065 12631 4123 12637
rect 4065 12597 4077 12631
rect 4111 12628 4123 12631
rect 4246 12628 4252 12640
rect 4111 12600 4252 12628
rect 4111 12597 4123 12600
rect 4065 12591 4123 12597
rect 4246 12588 4252 12600
rect 4304 12588 4310 12640
rect 4798 12628 4804 12640
rect 4759 12600 4804 12628
rect 4798 12588 4804 12600
rect 4856 12588 4862 12640
rect 4890 12588 4896 12640
rect 4948 12628 4954 12640
rect 6365 12631 6423 12637
rect 6365 12628 6377 12631
rect 4948 12600 6377 12628
rect 4948 12588 4954 12600
rect 6365 12597 6377 12600
rect 6411 12597 6423 12631
rect 8294 12628 8300 12640
rect 8255 12600 8300 12628
rect 6365 12591 6423 12597
rect 8294 12588 8300 12600
rect 8352 12588 8358 12640
rect 8754 12588 8760 12640
rect 8812 12628 8818 12640
rect 13740 12628 13768 12668
rect 8812 12600 13768 12628
rect 8812 12588 8818 12600
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14093 12631 14151 12637
rect 14093 12628 14105 12631
rect 13872 12600 14105 12628
rect 13872 12588 13878 12600
rect 14093 12597 14105 12600
rect 14139 12597 14151 12631
rect 14200 12628 14228 12668
rect 15672 12640 15700 12736
rect 16853 12733 16865 12736
rect 16899 12764 16911 12767
rect 17865 12767 17923 12773
rect 17865 12764 17877 12767
rect 16899 12736 17877 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17865 12733 17877 12736
rect 17911 12733 17923 12767
rect 20530 12764 20536 12776
rect 20491 12736 20536 12764
rect 17865 12727 17923 12733
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 19521 12699 19579 12705
rect 19521 12665 19533 12699
rect 19567 12696 19579 12699
rect 20070 12696 20076 12708
rect 19567 12668 20076 12696
rect 19567 12665 19579 12668
rect 19521 12659 19579 12665
rect 20070 12656 20076 12668
rect 20128 12656 20134 12708
rect 14826 12628 14832 12640
rect 14200 12600 14832 12628
rect 14093 12591 14151 12597
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 15654 12588 15660 12640
rect 15712 12628 15718 12640
rect 15749 12631 15807 12637
rect 15749 12628 15761 12631
rect 15712 12600 15761 12628
rect 15712 12588 15718 12600
rect 15749 12597 15761 12600
rect 15795 12597 15807 12631
rect 15749 12591 15807 12597
rect 17589 12631 17647 12637
rect 17589 12597 17601 12631
rect 17635 12628 17647 12631
rect 18046 12628 18052 12640
rect 17635 12600 18052 12628
rect 17635 12597 17647 12600
rect 17589 12591 17647 12597
rect 18046 12588 18052 12600
rect 18104 12588 18110 12640
rect 18138 12588 18144 12640
rect 18196 12628 18202 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 18196 12600 19257 12628
rect 18196 12588 18202 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19245 12591 19303 12597
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 3878 12424 3884 12436
rect 3839 12396 3884 12424
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 5534 12384 5540 12436
rect 5592 12384 5598 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 6086 12424 6092 12436
rect 5868 12396 6092 12424
rect 5868 12384 5874 12396
rect 6086 12384 6092 12396
rect 6144 12384 6150 12436
rect 6822 12384 6828 12436
rect 6880 12424 6886 12436
rect 6917 12427 6975 12433
rect 6917 12424 6929 12427
rect 6880 12396 6929 12424
rect 6880 12384 6886 12396
rect 6917 12393 6929 12396
rect 6963 12393 6975 12427
rect 6917 12387 6975 12393
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8481 12427 8539 12433
rect 8481 12424 8493 12427
rect 8076 12396 8493 12424
rect 8076 12384 8082 12396
rect 8481 12393 8493 12396
rect 8527 12424 8539 12427
rect 8938 12424 8944 12436
rect 8527 12396 8944 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 8938 12384 8944 12396
rect 8996 12384 9002 12436
rect 9214 12424 9220 12436
rect 9175 12396 9220 12424
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 11514 12384 11520 12436
rect 11572 12424 11578 12436
rect 12253 12427 12311 12433
rect 12253 12424 12265 12427
rect 11572 12396 12265 12424
rect 11572 12384 11578 12396
rect 12253 12393 12265 12396
rect 12299 12393 12311 12427
rect 12253 12387 12311 12393
rect 12618 12384 12624 12436
rect 12676 12424 12682 12436
rect 13630 12424 13636 12436
rect 12676 12396 13636 12424
rect 12676 12384 12682 12396
rect 13630 12384 13636 12396
rect 13688 12424 13694 12436
rect 14921 12427 14979 12433
rect 14921 12424 14933 12427
rect 13688 12396 14933 12424
rect 13688 12384 13694 12396
rect 14921 12393 14933 12396
rect 14967 12393 14979 12427
rect 18598 12424 18604 12436
rect 14921 12387 14979 12393
rect 15672 12396 18604 12424
rect 2958 12316 2964 12368
rect 3016 12356 3022 12368
rect 5261 12359 5319 12365
rect 5261 12356 5273 12359
rect 3016 12328 5273 12356
rect 3016 12316 3022 12328
rect 5261 12325 5273 12328
rect 5307 12325 5319 12359
rect 5552 12356 5580 12384
rect 5626 12356 5632 12368
rect 5552 12328 5632 12356
rect 5261 12319 5319 12325
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 5718 12316 5724 12368
rect 5776 12356 5782 12368
rect 6546 12356 6552 12368
rect 5776 12328 6552 12356
rect 5776 12316 5782 12328
rect 6546 12316 6552 12328
rect 6604 12316 6610 12368
rect 12802 12316 12808 12368
rect 12860 12356 12866 12368
rect 12897 12359 12955 12365
rect 12897 12356 12909 12359
rect 12860 12328 12909 12356
rect 12860 12316 12866 12328
rect 12897 12325 12909 12328
rect 12943 12356 12955 12359
rect 13814 12356 13820 12368
rect 12943 12328 13820 12356
rect 12943 12325 12955 12328
rect 12897 12319 12955 12325
rect 13814 12316 13820 12328
rect 13872 12316 13878 12368
rect 14274 12316 14280 12368
rect 14332 12356 14338 12368
rect 15672 12356 15700 12396
rect 18598 12384 18604 12396
rect 18656 12384 18662 12436
rect 19702 12424 19708 12436
rect 19663 12396 19708 12424
rect 19702 12384 19708 12396
rect 19760 12384 19766 12436
rect 20533 12427 20591 12433
rect 20533 12393 20545 12427
rect 20579 12424 20591 12427
rect 20622 12424 20628 12436
rect 20579 12396 20628 12424
rect 20579 12393 20591 12396
rect 20533 12387 20591 12393
rect 20622 12384 20628 12396
rect 20680 12384 20686 12436
rect 14332 12328 15700 12356
rect 14332 12316 14338 12328
rect 16942 12316 16948 12368
rect 17000 12356 17006 12368
rect 17000 12328 19334 12356
rect 17000 12316 17006 12328
rect 1210 12248 1216 12300
rect 1268 12288 1274 12300
rect 1949 12291 2007 12297
rect 1949 12288 1961 12291
rect 1268 12260 1961 12288
rect 1268 12248 1274 12260
rect 1949 12257 1961 12260
rect 1995 12257 2007 12291
rect 1949 12251 2007 12257
rect 2498 12248 2504 12300
rect 2556 12288 2562 12300
rect 3053 12291 3111 12297
rect 3053 12288 3065 12291
rect 2556 12260 3065 12288
rect 2556 12248 2562 12260
rect 3053 12257 3065 12260
rect 3099 12257 3111 12291
rect 4430 12288 4436 12300
rect 4391 12260 4436 12288
rect 3053 12251 3111 12257
rect 4430 12248 4436 12260
rect 4488 12248 4494 12300
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 7561 12291 7619 12297
rect 7561 12257 7573 12291
rect 7607 12288 7619 12291
rect 7742 12288 7748 12300
rect 7607 12260 7748 12288
rect 7607 12257 7619 12260
rect 7561 12251 7619 12257
rect 7742 12248 7748 12260
rect 7800 12248 7806 12300
rect 10520 12260 11008 12288
rect 2222 12220 2228 12232
rect 2183 12192 2228 12220
rect 2222 12180 2228 12192
rect 2280 12220 2286 12232
rect 2961 12223 3019 12229
rect 2280 12192 2774 12220
rect 2280 12180 2286 12192
rect 2746 12152 2774 12192
rect 2961 12189 2973 12223
rect 3007 12220 3019 12223
rect 3234 12220 3240 12232
rect 3007 12192 3240 12220
rect 3007 12189 3019 12192
rect 2961 12183 3019 12189
rect 3234 12180 3240 12192
rect 3292 12180 3298 12232
rect 4062 12180 4068 12232
rect 4120 12220 4126 12232
rect 6457 12223 6515 12229
rect 6457 12220 6469 12223
rect 4120 12192 6469 12220
rect 4120 12180 4126 12192
rect 6457 12189 6469 12192
rect 6503 12189 6515 12223
rect 7392 12220 7420 12248
rect 8113 12223 8171 12229
rect 8113 12220 8125 12223
rect 7392 12192 8125 12220
rect 6457 12183 6515 12189
rect 8113 12189 8125 12192
rect 8159 12189 8171 12223
rect 10520 12220 10548 12260
rect 8113 12183 8171 12189
rect 8220 12192 10548 12220
rect 10597 12223 10655 12229
rect 5629 12155 5687 12161
rect 5629 12152 5641 12155
rect 2746 12124 5641 12152
rect 5629 12121 5641 12124
rect 5675 12121 5687 12155
rect 8220 12152 8248 12192
rect 10597 12189 10609 12223
rect 10643 12220 10655 12223
rect 10870 12220 10876 12232
rect 10643 12192 10876 12220
rect 10643 12189 10655 12192
rect 10597 12183 10655 12189
rect 10870 12180 10876 12192
rect 10928 12180 10934 12232
rect 10980 12220 11008 12260
rect 12406 12260 15792 12288
rect 12406 12220 12434 12260
rect 10980 12192 12434 12220
rect 13357 12223 13415 12229
rect 13357 12189 13369 12223
rect 13403 12220 13415 12223
rect 13998 12220 14004 12232
rect 13403 12192 14004 12220
rect 13403 12189 13415 12192
rect 13357 12183 13415 12189
rect 13998 12180 14004 12192
rect 14056 12180 14062 12232
rect 15654 12220 15660 12232
rect 14108 12192 15660 12220
rect 10318 12152 10324 12164
rect 10376 12161 10382 12164
rect 5629 12115 5687 12121
rect 6012 12124 8248 12152
rect 10288 12124 10324 12152
rect 2038 12044 2044 12096
rect 2096 12084 2102 12096
rect 2501 12087 2559 12093
rect 2501 12084 2513 12087
rect 2096 12056 2513 12084
rect 2096 12044 2102 12056
rect 2501 12053 2513 12056
rect 2547 12053 2559 12087
rect 2866 12084 2872 12096
rect 2827 12056 2872 12084
rect 2501 12047 2559 12053
rect 2866 12044 2872 12056
rect 2924 12044 2930 12096
rect 3142 12044 3148 12096
rect 3200 12084 3206 12096
rect 3418 12084 3424 12096
rect 3200 12056 3424 12084
rect 3200 12044 3206 12056
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 3510 12044 3516 12096
rect 3568 12084 3574 12096
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 3568 12056 4261 12084
rect 3568 12044 3574 12056
rect 4249 12053 4261 12056
rect 4295 12053 4307 12087
rect 4249 12047 4307 12053
rect 4338 12044 4344 12096
rect 4396 12084 4402 12096
rect 4396 12056 4441 12084
rect 4396 12044 4402 12056
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 4985 12087 5043 12093
rect 4985 12084 4997 12087
rect 4672 12056 4997 12084
rect 4672 12044 4678 12056
rect 4985 12053 4997 12056
rect 5031 12084 5043 12087
rect 6012 12084 6040 12124
rect 10318 12112 10324 12124
rect 10376 12115 10388 12161
rect 11118 12155 11176 12161
rect 11118 12152 11130 12155
rect 10428 12124 11130 12152
rect 10376 12112 10382 12115
rect 5031 12056 6040 12084
rect 7285 12087 7343 12093
rect 5031 12053 5043 12056
rect 4985 12047 5043 12053
rect 7285 12053 7297 12087
rect 7331 12084 7343 12087
rect 8018 12084 8024 12096
rect 7331 12056 8024 12084
rect 7331 12053 7343 12056
rect 7285 12047 7343 12053
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 9214 12044 9220 12096
rect 9272 12084 9278 12096
rect 10428 12084 10456 12124
rect 11118 12121 11130 12124
rect 11164 12121 11176 12155
rect 11118 12115 11176 12121
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 13538 12152 13544 12164
rect 12667 12124 13544 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 13538 12112 13544 12124
rect 13596 12152 13602 12164
rect 13722 12152 13728 12164
rect 13596 12124 13728 12152
rect 13596 12112 13602 12124
rect 13722 12112 13728 12124
rect 13780 12152 13786 12164
rect 14108 12161 14136 12192
rect 15654 12180 15660 12192
rect 15712 12180 15718 12232
rect 15764 12220 15792 12260
rect 16850 12248 16856 12300
rect 16908 12288 16914 12300
rect 17681 12291 17739 12297
rect 17681 12288 17693 12291
rect 16908 12260 17693 12288
rect 16908 12248 16914 12260
rect 17681 12257 17693 12260
rect 17727 12257 17739 12291
rect 19306 12288 19334 12328
rect 19518 12316 19524 12368
rect 19576 12356 19582 12368
rect 19576 12328 21128 12356
rect 19576 12316 19582 12328
rect 21100 12297 21128 12328
rect 19981 12291 20039 12297
rect 19981 12288 19993 12291
rect 19306 12260 19993 12288
rect 17681 12251 17739 12257
rect 19981 12257 19993 12260
rect 20027 12257 20039 12291
rect 19981 12251 20039 12257
rect 21085 12291 21143 12297
rect 21085 12257 21097 12291
rect 21131 12257 21143 12291
rect 21085 12251 21143 12257
rect 19521 12223 19579 12229
rect 15764 12192 19472 12220
rect 14093 12155 14151 12161
rect 14093 12152 14105 12155
rect 13780 12124 14105 12152
rect 13780 12112 13786 12124
rect 14093 12121 14105 12124
rect 14139 12121 14151 12155
rect 14093 12115 14151 12121
rect 15194 12112 15200 12164
rect 15252 12152 15258 12164
rect 15924 12155 15982 12161
rect 15924 12152 15936 12155
rect 15252 12124 15936 12152
rect 15252 12112 15258 12124
rect 15924 12121 15936 12124
rect 15970 12152 15982 12155
rect 16850 12152 16856 12164
rect 15970 12124 16856 12152
rect 15970 12121 15982 12124
rect 15924 12115 15982 12121
rect 16850 12112 16856 12124
rect 16908 12112 16914 12164
rect 18049 12155 18107 12161
rect 18049 12152 18061 12155
rect 17328 12124 18061 12152
rect 17328 12096 17356 12124
rect 18049 12121 18061 12124
rect 18095 12152 18107 12155
rect 18417 12155 18475 12161
rect 18417 12152 18429 12155
rect 18095 12124 18429 12152
rect 18095 12121 18107 12124
rect 18049 12115 18107 12121
rect 18417 12121 18429 12124
rect 18463 12152 18475 12155
rect 18785 12155 18843 12161
rect 18785 12152 18797 12155
rect 18463 12124 18797 12152
rect 18463 12121 18475 12124
rect 18417 12115 18475 12121
rect 18785 12121 18797 12124
rect 18831 12121 18843 12155
rect 19444 12152 19472 12192
rect 19521 12189 19533 12223
rect 19567 12220 19579 12223
rect 21174 12220 21180 12232
rect 19567 12192 21180 12220
rect 19567 12189 19579 12192
rect 19521 12183 19579 12189
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 19978 12152 19984 12164
rect 19444 12124 19984 12152
rect 18785 12115 18843 12121
rect 19978 12112 19984 12124
rect 20036 12112 20042 12164
rect 20165 12155 20223 12161
rect 20165 12121 20177 12155
rect 20211 12152 20223 12155
rect 20530 12152 20536 12164
rect 20211 12124 20536 12152
rect 20211 12121 20223 12124
rect 20165 12115 20223 12121
rect 9272 12056 10456 12084
rect 13633 12087 13691 12093
rect 9272 12044 9278 12056
rect 13633 12053 13645 12087
rect 13679 12084 13691 12087
rect 14274 12084 14280 12096
rect 13679 12056 14280 12084
rect 13679 12053 13691 12056
rect 13633 12047 13691 12053
rect 14274 12044 14280 12056
rect 14332 12044 14338 12096
rect 14458 12084 14464 12096
rect 14419 12056 14464 12084
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 15378 12084 15384 12096
rect 15339 12056 15384 12084
rect 15378 12044 15384 12056
rect 15436 12044 15442 12096
rect 17034 12084 17040 12096
rect 16995 12056 17040 12084
rect 17034 12044 17040 12056
rect 17092 12044 17098 12096
rect 17310 12084 17316 12096
rect 17271 12056 17316 12084
rect 17310 12044 17316 12056
rect 17368 12044 17374 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 20180 12084 20208 12115
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 20901 12155 20959 12161
rect 20901 12121 20913 12155
rect 20947 12152 20959 12155
rect 21542 12152 21548 12164
rect 20947 12124 21548 12152
rect 20947 12121 20959 12124
rect 20901 12115 20959 12121
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 18196 12056 20208 12084
rect 20993 12087 21051 12093
rect 18196 12044 18202 12056
rect 20993 12053 21005 12087
rect 21039 12084 21051 12087
rect 21266 12084 21272 12096
rect 21039 12056 21272 12084
rect 21039 12053 21051 12056
rect 20993 12047 21051 12053
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 3510 11880 3516 11892
rect 3471 11852 3516 11880
rect 3510 11840 3516 11852
rect 3568 11840 3574 11892
rect 4246 11880 4252 11892
rect 4207 11852 4252 11880
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 4338 11840 4344 11892
rect 4396 11880 4402 11892
rect 5261 11883 5319 11889
rect 5261 11880 5273 11883
rect 4396 11852 5273 11880
rect 4396 11840 4402 11852
rect 5261 11849 5273 11852
rect 5307 11849 5319 11883
rect 7282 11880 7288 11892
rect 7243 11852 7288 11880
rect 5261 11843 5319 11849
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9493 11883 9551 11889
rect 9493 11880 9505 11883
rect 9180 11852 9505 11880
rect 9180 11840 9186 11852
rect 9493 11849 9505 11852
rect 9539 11849 9551 11883
rect 13170 11880 13176 11892
rect 13131 11852 13176 11880
rect 9493 11843 9551 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 15654 11840 15660 11892
rect 15712 11880 15718 11892
rect 15749 11883 15807 11889
rect 15749 11880 15761 11883
rect 15712 11852 15761 11880
rect 15712 11840 15718 11852
rect 15749 11849 15761 11852
rect 15795 11849 15807 11883
rect 15749 11843 15807 11849
rect 16945 11883 17003 11889
rect 16945 11849 16957 11883
rect 16991 11880 17003 11883
rect 19705 11883 19763 11889
rect 16991 11852 19288 11880
rect 16991 11849 17003 11852
rect 16945 11843 17003 11849
rect 3145 11815 3203 11821
rect 3145 11781 3157 11815
rect 3191 11812 3203 11815
rect 3970 11812 3976 11824
rect 3191 11784 3976 11812
rect 3191 11781 3203 11784
rect 3145 11775 3203 11781
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 4157 11815 4215 11821
rect 4157 11781 4169 11815
rect 4203 11812 4215 11815
rect 6454 11812 6460 11824
rect 4203 11784 6460 11812
rect 4203 11781 4215 11784
rect 4157 11775 4215 11781
rect 6454 11772 6460 11784
rect 6512 11772 6518 11824
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 7466 11812 7472 11824
rect 7239 11784 7472 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 7466 11772 7472 11784
rect 7524 11772 7530 11824
rect 10594 11772 10600 11824
rect 10652 11821 10658 11824
rect 10652 11812 10664 11821
rect 10652 11784 10697 11812
rect 10652 11775 10664 11784
rect 10652 11772 10658 11775
rect 11054 11772 11060 11824
rect 11112 11812 11118 11824
rect 12038 11815 12096 11821
rect 12038 11812 12050 11815
rect 11112 11784 12050 11812
rect 11112 11772 11118 11784
rect 12038 11781 12050 11784
rect 12084 11781 12096 11815
rect 12038 11775 12096 11781
rect 12158 11772 12164 11824
rect 12216 11812 12222 11824
rect 13262 11812 13268 11824
rect 12216 11784 13268 11812
rect 12216 11772 12222 11784
rect 13262 11772 13268 11784
rect 13320 11772 13326 11824
rect 1946 11744 1952 11756
rect 1907 11716 1952 11744
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2130 11744 2136 11756
rect 2056 11716 2136 11744
rect 2056 11676 2084 11716
rect 2130 11704 2136 11716
rect 2188 11704 2194 11756
rect 4062 11744 4068 11756
rect 2746 11716 4068 11744
rect 2222 11676 2228 11688
rect 1964 11648 2084 11676
rect 2183 11648 2228 11676
rect 1964 11620 1992 11648
rect 2222 11636 2228 11648
rect 2280 11676 2286 11688
rect 2746 11676 2774 11716
rect 4062 11704 4068 11716
rect 4120 11704 4126 11756
rect 5626 11744 5632 11756
rect 5587 11716 5632 11744
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 5721 11747 5779 11753
rect 5721 11713 5733 11747
rect 5767 11744 5779 11747
rect 8110 11744 8116 11756
rect 5767 11716 8116 11744
rect 5767 11713 5779 11716
rect 5721 11707 5779 11713
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 8938 11704 8944 11756
rect 8996 11744 9002 11756
rect 13556 11744 13584 11840
rect 14200 11784 19196 11812
rect 14093 11747 14151 11753
rect 14093 11744 14105 11747
rect 8996 11716 13512 11744
rect 13556 11716 14105 11744
rect 8996 11704 9002 11716
rect 2280 11648 2774 11676
rect 2961 11679 3019 11685
rect 2280 11636 2286 11648
rect 2961 11645 2973 11679
rect 3007 11645 3019 11679
rect 2961 11639 3019 11645
rect 3053 11679 3111 11685
rect 3053 11645 3065 11679
rect 3099 11676 3111 11679
rect 4338 11676 4344 11688
rect 3099 11648 4344 11676
rect 3099 11645 3111 11648
rect 3053 11639 3111 11645
rect 1946 11568 1952 11620
rect 2004 11568 2010 11620
rect 2976 11540 3004 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4433 11679 4491 11685
rect 4433 11645 4445 11679
rect 4479 11676 4491 11679
rect 4614 11676 4620 11688
rect 4479 11648 4620 11676
rect 4479 11645 4491 11648
rect 4433 11639 4491 11645
rect 4614 11636 4620 11648
rect 4672 11636 4678 11688
rect 4893 11679 4951 11685
rect 4893 11645 4905 11679
rect 4939 11676 4951 11679
rect 5810 11676 5816 11688
rect 4939 11648 5816 11676
rect 4939 11645 4951 11648
rect 4893 11639 4951 11645
rect 3234 11568 3240 11620
rect 3292 11608 3298 11620
rect 3789 11611 3847 11617
rect 3789 11608 3801 11611
rect 3292 11580 3801 11608
rect 3292 11568 3298 11580
rect 3789 11577 3801 11580
rect 3835 11577 3847 11611
rect 3789 11571 3847 11577
rect 4908 11540 4936 11639
rect 5810 11636 5816 11648
rect 5868 11636 5874 11688
rect 6638 11676 6644 11688
rect 6599 11648 6644 11676
rect 6638 11636 6644 11648
rect 6696 11636 6702 11688
rect 7101 11679 7159 11685
rect 7101 11645 7113 11679
rect 7147 11676 7159 11679
rect 10870 11676 10876 11688
rect 7147 11648 9904 11676
rect 10831 11648 10876 11676
rect 7147 11645 7159 11648
rect 7101 11639 7159 11645
rect 7653 11611 7711 11617
rect 7653 11577 7665 11611
rect 7699 11608 7711 11611
rect 8386 11608 8392 11620
rect 7699 11580 8392 11608
rect 7699 11577 7711 11580
rect 7653 11571 7711 11577
rect 8386 11568 8392 11580
rect 8444 11568 8450 11620
rect 8757 11611 8815 11617
rect 8757 11577 8769 11611
rect 8803 11608 8815 11611
rect 9398 11608 9404 11620
rect 8803 11580 9404 11608
rect 8803 11577 8815 11580
rect 8757 11571 8815 11577
rect 9398 11568 9404 11580
rect 9456 11568 9462 11620
rect 2976 11512 4936 11540
rect 7374 11500 7380 11552
rect 7432 11540 7438 11552
rect 7742 11540 7748 11552
rect 7432 11512 7748 11540
rect 7432 11500 7438 11512
rect 7742 11500 7748 11512
rect 7800 11540 7806 11552
rect 7929 11543 7987 11549
rect 7929 11540 7941 11543
rect 7800 11512 7941 11540
rect 7800 11500 7806 11512
rect 7929 11509 7941 11512
rect 7975 11509 7987 11543
rect 7929 11503 7987 11509
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8297 11543 8355 11549
rect 8297 11540 8309 11543
rect 8260 11512 8309 11540
rect 8260 11500 8266 11512
rect 8297 11509 8309 11512
rect 8343 11509 8355 11543
rect 8297 11503 8355 11509
rect 9125 11543 9183 11549
rect 9125 11509 9137 11543
rect 9171 11540 9183 11543
rect 9490 11540 9496 11552
rect 9171 11512 9496 11540
rect 9171 11509 9183 11512
rect 9125 11503 9183 11509
rect 9490 11500 9496 11512
rect 9548 11500 9554 11552
rect 9876 11540 9904 11648
rect 10870 11636 10876 11648
rect 10928 11676 10934 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 10928 11648 11805 11676
rect 10928 11636 10934 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 13484 11676 13512 11716
rect 14093 11713 14105 11716
rect 14139 11713 14151 11747
rect 14093 11707 14151 11713
rect 14200 11676 14228 11784
rect 14366 11753 14372 11756
rect 14360 11744 14372 11753
rect 14279 11716 14372 11744
rect 14360 11707 14372 11716
rect 14424 11744 14430 11756
rect 14826 11744 14832 11756
rect 14424 11716 14832 11744
rect 14366 11704 14372 11707
rect 14424 11704 14430 11716
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 16301 11747 16359 11753
rect 16301 11713 16313 11747
rect 16347 11744 16359 11747
rect 18046 11744 18052 11756
rect 16347 11716 18052 11744
rect 16347 11713 16359 11716
rect 16301 11707 16359 11713
rect 18046 11704 18052 11716
rect 18104 11704 18110 11756
rect 18230 11753 18236 11756
rect 18224 11707 18236 11753
rect 18288 11744 18294 11756
rect 18288 11716 18324 11744
rect 18230 11704 18236 11707
rect 18288 11704 18294 11716
rect 13484 11648 14228 11676
rect 11793 11639 11851 11645
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17957 11679 18015 11685
rect 17957 11676 17969 11679
rect 17368 11648 17969 11676
rect 17368 11636 17374 11648
rect 17957 11645 17969 11648
rect 18003 11645 18015 11679
rect 19168 11676 19196 11784
rect 19260 11744 19288 11852
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 19794 11880 19800 11892
rect 19751 11852 19800 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 19978 11840 19984 11892
rect 20036 11880 20042 11892
rect 20073 11883 20131 11889
rect 20073 11880 20085 11883
rect 20036 11852 20085 11880
rect 20036 11840 20042 11852
rect 20073 11849 20085 11852
rect 20119 11849 20131 11883
rect 20073 11843 20131 11849
rect 20809 11883 20867 11889
rect 20809 11849 20821 11883
rect 20855 11880 20867 11883
rect 20898 11880 20904 11892
rect 20855 11852 20904 11880
rect 20855 11849 20867 11852
rect 20809 11843 20867 11849
rect 20898 11840 20904 11852
rect 20956 11840 20962 11892
rect 21266 11880 21272 11892
rect 21227 11852 21272 11880
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 20162 11744 20168 11756
rect 19260 11716 20168 11744
rect 20162 11704 20168 11716
rect 20220 11704 20226 11756
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11744 20959 11747
rect 21450 11744 21456 11756
rect 20947 11716 21456 11744
rect 20947 11713 20959 11716
rect 20901 11707 20959 11713
rect 21450 11704 21456 11716
rect 21508 11704 21514 11756
rect 20717 11679 20775 11685
rect 19168 11648 20576 11676
rect 17957 11639 18015 11645
rect 15194 11568 15200 11620
rect 15252 11608 15258 11620
rect 15378 11608 15384 11620
rect 15252 11580 15384 11608
rect 15252 11568 15258 11580
rect 15378 11568 15384 11580
rect 15436 11608 15442 11620
rect 16482 11608 16488 11620
rect 15436 11580 16488 11608
rect 15436 11568 15442 11580
rect 16482 11568 16488 11580
rect 16540 11568 16546 11620
rect 17221 11611 17279 11617
rect 17221 11577 17233 11611
rect 17267 11608 17279 11611
rect 19337 11611 19395 11617
rect 17267 11580 18000 11608
rect 17267 11577 17279 11580
rect 17221 11571 17279 11577
rect 11054 11540 11060 11552
rect 9876 11512 11060 11540
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 15470 11540 15476 11552
rect 15431 11512 15476 11540
rect 15470 11500 15476 11512
rect 15528 11500 15534 11552
rect 17310 11500 17316 11552
rect 17368 11540 17374 11552
rect 17589 11543 17647 11549
rect 17589 11540 17601 11543
rect 17368 11512 17601 11540
rect 17368 11500 17374 11512
rect 17589 11509 17601 11512
rect 17635 11509 17647 11543
rect 17972 11540 18000 11580
rect 19337 11577 19349 11611
rect 19383 11608 19395 11611
rect 19794 11608 19800 11620
rect 19383 11580 19800 11608
rect 19383 11577 19395 11580
rect 19337 11571 19395 11577
rect 19794 11568 19800 11580
rect 19852 11608 19858 11620
rect 20438 11608 20444 11620
rect 19852 11580 20444 11608
rect 19852 11568 19858 11580
rect 20438 11568 20444 11580
rect 20496 11568 20502 11620
rect 19518 11540 19524 11552
rect 17972 11512 19524 11540
rect 17589 11503 17647 11509
rect 19518 11500 19524 11512
rect 19576 11500 19582 11552
rect 20548 11540 20576 11648
rect 20717 11645 20729 11679
rect 20763 11645 20775 11679
rect 20717 11639 20775 11645
rect 20732 11608 20760 11639
rect 20898 11608 20904 11620
rect 20732 11580 20904 11608
rect 20898 11568 20904 11580
rect 20956 11568 20962 11620
rect 21082 11540 21088 11552
rect 20548 11512 21088 11540
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1673 11339 1731 11345
rect 1673 11305 1685 11339
rect 1719 11336 1731 11339
rect 1854 11336 1860 11348
rect 1719 11308 1860 11336
rect 1719 11305 1731 11308
rect 1673 11299 1731 11305
rect 1854 11296 1860 11308
rect 1912 11296 1918 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 5166 11336 5172 11348
rect 4019 11308 5172 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 5166 11296 5172 11308
rect 5224 11296 5230 11348
rect 6914 11336 6920 11348
rect 5276 11308 6920 11336
rect 1946 11228 1952 11280
rect 2004 11268 2010 11280
rect 2961 11271 3019 11277
rect 2004 11240 2268 11268
rect 2004 11228 2010 11240
rect 2240 11212 2268 11240
rect 2961 11237 2973 11271
rect 3007 11268 3019 11271
rect 5276 11268 5304 11308
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 9674 11336 9680 11348
rect 9263 11308 9680 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10226 11296 10232 11348
rect 10284 11336 10290 11348
rect 11698 11336 11704 11348
rect 10284 11308 11704 11336
rect 10284 11296 10290 11308
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 13081 11339 13139 11345
rect 13081 11305 13093 11339
rect 13127 11336 13139 11339
rect 13538 11336 13544 11348
rect 13127 11308 13544 11336
rect 13127 11305 13139 11308
rect 13081 11299 13139 11305
rect 3007 11240 5304 11268
rect 5353 11271 5411 11277
rect 3007 11237 3019 11240
rect 2961 11231 3019 11237
rect 5353 11237 5365 11271
rect 5399 11268 5411 11271
rect 12618 11268 12624 11280
rect 5399 11240 6132 11268
rect 5399 11237 5411 11240
rect 5353 11231 5411 11237
rect 2222 11160 2228 11212
rect 2280 11200 2286 11212
rect 2280 11172 2325 11200
rect 2280 11160 2286 11172
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 4614 11200 4620 11212
rect 2556 11172 4620 11200
rect 2556 11160 2562 11172
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 5166 11200 5172 11212
rect 4847 11172 5172 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 5166 11160 5172 11172
rect 5224 11200 5230 11212
rect 5718 11200 5724 11212
rect 5224 11172 5724 11200
rect 5224 11160 5230 11172
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6104 11209 6132 11240
rect 10612 11240 12624 11268
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 6181 11203 6239 11209
rect 6181 11169 6193 11203
rect 6227 11169 6239 11203
rect 6181 11163 6239 11169
rect 7285 11203 7343 11209
rect 7285 11169 7297 11203
rect 7331 11200 7343 11203
rect 8018 11200 8024 11212
rect 7331 11172 8024 11200
rect 7331 11169 7343 11172
rect 7285 11163 7343 11169
rect 2038 11132 2044 11144
rect 1999 11104 2044 11132
rect 2038 11092 2044 11104
rect 2096 11092 2102 11144
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 2958 11132 2964 11144
rect 2823 11104 2964 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3234 11132 3240 11144
rect 3068 11104 3240 11132
rect 2133 11067 2191 11073
rect 2133 11033 2145 11067
rect 2179 11064 2191 11067
rect 3068 11064 3096 11104
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 3786 11132 3792 11144
rect 3747 11104 3792 11132
rect 3786 11092 3792 11104
rect 3844 11132 3850 11144
rect 4430 11132 4436 11144
rect 3844 11104 4436 11132
rect 3844 11092 3850 11104
rect 4430 11092 4436 11104
rect 4488 11092 4494 11144
rect 4982 11132 4988 11144
rect 4632 11104 4988 11132
rect 2179 11036 3096 11064
rect 4341 11067 4399 11073
rect 2179 11033 2191 11036
rect 2133 11027 2191 11033
rect 4341 11033 4353 11067
rect 4387 11064 4399 11067
rect 4632 11064 4660 11104
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5994 11132 6000 11144
rect 5955 11104 6000 11132
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 4387 11036 4660 11064
rect 4387 11033 4399 11036
rect 4341 11027 4399 11033
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4764 11036 4905 11064
rect 4764 11024 4770 11036
rect 4893 11033 4905 11036
rect 4939 11064 4951 11067
rect 5350 11064 5356 11076
rect 4939 11036 5356 11064
rect 4939 11033 4951 11036
rect 4893 11027 4951 11033
rect 5350 11024 5356 11036
rect 5408 11024 5414 11076
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 6196 11064 6224 11163
rect 8018 11160 8024 11172
rect 8076 11160 8082 11212
rect 8481 11203 8539 11209
rect 8481 11169 8493 11203
rect 8527 11200 8539 11203
rect 10612 11200 10640 11240
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 8527 11172 9076 11200
rect 8527 11169 8539 11172
rect 8481 11163 8539 11169
rect 8772 11144 8800 11172
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6696 11104 7021 11132
rect 6696 11092 6702 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7466 11092 7472 11144
rect 7524 11132 7530 11144
rect 8202 11132 8208 11144
rect 7524 11104 8208 11132
rect 7524 11092 7530 11104
rect 8202 11092 8208 11104
rect 8260 11092 8266 11144
rect 8294 11092 8300 11144
rect 8352 11132 8358 11144
rect 8570 11132 8576 11144
rect 8352 11104 8576 11132
rect 8352 11092 8358 11104
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8754 11092 8760 11144
rect 8812 11092 8818 11144
rect 7101 11067 7159 11073
rect 7101 11064 7113 11067
rect 5776 11036 6224 11064
rect 6840 11036 7113 11064
rect 5776 11024 5782 11036
rect 6840 11008 6868 11036
rect 7101 11033 7113 11036
rect 7147 11064 7159 11067
rect 8662 11064 8668 11076
rect 7147 11036 8668 11064
rect 7147 11033 7159 11036
rect 7101 11027 7159 11033
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 9048 11064 9076 11172
rect 10520 11172 10640 11200
rect 9122 11092 9128 11144
rect 9180 11132 9186 11144
rect 10330 11135 10388 11141
rect 10330 11132 10342 11135
rect 9180 11104 10342 11132
rect 9180 11092 9186 11104
rect 10330 11101 10342 11104
rect 10376 11101 10388 11135
rect 10330 11095 10388 11101
rect 10520 11064 10548 11172
rect 11054 11160 11060 11212
rect 11112 11200 11118 11212
rect 12526 11200 12532 11212
rect 11112 11172 12434 11200
rect 12487 11172 12532 11200
rect 11112 11160 11118 11172
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10778 11132 10784 11144
rect 10643 11104 10784 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10778 11092 10784 11104
rect 10836 11092 10842 11144
rect 12066 11132 12072 11144
rect 12027 11104 12072 11132
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12406 11132 12434 11172
rect 12526 11160 12532 11172
rect 12584 11200 12590 11212
rect 12894 11200 12900 11212
rect 12584 11172 12900 11200
rect 12584 11160 12590 11172
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 12618 11132 12624 11144
rect 12406 11104 12624 11132
rect 12618 11092 12624 11104
rect 12676 11092 12682 11144
rect 11882 11064 11888 11076
rect 9048 11036 10548 11064
rect 10612 11036 11888 11064
rect 3234 10996 3240 11008
rect 3195 10968 3240 10996
rect 3234 10956 3240 10968
rect 3292 10956 3298 11008
rect 5626 10996 5632 11008
rect 5587 10968 5632 10996
rect 5626 10956 5632 10968
rect 5684 10956 5690 11008
rect 6638 10996 6644 11008
rect 6599 10968 6644 10996
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 6822 10956 6828 11008
rect 6880 10956 6886 11008
rect 7834 10996 7840 11008
rect 7795 10968 7840 10996
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 8110 10956 8116 11008
rect 8168 10996 8174 11008
rect 8297 10999 8355 11005
rect 8297 10996 8309 10999
rect 8168 10968 8309 10996
rect 8168 10956 8174 10968
rect 8297 10965 8309 10968
rect 8343 10996 8355 10999
rect 10612 10996 10640 11036
rect 11882 11024 11888 11036
rect 11940 11024 11946 11076
rect 8343 10968 10640 10996
rect 8343 10965 8355 10968
rect 8297 10959 8355 10965
rect 10778 10956 10784 11008
rect 10836 10996 10842 11008
rect 11057 10999 11115 11005
rect 11057 10996 11069 10999
rect 10836 10968 11069 10996
rect 10836 10956 10842 10968
rect 11057 10965 11069 10968
rect 11103 10996 11115 10999
rect 11238 10996 11244 11008
rect 11103 10968 11244 10996
rect 11103 10965 11115 10968
rect 11057 10959 11115 10965
rect 11238 10956 11244 10968
rect 11296 10996 11302 11008
rect 11333 10999 11391 11005
rect 11333 10996 11345 10999
rect 11296 10968 11345 10996
rect 11296 10956 11302 10968
rect 11333 10965 11345 10968
rect 11379 10996 11391 10999
rect 13096 10996 13124 11299
rect 13538 11296 13544 11308
rect 13596 11336 13602 11348
rect 14093 11339 14151 11345
rect 14093 11336 14105 11339
rect 13596 11308 14105 11336
rect 13596 11296 13602 11308
rect 14093 11305 14105 11308
rect 14139 11336 14151 11339
rect 14829 11339 14887 11345
rect 14829 11336 14841 11339
rect 14139 11308 14841 11336
rect 14139 11305 14151 11308
rect 14093 11299 14151 11305
rect 14829 11305 14841 11308
rect 14875 11336 14887 11339
rect 14918 11336 14924 11348
rect 14875 11308 14924 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 15289 11339 15347 11345
rect 15289 11305 15301 11339
rect 15335 11336 15347 11339
rect 18966 11336 18972 11348
rect 15335 11308 18972 11336
rect 15335 11305 15347 11308
rect 15289 11299 15347 11305
rect 18966 11296 18972 11308
rect 19024 11296 19030 11348
rect 21266 11336 21272 11348
rect 19812 11308 21272 11336
rect 14553 11271 14611 11277
rect 14553 11237 14565 11271
rect 14599 11268 14611 11271
rect 15378 11268 15384 11280
rect 14599 11240 15384 11268
rect 14599 11237 14611 11240
rect 14553 11231 14611 11237
rect 15378 11228 15384 11240
rect 15436 11228 15442 11280
rect 16574 11228 16580 11280
rect 16632 11268 16638 11280
rect 16945 11271 17003 11277
rect 16945 11268 16957 11271
rect 16632 11240 16957 11268
rect 16632 11228 16638 11240
rect 16945 11237 16957 11240
rect 16991 11237 17003 11271
rect 16945 11231 17003 11237
rect 18598 11228 18604 11280
rect 18656 11268 18662 11280
rect 18693 11271 18751 11277
rect 18693 11268 18705 11271
rect 18656 11240 18705 11268
rect 18656 11228 18662 11240
rect 18693 11237 18705 11240
rect 18739 11237 18751 11271
rect 18693 11231 18751 11237
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 19518 11268 19524 11280
rect 19475 11240 19524 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 19518 11228 19524 11240
rect 19576 11228 19582 11280
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 14976 11172 15577 11200
rect 14976 11160 14982 11172
rect 15565 11169 15577 11172
rect 15611 11169 15623 11203
rect 15565 11163 15623 11169
rect 15010 11092 15016 11144
rect 15068 11132 15074 11144
rect 15821 11135 15879 11141
rect 15821 11132 15833 11135
rect 15068 11104 15833 11132
rect 15068 11092 15074 11104
rect 15821 11101 15833 11104
rect 15867 11101 15879 11135
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 15821 11095 15879 11101
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 17569 11135 17627 11141
rect 17569 11132 17581 11135
rect 17460 11104 17581 11132
rect 17460 11092 17466 11104
rect 17569 11101 17581 11104
rect 17615 11101 17627 11135
rect 17569 11095 17627 11101
rect 18046 11092 18052 11144
rect 18104 11132 18110 11144
rect 19812 11132 19840 11308
rect 21266 11296 21272 11308
rect 21324 11296 21330 11348
rect 18104 11104 19840 11132
rect 20809 11135 20867 11141
rect 18104 11092 18110 11104
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 20990 11132 20996 11144
rect 20855 11104 20996 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 21284 11141 21312 11296
rect 21269 11135 21327 11141
rect 21269 11101 21281 11135
rect 21315 11101 21327 11135
rect 21269 11095 21327 11101
rect 13262 11024 13268 11076
rect 13320 11064 13326 11076
rect 20564 11067 20622 11073
rect 13320 11036 20484 11064
rect 13320 11024 13326 11036
rect 13354 10996 13360 11008
rect 11379 10968 13124 10996
rect 13315 10968 13360 10996
rect 11379 10965 11391 10968
rect 11333 10959 11391 10965
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 20456 10996 20484 11036
rect 20564 11033 20576 11067
rect 20610 11064 20622 11067
rect 20898 11064 20904 11076
rect 20610 11036 20904 11064
rect 20610 11033 20622 11036
rect 20564 11027 20622 11033
rect 20898 11024 20904 11036
rect 20956 11024 20962 11076
rect 21085 11067 21143 11073
rect 21085 11064 21097 11067
rect 21008 11036 21097 11064
rect 21008 10996 21036 11036
rect 21085 11033 21097 11036
rect 21131 11033 21143 11067
rect 21085 11027 21143 11033
rect 20456 10968 21036 10996
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 2501 10795 2559 10801
rect 2501 10792 2513 10795
rect 2464 10764 2513 10792
rect 2464 10752 2470 10764
rect 2501 10761 2513 10764
rect 2547 10761 2559 10795
rect 2682 10792 2688 10804
rect 2501 10755 2559 10761
rect 2608 10764 2688 10792
rect 2130 10684 2136 10736
rect 2188 10724 2194 10736
rect 2608 10724 2636 10764
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 3878 10792 3884 10804
rect 3839 10764 3884 10792
rect 3878 10752 3884 10764
rect 3936 10752 3942 10804
rect 4430 10752 4436 10804
rect 4488 10792 4494 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4488 10764 4537 10792
rect 4488 10752 4494 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5442 10792 5448 10804
rect 5031 10764 5448 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 2188 10696 2636 10724
rect 2746 10696 4016 10724
rect 2188 10684 2194 10696
rect 2746 10668 2774 10696
rect 1762 10616 1768 10668
rect 1820 10656 1826 10668
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1820 10628 1961 10656
rect 1820 10616 1826 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2225 10659 2283 10665
rect 2225 10625 2237 10659
rect 2271 10656 2283 10659
rect 2746 10656 2780 10668
rect 2271 10628 2780 10656
rect 2271 10625 2283 10628
rect 2225 10619 2283 10625
rect 2774 10616 2780 10628
rect 2832 10616 2838 10668
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3418 10656 3424 10668
rect 2915 10628 3424 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 3418 10616 3424 10628
rect 3476 10616 3482 10668
rect 3988 10656 4016 10696
rect 4246 10684 4252 10736
rect 4304 10724 4310 10736
rect 5000 10724 5028 10755
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 6638 10752 6644 10804
rect 6696 10792 6702 10804
rect 6825 10795 6883 10801
rect 6825 10792 6837 10795
rect 6696 10764 6837 10792
rect 6696 10752 6702 10764
rect 6825 10761 6837 10764
rect 6871 10761 6883 10795
rect 6825 10755 6883 10761
rect 7469 10795 7527 10801
rect 7469 10761 7481 10795
rect 7515 10792 7527 10795
rect 7558 10792 7564 10804
rect 7515 10764 7564 10792
rect 7515 10761 7527 10764
rect 7469 10755 7527 10761
rect 7558 10752 7564 10764
rect 7616 10752 7622 10804
rect 7929 10795 7987 10801
rect 7929 10761 7941 10795
rect 7975 10792 7987 10795
rect 8202 10792 8208 10804
rect 7975 10764 8208 10792
rect 7975 10761 7987 10764
rect 7929 10755 7987 10761
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 8478 10752 8484 10804
rect 8536 10792 8542 10804
rect 9214 10792 9220 10804
rect 8536 10764 9220 10792
rect 8536 10752 8542 10764
rect 9214 10752 9220 10764
rect 9272 10752 9278 10804
rect 10318 10752 10324 10804
rect 10376 10792 10382 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 10376 10764 11529 10792
rect 10376 10752 10382 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 14918 10792 14924 10804
rect 14879 10764 14924 10792
rect 11517 10755 11575 10761
rect 14918 10752 14924 10764
rect 14976 10792 14982 10804
rect 15473 10795 15531 10801
rect 15473 10792 15485 10795
rect 14976 10764 15485 10792
rect 14976 10752 14982 10764
rect 15473 10761 15485 10764
rect 15519 10792 15531 10795
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15519 10764 15853 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 15841 10761 15853 10764
rect 15887 10792 15899 10795
rect 16209 10795 16267 10801
rect 16209 10792 16221 10795
rect 15887 10764 16221 10792
rect 15887 10761 15899 10764
rect 15841 10755 15899 10761
rect 16209 10761 16221 10764
rect 16255 10792 16267 10795
rect 17129 10795 17187 10801
rect 17129 10792 17141 10795
rect 16255 10764 17141 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 17129 10761 17141 10764
rect 17175 10792 17187 10795
rect 17310 10792 17316 10804
rect 17175 10764 17316 10792
rect 17175 10761 17187 10764
rect 17129 10755 17187 10761
rect 17310 10752 17316 10764
rect 17368 10792 17374 10804
rect 17497 10795 17555 10801
rect 17497 10792 17509 10795
rect 17368 10764 17509 10792
rect 17368 10752 17374 10764
rect 17497 10761 17509 10764
rect 17543 10761 17555 10795
rect 17497 10755 17555 10761
rect 4304 10696 5028 10724
rect 4304 10684 4310 10696
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 8110 10724 8116 10736
rect 5868 10696 8116 10724
rect 5868 10684 5874 10696
rect 8110 10684 8116 10696
rect 8168 10684 8174 10736
rect 8570 10724 8576 10736
rect 8312 10696 8576 10724
rect 4890 10656 4896 10668
rect 3988 10628 4896 10656
rect 4890 10616 4896 10628
rect 4948 10616 4954 10668
rect 5442 10656 5448 10668
rect 5403 10628 5448 10656
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 7837 10659 7895 10665
rect 5552 10628 7420 10656
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 2961 10591 3019 10597
rect 2961 10588 2973 10591
rect 2464 10560 2973 10588
rect 2464 10548 2470 10560
rect 2961 10557 2973 10560
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 3053 10591 3111 10597
rect 3053 10557 3065 10591
rect 3099 10557 3111 10591
rect 3970 10588 3976 10600
rect 3931 10560 3976 10588
rect 3053 10551 3111 10557
rect 2498 10480 2504 10532
rect 2556 10520 2562 10532
rect 2682 10520 2688 10532
rect 2556 10492 2688 10520
rect 2556 10480 2562 10492
rect 2682 10480 2688 10492
rect 2740 10520 2746 10532
rect 3068 10520 3096 10551
rect 3970 10548 3976 10560
rect 4028 10548 4034 10600
rect 4062 10548 4068 10600
rect 4120 10588 4126 10600
rect 4120 10560 4165 10588
rect 4120 10548 4126 10560
rect 4614 10548 4620 10600
rect 4672 10588 4678 10600
rect 5552 10588 5580 10628
rect 4672 10560 5580 10588
rect 6641 10591 6699 10597
rect 4672 10548 4678 10560
rect 6641 10557 6653 10591
rect 6687 10557 6699 10591
rect 6641 10551 6699 10557
rect 6733 10591 6791 10597
rect 6733 10557 6745 10591
rect 6779 10588 6791 10591
rect 7282 10588 7288 10600
rect 6779 10560 7288 10588
rect 6779 10557 6791 10560
rect 6733 10551 6791 10557
rect 2740 10492 3096 10520
rect 6656 10520 6684 10551
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7392 10588 7420 10628
rect 7837 10625 7849 10659
rect 7883 10656 7895 10659
rect 8312 10656 8340 10696
rect 8570 10684 8576 10696
rect 8628 10684 8634 10736
rect 8754 10724 8760 10736
rect 8715 10696 8760 10724
rect 8754 10684 8760 10696
rect 8812 10684 8818 10736
rect 11238 10684 11244 10736
rect 11296 10724 11302 10736
rect 11296 10696 12940 10724
rect 11296 10684 11302 10696
rect 7883 10628 8340 10656
rect 7883 10625 7895 10628
rect 7837 10619 7895 10625
rect 8110 10588 8116 10600
rect 7392 10560 7972 10588
rect 8071 10560 8116 10588
rect 7558 10520 7564 10532
rect 6656 10492 7564 10520
rect 2740 10480 2746 10492
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 2958 10412 2964 10464
rect 3016 10452 3022 10464
rect 3513 10455 3571 10461
rect 3513 10452 3525 10455
rect 3016 10424 3525 10452
rect 3016 10412 3022 10424
rect 3513 10421 3525 10424
rect 3559 10421 3571 10455
rect 5258 10452 5264 10464
rect 5219 10424 5264 10452
rect 3513 10415 3571 10421
rect 5258 10412 5264 10424
rect 5316 10412 5322 10464
rect 5350 10412 5356 10464
rect 5408 10452 5414 10464
rect 5810 10452 5816 10464
rect 5408 10424 5816 10452
rect 5408 10412 5414 10424
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 7098 10412 7104 10464
rect 7156 10452 7162 10464
rect 7193 10455 7251 10461
rect 7193 10452 7205 10455
rect 7156 10424 7205 10452
rect 7156 10412 7162 10424
rect 7193 10421 7205 10424
rect 7239 10421 7251 10455
rect 7944 10452 7972 10560
rect 8110 10548 8116 10560
rect 8168 10548 8174 10600
rect 8478 10548 8484 10600
rect 8536 10588 8542 10600
rect 8772 10588 8800 10684
rect 10341 10659 10399 10665
rect 10341 10625 10353 10659
rect 10387 10656 10399 10659
rect 10502 10656 10508 10668
rect 10387 10628 10508 10656
rect 10387 10625 10399 10628
rect 10341 10619 10399 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 12618 10616 12624 10668
rect 12676 10665 12682 10668
rect 12912 10665 12940 10696
rect 12676 10656 12688 10665
rect 12897 10659 12955 10665
rect 12676 10628 12721 10656
rect 12676 10619 12688 10628
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13265 10659 13323 10665
rect 13265 10656 13277 10659
rect 12943 10628 13277 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13265 10625 13277 10628
rect 13311 10625 13323 10659
rect 13265 10619 13323 10625
rect 12676 10616 12682 10619
rect 13354 10616 13360 10668
rect 13412 10656 13418 10668
rect 13521 10659 13579 10665
rect 13521 10656 13533 10659
rect 13412 10628 13533 10656
rect 13412 10616 13418 10628
rect 13521 10625 13533 10628
rect 13567 10625 13579 10659
rect 17512 10656 17540 10755
rect 17678 10752 17684 10804
rect 17736 10792 17742 10804
rect 17862 10792 17868 10804
rect 17736 10764 17868 10792
rect 17736 10752 17742 10764
rect 17862 10752 17868 10764
rect 17920 10792 17926 10804
rect 19245 10795 19303 10801
rect 19245 10792 19257 10795
rect 17920 10764 19257 10792
rect 17920 10752 17926 10764
rect 19245 10761 19257 10764
rect 19291 10761 19303 10795
rect 20898 10792 20904 10804
rect 20859 10764 20904 10792
rect 19245 10755 19303 10761
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 21174 10792 21180 10804
rect 21135 10764 21180 10792
rect 21174 10752 21180 10764
rect 21232 10752 21238 10804
rect 17770 10684 17776 10736
rect 17828 10724 17834 10736
rect 19794 10733 19800 10736
rect 18110 10727 18168 10733
rect 18110 10724 18122 10727
rect 17828 10696 18122 10724
rect 17828 10684 17834 10696
rect 18110 10693 18122 10696
rect 18156 10693 18168 10727
rect 19788 10724 19800 10733
rect 19755 10696 19800 10724
rect 18110 10687 18168 10693
rect 19788 10687 19800 10696
rect 19794 10684 19800 10687
rect 19852 10684 19858 10736
rect 17678 10656 17684 10668
rect 17512 10628 17684 10656
rect 13521 10619 13579 10625
rect 17678 10616 17684 10628
rect 17736 10656 17742 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17736 10628 17877 10656
rect 17736 10616 17742 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 20714 10656 20720 10668
rect 17865 10619 17923 10625
rect 19536 10628 20720 10656
rect 8536 10560 8800 10588
rect 10597 10591 10655 10597
rect 8536 10548 8542 10560
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 13372 10588 13400 10616
rect 19536 10597 19564 10628
rect 20714 10616 20720 10628
rect 20772 10656 20778 10668
rect 20990 10656 20996 10668
rect 20772 10628 20996 10656
rect 20772 10616 20778 10628
rect 20990 10616 20996 10628
rect 21048 10616 21054 10668
rect 21358 10656 21364 10668
rect 21319 10628 21364 10656
rect 21358 10616 21364 10628
rect 21416 10616 21422 10668
rect 10597 10551 10655 10557
rect 13280 10560 13400 10588
rect 19521 10591 19579 10597
rect 10410 10452 10416 10464
rect 7944 10424 10416 10452
rect 7193 10415 7251 10421
rect 10410 10412 10416 10424
rect 10468 10412 10474 10464
rect 10612 10452 10640 10551
rect 10686 10480 10692 10532
rect 10744 10520 10750 10532
rect 10744 10492 11376 10520
rect 10744 10480 10750 10492
rect 10965 10455 11023 10461
rect 10965 10452 10977 10455
rect 10612 10424 10977 10452
rect 10965 10421 10977 10424
rect 11011 10452 11023 10455
rect 11238 10452 11244 10464
rect 11011 10424 11244 10452
rect 11011 10421 11023 10424
rect 10965 10415 11023 10421
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11348 10452 11376 10492
rect 13280 10452 13308 10560
rect 19521 10557 19533 10591
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 14645 10523 14703 10529
rect 14645 10489 14657 10523
rect 14691 10520 14703 10523
rect 17126 10520 17132 10532
rect 14691 10492 17132 10520
rect 14691 10489 14703 10492
rect 14645 10483 14703 10489
rect 17126 10480 17132 10492
rect 17184 10480 17190 10532
rect 11348 10424 13308 10452
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 16853 10455 16911 10461
rect 16853 10452 16865 10455
rect 14332 10424 16865 10452
rect 14332 10412 14338 10424
rect 16853 10421 16865 10424
rect 16899 10452 16911 10455
rect 17586 10452 17592 10464
rect 16899 10424 17592 10452
rect 16899 10421 16911 10424
rect 16853 10415 16911 10421
rect 17586 10412 17592 10424
rect 17644 10452 17650 10464
rect 19518 10452 19524 10464
rect 17644 10424 19524 10452
rect 17644 10412 17650 10424
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 5258 10248 5264 10260
rect 1452 10220 5264 10248
rect 1452 10208 1458 10220
rect 5258 10208 5264 10220
rect 5316 10208 5322 10260
rect 6549 10251 6607 10257
rect 6549 10217 6561 10251
rect 6595 10248 6607 10251
rect 6822 10248 6828 10260
rect 6595 10220 6828 10248
rect 6595 10217 6607 10220
rect 6549 10211 6607 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7282 10248 7288 10260
rect 7243 10220 7288 10248
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8018 10208 8024 10260
rect 8076 10248 8082 10260
rect 13814 10248 13820 10260
rect 8076 10220 13820 10248
rect 8076 10208 8082 10220
rect 13814 10208 13820 10220
rect 13872 10208 13878 10260
rect 14645 10251 14703 10257
rect 14645 10217 14657 10251
rect 14691 10248 14703 10251
rect 17678 10248 17684 10260
rect 14691 10220 17540 10248
rect 17639 10220 17684 10248
rect 14691 10217 14703 10220
rect 14645 10211 14703 10217
rect 3326 10180 3332 10192
rect 2746 10152 3332 10180
rect 1670 10072 1676 10124
rect 1728 10112 1734 10124
rect 1949 10115 2007 10121
rect 1949 10112 1961 10115
rect 1728 10084 1961 10112
rect 1728 10072 1734 10084
rect 1949 10081 1961 10084
rect 1995 10081 2007 10115
rect 1949 10075 2007 10081
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 2222 10004 2228 10016
rect 2280 10044 2286 10056
rect 2746 10044 2774 10152
rect 3326 10140 3332 10152
rect 3384 10140 3390 10192
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 4338 10180 4344 10192
rect 3752 10152 4344 10180
rect 3752 10140 3758 10152
rect 4338 10140 4344 10152
rect 4396 10140 4402 10192
rect 4798 10140 4804 10192
rect 4856 10180 4862 10192
rect 6914 10180 6920 10192
rect 4856 10152 6920 10180
rect 4856 10140 4862 10152
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 8297 10183 8355 10189
rect 8297 10180 8309 10183
rect 8168 10152 8309 10180
rect 8168 10140 8174 10152
rect 8297 10149 8309 10152
rect 8343 10149 8355 10183
rect 8297 10143 8355 10149
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 10781 10183 10839 10189
rect 10781 10180 10793 10183
rect 10744 10152 10793 10180
rect 10744 10140 10750 10152
rect 10781 10149 10793 10152
rect 10827 10149 10839 10183
rect 15654 10180 15660 10192
rect 10781 10143 10839 10149
rect 11532 10152 12204 10180
rect 15615 10152 15660 10180
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10081 3203 10115
rect 3145 10075 3203 10081
rect 2280 10016 2774 10044
rect 2280 10004 2286 10016
rect 3050 10004 3056 10056
rect 3108 10004 3114 10056
rect 3160 10044 3188 10075
rect 3418 10072 3424 10124
rect 3476 10112 3482 10124
rect 3789 10115 3847 10121
rect 3789 10112 3801 10115
rect 3476 10084 3801 10112
rect 3476 10072 3482 10084
rect 3789 10081 3801 10084
rect 3835 10081 3847 10115
rect 3789 10075 3847 10081
rect 5077 10115 5135 10121
rect 5077 10081 5089 10115
rect 5123 10112 5135 10115
rect 5258 10112 5264 10124
rect 5123 10084 5264 10112
rect 5123 10081 5135 10084
rect 5077 10075 5135 10081
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 7929 10115 7987 10121
rect 7929 10081 7941 10115
rect 7975 10112 7987 10115
rect 8202 10112 8208 10124
rect 7975 10084 8208 10112
rect 7975 10081 7987 10084
rect 7929 10075 7987 10081
rect 8202 10072 8208 10084
rect 8260 10112 8266 10124
rect 9306 10112 9312 10124
rect 8260 10084 9312 10112
rect 8260 10072 8266 10084
rect 9306 10072 9312 10084
rect 9364 10072 9370 10124
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11532 10112 11560 10152
rect 10468 10084 11560 10112
rect 11609 10115 11667 10121
rect 10468 10072 10474 10084
rect 11609 10081 11621 10115
rect 11655 10112 11667 10115
rect 11790 10112 11796 10124
rect 11655 10084 11796 10112
rect 11655 10081 11667 10084
rect 11609 10075 11667 10081
rect 11790 10072 11796 10084
rect 11848 10072 11854 10124
rect 12176 10112 12204 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 17512 10180 17540 10220
rect 17678 10208 17684 10220
rect 17736 10208 17742 10260
rect 19521 10251 19579 10257
rect 19521 10217 19533 10251
rect 19567 10248 19579 10251
rect 19610 10248 19616 10260
rect 19567 10220 19616 10248
rect 19567 10217 19579 10220
rect 19521 10211 19579 10217
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 17512 10152 20576 10180
rect 15672 10112 15700 10140
rect 20548 10124 20576 10152
rect 12176 10084 12296 10112
rect 15672 10084 16160 10112
rect 3510 10044 3516 10056
rect 3160 10016 3516 10044
rect 3510 10004 3516 10016
rect 3568 10004 3574 10056
rect 8110 10004 8116 10056
rect 8168 10044 8174 10056
rect 9401 10047 9459 10053
rect 8168 10016 9168 10044
rect 8168 10004 8174 10016
rect 3068 9976 3096 10004
rect 3234 9976 3240 9988
rect 3068 9948 3240 9976
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 4706 9936 4712 9988
rect 4764 9976 4770 9988
rect 4893 9979 4951 9985
rect 4893 9976 4905 9979
rect 4764 9948 4905 9976
rect 4764 9936 4770 9948
rect 4893 9945 4905 9948
rect 4939 9976 4951 9979
rect 7653 9979 7711 9985
rect 7653 9976 7665 9979
rect 4939 9948 7665 9976
rect 4939 9945 4951 9948
rect 4893 9939 4951 9945
rect 7653 9945 7665 9948
rect 7699 9945 7711 9979
rect 7653 9939 7711 9945
rect 7742 9936 7748 9988
rect 7800 9976 7806 9988
rect 7800 9948 9076 9976
rect 7800 9936 7806 9948
rect 9048 9920 9076 9948
rect 2498 9908 2504 9920
rect 2459 9880 2504 9908
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2832 9880 2881 9908
rect 2832 9868 2838 9880
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 2869 9871 2927 9877
rect 2961 9911 3019 9917
rect 2961 9877 2973 9911
rect 3007 9908 3019 9911
rect 3050 9908 3056 9920
rect 3007 9880 3056 9908
rect 3007 9877 3019 9880
rect 2961 9871 3019 9877
rect 3050 9868 3056 9880
rect 3108 9868 3114 9920
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 4798 9908 4804 9920
rect 4759 9880 4804 9908
rect 4798 9868 4804 9880
rect 4856 9868 4862 9920
rect 5350 9868 5356 9920
rect 5408 9908 5414 9920
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 5408 9880 5549 9908
rect 5408 9868 5414 9880
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 5537 9871 5595 9877
rect 5994 9868 6000 9920
rect 6052 9908 6058 9920
rect 6181 9911 6239 9917
rect 6181 9908 6193 9911
rect 6052 9880 6193 9908
rect 6052 9868 6058 9880
rect 6181 9877 6193 9880
rect 6227 9908 6239 9911
rect 6638 9908 6644 9920
rect 6227 9880 6644 9908
rect 6227 9877 6239 9880
rect 6181 9871 6239 9877
rect 6638 9868 6644 9880
rect 6696 9868 6702 9920
rect 6914 9908 6920 9920
rect 6875 9880 6920 9908
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 7098 9868 7104 9920
rect 7156 9908 7162 9920
rect 7926 9908 7932 9920
rect 7156 9880 7932 9908
rect 7156 9868 7162 9880
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9140 9908 9168 10016
rect 9401 10013 9413 10047
rect 9447 10044 9459 10047
rect 9490 10044 9496 10056
rect 9447 10016 9496 10044
rect 9447 10013 9459 10016
rect 9401 10007 9459 10013
rect 9490 10004 9496 10016
rect 9548 10004 9554 10056
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 11296 10016 12173 10044
rect 11296 10004 11302 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 9214 9936 9220 9988
rect 9272 9976 9278 9988
rect 9646 9979 9704 9985
rect 9646 9976 9658 9979
rect 9272 9948 9658 9976
rect 9272 9936 9278 9948
rect 9646 9945 9658 9948
rect 9692 9945 9704 9979
rect 12268 9976 12296 10084
rect 14185 10047 14243 10053
rect 14185 10013 14197 10047
rect 14231 10044 14243 10047
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 14231 10016 15393 10044
rect 14231 10013 14243 10016
rect 14185 10007 14243 10013
rect 15381 10013 15393 10016
rect 15427 10044 15439 10047
rect 15930 10044 15936 10056
rect 15427 10016 15936 10044
rect 15427 10013 15439 10016
rect 15381 10007 15439 10013
rect 15930 10004 15936 10016
rect 15988 10044 15994 10056
rect 16025 10047 16083 10053
rect 16025 10044 16037 10047
rect 15988 10016 16037 10044
rect 15988 10004 15994 10016
rect 16025 10013 16037 10016
rect 16071 10013 16083 10047
rect 16132 10044 16160 10084
rect 17954 10072 17960 10124
rect 18012 10112 18018 10124
rect 18012 10084 18736 10112
rect 18012 10072 18018 10084
rect 16281 10047 16339 10053
rect 16281 10044 16293 10047
rect 16132 10016 16293 10044
rect 16025 10007 16083 10013
rect 16281 10013 16293 10016
rect 16327 10013 16339 10047
rect 18414 10044 18420 10056
rect 18375 10016 18420 10044
rect 16281 10007 16339 10013
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 18708 10053 18736 10084
rect 19518 10072 19524 10124
rect 19576 10112 19582 10124
rect 20073 10115 20131 10121
rect 20073 10112 20085 10115
rect 19576 10084 20085 10112
rect 19576 10072 19582 10084
rect 20073 10081 20085 10084
rect 20119 10081 20131 10115
rect 20530 10112 20536 10124
rect 20443 10084 20536 10112
rect 20073 10075 20131 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 20809 10115 20867 10121
rect 20809 10081 20821 10115
rect 20855 10112 20867 10115
rect 21082 10112 21088 10124
rect 20855 10084 21088 10112
rect 20855 10081 20867 10084
rect 20809 10075 20867 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 18693 10047 18751 10053
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 18782 10044 18788 10056
rect 18739 10016 18788 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18782 10004 18788 10016
rect 18840 10004 18846 10056
rect 19889 10047 19947 10053
rect 19889 10013 19901 10047
rect 19935 10044 19947 10047
rect 20622 10044 20628 10056
rect 19935 10016 20628 10044
rect 19935 10013 19947 10016
rect 19889 10007 19947 10013
rect 20622 10004 20628 10016
rect 20680 10004 20686 10056
rect 12406 9979 12464 9985
rect 12406 9976 12418 9979
rect 9646 9939 9704 9945
rect 9784 9948 11376 9976
rect 12268 9948 12418 9976
rect 9784 9908 9812 9948
rect 11238 9908 11244 9920
rect 9140 9880 9812 9908
rect 11199 9880 11244 9908
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11348 9908 11376 9948
rect 12406 9945 12418 9948
rect 12452 9945 12464 9979
rect 14090 9976 14096 9988
rect 12406 9939 12464 9945
rect 13484 9948 14096 9976
rect 13484 9908 13512 9948
rect 14090 9936 14096 9948
rect 14148 9976 14154 9988
rect 14458 9976 14464 9988
rect 14148 9948 14464 9976
rect 14148 9936 14154 9948
rect 14458 9936 14464 9948
rect 14516 9936 14522 9988
rect 15013 9979 15071 9985
rect 15013 9945 15025 9979
rect 15059 9976 15071 9979
rect 20162 9976 20168 9988
rect 15059 9948 20168 9976
rect 15059 9945 15071 9948
rect 15013 9939 15071 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 11348 9880 13512 9908
rect 13541 9911 13599 9917
rect 13541 9877 13553 9911
rect 13587 9908 13599 9911
rect 13814 9908 13820 9920
rect 13587 9880 13820 9908
rect 13587 9877 13599 9880
rect 13541 9871 13599 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 17402 9908 17408 9920
rect 17363 9880 17408 9908
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 17586 9868 17592 9920
rect 17644 9908 17650 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 17644 9880 18245 9908
rect 17644 9868 17650 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18233 9871 18291 9877
rect 18877 9911 18935 9917
rect 18877 9877 18889 9911
rect 18923 9908 18935 9911
rect 19794 9908 19800 9920
rect 18923 9880 19800 9908
rect 18923 9877 18935 9880
rect 18877 9871 18935 9877
rect 19794 9868 19800 9880
rect 19852 9868 19858 9920
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20036 9880 20081 9908
rect 20036 9868 20042 9880
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 2406 9704 2412 9716
rect 2367 9676 2412 9704
rect 2406 9664 2412 9676
rect 2464 9664 2470 9716
rect 3878 9704 3884 9716
rect 2700 9676 3884 9704
rect 2038 9568 2044 9580
rect 1951 9540 2044 9568
rect 2038 9528 2044 9540
rect 2096 9568 2102 9580
rect 2222 9568 2228 9580
rect 2096 9540 2228 9568
rect 2096 9528 2102 9540
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2406 9528 2412 9580
rect 2464 9568 2470 9580
rect 2700 9568 2728 9676
rect 3878 9664 3884 9676
rect 3936 9704 3942 9716
rect 3936 9676 4384 9704
rect 3936 9664 3942 9676
rect 3050 9596 3056 9648
rect 3108 9596 3114 9648
rect 3694 9596 3700 9648
rect 3752 9636 3758 9648
rect 4356 9645 4384 9676
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 7285 9707 7343 9713
rect 7285 9704 7297 9707
rect 6972 9676 7297 9704
rect 6972 9664 6978 9676
rect 7285 9673 7297 9676
rect 7331 9673 7343 9707
rect 7285 9667 7343 9673
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 8110 9704 8116 9716
rect 7616 9676 8116 9704
rect 7616 9664 7622 9676
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 9030 9664 9036 9716
rect 9088 9704 9094 9716
rect 9088 9676 16528 9704
rect 9088 9664 9094 9676
rect 4341 9639 4399 9645
rect 3752 9608 4292 9636
rect 3752 9596 3758 9608
rect 3068 9568 3096 9596
rect 3237 9571 3295 9577
rect 3237 9568 3249 9571
rect 2464 9540 2728 9568
rect 2884 9540 3249 9568
rect 2464 9528 2470 9540
rect 1857 9503 1915 9509
rect 1857 9469 1869 9503
rect 1903 9469 1915 9503
rect 1857 9463 1915 9469
rect 1949 9503 2007 9509
rect 1949 9469 1961 9503
rect 1995 9500 2007 9503
rect 2884 9500 2912 9540
rect 3237 9537 3249 9540
rect 3283 9568 3295 9571
rect 4154 9568 4160 9580
rect 3283 9540 4160 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 4154 9528 4160 9540
rect 4212 9528 4218 9580
rect 4264 9568 4292 9608
rect 4341 9605 4353 9639
rect 4387 9636 4399 9639
rect 4387 9608 4421 9636
rect 4387 9605 4399 9608
rect 4341 9599 4399 9605
rect 4890 9596 4896 9648
rect 4948 9636 4954 9648
rect 5902 9636 5908 9648
rect 4948 9608 5908 9636
rect 4948 9596 4954 9608
rect 5902 9596 5908 9608
rect 5960 9596 5966 9648
rect 6638 9596 6644 9648
rect 6696 9636 6702 9648
rect 7377 9639 7435 9645
rect 7377 9636 7389 9639
rect 6696 9608 7389 9636
rect 6696 9596 6702 9608
rect 7377 9605 7389 9608
rect 7423 9636 7435 9639
rect 8294 9636 8300 9648
rect 7423 9608 8300 9636
rect 7423 9605 7435 9608
rect 7377 9599 7435 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9306 9645 9312 9648
rect 9248 9639 9312 9645
rect 9248 9605 9260 9639
rect 9294 9605 9312 9639
rect 9248 9599 9312 9605
rect 9306 9596 9312 9599
rect 9364 9596 9370 9648
rect 9858 9596 9864 9648
rect 9916 9636 9922 9648
rect 10014 9639 10072 9645
rect 10014 9636 10026 9639
rect 9916 9608 10026 9636
rect 9916 9596 9922 9608
rect 10014 9605 10026 9608
rect 10060 9636 10072 9639
rect 10778 9636 10784 9648
rect 10060 9608 10784 9636
rect 10060 9605 10072 9608
rect 10014 9599 10072 9605
rect 10778 9596 10784 9608
rect 10836 9596 10842 9648
rect 11238 9596 11244 9648
rect 11296 9636 11302 9648
rect 11514 9636 11520 9648
rect 11296 9608 11520 9636
rect 11296 9596 11302 9608
rect 11514 9596 11520 9608
rect 11572 9636 11578 9648
rect 11572 9608 12112 9636
rect 11572 9596 11578 9608
rect 4433 9571 4491 9577
rect 4433 9568 4445 9571
rect 4264 9540 4445 9568
rect 4433 9537 4445 9540
rect 4479 9568 4491 9571
rect 4614 9568 4620 9580
rect 4479 9540 4620 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 5537 9571 5595 9577
rect 5537 9537 5549 9571
rect 5583 9568 5595 9571
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5583 9540 6377 9568
rect 5583 9537 5595 9540
rect 5537 9531 5595 9537
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 12084 9568 12112 9608
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 13050 9639 13108 9645
rect 13050 9636 13062 9639
rect 12492 9608 13062 9636
rect 12492 9596 12498 9608
rect 13050 9605 13062 9608
rect 13096 9636 13108 9639
rect 13722 9636 13728 9648
rect 13096 9608 13728 9636
rect 13096 9605 13108 9608
rect 13050 9599 13108 9605
rect 13722 9596 13728 9608
rect 13780 9596 13786 9648
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 15666 9639 15724 9645
rect 15666 9636 15678 9639
rect 13872 9608 15678 9636
rect 13872 9596 13878 9608
rect 15666 9605 15678 9608
rect 15712 9605 15724 9639
rect 16500 9636 16528 9676
rect 17402 9664 17408 9716
rect 17460 9704 17466 9716
rect 20990 9704 20996 9716
rect 17460 9676 20996 9704
rect 17460 9664 17466 9676
rect 20990 9664 20996 9676
rect 21048 9664 21054 9716
rect 15666 9599 15724 9605
rect 15764 9608 16436 9636
rect 16500 9608 20852 9636
rect 12805 9571 12863 9577
rect 12805 9568 12817 9571
rect 8720 9540 12020 9568
rect 12084 9540 12817 9568
rect 8720 9528 8726 9540
rect 3050 9500 3056 9512
rect 1995 9472 2912 9500
rect 3011 9472 3056 9500
rect 1995 9469 2007 9472
rect 1949 9463 2007 9469
rect 1872 9432 1900 9463
rect 3050 9460 3056 9472
rect 3108 9460 3114 9512
rect 3145 9503 3203 9509
rect 3145 9469 3157 9503
rect 3191 9500 3203 9503
rect 3326 9500 3332 9512
rect 3191 9472 3332 9500
rect 3191 9469 3203 9472
rect 3145 9463 3203 9469
rect 3326 9460 3332 9472
rect 3384 9500 3390 9512
rect 3970 9500 3976 9512
rect 3384 9472 3976 9500
rect 3384 9460 3390 9472
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4246 9500 4252 9512
rect 4207 9472 4252 9500
rect 4246 9460 4252 9472
rect 4304 9460 4310 9512
rect 5166 9460 5172 9512
rect 5224 9500 5230 9512
rect 5261 9503 5319 9509
rect 5261 9500 5273 9503
rect 5224 9472 5273 9500
rect 5224 9460 5230 9472
rect 5261 9469 5273 9472
rect 5307 9469 5319 9503
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 5261 9463 5319 9469
rect 2774 9432 2780 9444
rect 1872 9404 2780 9432
rect 2774 9392 2780 9404
rect 2832 9432 2838 9444
rect 4062 9432 4068 9444
rect 2832 9404 4068 9432
rect 2832 9392 2838 9404
rect 4062 9392 4068 9404
rect 4120 9392 4126 9444
rect 4522 9392 4528 9444
rect 4580 9432 4586 9444
rect 4801 9435 4859 9441
rect 4801 9432 4813 9435
rect 4580 9404 4813 9432
rect 4580 9392 4586 9404
rect 4801 9401 4813 9404
rect 4847 9401 4859 9435
rect 5276 9432 5304 9463
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6730 9500 6736 9512
rect 5868 9472 6736 9500
rect 5868 9460 5874 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7561 9503 7619 9509
rect 7561 9469 7573 9503
rect 7607 9500 7619 9503
rect 8294 9500 8300 9512
rect 7607 9472 8300 9500
rect 7607 9469 7619 9472
rect 7561 9463 7619 9469
rect 7576 9432 7604 9463
rect 8294 9460 8300 9472
rect 8352 9460 8358 9512
rect 9490 9500 9496 9512
rect 9451 9472 9496 9500
rect 9490 9460 9496 9472
rect 9548 9500 9554 9512
rect 9769 9503 9827 9509
rect 9769 9500 9781 9503
rect 9548 9472 9781 9500
rect 9548 9460 9554 9472
rect 9769 9469 9781 9472
rect 9815 9469 9827 9503
rect 9769 9463 9827 9469
rect 5276 9404 7604 9432
rect 4801 9395 4859 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 11149 9435 11207 9441
rect 11149 9432 11161 9435
rect 11112 9404 11161 9432
rect 11112 9392 11118 9404
rect 11149 9401 11161 9404
rect 11195 9401 11207 9435
rect 11149 9395 11207 9401
rect 3602 9364 3608 9376
rect 3563 9336 3608 9364
rect 3602 9324 3608 9336
rect 3660 9324 3666 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 5534 9364 5540 9376
rect 4028 9336 5540 9364
rect 4028 9324 4034 9336
rect 5534 9324 5540 9336
rect 5592 9324 5598 9376
rect 5905 9367 5963 9373
rect 5905 9333 5917 9367
rect 5951 9364 5963 9367
rect 6638 9364 6644 9376
rect 5951 9336 6644 9364
rect 5951 9333 5963 9336
rect 5905 9327 5963 9333
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 6917 9367 6975 9373
rect 6917 9364 6929 9367
rect 6788 9336 6929 9364
rect 6788 9324 6794 9336
rect 6917 9333 6929 9336
rect 6963 9333 6975 9367
rect 6917 9327 6975 9333
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 11238 9364 11244 9376
rect 8260 9336 11244 9364
rect 8260 9324 8266 9336
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 11514 9364 11520 9376
rect 11475 9336 11520 9364
rect 11514 9324 11520 9336
rect 11572 9324 11578 9376
rect 11992 9373 12020 9540
rect 12805 9537 12817 9540
rect 12851 9537 12863 9571
rect 15764 9568 15792 9608
rect 15930 9568 15936 9580
rect 12805 9531 12863 9537
rect 12912 9540 15792 9568
rect 15891 9540 15936 9568
rect 12529 9503 12587 9509
rect 12529 9469 12541 9503
rect 12575 9500 12587 9503
rect 12912 9500 12940 9540
rect 15930 9528 15936 9540
rect 15988 9568 15994 9580
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 15988 9540 16221 9568
rect 15988 9528 15994 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16408 9568 16436 9608
rect 17770 9568 17776 9580
rect 16408 9540 17776 9568
rect 16209 9531 16267 9537
rect 17770 9528 17776 9540
rect 17828 9528 17834 9580
rect 17862 9528 17868 9580
rect 17920 9568 17926 9580
rect 19070 9571 19128 9577
rect 19070 9568 19082 9571
rect 17920 9540 19082 9568
rect 17920 9528 17926 9540
rect 19070 9537 19082 9540
rect 19116 9537 19128 9571
rect 19070 9531 19128 9537
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 20162 9568 20168 9580
rect 19300 9540 19840 9568
rect 20123 9540 20168 9568
rect 19300 9528 19306 9540
rect 12575 9472 12940 9500
rect 16945 9503 17003 9509
rect 12575 9469 12587 9472
rect 12529 9463 12587 9469
rect 16945 9469 16957 9503
rect 16991 9500 17003 9503
rect 17954 9500 17960 9512
rect 16991 9472 17960 9500
rect 16991 9469 17003 9472
rect 16945 9463 17003 9469
rect 17954 9460 17960 9472
rect 18012 9460 18018 9512
rect 19337 9503 19395 9509
rect 19337 9469 19349 9503
rect 19383 9469 19395 9503
rect 19702 9500 19708 9512
rect 19663 9472 19708 9500
rect 19337 9463 19395 9469
rect 14090 9392 14096 9444
rect 14148 9432 14154 9444
rect 14185 9435 14243 9441
rect 14185 9432 14197 9435
rect 14148 9404 14197 9432
rect 14148 9392 14154 9404
rect 14185 9401 14197 9404
rect 14231 9401 14243 9435
rect 14550 9432 14556 9444
rect 14511 9404 14556 9432
rect 14185 9395 14243 9401
rect 14550 9392 14556 9404
rect 14608 9392 14614 9444
rect 19352 9432 19380 9463
rect 19702 9460 19708 9472
rect 19760 9460 19766 9512
rect 19812 9500 19840 9540
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20824 9577 20852 9608
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 20530 9500 20536 9512
rect 19812 9472 20536 9500
rect 20530 9460 20536 9472
rect 20588 9460 20594 9512
rect 20714 9432 20720 9444
rect 15948 9404 18092 9432
rect 19352 9404 20720 9432
rect 11977 9367 12035 9373
rect 11977 9333 11989 9367
rect 12023 9364 12035 9367
rect 14458 9364 14464 9376
rect 12023 9336 14464 9364
rect 12023 9333 12035 9336
rect 11977 9327 12035 9333
rect 14458 9324 14464 9336
rect 14516 9324 14522 9376
rect 14918 9324 14924 9376
rect 14976 9364 14982 9376
rect 15948 9364 15976 9404
rect 14976 9336 15976 9364
rect 14976 9324 14982 9336
rect 17034 9324 17040 9376
rect 17092 9364 17098 9376
rect 17313 9367 17371 9373
rect 17313 9364 17325 9367
rect 17092 9336 17325 9364
rect 17092 9324 17098 9336
rect 17313 9333 17325 9336
rect 17359 9364 17371 9367
rect 17494 9364 17500 9376
rect 17359 9336 17500 9364
rect 17359 9333 17371 9336
rect 17313 9327 17371 9333
rect 17494 9324 17500 9336
rect 17552 9324 17558 9376
rect 17862 9324 17868 9376
rect 17920 9364 17926 9376
rect 17957 9367 18015 9373
rect 17957 9364 17969 9367
rect 17920 9336 17969 9364
rect 17920 9324 17926 9336
rect 17957 9333 17969 9336
rect 18003 9333 18015 9367
rect 18064 9364 18092 9404
rect 20714 9392 20720 9404
rect 20772 9432 20778 9444
rect 21174 9432 21180 9444
rect 20772 9404 21180 9432
rect 20772 9392 20778 9404
rect 21174 9392 21180 9404
rect 21232 9392 21238 9444
rect 20073 9367 20131 9373
rect 20073 9364 20085 9367
rect 18064 9336 20085 9364
rect 17957 9327 18015 9333
rect 20073 9333 20085 9336
rect 20119 9333 20131 9367
rect 20073 9327 20131 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2593 9163 2651 9169
rect 2593 9129 2605 9163
rect 2639 9160 2651 9163
rect 2774 9160 2780 9172
rect 2639 9132 2780 9160
rect 2639 9129 2651 9132
rect 2593 9123 2651 9129
rect 2774 9120 2780 9132
rect 2832 9120 2838 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 5442 9160 5448 9172
rect 4019 9132 5448 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 5442 9120 5448 9132
rect 5500 9120 5506 9172
rect 10042 9160 10048 9172
rect 8680 9132 10048 9160
rect 2222 9052 2228 9104
rect 2280 9052 2286 9104
rect 3329 9095 3387 9101
rect 3329 9061 3341 9095
rect 3375 9092 3387 9095
rect 3878 9092 3884 9104
rect 3375 9064 3884 9092
rect 3375 9061 3387 9064
rect 3329 9055 3387 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4062 9052 4068 9104
rect 4120 9092 4126 9104
rect 4798 9092 4804 9104
rect 4120 9064 4804 9092
rect 4120 9052 4126 9064
rect 4798 9052 4804 9064
rect 4856 9052 4862 9104
rect 8680 9092 8708 9132
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10778 9160 10784 9172
rect 10739 9132 10784 9160
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 13722 9160 13728 9172
rect 10928 9132 13584 9160
rect 13683 9132 13728 9160
rect 10928 9120 10934 9132
rect 5460 9064 8708 9092
rect 13556 9092 13584 9132
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 15930 9160 15936 9172
rect 15764 9132 15936 9160
rect 15102 9092 15108 9104
rect 13556 9064 15108 9092
rect 1578 8984 1584 9036
rect 1636 9024 1642 9036
rect 1949 9027 2007 9033
rect 1949 9024 1961 9027
rect 1636 8996 1961 9024
rect 1636 8984 1642 8996
rect 1949 8993 1961 8996
rect 1995 8993 2007 9027
rect 2240 9024 2268 9052
rect 5460 9033 5488 9064
rect 15102 9052 15108 9064
rect 15160 9052 15166 9104
rect 4341 9027 4399 9033
rect 2240 8996 3832 9024
rect 1949 8987 2007 8993
rect 2130 8916 2136 8968
rect 2188 8956 2194 8968
rect 2225 8959 2283 8965
rect 2225 8956 2237 8959
rect 2188 8928 2237 8956
rect 2188 8916 2194 8928
rect 2225 8925 2237 8928
rect 2271 8925 2283 8959
rect 3142 8956 3148 8968
rect 3103 8928 3148 8956
rect 2225 8919 2283 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3804 8965 3832 8996
rect 4341 8993 4353 9027
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 5445 9027 5503 9033
rect 5445 8993 5457 9027
rect 5491 8993 5503 9027
rect 5445 8987 5503 8993
rect 5537 9027 5595 9033
rect 5537 8993 5549 9027
rect 5583 9024 5595 9027
rect 5626 9024 5632 9036
rect 5583 8996 5632 9024
rect 5583 8993 5595 8996
rect 5537 8987 5595 8993
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 4246 8956 4252 8968
rect 3835 8928 4252 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 1762 8848 1768 8900
rect 1820 8888 1826 8900
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 1820 8860 2697 8888
rect 1820 8848 1826 8860
rect 2685 8857 2697 8860
rect 2731 8857 2743 8891
rect 2685 8851 2743 8857
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 4356 8888 4384 8987
rect 5626 8984 5632 8996
rect 5684 8984 5690 9036
rect 6730 9024 6736 9036
rect 6691 8996 6736 9024
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 8202 9024 8208 9036
rect 8163 8996 8208 9024
rect 6825 8987 6883 8993
rect 4430 8916 4436 8968
rect 4488 8956 4494 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4488 8928 4629 8956
rect 4488 8916 4494 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 4617 8919 4675 8925
rect 5718 8916 5724 8968
rect 5776 8956 5782 8968
rect 6638 8956 6644 8968
rect 5776 8928 6500 8956
rect 6599 8928 6644 8956
rect 5776 8916 5782 8928
rect 5534 8888 5540 8900
rect 3108 8860 4108 8888
rect 4356 8860 5540 8888
rect 3108 8848 3114 8860
rect 2222 8780 2228 8832
rect 2280 8820 2286 8832
rect 3970 8820 3976 8832
rect 2280 8792 3976 8820
rect 2280 8780 2286 8792
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 4080 8820 4108 8860
rect 5534 8848 5540 8860
rect 5592 8848 5598 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 6472 8888 6500 8928
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 6840 8900 6868 8987
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 11698 8984 11704 9036
rect 11756 9024 11762 9036
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11756 8996 11989 9024
rect 11756 8984 11762 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 13814 8984 13820 9036
rect 13872 9024 13878 9036
rect 15764 9033 15792 9132
rect 15930 9120 15936 9132
rect 15988 9120 15994 9172
rect 16114 9120 16120 9172
rect 16172 9160 16178 9172
rect 17405 9163 17463 9169
rect 17405 9160 17417 9163
rect 16172 9132 17417 9160
rect 16172 9120 16178 9132
rect 17405 9129 17417 9132
rect 17451 9129 17463 9163
rect 17405 9123 17463 9129
rect 17770 9120 17776 9172
rect 17828 9160 17834 9172
rect 17828 9132 19932 9160
rect 17828 9120 17834 9132
rect 19904 9092 19932 9132
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20036 9132 20453 9160
rect 20036 9120 20042 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 21266 9092 21272 9104
rect 19904 9064 21272 9092
rect 21266 9052 21272 9064
rect 21324 9052 21330 9104
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13872 8996 14197 9024
rect 13872 8984 13878 8996
rect 14185 8993 14197 8996
rect 14231 9024 14243 9027
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14231 8996 14565 9024
rect 14231 8993 14243 8996
rect 14185 8987 14243 8993
rect 14553 8993 14565 8996
rect 14599 9024 14611 9027
rect 15749 9027 15807 9033
rect 15749 9024 15761 9027
rect 14599 8996 15761 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 15749 8993 15761 8996
rect 15795 8993 15807 9027
rect 17770 9024 17776 9036
rect 15749 8987 15807 8993
rect 17328 8996 17776 9024
rect 7929 8959 7987 8965
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8018 8956 8024 8968
rect 7975 8928 8024 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 9401 8959 9459 8965
rect 9401 8925 9413 8959
rect 9447 8956 9459 8959
rect 9490 8956 9496 8968
rect 9447 8928 9496 8956
rect 9447 8925 9459 8928
rect 9401 8919 9459 8925
rect 9490 8916 9496 8928
rect 9548 8956 9554 8968
rect 11514 8956 11520 8968
rect 9548 8928 11520 8956
rect 9548 8916 9554 8928
rect 6822 8888 6828 8900
rect 5675 8860 6316 8888
rect 6472 8860 6828 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 4338 8820 4344 8832
rect 4080 8792 4344 8820
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5718 8820 5724 8832
rect 5031 8792 5724 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5902 8780 5908 8832
rect 5960 8820 5966 8832
rect 6288 8829 6316 8860
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 9646 8891 9704 8897
rect 9646 8888 9658 8891
rect 8168 8860 9658 8888
rect 8168 8848 8174 8860
rect 9646 8857 9658 8860
rect 9692 8857 9704 8891
rect 10962 8888 10968 8900
rect 9646 8851 9704 8857
rect 10888 8860 10968 8888
rect 5997 8823 6055 8829
rect 5997 8820 6009 8823
rect 5960 8792 6009 8820
rect 5960 8780 5966 8792
rect 5997 8789 6009 8792
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8789 6331 8823
rect 6273 8783 6331 8789
rect 7098 8780 7104 8832
rect 7156 8820 7162 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 7156 8792 7573 8820
rect 7156 8780 7162 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 7742 8780 7748 8832
rect 7800 8820 7806 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7800 8792 8033 8820
rect 7800 8780 7806 8792
rect 8021 8789 8033 8792
rect 8067 8820 8079 8823
rect 8662 8820 8668 8832
rect 8067 8792 8668 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8662 8780 8668 8792
rect 8720 8820 8726 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8720 8792 8953 8820
rect 8720 8780 8726 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 10888 8820 10916 8860
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 11072 8832 11100 8928
rect 11514 8916 11520 8928
rect 11572 8956 11578 8968
rect 12345 8959 12403 8965
rect 12345 8956 12357 8959
rect 11572 8928 12357 8956
rect 11572 8916 11578 8928
rect 12345 8925 12357 8928
rect 12391 8925 12403 8959
rect 15286 8956 15292 8968
rect 15247 8928 15292 8956
rect 12345 8919 12403 8925
rect 15286 8916 15292 8928
rect 15344 8916 15350 8968
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 16005 8959 16063 8965
rect 16005 8956 16017 8959
rect 15528 8928 16017 8956
rect 15528 8916 15534 8928
rect 16005 8925 16017 8928
rect 16051 8925 16063 8959
rect 16005 8919 16063 8925
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 17328 8956 17356 8996
rect 17770 8984 17776 8996
rect 17828 8984 17834 9036
rect 19610 9024 19616 9036
rect 19571 8996 19616 9024
rect 19610 8984 19616 8996
rect 19668 8984 19674 9036
rect 19705 9027 19763 9033
rect 19705 8993 19717 9027
rect 19751 9024 19763 9027
rect 20806 9024 20812 9036
rect 19751 8996 20812 9024
rect 19751 8993 19763 8996
rect 19705 8987 19763 8993
rect 20806 8984 20812 8996
rect 20864 9024 20870 9036
rect 20901 9027 20959 9033
rect 20901 9024 20913 9027
rect 20864 8996 20913 9024
rect 20864 8984 20870 8996
rect 20901 8993 20913 8996
rect 20947 8993 20959 9027
rect 20901 8987 20959 8993
rect 20990 8984 20996 9036
rect 21048 9024 21054 9036
rect 21048 8996 21093 9024
rect 21048 8984 21054 8996
rect 16540 8928 17356 8956
rect 16540 8916 16546 8928
rect 17402 8916 17408 8968
rect 17460 8956 17466 8968
rect 18785 8959 18843 8965
rect 18785 8956 18797 8959
rect 17460 8928 18797 8956
rect 17460 8916 17466 8928
rect 18785 8925 18797 8928
rect 18831 8925 18843 8959
rect 18785 8919 18843 8925
rect 12590 8891 12648 8897
rect 12590 8888 12602 8891
rect 12360 8860 12602 8888
rect 12360 8832 12388 8860
rect 12590 8857 12602 8860
rect 12636 8857 12648 8891
rect 12590 8851 12648 8857
rect 15013 8891 15071 8897
rect 15013 8857 15025 8891
rect 15059 8888 15071 8891
rect 17862 8888 17868 8900
rect 15059 8860 17868 8888
rect 15059 8857 15071 8860
rect 15013 8851 15071 8857
rect 17862 8848 17868 8860
rect 17920 8848 17926 8900
rect 18518 8891 18576 8897
rect 18518 8888 18530 8891
rect 17972 8860 18530 8888
rect 11054 8820 11060 8832
rect 9088 8792 10916 8820
rect 11015 8792 11060 8820
rect 9088 8780 9094 8792
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 11701 8823 11759 8829
rect 11701 8789 11713 8823
rect 11747 8820 11759 8823
rect 12158 8820 12164 8832
rect 11747 8792 12164 8820
rect 11747 8789 11759 8792
rect 11701 8783 11759 8789
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12342 8780 12348 8832
rect 12400 8780 12406 8832
rect 12434 8780 12440 8832
rect 12492 8820 12498 8832
rect 15378 8820 15384 8832
rect 12492 8792 15384 8820
rect 12492 8780 12498 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15473 8823 15531 8829
rect 15473 8789 15485 8823
rect 15519 8820 15531 8823
rect 15746 8820 15752 8832
rect 15519 8792 15752 8820
rect 15519 8789 15531 8792
rect 15473 8783 15531 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16482 8820 16488 8832
rect 16264 8792 16488 8820
rect 16264 8780 16270 8792
rect 16482 8780 16488 8792
rect 16540 8780 16546 8832
rect 17034 8780 17040 8832
rect 17092 8820 17098 8832
rect 17129 8823 17187 8829
rect 17129 8820 17141 8823
rect 17092 8792 17141 8820
rect 17092 8780 17098 8792
rect 17129 8789 17141 8792
rect 17175 8789 17187 8823
rect 17129 8783 17187 8789
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17972 8820 18000 8860
rect 18518 8857 18530 8860
rect 18564 8857 18576 8891
rect 18966 8888 18972 8900
rect 18518 8851 18576 8857
rect 18616 8860 18972 8888
rect 17552 8792 18000 8820
rect 17552 8780 17558 8792
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18616 8820 18644 8860
rect 18966 8848 18972 8860
rect 19024 8888 19030 8900
rect 20809 8891 20867 8897
rect 20809 8888 20821 8891
rect 19024 8860 20821 8888
rect 19024 8848 19030 8860
rect 20809 8857 20821 8860
rect 20855 8857 20867 8891
rect 20809 8851 20867 8857
rect 18104 8792 18644 8820
rect 19797 8823 19855 8829
rect 18104 8780 18110 8792
rect 19797 8789 19809 8823
rect 19843 8820 19855 8823
rect 19978 8820 19984 8832
rect 19843 8792 19984 8820
rect 19843 8789 19855 8792
rect 19797 8783 19855 8789
rect 19978 8780 19984 8792
rect 20036 8780 20042 8832
rect 20162 8820 20168 8832
rect 20123 8792 20168 8820
rect 20162 8780 20168 8792
rect 20220 8780 20226 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2501 8619 2559 8625
rect 2501 8616 2513 8619
rect 2372 8588 2513 8616
rect 2372 8576 2378 8588
rect 2501 8585 2513 8588
rect 2547 8585 2559 8619
rect 2958 8616 2964 8628
rect 2919 8588 2964 8616
rect 2501 8579 2559 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4522 8616 4528 8628
rect 4483 8588 4528 8616
rect 4522 8576 4528 8588
rect 4580 8576 4586 8628
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5350 8576 5356 8628
rect 5408 8616 5414 8628
rect 7742 8616 7748 8628
rect 5408 8588 7748 8616
rect 5408 8576 5414 8588
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7892 8588 8033 8616
rect 7892 8576 7898 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 8481 8619 8539 8625
rect 8168 8588 8213 8616
rect 8168 8576 8174 8588
rect 8481 8585 8493 8619
rect 8527 8616 8539 8619
rect 8527 8588 12434 8616
rect 8527 8585 8539 8588
rect 8481 8579 8539 8585
rect 12406 8560 12434 8588
rect 12618 8576 12624 8628
rect 12676 8616 12682 8628
rect 12713 8619 12771 8625
rect 12713 8616 12725 8619
rect 12676 8588 12725 8616
rect 12676 8576 12682 8588
rect 12713 8585 12725 8588
rect 12759 8616 12771 8619
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 12759 8588 13461 8616
rect 12759 8585 12771 8588
rect 12713 8579 12771 8585
rect 13449 8585 13461 8588
rect 13495 8616 13507 8619
rect 13814 8616 13820 8628
rect 13495 8588 13820 8616
rect 13495 8585 13507 8588
rect 13449 8579 13507 8585
rect 13814 8576 13820 8588
rect 13872 8576 13878 8628
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15470 8616 15476 8628
rect 15252 8588 15476 8616
rect 15252 8576 15258 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 15841 8619 15899 8625
rect 15841 8585 15853 8619
rect 15887 8616 15899 8619
rect 15930 8616 15936 8628
rect 15887 8588 15936 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1636 8520 6776 8548
rect 1636 8508 1642 8520
rect 1946 8480 1952 8492
rect 1907 8452 1952 8480
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 2866 8480 2872 8492
rect 2827 8452 2872 8480
rect 2866 8440 2872 8452
rect 2924 8440 2930 8492
rect 6748 8480 6776 8520
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 9490 8548 9496 8560
rect 6880 8520 9496 8548
rect 6880 8508 6886 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 9950 8508 9956 8560
rect 10008 8548 10014 8560
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10008 8520 10793 8548
rect 10008 8508 10014 8520
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 10781 8511 10839 8517
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 11974 8548 11980 8560
rect 11020 8520 11376 8548
rect 11935 8520 11980 8548
rect 11020 8508 11026 8520
rect 6914 8480 6920 8492
rect 6748 8452 6920 8480
rect 6914 8440 6920 8452
rect 6972 8440 6978 8492
rect 8018 8440 8024 8492
rect 8076 8480 8082 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8076 8452 8769 8480
rect 8076 8440 8082 8452
rect 8757 8449 8769 8452
rect 8803 8480 8815 8483
rect 9030 8480 9036 8492
rect 8803 8452 9036 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 9030 8440 9036 8452
rect 9088 8440 9094 8492
rect 10045 8483 10103 8489
rect 10045 8449 10057 8483
rect 10091 8480 10103 8483
rect 11238 8480 11244 8492
rect 10091 8452 11244 8480
rect 10091 8449 10103 8452
rect 10045 8443 10103 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11348 8480 11376 8520
rect 11974 8508 11980 8520
rect 12032 8508 12038 8560
rect 12406 8520 12440 8560
rect 12434 8508 12440 8520
rect 12492 8508 12498 8560
rect 13081 8551 13139 8557
rect 13081 8517 13093 8551
rect 13127 8548 13139 8551
rect 15654 8548 15660 8560
rect 13127 8520 15660 8548
rect 13127 8517 13139 8520
rect 13081 8511 13139 8517
rect 15654 8508 15660 8520
rect 15712 8508 15718 8560
rect 12544 8480 12664 8484
rect 14918 8480 14924 8492
rect 11348 8456 14924 8480
rect 11348 8452 12572 8456
rect 12636 8452 14924 8456
rect 14918 8440 14924 8452
rect 14976 8440 14982 8492
rect 15194 8440 15200 8492
rect 15252 8489 15258 8492
rect 15252 8480 15264 8489
rect 15252 8452 15297 8480
rect 15252 8443 15264 8452
rect 15252 8440 15258 8443
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 15473 8483 15531 8489
rect 15473 8449 15485 8483
rect 15519 8480 15531 8483
rect 15856 8480 15884 8579
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 17405 8619 17463 8625
rect 17405 8585 17417 8619
rect 17451 8616 17463 8619
rect 18046 8616 18052 8628
rect 17451 8588 18052 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 18046 8576 18052 8588
rect 18104 8576 18110 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 19797 8619 19855 8625
rect 19797 8616 19809 8619
rect 18288 8588 19809 8616
rect 18288 8576 18294 8588
rect 19797 8585 19809 8588
rect 19843 8585 19855 8619
rect 19797 8579 19855 8585
rect 18874 8508 18880 8560
rect 18932 8548 18938 8560
rect 20910 8551 20968 8557
rect 20910 8548 20922 8551
rect 18932 8520 20922 8548
rect 18932 8508 18938 8520
rect 20910 8517 20922 8520
rect 20956 8517 20968 8551
rect 20910 8511 20968 8517
rect 15519 8452 15884 8480
rect 17221 8483 17279 8489
rect 15519 8449 15531 8452
rect 15473 8443 15531 8449
rect 17221 8449 17233 8483
rect 17267 8480 17279 8483
rect 17494 8480 17500 8492
rect 17267 8452 17500 8480
rect 17267 8449 17279 8452
rect 17221 8443 17279 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 17862 8480 17868 8492
rect 17727 8452 17868 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 17862 8440 17868 8452
rect 17920 8440 17926 8492
rect 18046 8440 18052 8492
rect 18104 8480 18110 8492
rect 18397 8483 18455 8489
rect 18397 8480 18409 8483
rect 18104 8452 18409 8480
rect 18104 8440 18110 8452
rect 18397 8449 18409 8452
rect 18443 8449 18455 8483
rect 21174 8480 21180 8492
rect 21135 8452 21180 8480
rect 18397 8443 18455 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2682 8372 2688 8424
rect 2740 8412 2746 8424
rect 3053 8415 3111 8421
rect 2740 8384 2912 8412
rect 2740 8372 2746 8384
rect 2884 8344 2912 8384
rect 3053 8381 3065 8415
rect 3099 8381 3111 8415
rect 3053 8375 3111 8381
rect 3068 8344 3096 8375
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 3200 8384 3525 8412
rect 3200 8372 3206 8384
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 4982 8412 4988 8424
rect 4895 8384 4988 8412
rect 3513 8375 3571 8381
rect 4982 8372 4988 8384
rect 5040 8372 5046 8424
rect 5166 8412 5172 8424
rect 5127 8384 5172 8412
rect 5166 8372 5172 8384
rect 5224 8372 5230 8424
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8412 6055 8415
rect 7558 8412 7564 8424
rect 6043 8384 7564 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 7558 8372 7564 8384
rect 7616 8372 7622 8424
rect 7929 8415 7987 8421
rect 7929 8381 7941 8415
rect 7975 8412 7987 8415
rect 10870 8412 10876 8424
rect 7975 8384 10876 8412
rect 7975 8381 7987 8384
rect 7929 8375 7987 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11330 8372 11336 8424
rect 11388 8412 11394 8424
rect 11974 8412 11980 8424
rect 11388 8384 11980 8412
rect 11388 8372 11394 8384
rect 11974 8372 11980 8384
rect 12032 8412 12038 8424
rect 15396 8412 15424 8440
rect 12032 8384 14136 8412
rect 15396 8384 16896 8412
rect 12032 8372 12038 8384
rect 2884 8316 3096 8344
rect 3878 8304 3884 8356
rect 3936 8344 3942 8356
rect 4062 8344 4068 8356
rect 3936 8316 4068 8344
rect 3936 8304 3942 8316
rect 4062 8304 4068 8316
rect 4120 8344 4126 8356
rect 4157 8347 4215 8353
rect 4157 8344 4169 8347
rect 4120 8316 4169 8344
rect 4120 8304 4126 8316
rect 4157 8313 4169 8316
rect 4203 8313 4215 8347
rect 5000 8344 5028 8372
rect 5629 8347 5687 8353
rect 5629 8344 5641 8347
rect 5000 8316 5641 8344
rect 4157 8307 4215 8313
rect 5629 8313 5641 8316
rect 5675 8344 5687 8347
rect 6457 8347 6515 8353
rect 5675 8316 6408 8344
rect 5675 8313 5687 8316
rect 5629 8307 5687 8313
rect 3510 8236 3516 8288
rect 3568 8276 3574 8288
rect 4614 8276 4620 8288
rect 3568 8248 4620 8276
rect 3568 8236 3574 8248
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 6380 8276 6408 8316
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 6546 8344 6552 8356
rect 6503 8316 6552 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6546 8304 6552 8316
rect 6604 8304 6610 8356
rect 6825 8347 6883 8353
rect 6825 8313 6837 8347
rect 6871 8344 6883 8347
rect 6914 8344 6920 8356
rect 6871 8316 6920 8344
rect 6871 8313 6883 8316
rect 6825 8307 6883 8313
rect 6914 8304 6920 8316
rect 6972 8304 6978 8356
rect 7469 8347 7527 8353
rect 7469 8313 7481 8347
rect 7515 8344 7527 8347
rect 7650 8344 7656 8356
rect 7515 8316 7656 8344
rect 7515 8313 7527 8316
rect 7469 8307 7527 8313
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 7760 8316 8616 8344
rect 7760 8276 7788 8316
rect 6380 8248 7788 8276
rect 8588 8276 8616 8316
rect 8662 8304 8668 8356
rect 8720 8344 8726 8356
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 8720 8316 9137 8344
rect 8720 8304 8726 8316
rect 9125 8313 9137 8316
rect 9171 8313 9183 8347
rect 9125 8307 9183 8313
rect 9677 8347 9735 8353
rect 9677 8313 9689 8347
rect 9723 8344 9735 8347
rect 10505 8347 10563 8353
rect 10505 8344 10517 8347
rect 9723 8316 10517 8344
rect 9723 8313 9735 8316
rect 9677 8307 9735 8313
rect 10505 8313 10517 8316
rect 10551 8344 10563 8347
rect 11054 8344 11060 8356
rect 10551 8316 11060 8344
rect 10551 8313 10563 8316
rect 10505 8307 10563 8313
rect 11054 8304 11060 8316
rect 11112 8344 11118 8356
rect 11517 8347 11575 8353
rect 11517 8344 11529 8347
rect 11112 8316 11529 8344
rect 11112 8304 11118 8316
rect 11517 8313 11529 8316
rect 11563 8344 11575 8347
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 11563 8316 12265 8344
rect 11563 8313 11575 8316
rect 11517 8307 11575 8313
rect 12253 8313 12265 8316
rect 12299 8344 12311 8347
rect 12434 8344 12440 8356
rect 12299 8316 12440 8344
rect 12299 8313 12311 8316
rect 12253 8307 12311 8313
rect 12434 8304 12440 8316
rect 12492 8344 12498 8356
rect 12618 8344 12624 8356
rect 12492 8316 12624 8344
rect 12492 8304 12498 8316
rect 12618 8304 12624 8316
rect 12676 8304 12682 8356
rect 14108 8353 14136 8384
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 15470 8304 15476 8356
rect 15528 8344 15534 8356
rect 15838 8344 15844 8356
rect 15528 8316 15844 8344
rect 15528 8304 15534 8316
rect 15838 8304 15844 8316
rect 15896 8344 15902 8356
rect 16114 8344 16120 8356
rect 15896 8316 16120 8344
rect 15896 8304 15902 8316
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16868 8344 16896 8384
rect 17402 8372 17408 8424
rect 17460 8412 17466 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 17460 8384 18153 8412
rect 17460 8372 17466 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 16868 8316 17724 8344
rect 15562 8276 15568 8288
rect 8588 8248 15568 8276
rect 15562 8236 15568 8248
rect 15620 8236 15626 8288
rect 16945 8279 17003 8285
rect 16945 8245 16957 8279
rect 16991 8276 17003 8279
rect 17402 8276 17408 8288
rect 16991 8248 17408 8276
rect 16991 8245 17003 8248
rect 16945 8239 17003 8245
rect 17402 8236 17408 8248
rect 17460 8236 17466 8288
rect 17696 8276 17724 8316
rect 17770 8304 17776 8356
rect 17828 8344 17834 8356
rect 17865 8347 17923 8353
rect 17865 8344 17877 8347
rect 17828 8316 17877 8344
rect 17828 8304 17834 8316
rect 17865 8313 17877 8316
rect 17911 8313 17923 8347
rect 17865 8307 17923 8313
rect 19058 8276 19064 8288
rect 17696 8248 19064 8276
rect 19058 8236 19064 8248
rect 19116 8236 19122 8288
rect 19521 8279 19579 8285
rect 19521 8245 19533 8279
rect 19567 8276 19579 8279
rect 19610 8276 19616 8288
rect 19567 8248 19616 8276
rect 19567 8245 19579 8248
rect 19521 8239 19579 8245
rect 19610 8236 19616 8248
rect 19668 8236 19674 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2225 8075 2283 8081
rect 2225 8041 2237 8075
rect 2271 8072 2283 8075
rect 2774 8072 2780 8084
rect 2271 8044 2780 8072
rect 2271 8041 2283 8044
rect 2225 8035 2283 8041
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4985 8075 5043 8081
rect 4985 8072 4997 8075
rect 4304 8044 4997 8072
rect 4304 8032 4310 8044
rect 4985 8041 4997 8044
rect 5031 8041 5043 8075
rect 4985 8035 5043 8041
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6822 8072 6828 8084
rect 6604 8044 6828 8072
rect 6604 8032 6610 8044
rect 6822 8032 6828 8044
rect 6880 8032 6886 8084
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8754 8072 8760 8084
rect 8352 8044 8760 8072
rect 8352 8032 8358 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9582 8072 9588 8084
rect 8987 8044 9588 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10100 8044 10609 8072
rect 10100 8032 10106 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 14642 8032 14648 8084
rect 14700 8072 14706 8084
rect 15013 8075 15071 8081
rect 15013 8072 15025 8075
rect 14700 8044 15025 8072
rect 14700 8032 14706 8044
rect 15013 8041 15025 8044
rect 15059 8041 15071 8075
rect 15013 8035 15071 8041
rect 15841 8075 15899 8081
rect 15841 8041 15853 8075
rect 15887 8072 15899 8075
rect 15930 8072 15936 8084
rect 15887 8044 15936 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 16577 8075 16635 8081
rect 16577 8041 16589 8075
rect 16623 8072 16635 8075
rect 16942 8072 16948 8084
rect 16623 8044 16948 8072
rect 16623 8041 16635 8044
rect 16577 8035 16635 8041
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 18046 8072 18052 8084
rect 17052 8044 18052 8072
rect 4709 8007 4767 8013
rect 2700 7976 4476 8004
rect 1670 7936 1676 7948
rect 1631 7908 1676 7936
rect 1670 7896 1676 7908
rect 1728 7896 1734 7948
rect 2700 7945 2728 7976
rect 2685 7939 2743 7945
rect 2685 7905 2697 7939
rect 2731 7905 2743 7939
rect 4338 7936 4344 7948
rect 2685 7899 2743 7905
rect 2792 7908 4344 7936
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7868 1823 7871
rect 2792 7868 2820 7908
rect 4338 7896 4344 7908
rect 4396 7896 4402 7948
rect 4448 7936 4476 7976
rect 4709 7973 4721 8007
rect 4755 8004 4767 8007
rect 4890 8004 4896 8016
rect 4755 7976 4896 8004
rect 4755 7973 4767 7976
rect 4709 7967 4767 7973
rect 4890 7964 4896 7976
rect 4948 7964 4954 8016
rect 7653 8007 7711 8013
rect 5460 7976 7604 8004
rect 5166 7936 5172 7948
rect 4448 7908 5172 7936
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 1811 7840 2820 7868
rect 2869 7871 2927 7877
rect 1811 7837 1823 7840
rect 1765 7831 1823 7837
rect 2869 7837 2881 7871
rect 2915 7868 2927 7871
rect 3142 7868 3148 7880
rect 2915 7840 3148 7868
rect 2915 7837 2927 7840
rect 2869 7831 2927 7837
rect 3142 7828 3148 7840
rect 3200 7828 3206 7880
rect 3970 7868 3976 7880
rect 3931 7840 3976 7868
rect 3970 7828 3976 7840
rect 4028 7828 4034 7880
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7868 4307 7871
rect 4430 7868 4436 7880
rect 4295 7840 4436 7868
rect 4295 7837 4307 7840
rect 4249 7831 4307 7837
rect 4430 7828 4436 7840
rect 4488 7868 4494 7880
rect 5460 7868 5488 7976
rect 5537 7939 5595 7945
rect 5537 7905 5549 7939
rect 5583 7905 5595 7939
rect 5718 7936 5724 7948
rect 5679 7908 5724 7936
rect 5537 7899 5595 7905
rect 4488 7840 5488 7868
rect 5552 7868 5580 7899
rect 5718 7896 5724 7908
rect 5776 7896 5782 7948
rect 7098 7936 7104 7948
rect 7059 7908 7104 7936
rect 7098 7896 7104 7908
rect 7156 7896 7162 7948
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7905 7343 7939
rect 7576 7936 7604 7976
rect 7653 7973 7665 8007
rect 7699 8004 7711 8007
rect 7742 8004 7748 8016
rect 7699 7976 7748 8004
rect 7699 7973 7711 7976
rect 7653 7967 7711 7973
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 9030 7964 9036 8016
rect 9088 8004 9094 8016
rect 9214 8004 9220 8016
rect 9088 7976 9220 8004
rect 9088 7964 9094 7976
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 12860 7976 13001 8004
rect 12860 7964 12866 7976
rect 12989 7973 13001 7976
rect 13035 8004 13047 8007
rect 17052 8004 17080 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 18693 8075 18751 8081
rect 18693 8041 18705 8075
rect 18739 8072 18751 8075
rect 18782 8072 18788 8084
rect 18739 8044 18788 8072
rect 18739 8041 18751 8044
rect 18693 8035 18751 8041
rect 18782 8032 18788 8044
rect 18840 8032 18846 8084
rect 13035 7976 17080 8004
rect 13035 7973 13047 7976
rect 12989 7967 13047 7973
rect 17954 7964 17960 8016
rect 18012 8004 18018 8016
rect 19981 8007 20039 8013
rect 19981 8004 19993 8007
rect 18012 7976 19993 8004
rect 18012 7964 18018 7976
rect 19981 7973 19993 7976
rect 20027 7973 20039 8007
rect 19981 7967 20039 7973
rect 8294 7936 8300 7948
rect 7576 7908 8300 7936
rect 7285 7899 7343 7905
rect 7300 7868 7328 7899
rect 8294 7896 8300 7908
rect 8352 7936 8358 7948
rect 8352 7908 9352 7936
rect 8352 7896 8358 7908
rect 7834 7868 7840 7880
rect 5552 7840 7236 7868
rect 7300 7840 7840 7868
rect 4488 7828 4494 7840
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2777 7803 2835 7809
rect 2777 7800 2789 7803
rect 2188 7772 2789 7800
rect 2188 7760 2194 7772
rect 2777 7769 2789 7772
rect 2823 7769 2835 7803
rect 2777 7763 2835 7769
rect 3418 7760 3424 7812
rect 3476 7800 3482 7812
rect 3476 7772 6684 7800
rect 3476 7760 3482 7772
rect 1854 7692 1860 7744
rect 1912 7732 1918 7744
rect 3234 7732 3240 7744
rect 1912 7704 1957 7732
rect 3195 7704 3240 7732
rect 1912 7692 1918 7704
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 3384 7704 3801 7732
rect 3384 7692 3390 7704
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 5813 7735 5871 7741
rect 5813 7701 5825 7735
rect 5859 7732 5871 7735
rect 5994 7732 6000 7744
rect 5859 7704 6000 7732
rect 5859 7701 5871 7704
rect 5813 7695 5871 7701
rect 5994 7692 6000 7704
rect 6052 7692 6058 7744
rect 6181 7735 6239 7741
rect 6181 7701 6193 7735
rect 6227 7732 6239 7735
rect 6546 7732 6552 7744
rect 6227 7704 6552 7732
rect 6227 7701 6239 7704
rect 6181 7695 6239 7701
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6656 7741 6684 7772
rect 6641 7735 6699 7741
rect 6641 7701 6653 7735
rect 6687 7701 6699 7735
rect 7006 7732 7012 7744
rect 6967 7704 7012 7732
rect 6641 7695 6699 7701
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7208 7732 7236 7840
rect 7834 7828 7840 7840
rect 7892 7828 7898 7880
rect 9214 7868 9220 7880
rect 7944 7840 9220 7868
rect 7944 7732 7972 7840
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 9324 7868 9352 7908
rect 18414 7896 18420 7948
rect 18472 7936 18478 7948
rect 19242 7936 19248 7948
rect 18472 7908 19248 7936
rect 18472 7896 18478 7908
rect 19242 7896 19248 7908
rect 19300 7896 19306 7948
rect 19794 7896 19800 7948
rect 19852 7936 19858 7948
rect 20441 7939 20499 7945
rect 20441 7936 20453 7939
rect 19852 7908 20453 7936
rect 19852 7896 19858 7908
rect 20441 7905 20453 7908
rect 20487 7905 20499 7939
rect 20441 7899 20499 7905
rect 20533 7939 20591 7945
rect 20533 7905 20545 7939
rect 20579 7905 20591 7939
rect 20533 7899 20591 7905
rect 9324 7840 9444 7868
rect 8021 7803 8079 7809
rect 8021 7769 8033 7803
rect 8067 7800 8079 7803
rect 9306 7800 9312 7812
rect 8067 7772 9312 7800
rect 8067 7769 8079 7772
rect 8021 7763 8079 7769
rect 9306 7760 9312 7772
rect 9364 7760 9370 7812
rect 7208 7704 7972 7732
rect 8113 7735 8171 7741
rect 8113 7701 8125 7735
rect 8159 7732 8171 7735
rect 9122 7732 9128 7744
rect 8159 7704 9128 7732
rect 8159 7701 8171 7704
rect 8113 7695 8171 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9416 7732 9444 7840
rect 10042 7828 10048 7880
rect 10100 7877 10106 7880
rect 10100 7868 10112 7877
rect 10321 7871 10379 7877
rect 10100 7840 10145 7868
rect 10100 7831 10112 7840
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 10367 7840 11989 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 11977 7837 11989 7840
rect 12023 7868 12035 7871
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 12023 7840 12265 7868
rect 12023 7837 12035 7840
rect 11977 7831 12035 7837
rect 12253 7837 12265 7840
rect 12299 7868 12311 7871
rect 12342 7868 12348 7880
rect 12299 7840 12348 7868
rect 12299 7837 12311 7840
rect 12253 7831 12311 7837
rect 10100 7828 10106 7831
rect 12342 7828 12348 7840
rect 12400 7868 12406 7880
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 12400 7840 13645 7868
rect 12400 7828 12406 7840
rect 13633 7837 13645 7840
rect 13679 7837 13691 7871
rect 13633 7831 13691 7837
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 16942 7868 16948 7880
rect 15160 7840 16948 7868
rect 15160 7828 15166 7840
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 17402 7828 17408 7880
rect 17460 7868 17466 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17460 7840 17969 7868
rect 17460 7828 17466 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18506 7868 18512 7880
rect 18104 7840 18512 7868
rect 18104 7828 18110 7840
rect 18506 7828 18512 7840
rect 18564 7828 18570 7880
rect 18690 7828 18696 7880
rect 18748 7868 18754 7880
rect 19886 7868 19892 7880
rect 18748 7840 19892 7868
rect 18748 7828 18754 7840
rect 19886 7828 19892 7840
rect 19944 7868 19950 7880
rect 20548 7868 20576 7899
rect 21266 7868 21272 7880
rect 19944 7840 20576 7868
rect 21227 7840 21272 7868
rect 19944 7828 19950 7840
rect 21266 7828 21272 7840
rect 21324 7828 21330 7880
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 11710 7803 11768 7809
rect 11710 7800 11722 7803
rect 9640 7772 11722 7800
rect 9640 7760 9646 7772
rect 11710 7769 11722 7772
rect 11756 7769 11768 7803
rect 11710 7763 11768 7769
rect 13357 7803 13415 7809
rect 13357 7769 13369 7803
rect 13403 7800 13415 7803
rect 15286 7800 15292 7812
rect 13403 7772 15292 7800
rect 13403 7769 13415 7772
rect 13357 7763 13415 7769
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 15654 7760 15660 7812
rect 15712 7800 15718 7812
rect 17712 7803 17770 7809
rect 15712 7772 17632 7800
rect 15712 7760 15718 7772
rect 10686 7732 10692 7744
rect 9416 7704 10692 7732
rect 10686 7692 10692 7704
rect 10744 7692 10750 7744
rect 12158 7692 12164 7744
rect 12216 7732 12222 7744
rect 13722 7732 13728 7744
rect 12216 7704 13728 7732
rect 12216 7692 12222 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 14274 7732 14280 7744
rect 14235 7704 14280 7732
rect 14274 7692 14280 7704
rect 14332 7692 14338 7744
rect 14642 7732 14648 7744
rect 14603 7704 14648 7732
rect 14642 7692 14648 7704
rect 14700 7692 14706 7744
rect 15470 7732 15476 7744
rect 15431 7704 15476 7732
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16206 7732 16212 7744
rect 16167 7704 16212 7732
rect 16206 7692 16212 7704
rect 16264 7692 16270 7744
rect 17604 7732 17632 7772
rect 17712 7769 17724 7803
rect 17758 7800 17770 7803
rect 18064 7800 18092 7828
rect 18782 7800 18788 7812
rect 17758 7772 18092 7800
rect 18136 7772 18788 7800
rect 17758 7769 17770 7772
rect 17712 7763 17770 7769
rect 18136 7732 18164 7772
rect 18782 7760 18788 7772
rect 18840 7760 18846 7812
rect 19610 7800 19616 7812
rect 19523 7772 19616 7800
rect 19610 7760 19616 7772
rect 19668 7800 19674 7812
rect 20070 7800 20076 7812
rect 19668 7772 20076 7800
rect 19668 7760 19674 7772
rect 20070 7760 20076 7772
rect 20128 7760 20134 7812
rect 20349 7803 20407 7809
rect 20349 7769 20361 7803
rect 20395 7800 20407 7803
rect 20438 7800 20444 7812
rect 20395 7772 20444 7800
rect 20395 7769 20407 7772
rect 20349 7763 20407 7769
rect 20438 7760 20444 7772
rect 20496 7760 20502 7812
rect 21082 7800 21088 7812
rect 21043 7772 21088 7800
rect 21082 7760 21088 7772
rect 21140 7760 21146 7812
rect 17604 7704 18164 7732
rect 18325 7735 18383 7741
rect 18325 7701 18337 7735
rect 18371 7732 18383 7735
rect 18690 7732 18696 7744
rect 18371 7704 18696 7732
rect 18371 7701 18383 7704
rect 18325 7695 18383 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 19521 7735 19579 7741
rect 19521 7701 19533 7735
rect 19567 7732 19579 7735
rect 20714 7732 20720 7744
rect 19567 7704 20720 7732
rect 19567 7701 19579 7704
rect 19521 7695 19579 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1578 7528 1584 7540
rect 1539 7500 1584 7528
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2498 7528 2504 7540
rect 2363 7500 2504 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 3329 7531 3387 7537
rect 3329 7497 3341 7531
rect 3375 7528 3387 7531
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3375 7500 3985 7528
rect 3375 7497 3387 7500
rect 3329 7491 3387 7497
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 4338 7528 4344 7540
rect 4299 7500 4344 7528
rect 3973 7491 4031 7497
rect 4338 7488 4344 7500
rect 4396 7528 4402 7540
rect 5442 7528 5448 7540
rect 4396 7500 5448 7528
rect 4396 7488 4402 7500
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5994 7528 6000 7540
rect 5955 7500 6000 7528
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 10870 7528 10876 7540
rect 6104 7500 10876 7528
rect 3050 7460 3056 7472
rect 1504 7432 3056 7460
rect 1504 7404 1532 7432
rect 3050 7420 3056 7432
rect 3108 7420 3114 7472
rect 3234 7420 3240 7472
rect 3292 7460 3298 7472
rect 5629 7463 5687 7469
rect 5629 7460 5641 7463
rect 3292 7432 5641 7460
rect 3292 7420 3298 7432
rect 5629 7429 5641 7432
rect 5675 7429 5687 7463
rect 5629 7423 5687 7429
rect 1486 7392 1492 7404
rect 1447 7364 1492 7392
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 3418 7392 3424 7404
rect 3379 7364 3424 7392
rect 3418 7352 3424 7364
rect 3476 7352 3482 7404
rect 6104 7392 6132 7500
rect 10870 7488 10876 7500
rect 10928 7488 10934 7540
rect 15381 7531 15439 7537
rect 15381 7497 15393 7531
rect 15427 7528 15439 7531
rect 15930 7528 15936 7540
rect 15427 7500 15936 7528
rect 15427 7497 15439 7500
rect 15381 7491 15439 7497
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 16301 7531 16359 7537
rect 16301 7497 16313 7531
rect 16347 7528 16359 7531
rect 18049 7531 18107 7537
rect 16347 7500 18000 7528
rect 16347 7497 16359 7500
rect 16301 7491 16359 7497
rect 7374 7460 7380 7472
rect 7287 7432 7380 7460
rect 7374 7420 7380 7432
rect 7432 7460 7438 7472
rect 12250 7460 12256 7472
rect 7432 7432 12256 7460
rect 7432 7420 7438 7432
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 12342 7420 12348 7472
rect 12400 7460 12406 7472
rect 12434 7460 12440 7472
rect 12400 7432 12440 7460
rect 12400 7420 12406 7432
rect 12434 7420 12440 7432
rect 12492 7460 12498 7472
rect 13173 7463 13231 7469
rect 13173 7460 13185 7463
rect 12492 7432 13185 7460
rect 12492 7420 12498 7432
rect 7926 7392 7932 7404
rect 3620 7364 6132 7392
rect 7887 7364 7932 7392
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7293 2099 7327
rect 2222 7324 2228 7336
rect 2183 7296 2228 7324
rect 2041 7287 2099 7293
rect 2056 7256 2084 7287
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 3620 7333 3648 7364
rect 7926 7352 7932 7364
rect 7984 7352 7990 7404
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8352 7364 8493 7392
rect 8352 7352 8358 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8481 7355 8539 7361
rect 9214 7352 9220 7404
rect 9272 7392 9278 7404
rect 10514 7395 10572 7401
rect 10514 7392 10526 7395
rect 9272 7364 10526 7392
rect 9272 7352 9278 7364
rect 10514 7361 10526 7364
rect 10560 7361 10572 7395
rect 10514 7355 10572 7361
rect 12618 7352 12624 7404
rect 12676 7401 12682 7404
rect 12912 7401 12940 7432
rect 13173 7429 13185 7432
rect 13219 7460 13231 7463
rect 15948 7460 15976 7488
rect 16942 7469 16948 7472
rect 16936 7460 16948 7469
rect 13219 7432 13676 7460
rect 15948 7432 16712 7460
rect 16903 7432 16948 7460
rect 13219 7429 13231 7432
rect 13173 7423 13231 7429
rect 13648 7404 13676 7432
rect 12676 7392 12688 7401
rect 12897 7395 12955 7401
rect 12676 7364 12721 7392
rect 12676 7355 12688 7364
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 13630 7392 13636 7404
rect 13543 7364 13636 7392
rect 12897 7355 12955 7361
rect 12676 7352 12682 7355
rect 13630 7352 13636 7364
rect 13688 7352 13694 7404
rect 13900 7395 13958 7401
rect 13900 7392 13912 7395
rect 13740 7364 13912 7392
rect 3605 7327 3663 7333
rect 3605 7324 3617 7327
rect 2746 7296 3617 7324
rect 2746 7256 2774 7296
rect 3605 7293 3617 7296
rect 3651 7293 3663 7327
rect 3605 7287 3663 7293
rect 4062 7284 4068 7336
rect 4120 7324 4126 7336
rect 4433 7327 4491 7333
rect 4433 7324 4445 7327
rect 4120 7296 4445 7324
rect 4120 7284 4126 7296
rect 4433 7293 4445 7296
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5353 7327 5411 7333
rect 4672 7296 5304 7324
rect 4672 7284 4678 7296
rect 2056 7228 2774 7256
rect 2682 7188 2688 7200
rect 2643 7160 2688 7188
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 2958 7188 2964 7200
rect 2919 7160 2964 7188
rect 2958 7148 2964 7160
rect 3016 7148 3022 7200
rect 3234 7148 3240 7200
rect 3292 7188 3298 7200
rect 3970 7188 3976 7200
rect 3292 7160 3976 7188
rect 3292 7148 3298 7160
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 5276 7188 5304 7296
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5353 7287 5411 7293
rect 5368 7256 5396 7287
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 9766 7324 9772 7336
rect 5644 7296 9772 7324
rect 5644 7268 5672 7296
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 13740 7324 13768 7364
rect 13900 7361 13912 7364
rect 13946 7392 13958 7395
rect 15194 7392 15200 7404
rect 13946 7364 15200 7392
rect 13946 7361 13958 7364
rect 13900 7355 13958 7361
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 16117 7395 16175 7401
rect 16117 7361 16129 7395
rect 16163 7392 16175 7395
rect 16206 7392 16212 7404
rect 16163 7364 16212 7392
rect 16163 7361 16175 7364
rect 16117 7355 16175 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16684 7401 16712 7432
rect 16936 7423 16948 7432
rect 17000 7460 17006 7472
rect 17126 7460 17132 7472
rect 17000 7432 17132 7460
rect 16942 7420 16948 7423
rect 17000 7420 17006 7432
rect 17126 7420 17132 7432
rect 17184 7420 17190 7472
rect 17972 7460 18000 7500
rect 18049 7497 18061 7531
rect 18095 7528 18107 7531
rect 18138 7528 18144 7540
rect 18095 7500 18144 7528
rect 18095 7497 18107 7500
rect 18049 7491 18107 7497
rect 18138 7488 18144 7500
rect 18196 7528 18202 7540
rect 18874 7528 18880 7540
rect 18196 7500 18880 7528
rect 18196 7488 18202 7500
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19116 7500 19257 7528
rect 19116 7488 19122 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 19613 7531 19671 7537
rect 19613 7497 19625 7531
rect 19659 7528 19671 7531
rect 21358 7528 21364 7540
rect 19659 7500 21364 7528
rect 19659 7497 19671 7500
rect 19613 7491 19671 7497
rect 21358 7488 21364 7500
rect 21416 7488 21422 7540
rect 19150 7460 19156 7472
rect 17972 7432 19012 7460
rect 19111 7432 19156 7460
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 17494 7352 17500 7404
rect 17552 7392 17558 7404
rect 18690 7392 18696 7404
rect 17552 7364 18696 7392
rect 17552 7352 17558 7364
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 18984 7392 19012 7432
rect 19150 7420 19156 7432
rect 19208 7420 19214 7472
rect 19794 7420 19800 7472
rect 19852 7460 19858 7472
rect 19889 7463 19947 7469
rect 19889 7460 19901 7463
rect 19852 7432 19901 7460
rect 19852 7420 19858 7432
rect 19889 7429 19901 7432
rect 19935 7429 19947 7463
rect 20070 7460 20076 7472
rect 20031 7432 20076 7460
rect 19889 7423 19947 7429
rect 20070 7420 20076 7432
rect 20128 7420 20134 7472
rect 18984 7364 19196 7392
rect 10827 7296 11100 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 5626 7256 5632 7268
rect 5368 7228 5632 7256
rect 5626 7216 5632 7228
rect 5684 7216 5690 7268
rect 7834 7256 7840 7268
rect 5736 7228 7840 7256
rect 5736 7188 5764 7228
rect 7834 7216 7840 7228
rect 7892 7216 7898 7268
rect 8294 7216 8300 7268
rect 8352 7256 8358 7268
rect 8849 7259 8907 7265
rect 8849 7256 8861 7259
rect 8352 7228 8861 7256
rect 8352 7216 8358 7228
rect 8849 7225 8861 7228
rect 8895 7225 8907 7259
rect 8849 7219 8907 7225
rect 11072 7200 11100 7296
rect 13648 7296 13768 7324
rect 5276 7160 5764 7188
rect 5994 7148 6000 7200
rect 6052 7188 6058 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 6052 7160 6377 7188
rect 6052 7148 6058 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 7009 7191 7067 7197
rect 7009 7157 7021 7191
rect 7055 7188 7067 7191
rect 7190 7188 7196 7200
rect 7055 7160 7196 7188
rect 7055 7157 7067 7160
rect 7009 7151 7067 7157
rect 7190 7148 7196 7160
rect 7248 7148 7254 7200
rect 7926 7148 7932 7200
rect 7984 7188 7990 7200
rect 8113 7191 8171 7197
rect 8113 7188 8125 7191
rect 7984 7160 8125 7188
rect 7984 7148 7990 7160
rect 8113 7157 8125 7160
rect 8159 7157 8171 7191
rect 8113 7151 8171 7157
rect 8754 7148 8760 7200
rect 8812 7188 8818 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 8812 7160 9413 7188
rect 8812 7148 8818 7160
rect 9401 7157 9413 7160
rect 9447 7188 9459 7191
rect 10042 7188 10048 7200
rect 9447 7160 10048 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 10042 7148 10048 7160
rect 10100 7148 10106 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11517 7191 11575 7197
rect 11517 7157 11529 7191
rect 11563 7188 11575 7191
rect 12158 7188 12164 7200
rect 11563 7160 12164 7188
rect 11563 7157 11575 7160
rect 11517 7151 11575 7157
rect 12158 7148 12164 7160
rect 12216 7148 12222 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 13648 7188 13676 7296
rect 15212 7256 15240 7352
rect 15562 7284 15568 7336
rect 15620 7324 15626 7336
rect 18322 7324 18328 7336
rect 15620 7296 16068 7324
rect 18283 7296 18328 7324
rect 15620 7284 15626 7296
rect 15212 7228 15792 7256
rect 15010 7188 15016 7200
rect 12308 7160 13676 7188
rect 14971 7160 15016 7188
rect 12308 7148 12314 7160
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 15764 7197 15792 7228
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7188 15807 7191
rect 15930 7188 15936 7200
rect 15795 7160 15936 7188
rect 15795 7157 15807 7160
rect 15749 7151 15807 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16040 7188 16068 7296
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 18874 7284 18880 7336
rect 18932 7324 18938 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18932 7296 18981 7324
rect 18932 7284 18938 7296
rect 18969 7293 18981 7296
rect 19015 7293 19027 7327
rect 19168 7324 19196 7364
rect 19242 7352 19248 7404
rect 19300 7392 19306 7404
rect 20530 7392 20536 7404
rect 19300 7364 20536 7392
rect 19300 7352 19306 7364
rect 20530 7352 20536 7364
rect 20588 7352 20594 7404
rect 21450 7392 21456 7404
rect 20640 7364 21456 7392
rect 20640 7324 20668 7364
rect 21450 7352 21456 7364
rect 21508 7352 21514 7404
rect 19168 7296 20668 7324
rect 20809 7327 20867 7333
rect 18969 7287 19027 7293
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 20824 7256 20852 7287
rect 19306 7228 20852 7256
rect 19306 7188 19334 7228
rect 16040 7160 19334 7188
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2130 6984 2136 6996
rect 2091 6956 2136 6984
rect 2130 6944 2136 6956
rect 2188 6944 2194 6996
rect 2222 6944 2228 6996
rect 2280 6984 2286 6996
rect 2409 6987 2467 6993
rect 2409 6984 2421 6987
rect 2280 6956 2421 6984
rect 2280 6944 2286 6956
rect 2409 6953 2421 6956
rect 2455 6953 2467 6987
rect 2409 6947 2467 6953
rect 2498 6944 2504 6996
rect 2556 6984 2562 6996
rect 4890 6984 4896 6996
rect 2556 6956 4896 6984
rect 2556 6944 2562 6956
rect 4890 6944 4896 6956
rect 4948 6944 4954 6996
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 6914 6984 6920 6996
rect 5224 6956 6920 6984
rect 5224 6944 5230 6956
rect 6914 6944 6920 6956
rect 6972 6944 6978 6996
rect 7006 6944 7012 6996
rect 7064 6984 7070 6996
rect 7469 6987 7527 6993
rect 7469 6984 7481 6987
rect 7064 6956 7481 6984
rect 7064 6944 7070 6956
rect 7469 6953 7481 6956
rect 7515 6953 7527 6987
rect 7469 6947 7527 6953
rect 8018 6944 8024 6996
rect 8076 6984 8082 6996
rect 8478 6984 8484 6996
rect 8076 6956 8484 6984
rect 8076 6944 8082 6956
rect 8478 6944 8484 6956
rect 8536 6944 8542 6996
rect 9214 6984 9220 6996
rect 9175 6956 9220 6984
rect 9214 6944 9220 6956
rect 9272 6944 9278 6996
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10594 6984 10600 6996
rect 9916 6956 10600 6984
rect 9916 6944 9922 6956
rect 10594 6944 10600 6956
rect 10652 6984 10658 6996
rect 12250 6984 12256 6996
rect 10652 6956 12256 6984
rect 10652 6944 10658 6956
rect 12250 6944 12256 6956
rect 12308 6944 12314 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12802 6984 12808 6996
rect 12400 6956 12808 6984
rect 12400 6944 12406 6956
rect 12802 6944 12808 6956
rect 12860 6944 12866 6996
rect 18877 6987 18935 6993
rect 18340 6956 18552 6984
rect 2774 6876 2780 6928
rect 2832 6876 2838 6928
rect 4614 6876 4620 6928
rect 4672 6876 4678 6928
rect 7374 6916 7380 6928
rect 6656 6888 7380 6916
rect 2792 6848 2820 6876
rect 1964 6820 2820 6848
rect 3053 6851 3111 6857
rect 1486 6780 1492 6792
rect 1447 6752 1492 6780
rect 1486 6740 1492 6752
rect 1544 6740 1550 6792
rect 1964 6789 1992 6820
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 4632 6848 4660 6876
rect 3099 6820 4660 6848
rect 4801 6851 4859 6857
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 4801 6817 4813 6851
rect 4847 6848 4859 6851
rect 5810 6848 5816 6860
rect 4847 6820 5816 6848
rect 4847 6817 4859 6820
rect 4801 6811 4859 6817
rect 5810 6808 5816 6820
rect 5868 6808 5874 6860
rect 6656 6857 6684 6888
rect 7374 6876 7380 6888
rect 7432 6876 7438 6928
rect 12069 6919 12127 6925
rect 12069 6885 12081 6919
rect 12115 6885 12127 6919
rect 12069 6879 12127 6885
rect 6641 6851 6699 6857
rect 6641 6817 6653 6851
rect 6687 6817 6699 6851
rect 6641 6811 6699 6817
rect 7466 6808 7472 6860
rect 7524 6808 7530 6860
rect 8113 6851 8171 6857
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8202 6848 8208 6860
rect 8159 6820 8208 6848
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8202 6808 8208 6820
rect 8260 6808 8266 6860
rect 12084 6848 12112 6879
rect 10520 6820 12112 6848
rect 13449 6851 13507 6857
rect 1949 6783 2007 6789
rect 1949 6749 1961 6783
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 2774 6740 2780 6792
rect 2832 6780 2838 6792
rect 3326 6780 3332 6792
rect 2832 6752 3332 6780
rect 2832 6740 2838 6752
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5350 6780 5356 6792
rect 4663 6752 5356 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 5350 6740 5356 6752
rect 5408 6740 5414 6792
rect 5629 6783 5687 6789
rect 5629 6749 5641 6783
rect 5675 6780 5687 6783
rect 5994 6780 6000 6792
rect 5675 6752 6000 6780
rect 5675 6749 5687 6752
rect 5629 6743 5687 6749
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 7484 6780 7512 6808
rect 6196 6752 7512 6780
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1719 6684 5672 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3234 6644 3240 6656
rect 2915 6616 3240 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3234 6604 3240 6616
rect 3292 6644 3298 6656
rect 3418 6644 3424 6656
rect 3292 6616 3424 6644
rect 3292 6604 3298 6616
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3881 6647 3939 6653
rect 3881 6613 3893 6647
rect 3927 6644 3939 6647
rect 3970 6644 3976 6656
rect 3927 6616 3976 6644
rect 3927 6613 3939 6616
rect 3881 6607 3939 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4525 6647 4583 6653
rect 4525 6613 4537 6647
rect 4571 6644 4583 6647
rect 4614 6644 4620 6656
rect 4571 6616 4620 6644
rect 4571 6613 4583 6616
rect 4525 6607 4583 6613
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5166 6644 5172 6656
rect 5127 6616 5172 6644
rect 5166 6604 5172 6616
rect 5224 6604 5230 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5537 6647 5595 6653
rect 5537 6644 5549 6647
rect 5316 6616 5549 6644
rect 5316 6604 5322 6616
rect 5537 6613 5549 6616
rect 5583 6613 5595 6647
rect 5644 6644 5672 6684
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 6196 6712 6224 6752
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 7892 6752 9674 6780
rect 7892 6740 7898 6752
rect 5776 6684 6224 6712
rect 6733 6715 6791 6721
rect 5776 6672 5782 6684
rect 6733 6681 6745 6715
rect 6779 6712 6791 6715
rect 7466 6712 7472 6724
rect 6779 6684 7472 6712
rect 6779 6681 6791 6684
rect 6733 6675 6791 6681
rect 7466 6672 7472 6684
rect 7524 6672 7530 6724
rect 7742 6672 7748 6724
rect 7800 6712 7806 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 7800 6684 7941 6712
rect 7800 6672 7806 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 9646 6712 9674 6752
rect 9766 6740 9772 6792
rect 9824 6780 9830 6792
rect 10330 6783 10388 6789
rect 10330 6780 10342 6783
rect 9824 6752 10342 6780
rect 9824 6740 9830 6752
rect 10330 6749 10342 6752
rect 10376 6780 10388 6783
rect 10520 6780 10548 6820
rect 13449 6817 13461 6851
rect 13495 6848 13507 6851
rect 13630 6848 13636 6860
rect 13495 6820 13636 6848
rect 13495 6817 13507 6820
rect 13449 6811 13507 6817
rect 13630 6808 13636 6820
rect 13688 6848 13694 6860
rect 14093 6851 14151 6857
rect 14093 6848 14105 6851
rect 13688 6820 14105 6848
rect 13688 6808 13694 6820
rect 14093 6817 14105 6820
rect 14139 6848 14151 6851
rect 14553 6851 14611 6857
rect 14553 6848 14565 6851
rect 14139 6820 14565 6848
rect 14139 6817 14151 6820
rect 14093 6811 14151 6817
rect 14553 6817 14565 6820
rect 14599 6817 14611 6851
rect 14553 6811 14611 6817
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6848 17647 6851
rect 18046 6848 18052 6860
rect 17635 6820 18052 6848
rect 17635 6817 17647 6820
rect 17589 6811 17647 6817
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 18233 6851 18291 6857
rect 18233 6817 18245 6851
rect 18279 6848 18291 6851
rect 18340 6848 18368 6956
rect 18524 6916 18552 6956
rect 18877 6953 18889 6987
rect 18923 6984 18935 6987
rect 20346 6984 20352 6996
rect 18923 6956 20352 6984
rect 18923 6953 18935 6956
rect 18877 6947 18935 6953
rect 20346 6944 20352 6956
rect 20404 6944 20410 6996
rect 18524 6888 19334 6916
rect 18279 6820 18368 6848
rect 19306 6848 19334 6888
rect 19426 6848 19432 6860
rect 19306 6820 19432 6848
rect 18279 6817 18291 6820
rect 18233 6811 18291 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 19610 6848 19616 6860
rect 19571 6820 19616 6848
rect 19610 6808 19616 6820
rect 19668 6808 19674 6860
rect 19797 6851 19855 6857
rect 19797 6817 19809 6851
rect 19843 6848 19855 6851
rect 20162 6848 20168 6860
rect 19843 6820 20168 6848
rect 19843 6817 19855 6820
rect 19797 6811 19855 6817
rect 20162 6808 20168 6820
rect 20220 6808 20226 6860
rect 20809 6851 20867 6857
rect 20809 6848 20821 6851
rect 20272 6820 20821 6848
rect 10376 6752 10548 6780
rect 10597 6783 10655 6789
rect 10376 6749 10388 6752
rect 10330 6743 10388 6749
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 11054 6780 11060 6792
rect 10643 6752 11060 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11054 6740 11060 6752
rect 11112 6740 11118 6792
rect 13182 6783 13240 6789
rect 13182 6780 13194 6783
rect 12268 6752 13194 6780
rect 10134 6712 10140 6724
rect 9646 6684 10140 6712
rect 7929 6675 7987 6681
rect 10134 6672 10140 6684
rect 10192 6672 10198 6724
rect 10244 6684 11376 6712
rect 6178 6644 6184 6656
rect 5644 6616 6184 6644
rect 5537 6607 5595 6613
rect 6178 6604 6184 6616
rect 6236 6604 6242 6656
rect 6825 6647 6883 6653
rect 6825 6613 6837 6647
rect 6871 6644 6883 6647
rect 7006 6644 7012 6656
rect 6871 6616 7012 6644
rect 6871 6613 6883 6616
rect 6825 6607 6883 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 7156 6616 7205 6644
rect 7156 6604 7162 6616
rect 7193 6613 7205 6616
rect 7239 6613 7251 6647
rect 7834 6644 7840 6656
rect 7795 6616 7840 6644
rect 7193 6607 7251 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10244 6644 10272 6684
rect 9824 6616 10272 6644
rect 10965 6647 11023 6653
rect 9824 6604 9830 6616
rect 10965 6613 10977 6647
rect 11011 6644 11023 6647
rect 11054 6644 11060 6656
rect 11011 6616 11060 6644
rect 11011 6613 11023 6616
rect 10965 6607 11023 6613
rect 11054 6604 11060 6616
rect 11112 6644 11118 6656
rect 11241 6647 11299 6653
rect 11241 6644 11253 6647
rect 11112 6616 11253 6644
rect 11112 6604 11118 6616
rect 11241 6613 11253 6616
rect 11287 6613 11299 6647
rect 11348 6644 11376 6684
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 11848 6684 11893 6712
rect 11848 6672 11854 6684
rect 12268 6644 12296 6752
rect 13182 6749 13194 6752
rect 13228 6749 13240 6783
rect 13182 6743 13240 6749
rect 13814 6740 13820 6792
rect 13872 6780 13878 6792
rect 14826 6789 14832 6792
rect 14820 6780 14832 6789
rect 13872 6752 14832 6780
rect 13872 6740 13878 6752
rect 14820 6743 14832 6752
rect 14826 6740 14832 6743
rect 14884 6740 14890 6792
rect 15286 6740 15292 6792
rect 15344 6780 15350 6792
rect 16669 6783 16727 6789
rect 16669 6780 16681 6783
rect 15344 6752 16681 6780
rect 15344 6740 15350 6752
rect 16669 6749 16681 6752
rect 16715 6780 16727 6783
rect 17313 6783 17371 6789
rect 16715 6752 17264 6780
rect 16715 6749 16727 6752
rect 16669 6743 16727 6749
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 15252 6684 16528 6712
rect 15252 6672 15258 6684
rect 11348 6616 12296 6644
rect 15933 6647 15991 6653
rect 11241 6607 11299 6613
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 16022 6644 16028 6656
rect 15979 6616 16028 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 16022 6604 16028 6616
rect 16080 6604 16086 6656
rect 16500 6653 16528 6684
rect 16485 6647 16543 6653
rect 16485 6613 16497 6647
rect 16531 6613 16543 6647
rect 16942 6644 16948 6656
rect 16903 6616 16948 6644
rect 16485 6607 16543 6613
rect 16942 6604 16948 6616
rect 17000 6604 17006 6656
rect 17236 6644 17264 6752
rect 17313 6749 17325 6783
rect 17359 6780 17371 6783
rect 18322 6780 18328 6792
rect 17359 6752 18328 6780
rect 17359 6749 17371 6752
rect 17313 6743 17371 6749
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 18782 6740 18788 6792
rect 18840 6780 18846 6792
rect 20272 6780 20300 6820
rect 20809 6817 20821 6820
rect 20855 6817 20867 6851
rect 20809 6811 20867 6817
rect 18840 6752 20300 6780
rect 20533 6783 20591 6789
rect 18840 6740 18846 6752
rect 20533 6749 20545 6783
rect 20579 6749 20591 6783
rect 20533 6743 20591 6749
rect 17405 6715 17463 6721
rect 17405 6681 17417 6715
rect 17451 6712 17463 6715
rect 17954 6712 17960 6724
rect 17451 6684 17960 6712
rect 17451 6681 17463 6684
rect 17405 6675 17463 6681
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 18598 6712 18604 6724
rect 18064 6684 18604 6712
rect 18064 6644 18092 6684
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 19610 6672 19616 6724
rect 19668 6712 19674 6724
rect 19889 6715 19947 6721
rect 19889 6712 19901 6715
rect 19668 6684 19901 6712
rect 19668 6672 19674 6684
rect 19889 6681 19901 6684
rect 19935 6681 19947 6715
rect 20548 6712 20576 6743
rect 19889 6675 19947 6681
rect 20088 6684 20576 6712
rect 18414 6644 18420 6656
rect 17236 6616 18092 6644
rect 18375 6616 18420 6644
rect 18414 6604 18420 6616
rect 18472 6604 18478 6656
rect 18509 6647 18567 6653
rect 18509 6613 18521 6647
rect 18555 6644 18567 6647
rect 18782 6644 18788 6656
rect 18555 6616 18788 6644
rect 18555 6613 18567 6616
rect 18509 6607 18567 6613
rect 18782 6604 18788 6616
rect 18840 6604 18846 6656
rect 19242 6604 19248 6656
rect 19300 6644 19306 6656
rect 20088 6644 20116 6684
rect 20254 6644 20260 6656
rect 19300 6616 20116 6644
rect 20215 6616 20260 6644
rect 19300 6604 19306 6616
rect 20254 6604 20260 6616
rect 20312 6604 20318 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 2590 6440 2596 6452
rect 2551 6412 2596 6440
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 3053 6443 3111 6449
rect 3053 6440 3065 6443
rect 3016 6412 3065 6440
rect 3016 6400 3022 6412
rect 3053 6409 3065 6412
rect 3099 6409 3111 6443
rect 3053 6403 3111 6409
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 4341 6443 4399 6449
rect 3384 6412 4292 6440
rect 3384 6400 3390 6412
rect 1857 6375 1915 6381
rect 1857 6341 1869 6375
rect 1903 6372 1915 6375
rect 2774 6372 2780 6384
rect 1903 6344 2780 6372
rect 1903 6341 1915 6344
rect 1857 6335 1915 6341
rect 2774 6332 2780 6344
rect 2832 6332 2838 6384
rect 4264 6372 4292 6412
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 5258 6440 5264 6452
rect 4387 6412 5264 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 5258 6400 5264 6412
rect 5316 6400 5322 6452
rect 12618 6440 12624 6452
rect 5552 6412 12624 6440
rect 3068 6344 4200 6372
rect 4264 6344 4660 6372
rect 3068 6316 3096 6344
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1762 6236 1768 6248
rect 1723 6208 1768 6236
rect 1762 6196 1768 6208
rect 1820 6196 1826 6248
rect 1964 6236 1992 6267
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 2961 6307 3019 6313
rect 2961 6304 2973 6307
rect 2740 6276 2973 6304
rect 2740 6264 2746 6276
rect 2961 6273 2973 6276
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 4172 6313 4200 6344
rect 4632 6313 4660 6344
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3476 6276 3709 6304
rect 3476 6264 3482 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6273 4675 6307
rect 4617 6267 4675 6273
rect 3237 6239 3295 6245
rect 1964 6208 3188 6236
rect 2317 6171 2375 6177
rect 2317 6137 2329 6171
rect 2363 6168 2375 6171
rect 2866 6168 2872 6180
rect 2363 6140 2872 6168
rect 2363 6137 2375 6140
rect 2317 6131 2375 6137
rect 2866 6128 2872 6140
rect 2924 6128 2930 6180
rect 3160 6168 3188 6208
rect 3237 6205 3249 6239
rect 3283 6236 3295 6239
rect 5552 6236 5580 6412
rect 12618 6400 12624 6412
rect 12676 6440 12682 6452
rect 13449 6443 13507 6449
rect 13449 6440 13461 6443
rect 12676 6412 13461 6440
rect 12676 6400 12682 6412
rect 13449 6409 13461 6412
rect 13495 6409 13507 6443
rect 13449 6403 13507 6409
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 13725 6443 13783 6449
rect 13725 6440 13737 6443
rect 13688 6412 13737 6440
rect 13688 6400 13694 6412
rect 13725 6409 13737 6412
rect 13771 6409 13783 6443
rect 13725 6403 13783 6409
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 14884 6412 15117 6440
rect 14884 6400 14890 6412
rect 15105 6409 15117 6412
rect 15151 6409 15163 6443
rect 15105 6403 15163 6409
rect 15286 6400 15292 6452
rect 15344 6440 15350 6452
rect 15470 6440 15476 6452
rect 15344 6412 15476 6440
rect 15344 6400 15350 6412
rect 15470 6400 15476 6412
rect 15528 6400 15534 6452
rect 16298 6440 16304 6452
rect 16259 6412 16304 6440
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 16850 6400 16856 6452
rect 16908 6440 16914 6452
rect 16945 6443 17003 6449
rect 16945 6440 16957 6443
rect 16908 6412 16957 6440
rect 16908 6400 16914 6412
rect 16945 6409 16957 6412
rect 16991 6409 17003 6443
rect 16945 6403 17003 6409
rect 17405 6443 17463 6449
rect 17405 6409 17417 6443
rect 17451 6440 17463 6443
rect 18138 6440 18144 6452
rect 17451 6412 18144 6440
rect 17451 6409 17463 6412
rect 17405 6403 17463 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18414 6400 18420 6452
rect 18472 6440 18478 6452
rect 20625 6443 20683 6449
rect 20625 6440 20637 6443
rect 18472 6412 20637 6440
rect 18472 6400 18478 6412
rect 20625 6409 20637 6412
rect 20671 6409 20683 6443
rect 20625 6403 20683 6409
rect 20806 6400 20812 6452
rect 20864 6440 20870 6452
rect 21085 6443 21143 6449
rect 21085 6440 21097 6443
rect 20864 6412 21097 6440
rect 20864 6400 20870 6412
rect 21085 6409 21097 6412
rect 21131 6440 21143 6443
rect 21542 6440 21548 6452
rect 21131 6412 21548 6440
rect 21131 6409 21143 6412
rect 21085 6403 21143 6409
rect 21542 6400 21548 6412
rect 21600 6400 21606 6452
rect 5629 6375 5687 6381
rect 5629 6341 5641 6375
rect 5675 6372 5687 6375
rect 7006 6372 7012 6384
rect 5675 6344 7012 6372
rect 5675 6341 5687 6344
rect 5629 6335 5687 6341
rect 7006 6332 7012 6344
rect 7064 6372 7070 6384
rect 7282 6372 7288 6384
rect 7064 6344 7288 6372
rect 7064 6332 7070 6344
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 8570 6372 8576 6384
rect 7944 6344 8432 6372
rect 8531 6344 8576 6372
rect 5718 6304 5724 6316
rect 5679 6276 5724 6304
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6304 6607 6307
rect 6822 6304 6828 6316
rect 6595 6276 6828 6304
rect 6595 6273 6607 6276
rect 6549 6267 6607 6273
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7098 6264 7104 6316
rect 7156 6304 7162 6316
rect 7561 6307 7619 6313
rect 7561 6304 7573 6307
rect 7156 6276 7573 6304
rect 7156 6264 7162 6276
rect 7561 6273 7573 6276
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 5810 6236 5816 6248
rect 3283 6208 5580 6236
rect 5771 6208 5816 6236
rect 3283 6205 3295 6208
rect 3237 6199 3295 6205
rect 5810 6196 5816 6208
rect 5868 6196 5874 6248
rect 7374 6236 7380 6248
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7524 6208 7569 6236
rect 7524 6196 7530 6208
rect 3881 6171 3939 6177
rect 3160 6140 3464 6168
rect 3436 6100 3464 6140
rect 3881 6137 3893 6171
rect 3927 6168 3939 6171
rect 4338 6168 4344 6180
rect 3927 6140 4344 6168
rect 3927 6137 3939 6140
rect 3881 6131 3939 6137
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4798 6168 4804 6180
rect 4759 6140 4804 6168
rect 4798 6128 4804 6140
rect 4856 6128 4862 6180
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 7944 6177 7972 6344
rect 8404 6304 8432 6344
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 8754 6332 8760 6384
rect 8812 6372 8818 6384
rect 11790 6372 11796 6384
rect 8812 6344 11796 6372
rect 8812 6332 8818 6344
rect 11790 6332 11796 6344
rect 11848 6332 11854 6384
rect 12802 6332 12808 6384
rect 12860 6372 12866 6384
rect 17037 6375 17095 6381
rect 17037 6372 17049 6375
rect 12860 6344 17049 6372
rect 12860 6332 12866 6344
rect 17037 6341 17049 6344
rect 17083 6341 17095 6375
rect 17037 6335 17095 6341
rect 18046 6332 18052 6384
rect 18104 6372 18110 6384
rect 18325 6375 18383 6381
rect 18325 6372 18337 6375
rect 18104 6344 18337 6372
rect 18104 6332 18110 6344
rect 18325 6341 18337 6344
rect 18371 6341 18383 6375
rect 18325 6335 18383 6341
rect 19334 6332 19340 6384
rect 19392 6372 19398 6384
rect 19518 6372 19524 6384
rect 19392 6344 19524 6372
rect 19392 6332 19398 6344
rect 19518 6332 19524 6344
rect 19576 6372 19582 6384
rect 20082 6375 20140 6381
rect 20082 6372 20094 6375
rect 19576 6344 20094 6372
rect 19576 6332 19582 6344
rect 20082 6341 20094 6344
rect 20128 6341 20140 6375
rect 20082 6335 20140 6341
rect 20714 6332 20720 6384
rect 20772 6332 20778 6384
rect 9858 6304 9864 6316
rect 8404 6276 9076 6304
rect 9819 6276 9864 6304
rect 8018 6196 8024 6248
rect 8076 6236 8082 6248
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8076 6208 8309 6236
rect 8076 6196 8082 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8478 6236 8484 6248
rect 8439 6208 8484 6236
rect 8297 6199 8355 6205
rect 6365 6171 6423 6177
rect 6365 6168 6377 6171
rect 5500 6140 6377 6168
rect 5500 6128 5506 6140
rect 6365 6137 6377 6140
rect 6411 6137 6423 6171
rect 6365 6131 6423 6137
rect 7929 6171 7987 6177
rect 7929 6137 7941 6171
rect 7975 6137 7987 6171
rect 7929 6131 7987 6137
rect 4522 6100 4528 6112
rect 3436 6072 4528 6100
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 4890 6060 4896 6112
rect 4948 6100 4954 6112
rect 5261 6103 5319 6109
rect 5261 6100 5273 6103
rect 4948 6072 5273 6100
rect 4948 6060 4954 6072
rect 5261 6069 5273 6072
rect 5307 6069 5319 6103
rect 5261 6063 5319 6069
rect 6917 6103 6975 6109
rect 6917 6069 6929 6103
rect 6963 6100 6975 6103
rect 8018 6100 8024 6112
rect 6963 6072 8024 6100
rect 6963 6069 6975 6072
rect 6917 6063 6975 6069
rect 8018 6060 8024 6072
rect 8076 6060 8082 6112
rect 8312 6100 8340 6199
rect 8478 6196 8484 6208
rect 8536 6196 8542 6248
rect 8754 6128 8760 6180
rect 8812 6168 8818 6180
rect 8941 6171 8999 6177
rect 8941 6168 8953 6171
rect 8812 6140 8953 6168
rect 8812 6128 8818 6140
rect 8941 6137 8953 6140
rect 8987 6137 8999 6171
rect 9048 6168 9076 6276
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 10870 6264 10876 6316
rect 10928 6304 10934 6316
rect 12336 6308 12394 6313
rect 12268 6307 12394 6308
rect 12268 6304 12348 6307
rect 10928 6280 12348 6304
rect 10928 6276 12296 6280
rect 10928 6264 10934 6276
rect 12336 6273 12348 6280
rect 12382 6273 12394 6307
rect 12336 6267 12394 6273
rect 14550 6264 14556 6316
rect 14608 6304 14614 6316
rect 14645 6307 14703 6313
rect 14645 6304 14657 6307
rect 14608 6276 14657 6304
rect 14608 6264 14614 6276
rect 14645 6273 14657 6276
rect 14691 6273 14703 6307
rect 15286 6304 15292 6316
rect 15247 6276 15292 6304
rect 14645 6267 14703 6273
rect 15286 6264 15292 6276
rect 15344 6264 15350 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6273 15991 6307
rect 17126 6304 17132 6316
rect 15933 6267 15991 6273
rect 16868 6276 17132 6304
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 10686 6236 10692 6248
rect 9272 6208 10692 6236
rect 9272 6196 9278 6208
rect 10686 6196 10692 6208
rect 10744 6196 10750 6248
rect 11514 6196 11520 6248
rect 11572 6236 11578 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11572 6208 12081 6236
rect 11572 6196 11578 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 15654 6236 15660 6248
rect 15615 6208 15660 6236
rect 12069 6199 12127 6205
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15838 6236 15844 6248
rect 15799 6208 15844 6236
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 15948 6168 15976 6267
rect 16868 6245 16896 6276
rect 17126 6264 17132 6276
rect 17184 6264 17190 6316
rect 20530 6304 20536 6316
rect 18156 6276 20536 6304
rect 18156 6245 18184 6276
rect 20530 6264 20536 6276
rect 20588 6304 20594 6316
rect 20732 6304 20760 6332
rect 20588 6276 20760 6304
rect 20993 6307 21051 6313
rect 20588 6264 20594 6276
rect 20993 6273 21005 6307
rect 21039 6304 21051 6307
rect 21358 6304 21364 6316
rect 21039 6276 21364 6304
rect 21039 6273 21051 6276
rect 20993 6267 21051 6273
rect 21358 6264 21364 6276
rect 21416 6264 21422 6316
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6205 16911 6239
rect 16853 6199 16911 6205
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6205 18199 6239
rect 18141 6199 18199 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6205 18291 6239
rect 18233 6199 18291 6205
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 20714 6236 20720 6248
rect 20395 6208 20720 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 9048 6140 11652 6168
rect 8941 6131 8999 6137
rect 9214 6100 9220 6112
rect 8312 6072 9220 6100
rect 9214 6060 9220 6072
rect 9272 6060 9278 6112
rect 10229 6103 10287 6109
rect 10229 6069 10241 6103
rect 10275 6100 10287 6103
rect 10318 6100 10324 6112
rect 10275 6072 10324 6100
rect 10275 6069 10287 6072
rect 10229 6063 10287 6069
rect 10318 6060 10324 6072
rect 10376 6060 10382 6112
rect 10502 6100 10508 6112
rect 10463 6072 10508 6100
rect 10502 6060 10508 6072
rect 10560 6060 10566 6112
rect 10965 6103 11023 6109
rect 10965 6069 10977 6103
rect 11011 6100 11023 6103
rect 11054 6100 11060 6112
rect 11011 6072 11060 6100
rect 11011 6069 11023 6072
rect 10965 6063 11023 6069
rect 11054 6060 11060 6072
rect 11112 6100 11118 6112
rect 11514 6100 11520 6112
rect 11112 6072 11520 6100
rect 11112 6060 11118 6072
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 11624 6100 11652 6140
rect 13372 6140 15976 6168
rect 13372 6100 13400 6140
rect 16390 6128 16396 6180
rect 16448 6168 16454 6180
rect 16448 6140 17908 6168
rect 16448 6128 16454 6140
rect 11624 6072 13400 6100
rect 14369 6103 14427 6109
rect 14369 6069 14381 6103
rect 14415 6100 14427 6103
rect 14550 6100 14556 6112
rect 14415 6072 14556 6100
rect 14415 6069 14427 6072
rect 14369 6063 14427 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14829 6103 14887 6109
rect 14829 6069 14841 6103
rect 14875 6100 14887 6103
rect 17494 6100 17500 6112
rect 14875 6072 17500 6100
rect 14875 6069 14887 6072
rect 14829 6063 14887 6069
rect 17494 6060 17500 6072
rect 17552 6060 17558 6112
rect 17880 6100 17908 6140
rect 17954 6128 17960 6180
rect 18012 6168 18018 6180
rect 18248 6168 18276 6199
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 21082 6196 21088 6248
rect 21140 6236 21146 6248
rect 21177 6239 21235 6245
rect 21177 6236 21189 6239
rect 21140 6208 21189 6236
rect 21140 6196 21146 6208
rect 21177 6205 21189 6208
rect 21223 6205 21235 6239
rect 21177 6199 21235 6205
rect 18012 6140 18276 6168
rect 18693 6171 18751 6177
rect 18012 6128 18018 6140
rect 18693 6137 18705 6171
rect 18739 6168 18751 6171
rect 18739 6140 19380 6168
rect 18739 6137 18751 6140
rect 18693 6131 18751 6137
rect 18414 6100 18420 6112
rect 17880 6072 18420 6100
rect 18414 6060 18420 6072
rect 18472 6060 18478 6112
rect 18506 6060 18512 6112
rect 18564 6100 18570 6112
rect 18969 6103 19027 6109
rect 18969 6100 18981 6103
rect 18564 6072 18981 6100
rect 18564 6060 18570 6072
rect 18969 6069 18981 6072
rect 19015 6069 19027 6103
rect 19352 6100 19380 6140
rect 19978 6100 19984 6112
rect 19352 6072 19984 6100
rect 18969 6063 19027 6069
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1578 5856 1584 5908
rect 1636 5896 1642 5908
rect 3326 5896 3332 5908
rect 1636 5868 3332 5896
rect 1636 5856 1642 5868
rect 3326 5856 3332 5868
rect 3384 5856 3390 5908
rect 3786 5896 3792 5908
rect 3747 5868 3792 5896
rect 3786 5856 3792 5868
rect 3844 5856 3850 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4706 5896 4712 5908
rect 4667 5868 4712 5896
rect 4706 5856 4712 5868
rect 4764 5856 4770 5908
rect 5534 5856 5540 5908
rect 5592 5896 5598 5908
rect 5813 5899 5871 5905
rect 5813 5896 5825 5899
rect 5592 5868 5825 5896
rect 5592 5856 5598 5868
rect 5813 5865 5825 5868
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 7374 5856 7380 5908
rect 7432 5896 7438 5908
rect 7432 5868 14596 5896
rect 7432 5856 7438 5868
rect 3234 5788 3240 5840
rect 3292 5828 3298 5840
rect 6825 5831 6883 5837
rect 6825 5828 6837 5831
rect 3292 5800 6837 5828
rect 3292 5788 3298 5800
rect 6825 5797 6837 5800
rect 6871 5797 6883 5831
rect 6825 5791 6883 5797
rect 7282 5788 7288 5840
rect 7340 5828 7346 5840
rect 7929 5831 7987 5837
rect 7929 5828 7941 5831
rect 7340 5800 7941 5828
rect 7340 5788 7346 5800
rect 7929 5797 7941 5800
rect 7975 5828 7987 5831
rect 8110 5828 8116 5840
rect 7975 5800 8116 5828
rect 7975 5797 7987 5800
rect 7929 5791 7987 5797
rect 8110 5788 8116 5800
rect 8168 5788 8174 5840
rect 9122 5788 9128 5840
rect 9180 5828 9186 5840
rect 9217 5831 9275 5837
rect 9217 5828 9229 5831
rect 9180 5800 9229 5828
rect 9180 5788 9186 5800
rect 9217 5797 9229 5800
rect 9263 5797 9275 5831
rect 9582 5828 9588 5840
rect 9543 5800 9588 5828
rect 9217 5791 9275 5797
rect 9582 5788 9588 5800
rect 9640 5788 9646 5840
rect 10962 5788 10968 5840
rect 11020 5828 11026 5840
rect 13078 5828 13084 5840
rect 11020 5800 13084 5828
rect 11020 5788 11026 5800
rect 13078 5788 13084 5800
rect 13136 5828 13142 5840
rect 13814 5828 13820 5840
rect 13136 5800 13820 5828
rect 13136 5788 13142 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 1857 5763 1915 5769
rect 1857 5729 1869 5763
rect 1903 5729 1915 5763
rect 1857 5723 1915 5729
rect 1949 5763 2007 5769
rect 1949 5729 1961 5763
rect 1995 5760 2007 5763
rect 2774 5760 2780 5772
rect 1995 5732 2780 5760
rect 1995 5729 2007 5732
rect 1949 5723 2007 5729
rect 1872 5692 1900 5723
rect 2774 5720 2780 5732
rect 2832 5720 2838 5772
rect 3326 5760 3332 5772
rect 3287 5732 3332 5760
rect 3326 5720 3332 5732
rect 3384 5720 3390 5772
rect 3510 5720 3516 5772
rect 3568 5760 3574 5772
rect 6457 5763 6515 5769
rect 3568 5732 4936 5760
rect 3568 5720 3574 5732
rect 2590 5692 2596 5704
rect 1872 5664 2596 5692
rect 2590 5652 2596 5664
rect 2648 5652 2654 5704
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3200 5664 3985 5692
rect 3200 5652 3206 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4430 5692 4436 5704
rect 4120 5664 4436 5692
rect 4120 5652 4126 5664
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4908 5701 4936 5732
rect 6457 5729 6469 5763
rect 6503 5760 6515 5763
rect 6914 5760 6920 5772
rect 6503 5732 6920 5760
rect 6503 5729 6515 5732
rect 6457 5723 6515 5729
rect 6914 5720 6920 5732
rect 6972 5760 6978 5772
rect 9766 5760 9772 5772
rect 6972 5732 8156 5760
rect 6972 5720 6978 5732
rect 4893 5695 4951 5701
rect 4893 5661 4905 5695
rect 4939 5692 4951 5695
rect 5074 5692 5080 5704
rect 4939 5664 5080 5692
rect 4939 5661 4951 5664
rect 4893 5655 4951 5661
rect 5074 5652 5080 5664
rect 5132 5652 5138 5704
rect 5718 5652 5724 5704
rect 5776 5692 5782 5704
rect 6730 5692 6736 5704
rect 5776 5664 6736 5692
rect 5776 5652 5782 5664
rect 6730 5652 6736 5664
rect 6788 5692 6794 5704
rect 7009 5695 7067 5701
rect 7009 5692 7021 5695
rect 6788 5664 7021 5692
rect 6788 5652 6794 5664
rect 7009 5661 7021 5664
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 8128 5688 8156 5732
rect 8312 5732 9772 5760
rect 8312 5688 8340 5732
rect 9766 5720 9772 5732
rect 9824 5720 9830 5772
rect 12158 5760 12164 5772
rect 12119 5732 12164 5760
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 8128 5660 8340 5688
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8444 5664 8489 5692
rect 8444 5652 8450 5664
rect 9398 5652 9404 5704
rect 9456 5692 9462 5704
rect 10965 5695 11023 5701
rect 10965 5692 10977 5695
rect 9456 5664 10977 5692
rect 9456 5652 9462 5664
rect 10965 5661 10977 5664
rect 11011 5692 11023 5695
rect 11054 5692 11060 5704
rect 11011 5664 11060 5692
rect 11011 5661 11023 5664
rect 10965 5655 11023 5661
rect 11054 5652 11060 5664
rect 11112 5692 11118 5704
rect 11241 5695 11299 5701
rect 11241 5692 11253 5695
rect 11112 5664 11253 5692
rect 11112 5652 11118 5664
rect 11241 5661 11253 5664
rect 11287 5661 11299 5695
rect 11241 5655 11299 5661
rect 13265 5695 13323 5701
rect 13265 5661 13277 5695
rect 13311 5692 13323 5695
rect 13725 5695 13783 5701
rect 13725 5692 13737 5695
rect 13311 5664 13737 5692
rect 13311 5661 13323 5664
rect 13265 5655 13323 5661
rect 13725 5661 13737 5664
rect 13771 5692 13783 5695
rect 14458 5692 14464 5704
rect 13771 5664 14464 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 14568 5692 14596 5868
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 15344 5868 15608 5896
rect 15344 5856 15350 5868
rect 15580 5828 15608 5868
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15712 5868 16129 5896
rect 15712 5856 15718 5868
rect 16117 5865 16129 5868
rect 16163 5896 16175 5899
rect 17678 5896 17684 5908
rect 16163 5868 17684 5896
rect 16163 5865 16175 5868
rect 16117 5859 16175 5865
rect 17678 5856 17684 5868
rect 17736 5856 17742 5908
rect 17957 5899 18015 5905
rect 17957 5865 17969 5899
rect 18003 5896 18015 5899
rect 20898 5896 20904 5908
rect 18003 5868 20904 5896
rect 18003 5865 18015 5868
rect 17957 5859 18015 5865
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 16206 5828 16212 5840
rect 15580 5800 16212 5828
rect 16206 5788 16212 5800
rect 16264 5788 16270 5840
rect 19337 5831 19395 5837
rect 19337 5797 19349 5831
rect 19383 5828 19395 5831
rect 19702 5828 19708 5840
rect 19383 5800 19708 5828
rect 19383 5797 19395 5800
rect 19337 5791 19395 5797
rect 19702 5788 19708 5800
rect 19760 5788 19766 5840
rect 20990 5788 20996 5840
rect 21048 5828 21054 5840
rect 21085 5831 21143 5837
rect 21085 5828 21097 5831
rect 21048 5800 21097 5828
rect 21048 5788 21054 5800
rect 21085 5797 21097 5800
rect 21131 5797 21143 5831
rect 21085 5791 21143 5797
rect 15562 5692 15568 5704
rect 14568 5664 15424 5692
rect 15523 5664 15568 5692
rect 3053 5627 3111 5633
rect 3053 5593 3065 5627
rect 3099 5624 3111 5627
rect 3786 5624 3792 5636
rect 3099 5596 3792 5624
rect 3099 5593 3111 5596
rect 3053 5587 3111 5593
rect 3786 5584 3792 5596
rect 3844 5584 3850 5636
rect 6178 5624 6184 5636
rect 4356 5596 5488 5624
rect 6139 5596 6184 5624
rect 2038 5516 2044 5568
rect 2096 5556 2102 5568
rect 2406 5556 2412 5568
rect 2096 5528 2141 5556
rect 2367 5528 2412 5556
rect 2096 5516 2102 5528
rect 2406 5516 2412 5528
rect 2464 5516 2470 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 3145 5559 3203 5565
rect 3145 5525 3157 5559
rect 3191 5556 3203 5559
rect 4356 5556 4384 5596
rect 5460 5568 5488 5596
rect 6178 5584 6184 5596
rect 6236 5584 6242 5636
rect 7561 5627 7619 5633
rect 7561 5593 7573 5627
rect 7607 5624 7619 5627
rect 8938 5624 8944 5636
rect 7607 5596 8944 5624
rect 7607 5593 7619 5596
rect 7561 5587 7619 5593
rect 8938 5584 8944 5596
rect 8996 5584 9002 5636
rect 10042 5584 10048 5636
rect 10100 5624 10106 5636
rect 10698 5627 10756 5633
rect 10698 5624 10710 5627
rect 10100 5596 10710 5624
rect 10100 5584 10106 5596
rect 10698 5593 10710 5596
rect 10744 5593 10756 5627
rect 10698 5587 10756 5593
rect 14366 5584 14372 5636
rect 14424 5624 14430 5636
rect 15298 5627 15356 5633
rect 15298 5624 15310 5627
rect 14424 5596 15310 5624
rect 14424 5584 14430 5596
rect 15298 5593 15310 5596
rect 15344 5593 15356 5627
rect 15396 5624 15424 5664
rect 15562 5652 15568 5664
rect 15620 5692 15626 5704
rect 17402 5692 17408 5704
rect 15620 5664 17408 5692
rect 15620 5652 15626 5664
rect 17402 5652 17408 5664
rect 17460 5692 17466 5704
rect 17497 5695 17555 5701
rect 17497 5692 17509 5695
rect 17460 5664 17509 5692
rect 17460 5652 17466 5664
rect 17497 5661 17509 5664
rect 17543 5661 17555 5695
rect 17770 5692 17776 5704
rect 17731 5664 17776 5692
rect 17497 5655 17555 5661
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18874 5701 18880 5704
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 18869 5692 18880 5701
rect 18279 5664 18736 5692
rect 18835 5664 18880 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 17126 5624 17132 5636
rect 15396 5596 17132 5624
rect 15298 5587 15356 5593
rect 17126 5584 17132 5596
rect 17184 5624 17190 5636
rect 17230 5627 17288 5633
rect 17230 5624 17242 5627
rect 17184 5596 17242 5624
rect 17184 5584 17190 5596
rect 17230 5593 17242 5596
rect 17276 5624 17288 5627
rect 17678 5624 17684 5636
rect 17276 5596 17684 5624
rect 17276 5593 17288 5596
rect 17230 5587 17288 5593
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 3191 5528 4384 5556
rect 3191 5525 3203 5528
rect 3145 5519 3203 5525
rect 4430 5516 4436 5568
rect 4488 5556 4494 5568
rect 4706 5556 4712 5568
rect 4488 5528 4712 5556
rect 4488 5516 4494 5528
rect 4706 5516 4712 5528
rect 4764 5516 4770 5568
rect 5350 5556 5356 5568
rect 5311 5528 5356 5556
rect 5350 5516 5356 5528
rect 5408 5516 5414 5568
rect 5442 5516 5448 5568
rect 5500 5556 5506 5568
rect 6273 5559 6331 5565
rect 6273 5556 6285 5559
rect 5500 5528 6285 5556
rect 5500 5516 5506 5528
rect 6273 5525 6285 5528
rect 6319 5556 6331 5559
rect 7374 5556 7380 5568
rect 6319 5528 7380 5556
rect 6319 5525 6331 5528
rect 6273 5519 6331 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8260 5528 8305 5556
rect 8260 5516 8266 5528
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 10226 5556 10232 5568
rect 8812 5528 10232 5556
rect 8812 5516 8818 5528
rect 10226 5516 10232 5528
rect 10284 5516 10290 5568
rect 11609 5559 11667 5565
rect 11609 5525 11621 5559
rect 11655 5556 11667 5559
rect 11698 5556 11704 5568
rect 11655 5528 11704 5556
rect 11655 5525 11667 5528
rect 11609 5519 11667 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12713 5559 12771 5565
rect 12713 5525 12725 5559
rect 12759 5556 12771 5559
rect 12894 5556 12900 5568
rect 12759 5528 12900 5556
rect 12759 5525 12771 5528
rect 12713 5519 12771 5525
rect 12894 5516 12900 5528
rect 12952 5516 12958 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13630 5556 13636 5568
rect 13587 5528 13636 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 14182 5556 14188 5568
rect 14143 5528 14188 5556
rect 14182 5516 14188 5528
rect 14240 5516 14246 5568
rect 16850 5516 16856 5568
rect 16908 5556 16914 5568
rect 17034 5556 17040 5568
rect 16908 5528 17040 5556
rect 16908 5516 16914 5528
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5556 18475 5559
rect 18506 5556 18512 5568
rect 18463 5528 18512 5556
rect 18463 5525 18475 5528
rect 18417 5519 18475 5525
rect 18506 5516 18512 5528
rect 18564 5516 18570 5568
rect 18708 5565 18736 5664
rect 18869 5655 18880 5664
rect 18874 5652 18880 5655
rect 18932 5652 18938 5704
rect 20162 5652 20168 5704
rect 20220 5692 20226 5704
rect 20714 5692 20720 5704
rect 20220 5664 20576 5692
rect 20675 5664 20720 5692
rect 20220 5652 20226 5664
rect 20438 5624 20444 5636
rect 20496 5633 20502 5636
rect 20408 5596 20444 5624
rect 20438 5584 20444 5596
rect 20496 5587 20508 5633
rect 20548 5624 20576 5664
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 21269 5627 21327 5633
rect 21269 5624 21281 5627
rect 20548 5596 21281 5624
rect 21269 5593 21281 5596
rect 21315 5593 21327 5627
rect 21269 5587 21327 5593
rect 20496 5584 20502 5587
rect 18693 5559 18751 5565
rect 18693 5525 18705 5559
rect 18739 5525 18751 5559
rect 18693 5519 18751 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 2038 5312 2044 5364
rect 2096 5352 2102 5364
rect 3237 5355 3295 5361
rect 3237 5352 3249 5355
rect 2096 5324 3249 5352
rect 2096 5312 2102 5324
rect 3237 5321 3249 5324
rect 3283 5321 3295 5355
rect 3237 5315 3295 5321
rect 4154 5312 4160 5364
rect 4212 5352 4218 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4212 5324 4261 5352
rect 4212 5312 4218 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 4249 5315 4307 5321
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 4890 5352 4896 5364
rect 4387 5324 4896 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 4890 5312 4896 5324
rect 4948 5312 4954 5364
rect 5350 5352 5356 5364
rect 5311 5324 5356 5352
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 6365 5355 6423 5361
rect 6365 5352 6377 5355
rect 5460 5324 6377 5352
rect 1486 5284 1492 5296
rect 1447 5256 1492 5284
rect 1486 5244 1492 5256
rect 1544 5244 1550 5296
rect 2498 5244 2504 5296
rect 2556 5284 2562 5296
rect 2593 5287 2651 5293
rect 2593 5284 2605 5287
rect 2556 5256 2605 5284
rect 2556 5244 2562 5256
rect 2593 5253 2605 5256
rect 2639 5253 2651 5287
rect 2593 5247 2651 5253
rect 2774 5244 2780 5296
rect 2832 5284 2838 5296
rect 3786 5284 3792 5296
rect 2832 5256 3792 5284
rect 2832 5244 2838 5256
rect 3786 5244 3792 5256
rect 3844 5244 3850 5296
rect 4522 5244 4528 5296
rect 4580 5284 4586 5296
rect 5460 5284 5488 5324
rect 6365 5321 6377 5324
rect 6411 5321 6423 5355
rect 6365 5315 6423 5321
rect 6914 5312 6920 5364
rect 6972 5352 6978 5364
rect 7561 5355 7619 5361
rect 7561 5352 7573 5355
rect 6972 5324 7573 5352
rect 6972 5312 6978 5324
rect 7561 5321 7573 5324
rect 7607 5321 7619 5355
rect 7561 5315 7619 5321
rect 8297 5355 8355 5361
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 10962 5352 10968 5364
rect 8343 5324 10968 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11054 5312 11060 5364
rect 11112 5352 11118 5364
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 11112 5324 11529 5352
rect 11112 5312 11118 5324
rect 11517 5321 11529 5324
rect 11563 5352 11575 5355
rect 11790 5352 11796 5364
rect 11563 5324 11796 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 11790 5312 11796 5324
rect 11848 5352 11854 5364
rect 11885 5355 11943 5361
rect 11885 5352 11897 5355
rect 11848 5324 11897 5352
rect 11848 5312 11854 5324
rect 11885 5321 11897 5324
rect 11931 5321 11943 5355
rect 11885 5315 11943 5321
rect 14642 5312 14648 5364
rect 14700 5352 14706 5364
rect 16758 5352 16764 5364
rect 14700 5324 16764 5352
rect 14700 5312 14706 5324
rect 16758 5312 16764 5324
rect 16816 5312 16822 5364
rect 16853 5355 16911 5361
rect 16853 5321 16865 5355
rect 16899 5352 16911 5355
rect 16899 5324 17080 5352
rect 16899 5321 16911 5324
rect 16853 5315 16911 5321
rect 5810 5284 5816 5296
rect 4580 5256 5488 5284
rect 5644 5256 5816 5284
rect 4580 5244 4586 5256
rect 4982 5216 4988 5228
rect 2746 5188 4988 5216
rect 2314 5148 2320 5160
rect 2275 5120 2320 5148
rect 2314 5108 2320 5120
rect 2372 5108 2378 5160
rect 2501 5151 2559 5157
rect 2501 5117 2513 5151
rect 2547 5117 2559 5151
rect 2501 5111 2559 5117
rect 2222 5040 2228 5092
rect 2280 5080 2286 5092
rect 2516 5080 2544 5111
rect 2280 5052 2544 5080
rect 2280 5040 2286 5052
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 2746 5012 2774 5188
rect 4982 5176 4988 5188
rect 5040 5216 5046 5228
rect 5445 5219 5503 5225
rect 5445 5216 5457 5219
rect 5040 5188 5457 5216
rect 5040 5176 5046 5188
rect 5445 5185 5457 5188
rect 5491 5185 5503 5219
rect 5445 5179 5503 5185
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4614 5148 4620 5160
rect 4203 5120 4620 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 5644 5157 5672 5256
rect 5810 5244 5816 5256
rect 5868 5284 5874 5296
rect 12342 5284 12348 5296
rect 5868 5256 12348 5284
rect 5868 5244 5874 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 13572 5287 13630 5293
rect 13572 5284 13584 5287
rect 13372 5256 13584 5284
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6730 5216 6736 5228
rect 6595 5188 6736 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7098 5216 7104 5228
rect 7059 5188 7104 5216
rect 7098 5176 7104 5188
rect 7156 5176 7162 5228
rect 7190 5176 7196 5228
rect 7248 5216 7254 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7248 5188 7757 5216
rect 7248 5176 7254 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 8110 5216 8116 5228
rect 8071 5188 8116 5216
rect 7745 5179 7803 5185
rect 8110 5176 8116 5188
rect 8168 5176 8174 5228
rect 8570 5216 8576 5228
rect 8531 5188 8576 5216
rect 8570 5176 8576 5188
rect 8628 5176 8634 5228
rect 8938 5176 8944 5228
rect 8996 5216 9002 5228
rect 9398 5216 9404 5228
rect 8996 5188 9404 5216
rect 8996 5176 9002 5188
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9657 5219 9715 5225
rect 9657 5216 9669 5219
rect 9508 5188 9669 5216
rect 5629 5151 5687 5157
rect 5629 5117 5641 5151
rect 5675 5117 5687 5151
rect 9508 5148 9536 5188
rect 9657 5185 9669 5188
rect 9703 5185 9715 5219
rect 9657 5179 9715 5185
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 13372 5216 13400 5256
rect 13572 5253 13584 5256
rect 13618 5284 13630 5287
rect 14182 5284 14188 5296
rect 13618 5256 14188 5284
rect 13618 5253 13630 5256
rect 13572 5247 13630 5253
rect 14182 5244 14188 5256
rect 14240 5244 14246 5296
rect 14274 5244 14280 5296
rect 14332 5284 14338 5296
rect 14332 5256 14872 5284
rect 14332 5244 14338 5256
rect 10100 5188 13400 5216
rect 14369 5219 14427 5225
rect 10100 5176 10106 5188
rect 14369 5185 14381 5219
rect 14415 5216 14427 5219
rect 14642 5216 14648 5228
rect 14415 5188 14648 5216
rect 14415 5185 14427 5188
rect 14369 5179 14427 5185
rect 14642 5176 14648 5188
rect 14700 5176 14706 5228
rect 14844 5225 14872 5256
rect 14829 5219 14887 5225
rect 14829 5185 14841 5219
rect 14875 5185 14887 5219
rect 14829 5179 14887 5185
rect 5629 5111 5687 5117
rect 8588 5120 9536 5148
rect 8588 5092 8616 5120
rect 3786 5040 3792 5092
rect 3844 5080 3850 5092
rect 7742 5080 7748 5092
rect 3844 5052 7748 5080
rect 3844 5040 3850 5052
rect 7742 5040 7748 5052
rect 7800 5080 7806 5092
rect 8110 5080 8116 5092
rect 7800 5052 8116 5080
rect 7800 5040 7806 5052
rect 8110 5040 8116 5052
rect 8168 5040 8174 5092
rect 8570 5040 8576 5092
rect 8628 5040 8634 5092
rect 8757 5083 8815 5089
rect 8757 5049 8769 5083
rect 8803 5080 8815 5083
rect 9214 5080 9220 5092
rect 8803 5052 9220 5080
rect 8803 5049 8815 5052
rect 8757 5043 8815 5049
rect 9214 5040 9220 5052
rect 9272 5040 9278 5092
rect 2958 5012 2964 5024
rect 1627 4984 2774 5012
rect 2919 4984 2964 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 2958 4972 2964 4984
rect 3016 4972 3022 5024
rect 4706 5012 4712 5024
rect 4667 4984 4712 5012
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 4985 5015 5043 5021
rect 4985 5012 4997 5015
rect 4948 4984 4997 5012
rect 4948 4972 4954 4984
rect 4985 4981 4997 4984
rect 5031 4981 5043 5015
rect 4985 4975 5043 4981
rect 7285 5015 7343 5021
rect 7285 4981 7297 5015
rect 7331 5012 7343 5015
rect 7374 5012 7380 5024
rect 7331 4984 7380 5012
rect 7331 4981 7343 4984
rect 7285 4975 7343 4981
rect 7374 4972 7380 4984
rect 7432 4972 7438 5024
rect 9122 5012 9128 5024
rect 9083 4984 9128 5012
rect 9122 4972 9128 4984
rect 9180 4972 9186 5024
rect 9416 5012 9444 5120
rect 12342 5108 12348 5160
rect 12400 5148 12406 5160
rect 12618 5148 12624 5160
rect 12400 5120 12624 5148
rect 12400 5108 12406 5120
rect 12452 5089 12480 5120
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 13817 5151 13875 5157
rect 13817 5117 13829 5151
rect 13863 5117 13875 5151
rect 14844 5148 14872 5179
rect 15378 5176 15384 5228
rect 15436 5216 15442 5228
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15436 5188 15485 5216
rect 15436 5176 15442 5188
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15746 5216 15752 5228
rect 15707 5188 15752 5216
rect 15473 5179 15531 5185
rect 15488 5148 15516 5179
rect 15746 5176 15752 5188
rect 15804 5176 15810 5228
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5216 16727 5219
rect 16942 5216 16948 5228
rect 16715 5188 16948 5216
rect 16715 5185 16727 5188
rect 16669 5179 16727 5185
rect 16942 5176 16948 5188
rect 17000 5176 17006 5228
rect 17052 5216 17080 5324
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17310 5352 17316 5364
rect 17184 5324 17316 5352
rect 17184 5312 17190 5324
rect 17310 5312 17316 5324
rect 17368 5352 17374 5364
rect 19702 5352 19708 5364
rect 17368 5324 19708 5352
rect 17368 5312 17374 5324
rect 19702 5312 19708 5324
rect 19760 5312 19766 5364
rect 19978 5352 19984 5364
rect 19939 5324 19984 5352
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 20346 5352 20352 5364
rect 20307 5324 20352 5352
rect 20346 5312 20352 5324
rect 20404 5312 20410 5364
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 21085 5355 21143 5361
rect 21085 5321 21097 5355
rect 21131 5352 21143 5355
rect 21450 5352 21456 5364
rect 21131 5324 21456 5352
rect 21131 5321 21143 5324
rect 21085 5315 21143 5321
rect 21450 5312 21456 5324
rect 21508 5312 21514 5364
rect 18414 5244 18420 5296
rect 18472 5284 18478 5296
rect 20993 5287 21051 5293
rect 20993 5284 21005 5287
rect 18472 5256 21005 5284
rect 18472 5244 18478 5256
rect 20993 5253 21005 5256
rect 21039 5253 21051 5287
rect 20993 5247 21051 5253
rect 17129 5219 17187 5225
rect 17129 5216 17141 5219
rect 17052 5188 17141 5216
rect 17129 5185 17141 5188
rect 17175 5185 17187 5219
rect 17586 5216 17592 5228
rect 17547 5188 17592 5216
rect 17129 5179 17187 5185
rect 17586 5176 17592 5188
rect 17644 5176 17650 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 17736 5188 18337 5216
rect 17736 5176 17742 5188
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18874 5216 18880 5228
rect 18835 5188 18880 5216
rect 18325 5179 18383 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 18598 5148 18604 5160
rect 14844 5120 15424 5148
rect 15488 5120 18604 5148
rect 13817 5111 13875 5117
rect 12437 5083 12495 5089
rect 10612 5052 11192 5080
rect 10612 5012 10640 5052
rect 10778 5012 10784 5024
rect 9416 4984 10640 5012
rect 10739 4984 10784 5012
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 11164 5021 11192 5052
rect 12437 5049 12449 5083
rect 12483 5049 12495 5083
rect 12437 5043 12495 5049
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11330 5012 11336 5024
rect 11195 4984 11336 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 13832 5012 13860 5111
rect 14274 5040 14280 5092
rect 14332 5080 14338 5092
rect 15289 5083 15347 5089
rect 15289 5080 15301 5083
rect 14332 5052 15301 5080
rect 14332 5040 14338 5052
rect 15289 5049 15301 5052
rect 15335 5049 15347 5083
rect 15396 5080 15424 5120
rect 18598 5108 18604 5120
rect 18656 5108 18662 5160
rect 19702 5148 19708 5160
rect 19663 5120 19708 5148
rect 19702 5108 19708 5120
rect 19760 5108 19766 5160
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5148 19947 5151
rect 20622 5148 20628 5160
rect 19935 5120 20628 5148
rect 19935 5117 19947 5120
rect 19889 5111 19947 5117
rect 20622 5108 20628 5120
rect 20680 5108 20686 5160
rect 21174 5148 21180 5160
rect 21135 5120 21180 5148
rect 21174 5108 21180 5120
rect 21232 5108 21238 5160
rect 18509 5083 18567 5089
rect 15396 5052 18000 5080
rect 15289 5043 15347 5049
rect 17972 5024 18000 5052
rect 18509 5049 18521 5083
rect 18555 5080 18567 5083
rect 20254 5080 20260 5092
rect 18555 5052 20260 5080
rect 18555 5049 18567 5052
rect 18509 5043 18567 5049
rect 20254 5040 20260 5052
rect 20312 5040 20318 5092
rect 11848 4984 13860 5012
rect 14553 5015 14611 5021
rect 11848 4972 11854 4984
rect 14553 4981 14565 5015
rect 14599 5012 14611 5015
rect 14918 5012 14924 5024
rect 14599 4984 14924 5012
rect 14599 4981 14611 4984
rect 14553 4975 14611 4981
rect 14918 4972 14924 4984
rect 14976 4972 14982 5024
rect 15013 5015 15071 5021
rect 15013 4981 15025 5015
rect 15059 5012 15071 5015
rect 15746 5012 15752 5024
rect 15059 4984 15752 5012
rect 15059 4981 15071 4984
rect 15013 4975 15071 4981
rect 15746 4972 15752 4984
rect 15804 4972 15810 5024
rect 15933 5015 15991 5021
rect 15933 4981 15945 5015
rect 15979 5012 15991 5015
rect 16022 5012 16028 5024
rect 15979 4984 16028 5012
rect 15979 4981 15991 4984
rect 15933 4975 15991 4981
rect 16022 4972 16028 4984
rect 16080 4972 16086 5024
rect 16301 5015 16359 5021
rect 16301 4981 16313 5015
rect 16347 5012 16359 5015
rect 16390 5012 16396 5024
rect 16347 4984 16396 5012
rect 16347 4981 16359 4984
rect 16301 4975 16359 4981
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 17313 5015 17371 5021
rect 17313 4981 17325 5015
rect 17359 5012 17371 5015
rect 17402 5012 17408 5024
rect 17359 4984 17408 5012
rect 17359 4981 17371 4984
rect 17313 4975 17371 4981
rect 17402 4972 17408 4984
rect 17460 4972 17466 5024
rect 17586 4972 17592 5024
rect 17644 5012 17650 5024
rect 17773 5015 17831 5021
rect 17773 5012 17785 5015
rect 17644 4984 17785 5012
rect 17644 4972 17650 4984
rect 17773 4981 17785 4984
rect 17819 4981 17831 5015
rect 17773 4975 17831 4981
rect 17954 4972 17960 5024
rect 18012 4972 18018 5024
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 18840 4984 19073 5012
rect 18840 4972 18846 4984
rect 19061 4981 19073 4984
rect 19107 4981 19119 5015
rect 19061 4975 19119 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 3234 4808 3240 4820
rect 3195 4780 3240 4808
rect 3234 4768 3240 4780
rect 3292 4768 3298 4820
rect 3973 4811 4031 4817
rect 3973 4777 3985 4811
rect 4019 4808 4031 4811
rect 5534 4808 5540 4820
rect 4019 4780 5540 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 6365 4811 6423 4817
rect 6365 4777 6377 4811
rect 6411 4808 6423 4811
rect 7098 4808 7104 4820
rect 6411 4780 7104 4808
rect 6411 4777 6423 4780
rect 6365 4771 6423 4777
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 7561 4811 7619 4817
rect 7561 4808 7573 4811
rect 7524 4780 7573 4808
rect 7524 4768 7530 4780
rect 7561 4777 7573 4780
rect 7607 4777 7619 4811
rect 7561 4771 7619 4777
rect 8110 4768 8116 4820
rect 8168 4808 8174 4820
rect 8938 4808 8944 4820
rect 8168 4780 8944 4808
rect 8168 4768 8174 4780
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9398 4768 9404 4820
rect 9456 4808 9462 4820
rect 9953 4811 10011 4817
rect 9953 4808 9965 4811
rect 9456 4780 9965 4808
rect 9456 4768 9462 4780
rect 9953 4777 9965 4780
rect 9999 4777 10011 4811
rect 10410 4808 10416 4820
rect 10371 4780 10416 4808
rect 9953 4771 10011 4777
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 14734 4808 14740 4820
rect 10888 4780 12434 4808
rect 3878 4740 3884 4752
rect 2240 4712 3884 4740
rect 1946 4672 1952 4684
rect 1907 4644 1952 4672
rect 1946 4632 1952 4644
rect 2004 4632 2010 4684
rect 2240 4616 2268 4712
rect 3878 4700 3884 4712
rect 3936 4700 3942 4752
rect 4706 4700 4712 4752
rect 4764 4740 4770 4752
rect 7285 4743 7343 4749
rect 4764 4712 5948 4740
rect 4764 4700 4770 4712
rect 2685 4675 2743 4681
rect 2685 4641 2697 4675
rect 2731 4672 2743 4675
rect 3694 4672 3700 4684
rect 2731 4644 3700 4672
rect 2731 4641 2743 4644
rect 2685 4635 2743 4641
rect 3694 4632 3700 4644
rect 3752 4632 3758 4684
rect 4614 4672 4620 4684
rect 4575 4644 4620 4672
rect 4614 4632 4620 4644
rect 4672 4632 4678 4684
rect 4801 4675 4859 4681
rect 4801 4641 4813 4675
rect 4847 4672 4859 4675
rect 5166 4672 5172 4684
rect 4847 4644 5172 4672
rect 4847 4641 4859 4644
rect 4801 4635 4859 4641
rect 5166 4632 5172 4644
rect 5224 4632 5230 4684
rect 5920 4681 5948 4712
rect 6472 4712 7236 4740
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4641 5871 4675
rect 5813 4635 5871 4641
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 2406 4564 2412 4616
rect 2464 4604 2470 4616
rect 2869 4607 2927 4613
rect 2869 4604 2881 4607
rect 2464 4576 2881 4604
rect 2464 4564 2470 4576
rect 2869 4573 2881 4576
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3789 4607 3847 4613
rect 3789 4604 3801 4607
rect 3292 4576 3801 4604
rect 3292 4564 3298 4576
rect 3789 4573 3801 4576
rect 3835 4573 3847 4607
rect 4890 4604 4896 4616
rect 4851 4576 4896 4604
rect 3789 4567 3847 4573
rect 4890 4564 4896 4576
rect 4948 4564 4954 4616
rect 5828 4604 5856 4635
rect 6472 4604 6500 4712
rect 6546 4632 6552 4684
rect 6604 4672 6610 4684
rect 7208 4672 7236 4712
rect 7285 4709 7297 4743
rect 7331 4740 7343 4743
rect 9582 4740 9588 4752
rect 7331 4712 9588 4740
rect 7331 4709 7343 4712
rect 7285 4703 7343 4709
rect 9582 4700 9588 4712
rect 9640 4700 9646 4752
rect 9677 4743 9735 4749
rect 9677 4709 9689 4743
rect 9723 4740 9735 4743
rect 10888 4740 10916 4780
rect 9723 4712 10916 4740
rect 12406 4740 12434 4780
rect 12728 4780 14740 4808
rect 12728 4740 12756 4780
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 14829 4811 14887 4817
rect 14829 4777 14841 4811
rect 14875 4808 14887 4811
rect 14918 4808 14924 4820
rect 14875 4780 14924 4808
rect 14875 4777 14887 4780
rect 14829 4771 14887 4777
rect 14918 4768 14924 4780
rect 14976 4768 14982 4820
rect 15102 4808 15108 4820
rect 15063 4780 15108 4808
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 19702 4808 19708 4820
rect 15488 4780 19708 4808
rect 12406 4712 12756 4740
rect 9723 4709 9735 4712
rect 9677 4703 9735 4709
rect 9125 4675 9183 4681
rect 6604 4644 6868 4672
rect 7208 4644 9076 4672
rect 6604 4632 6610 4644
rect 6840 4613 6868 4644
rect 5828 4576 6500 4604
rect 6825 4607 6883 4613
rect 6825 4573 6837 4607
rect 6871 4573 6883 4607
rect 6825 4567 6883 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7101 4567 7159 4573
rect 2777 4539 2835 4545
rect 2777 4505 2789 4539
rect 2823 4536 2835 4539
rect 4798 4536 4804 4548
rect 2823 4508 4804 4536
rect 2823 4505 2835 4508
rect 2777 4499 2835 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 5997 4539 6055 4545
rect 5997 4536 6009 4539
rect 5276 4508 6009 4536
rect 1762 4428 1768 4480
rect 1820 4468 1826 4480
rect 5166 4468 5172 4480
rect 1820 4440 5172 4468
rect 1820 4428 1826 4440
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 5276 4477 5304 4508
rect 5997 4505 6009 4508
rect 6043 4505 6055 4539
rect 5997 4499 6055 4505
rect 6546 4496 6552 4548
rect 6604 4536 6610 4548
rect 7116 4536 7144 4567
rect 7558 4564 7564 4616
rect 7616 4604 7622 4616
rect 7745 4607 7803 4613
rect 7745 4604 7757 4607
rect 7616 4576 7757 4604
rect 7616 4564 7622 4576
rect 7745 4573 7757 4576
rect 7791 4573 7803 4607
rect 7745 4567 7803 4573
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8389 4607 8447 4613
rect 8389 4604 8401 4607
rect 8076 4576 8401 4604
rect 8076 4564 8082 4576
rect 8389 4573 8401 4576
rect 8435 4573 8447 4607
rect 9048 4604 9076 4644
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 10594 4672 10600 4684
rect 9171 4644 10600 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 11790 4672 11796 4684
rect 11751 4644 11796 4672
rect 11790 4632 11796 4644
rect 11848 4672 11854 4684
rect 15378 4672 15384 4684
rect 11848 4644 12434 4672
rect 11848 4632 11854 4644
rect 11537 4607 11595 4613
rect 9048 4576 9720 4604
rect 8389 4567 8447 4573
rect 6604 4508 7144 4536
rect 6604 4496 6610 4508
rect 7834 4496 7840 4548
rect 7892 4536 7898 4548
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 7892 4508 9321 4536
rect 7892 4496 7898 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9309 4499 9367 4505
rect 5261 4471 5319 4477
rect 5261 4437 5273 4471
rect 5307 4437 5319 4471
rect 5261 4431 5319 4437
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5626 4468 5632 4480
rect 5408 4440 5632 4468
rect 5408 4428 5414 4440
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 6638 4468 6644 4480
rect 6599 4440 6644 4468
rect 6638 4428 6644 4440
rect 6696 4428 6702 4480
rect 6730 4428 6736 4480
rect 6788 4468 6794 4480
rect 8205 4471 8263 4477
rect 8205 4468 8217 4471
rect 6788 4440 8217 4468
rect 6788 4428 6794 4440
rect 8205 4437 8217 4440
rect 8251 4437 8263 4471
rect 8205 4431 8263 4437
rect 8938 4428 8944 4480
rect 8996 4468 9002 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8996 4440 9229 4468
rect 8996 4428 9002 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9692 4468 9720 4576
rect 11537 4573 11549 4607
rect 11583 4604 11595 4607
rect 11698 4604 11704 4616
rect 11583 4576 11704 4604
rect 11583 4573 11595 4576
rect 11537 4567 11595 4573
rect 11698 4564 11704 4576
rect 11756 4564 11762 4616
rect 12406 4604 12434 4644
rect 14384 4644 15384 4672
rect 14384 4613 14412 4644
rect 15378 4632 15384 4644
rect 15436 4632 15442 4684
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 12406 4576 13645 4604
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4604 14703 4607
rect 15488 4604 15516 4780
rect 19702 4768 19708 4780
rect 19760 4768 19766 4820
rect 20162 4808 20168 4820
rect 19812 4780 20168 4808
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 19812 4740 19840 4780
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 21082 4740 21088 4752
rect 19475 4712 19840 4740
rect 21043 4712 21088 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 21082 4700 21088 4712
rect 21140 4700 21146 4752
rect 16390 4604 16396 4616
rect 14691 4576 15516 4604
rect 15580 4576 16396 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 10134 4496 10140 4548
rect 10192 4536 10198 4548
rect 10686 4536 10692 4548
rect 10192 4508 10692 4536
rect 10192 4496 10198 4508
rect 10686 4496 10692 4508
rect 10744 4536 10750 4548
rect 13366 4539 13424 4545
rect 13366 4536 13378 4539
rect 10744 4508 13378 4536
rect 10744 4496 10750 4508
rect 13366 4505 13378 4508
rect 13412 4505 13424 4539
rect 13648 4536 13676 4567
rect 15580 4548 15608 4576
rect 16390 4564 16396 4576
rect 16448 4604 16454 4616
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16448 4576 16497 4604
rect 16448 4564 16454 4576
rect 16485 4573 16497 4576
rect 16531 4604 16543 4607
rect 18233 4607 18291 4613
rect 18233 4604 18245 4607
rect 16531 4576 18245 4604
rect 16531 4573 16543 4576
rect 16485 4567 16543 4573
rect 18233 4573 18245 4576
rect 18279 4573 18291 4607
rect 18506 4604 18512 4616
rect 18467 4576 18512 4604
rect 18233 4567 18291 4573
rect 15562 4536 15568 4548
rect 13648 4508 15568 4536
rect 13366 4499 13424 4505
rect 15562 4496 15568 4508
rect 15620 4496 15626 4548
rect 15930 4496 15936 4548
rect 15988 4536 15994 4548
rect 16218 4539 16276 4545
rect 16218 4536 16230 4539
rect 15988 4508 16230 4536
rect 15988 4496 15994 4508
rect 16218 4505 16230 4508
rect 16264 4536 16276 4539
rect 17988 4539 18046 4545
rect 16264 4508 16896 4536
rect 16264 4505 16276 4508
rect 16218 4499 16276 4505
rect 9766 4468 9772 4480
rect 9692 4440 9772 4468
rect 9217 4431 9275 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 10928 4440 12265 4468
rect 10928 4428 10934 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 13722 4428 13728 4480
rect 13780 4468 13786 4480
rect 16868 4477 16896 4508
rect 17988 4505 18000 4539
rect 18034 4536 18046 4539
rect 18138 4536 18144 4548
rect 18034 4508 18144 4536
rect 18034 4505 18046 4508
rect 17988 4499 18046 4505
rect 18138 4496 18144 4508
rect 18196 4496 18202 4548
rect 18248 4536 18276 4567
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 20714 4604 20720 4616
rect 19904 4576 20720 4604
rect 19904 4548 19932 4576
rect 20714 4564 20720 4576
rect 20772 4604 20778 4616
rect 20809 4607 20867 4613
rect 20809 4604 20821 4607
rect 20772 4576 20821 4604
rect 20772 4564 20778 4576
rect 20809 4573 20821 4576
rect 20855 4573 20867 4607
rect 21266 4604 21272 4616
rect 21227 4576 21272 4604
rect 20809 4567 20867 4573
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 19886 4536 19892 4548
rect 18248 4508 19892 4536
rect 19886 4496 19892 4508
rect 19944 4496 19950 4548
rect 20564 4539 20622 4545
rect 20564 4505 20576 4539
rect 20610 4536 20622 4539
rect 21174 4536 21180 4548
rect 20610 4508 21180 4536
rect 20610 4505 20622 4508
rect 20564 4499 20622 4505
rect 21174 4496 21180 4508
rect 21232 4496 21238 4548
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 13780 4440 14197 4468
rect 13780 4428 13786 4440
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 14185 4431 14243 4437
rect 16853 4471 16911 4477
rect 16853 4437 16865 4471
rect 16899 4468 16911 4471
rect 17310 4468 17316 4480
rect 16899 4440 17316 4468
rect 16899 4437 16911 4440
rect 16853 4431 16911 4437
rect 17310 4428 17316 4440
rect 17368 4428 17374 4480
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 18693 4471 18751 4477
rect 18693 4468 18705 4471
rect 18472 4440 18705 4468
rect 18472 4428 18478 4440
rect 18693 4437 18705 4440
rect 18739 4437 18751 4471
rect 18693 4431 18751 4437
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 1578 4264 1584 4276
rect 1539 4236 1584 4264
rect 1578 4224 1584 4236
rect 1636 4224 1642 4276
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3016 4236 3801 4264
rect 3016 4224 3022 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 3789 4227 3847 4233
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 5997 4267 6055 4273
rect 4672 4236 5580 4264
rect 4672 4224 4678 4236
rect 3050 4156 3056 4208
rect 3108 4196 3114 4208
rect 3237 4199 3295 4205
rect 3237 4196 3249 4199
rect 3108 4168 3249 4196
rect 3108 4156 3114 4168
rect 3237 4165 3249 4168
rect 3283 4196 3295 4199
rect 3510 4196 3516 4208
rect 3283 4168 3516 4196
rect 3283 4165 3295 4168
rect 3237 4159 3295 4165
rect 3510 4156 3516 4168
rect 3568 4156 3574 4208
rect 3881 4199 3939 4205
rect 3881 4165 3893 4199
rect 3927 4196 3939 4199
rect 4246 4196 4252 4208
rect 3927 4168 4252 4196
rect 3927 4165 3939 4168
rect 3881 4159 3939 4165
rect 4246 4156 4252 4168
rect 4304 4156 4310 4208
rect 5552 4196 5580 4236
rect 5997 4233 6009 4267
rect 6043 4264 6055 4267
rect 6546 4264 6552 4276
rect 6043 4236 6552 4264
rect 6043 4233 6055 4236
rect 5997 4227 6055 4233
rect 6546 4224 6552 4236
rect 6604 4224 6610 4276
rect 6914 4224 6920 4276
rect 6972 4264 6978 4276
rect 7558 4264 7564 4276
rect 6972 4236 7564 4264
rect 6972 4224 6978 4236
rect 7558 4224 7564 4236
rect 7616 4224 7622 4276
rect 7834 4264 7840 4276
rect 7795 4236 7840 4264
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 7944 4236 10640 4264
rect 7944 4196 7972 4236
rect 10612 4208 10640 4236
rect 11238 4224 11244 4276
rect 11296 4264 11302 4276
rect 11330 4264 11336 4276
rect 11296 4236 11336 4264
rect 11296 4224 11302 4236
rect 11330 4224 11336 4236
rect 11388 4224 11394 4276
rect 15746 4224 15752 4276
rect 15804 4264 15810 4276
rect 17497 4267 17555 4273
rect 17497 4264 17509 4267
rect 15804 4236 17509 4264
rect 15804 4224 15810 4236
rect 17497 4233 17509 4236
rect 17543 4264 17555 4267
rect 18046 4264 18052 4276
rect 17543 4236 18052 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 5552 4168 7972 4196
rect 8938 4156 8944 4208
rect 8996 4196 9002 4208
rect 8996 4168 9041 4196
rect 8996 4156 9002 4168
rect 10594 4156 10600 4208
rect 10652 4196 10658 4208
rect 10882 4199 10940 4205
rect 10882 4196 10894 4199
rect 10652 4168 10894 4196
rect 10652 4156 10658 4168
rect 10882 4165 10894 4168
rect 10928 4165 10940 4199
rect 10882 4159 10940 4165
rect 11701 4199 11759 4205
rect 11701 4165 11713 4199
rect 11747 4196 11759 4199
rect 12158 4196 12164 4208
rect 11747 4168 12164 4196
rect 11747 4165 11759 4168
rect 11701 4159 11759 4165
rect 12158 4156 12164 4168
rect 12216 4156 12222 4208
rect 13556 4168 13860 4196
rect 1394 4128 1400 4140
rect 1355 4100 1400 4128
rect 1394 4088 1400 4100
rect 1452 4088 1458 4140
rect 2498 4128 2504 4140
rect 2459 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4088 2562 4140
rect 2590 4088 2596 4140
rect 2648 4128 2654 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 2648 4100 4537 4128
rect 2648 4088 2654 4100
rect 4525 4097 4537 4100
rect 4571 4128 4583 4131
rect 4706 4128 4712 4140
rect 4571 4100 4712 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4706 4088 4712 4100
rect 4764 4088 4770 4140
rect 4893 4131 4951 4137
rect 4893 4097 4905 4131
rect 4939 4128 4951 4131
rect 4982 4128 4988 4140
rect 4939 4100 4988 4128
rect 4939 4097 4951 4100
rect 4893 4091 4951 4097
rect 4982 4088 4988 4100
rect 5040 4088 5046 4140
rect 5350 4128 5356 4140
rect 5311 4100 5356 4128
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5810 4128 5816 4140
rect 5771 4100 5816 4128
rect 5810 4088 5816 4100
rect 5868 4088 5874 4140
rect 5902 4088 5908 4140
rect 5960 4128 5966 4140
rect 6365 4131 6423 4137
rect 6365 4128 6377 4131
rect 5960 4100 6377 4128
rect 5960 4088 5966 4100
rect 6365 4097 6377 4100
rect 6411 4097 6423 4131
rect 7009 4131 7067 4137
rect 7009 4128 7021 4131
rect 6365 4091 6423 4097
rect 6564 4100 7021 4128
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4029 2375 4063
rect 2317 4023 2375 4029
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 2682 4060 2688 4072
rect 2455 4032 2688 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 2332 3992 2360 4023
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 3697 4063 3755 4069
rect 3697 4060 3709 4063
rect 2792 4032 3709 4060
rect 2792 3992 2820 4032
rect 3697 4029 3709 4032
rect 3743 4060 3755 4063
rect 6178 4060 6184 4072
rect 3743 4032 6184 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 2332 3964 2820 3992
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 4154 3992 4160 4004
rect 2915 3964 4160 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 4154 3952 4160 3964
rect 4212 3952 4218 4004
rect 5074 3992 5080 4004
rect 5035 3964 5080 3992
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 6564 4001 6592 4100
rect 7009 4097 7021 4100
rect 7055 4097 7067 4131
rect 7650 4128 7656 4140
rect 7611 4100 7656 4128
rect 7009 4091 7067 4097
rect 7650 4088 7656 4100
rect 7708 4088 7714 4140
rect 8294 4128 8300 4140
rect 8255 4100 8300 4128
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 11517 4131 11575 4137
rect 11517 4128 11529 4131
rect 8404 4100 11529 4128
rect 7098 4020 7104 4072
rect 7156 4060 7162 4072
rect 8404 4060 8432 4100
rect 11517 4097 11529 4100
rect 11563 4097 11575 4131
rect 12250 4128 12256 4140
rect 12211 4100 12256 4128
rect 11517 4091 11575 4097
rect 12250 4088 12256 4100
rect 12308 4088 12314 4140
rect 12805 4131 12863 4137
rect 12805 4097 12817 4131
rect 12851 4097 12863 4131
rect 12805 4091 12863 4097
rect 13265 4131 13323 4137
rect 13265 4097 13277 4131
rect 13311 4128 13323 4131
rect 13556 4128 13584 4168
rect 13722 4128 13728 4140
rect 13311 4100 13584 4128
rect 13683 4100 13728 4128
rect 13311 4097 13323 4100
rect 13265 4091 13323 4097
rect 7156 4032 8432 4060
rect 8665 4063 8723 4069
rect 7156 4020 7162 4032
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 8846 4060 8852 4072
rect 8807 4032 8852 4060
rect 8665 4023 8723 4029
rect 6549 3995 6607 4001
rect 5224 3964 5672 3992
rect 5224 3952 5230 3964
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 4338 3924 4344 3936
rect 4295 3896 4344 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 4338 3884 4344 3896
rect 4396 3884 4402 3936
rect 5534 3924 5540 3936
rect 5495 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5644 3924 5672 3964
rect 6549 3961 6561 3995
rect 6595 3961 6607 3995
rect 6549 3955 6607 3961
rect 7282 3952 7288 4004
rect 7340 3992 7346 4004
rect 8680 3992 8708 4023
rect 8846 4020 8852 4032
rect 8904 4020 8910 4072
rect 8938 4020 8944 4072
rect 8996 4060 9002 4072
rect 8996 4032 9904 4060
rect 8996 4020 9002 4032
rect 9306 3992 9312 4004
rect 7340 3964 8708 3992
rect 9267 3964 9312 3992
rect 7340 3952 7346 3964
rect 9306 3952 9312 3964
rect 9364 3952 9370 4004
rect 9766 3992 9772 4004
rect 9727 3964 9772 3992
rect 9766 3952 9772 3964
rect 9824 3952 9830 4004
rect 7098 3924 7104 3936
rect 5644 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7193 3927 7251 3933
rect 7193 3893 7205 3927
rect 7239 3924 7251 3927
rect 7742 3924 7748 3936
rect 7239 3896 7748 3924
rect 7239 3893 7251 3896
rect 7193 3887 7251 3893
rect 7742 3884 7748 3896
rect 7800 3884 7806 3936
rect 8110 3924 8116 3936
rect 8071 3896 8116 3924
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 9398 3924 9404 3936
rect 8904 3896 9404 3924
rect 8904 3884 8910 3896
rect 9398 3884 9404 3896
rect 9456 3924 9462 3936
rect 9582 3924 9588 3936
rect 9456 3896 9588 3924
rect 9456 3884 9462 3896
rect 9582 3884 9588 3896
rect 9640 3884 9646 3936
rect 9876 3924 9904 4032
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11790 4060 11796 4072
rect 11204 4032 11796 4060
rect 11204 4020 11210 4032
rect 11790 4020 11796 4032
rect 11848 4020 11854 4072
rect 12820 4060 12848 4091
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 13832 4128 13860 4168
rect 15194 4156 15200 4208
rect 15252 4156 15258 4208
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 19794 4196 19800 4208
rect 15436 4168 18184 4196
rect 15436 4156 15442 4168
rect 15212 4128 15240 4156
rect 18156 4140 18184 4168
rect 19720 4168 19800 4196
rect 13832 4100 15240 4128
rect 15286 4088 15292 4140
rect 15344 4137 15350 4140
rect 15344 4128 15356 4137
rect 15562 4128 15568 4140
rect 15344 4100 15389 4128
rect 15523 4100 15568 4128
rect 15344 4091 15356 4100
rect 15344 4088 15350 4091
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 15841 4131 15899 4137
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 16666 4128 16672 4140
rect 16627 4100 16672 4128
rect 15841 4091 15899 4097
rect 14274 4060 14280 4072
rect 12820 4032 14280 4060
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 13906 3992 13912 4004
rect 11164 3964 13768 3992
rect 13867 3964 13912 3992
rect 11164 3924 11192 3964
rect 9876 3896 11192 3924
rect 11882 3884 11888 3936
rect 11940 3924 11946 3936
rect 12069 3927 12127 3933
rect 12069 3924 12081 3927
rect 11940 3896 12081 3924
rect 11940 3884 11946 3896
rect 12069 3893 12081 3896
rect 12115 3893 12127 3927
rect 12986 3924 12992 3936
rect 12947 3896 12992 3924
rect 12069 3887 12127 3893
rect 12986 3884 12992 3896
rect 13044 3884 13050 3936
rect 13449 3927 13507 3933
rect 13449 3893 13461 3927
rect 13495 3924 13507 3927
rect 13538 3924 13544 3936
rect 13495 3896 13544 3924
rect 13495 3893 13507 3896
rect 13449 3887 13507 3893
rect 13538 3884 13544 3896
rect 13596 3884 13602 3936
rect 13740 3924 13768 3964
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 14185 3995 14243 4001
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 14366 3992 14372 4004
rect 14231 3964 14372 3992
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 14200 3924 14228 3955
rect 14366 3952 14372 3964
rect 14424 3952 14430 4004
rect 13740 3896 14228 3924
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 15856 3924 15884 4091
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 17494 4088 17500 4140
rect 17552 4128 17558 4140
rect 17589 4131 17647 4137
rect 17589 4128 17601 4131
rect 17552 4100 17601 4128
rect 17552 4088 17558 4100
rect 17589 4097 17601 4100
rect 17635 4097 17647 4131
rect 18138 4128 18144 4140
rect 18051 4100 18144 4128
rect 17589 4091 17647 4097
rect 18138 4088 18144 4100
rect 18196 4088 18202 4140
rect 19334 4128 19340 4140
rect 18708 4100 19340 4128
rect 17770 4060 17776 4072
rect 17731 4032 17776 4060
rect 17770 4020 17776 4032
rect 17828 4020 17834 4072
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16853 3995 16911 4001
rect 15988 3964 16528 3992
rect 15988 3952 15994 3964
rect 14332 3896 15884 3924
rect 16025 3927 16083 3933
rect 14332 3884 14338 3896
rect 16025 3893 16037 3927
rect 16071 3924 16083 3927
rect 16298 3924 16304 3936
rect 16071 3896 16304 3924
rect 16071 3893 16083 3896
rect 16025 3887 16083 3893
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16500 3924 16528 3964
rect 16853 3961 16865 3995
rect 16899 3992 16911 3995
rect 17862 3992 17868 4004
rect 16899 3964 17868 3992
rect 16899 3961 16911 3964
rect 16853 3955 16911 3961
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 18509 3995 18567 4001
rect 18509 3961 18521 3995
rect 18555 3992 18567 3995
rect 18708 3992 18736 4100
rect 19334 4088 19340 4100
rect 19392 4088 19398 4140
rect 19633 4131 19691 4137
rect 19633 4097 19645 4131
rect 19679 4128 19691 4131
rect 19720 4128 19748 4168
rect 19794 4156 19800 4168
rect 19852 4156 19858 4208
rect 20714 4196 20720 4208
rect 20675 4168 20720 4196
rect 20714 4156 20720 4168
rect 20772 4156 20778 4208
rect 19886 4128 19892 4140
rect 19679 4100 19748 4128
rect 19847 4100 19892 4128
rect 19679 4097 19691 4100
rect 19633 4091 19691 4097
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 20806 4128 20812 4140
rect 20767 4100 20812 4128
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 20530 4020 20536 4072
rect 20588 4060 20594 4072
rect 20901 4063 20959 4069
rect 20901 4060 20913 4063
rect 20588 4032 20913 4060
rect 20588 4020 20594 4032
rect 20901 4029 20913 4032
rect 20947 4029 20959 4063
rect 20901 4023 20959 4029
rect 18555 3964 18736 3992
rect 18555 3961 18567 3964
rect 18509 3955 18567 3961
rect 17129 3927 17187 3933
rect 17129 3924 17141 3927
rect 16500 3896 17141 3924
rect 17129 3893 17141 3896
rect 17175 3893 17187 3927
rect 17129 3887 17187 3893
rect 18598 3884 18604 3936
rect 18656 3924 18662 3936
rect 20349 3927 20407 3933
rect 20349 3924 20361 3927
rect 18656 3896 20361 3924
rect 18656 3884 18662 3896
rect 20349 3893 20361 3896
rect 20395 3893 20407 3927
rect 20349 3887 20407 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2498 3680 2504 3732
rect 2556 3720 2562 3732
rect 2593 3723 2651 3729
rect 2593 3720 2605 3723
rect 2556 3692 2605 3720
rect 2556 3680 2562 3692
rect 2593 3689 2605 3692
rect 2639 3689 2651 3723
rect 2593 3683 2651 3689
rect 2961 3723 3019 3729
rect 2961 3689 2973 3723
rect 3007 3720 3019 3723
rect 3007 3692 4752 3720
rect 3007 3689 3019 3692
rect 2961 3683 3019 3689
rect 3881 3655 3939 3661
rect 3881 3621 3893 3655
rect 3927 3621 3939 3655
rect 4724 3652 4752 3692
rect 4798 3680 4804 3732
rect 4856 3720 4862 3732
rect 4893 3723 4951 3729
rect 4893 3720 4905 3723
rect 4856 3692 4905 3720
rect 4856 3680 4862 3692
rect 4893 3689 4905 3692
rect 4939 3689 4951 3723
rect 4893 3683 4951 3689
rect 8113 3723 8171 3729
rect 8113 3689 8125 3723
rect 8159 3720 8171 3723
rect 13630 3720 13636 3732
rect 8159 3692 13636 3720
rect 8159 3689 8171 3692
rect 8113 3683 8171 3689
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 13725 3723 13783 3729
rect 13725 3689 13737 3723
rect 13771 3720 13783 3723
rect 14274 3720 14280 3732
rect 13771 3692 14280 3720
rect 13771 3689 13783 3692
rect 13725 3683 13783 3689
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 15565 3723 15623 3729
rect 14424 3692 14469 3720
rect 14424 3680 14430 3692
rect 15565 3689 15577 3723
rect 15611 3720 15623 3723
rect 16666 3720 16672 3732
rect 15611 3692 16672 3720
rect 15611 3689 15623 3692
rect 15565 3683 15623 3689
rect 16666 3680 16672 3692
rect 16724 3680 16730 3732
rect 17218 3680 17224 3732
rect 17276 3720 17282 3732
rect 17865 3723 17923 3729
rect 17865 3720 17877 3723
rect 17276 3692 17877 3720
rect 17276 3680 17282 3692
rect 17865 3689 17877 3692
rect 17911 3689 17923 3723
rect 17865 3683 17923 3689
rect 18138 3680 18144 3732
rect 18196 3720 18202 3732
rect 19610 3720 19616 3732
rect 18196 3692 19196 3720
rect 19571 3692 19616 3720
rect 18196 3680 18202 3692
rect 5074 3652 5080 3664
rect 4724 3624 5080 3652
rect 3881 3615 3939 3621
rect 2041 3587 2099 3593
rect 2041 3553 2053 3587
rect 2087 3584 2099 3587
rect 2314 3584 2320 3596
rect 2087 3556 2320 3584
rect 2087 3553 2099 3556
rect 2041 3547 2099 3553
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2133 3519 2191 3525
rect 2133 3485 2145 3519
rect 2179 3516 2191 3519
rect 3050 3516 3056 3528
rect 2179 3488 3056 3516
rect 2179 3485 2191 3488
rect 2133 3479 2191 3485
rect 3050 3476 3056 3488
rect 3108 3476 3114 3528
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3896 3516 3924 3615
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 5534 3612 5540 3664
rect 5592 3652 5598 3664
rect 10686 3652 10692 3664
rect 5592 3624 9444 3652
rect 10647 3624 10692 3652
rect 5592 3612 5598 3624
rect 9416 3596 9444 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 12529 3655 12587 3661
rect 12529 3621 12541 3655
rect 12575 3621 12587 3655
rect 12529 3615 12587 3621
rect 4338 3584 4344 3596
rect 4299 3556 4344 3584
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 4522 3584 4528 3596
rect 4483 3556 4528 3584
rect 4522 3544 4528 3556
rect 4580 3544 4586 3596
rect 4706 3544 4712 3596
rect 4764 3584 4770 3596
rect 5445 3587 5503 3593
rect 5445 3584 5457 3587
rect 4764 3556 5457 3584
rect 4764 3544 4770 3556
rect 5445 3553 5457 3556
rect 5491 3584 5503 3587
rect 5810 3584 5816 3596
rect 5491 3556 5816 3584
rect 5491 3553 5503 3556
rect 5445 3547 5503 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 5994 3544 6000 3596
rect 6052 3584 6058 3596
rect 6089 3587 6147 3593
rect 6089 3584 6101 3587
rect 6052 3556 6101 3584
rect 6052 3544 6058 3556
rect 6089 3553 6101 3556
rect 6135 3553 6147 3587
rect 8202 3584 8208 3596
rect 6089 3547 6147 3553
rect 7484 3556 8208 3584
rect 3283 3488 3924 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 4154 3476 4160 3528
rect 4212 3516 4218 3528
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4212 3488 4261 3516
rect 4212 3476 4218 3488
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3516 6423 3519
rect 6546 3516 6552 3528
rect 6411 3488 6552 3516
rect 6411 3485 6423 3488
rect 6365 3479 6423 3485
rect 6546 3476 6552 3488
rect 6604 3516 6610 3528
rect 6730 3516 6736 3528
rect 6604 3488 6736 3516
rect 6604 3476 6610 3488
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 7484 3525 7512 3556
rect 8202 3544 8208 3556
rect 8260 3544 8266 3596
rect 8754 3544 8760 3596
rect 8812 3584 8818 3596
rect 9398 3584 9404 3596
rect 8812 3556 9260 3584
rect 9311 3556 9404 3584
rect 8812 3544 8818 3556
rect 7009 3519 7067 3525
rect 7009 3485 7021 3519
rect 7055 3485 7067 3519
rect 7009 3479 7067 3485
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7926 3516 7932 3528
rect 7887 3488 7932 3516
rect 7469 3479 7527 3485
rect 1581 3451 1639 3457
rect 1581 3417 1593 3451
rect 1627 3448 1639 3451
rect 2225 3451 2283 3457
rect 2225 3448 2237 3451
rect 1627 3420 2237 3448
rect 1627 3417 1639 3420
rect 1581 3411 1639 3417
rect 2225 3417 2237 3420
rect 2271 3417 2283 3451
rect 7024 3448 7052 3479
rect 7926 3476 7932 3488
rect 7984 3476 7990 3528
rect 8573 3519 8631 3525
rect 8573 3485 8585 3519
rect 8619 3516 8631 3519
rect 8662 3516 8668 3528
rect 8619 3488 8668 3516
rect 8619 3485 8631 3488
rect 8573 3479 8631 3485
rect 8662 3476 8668 3488
rect 8720 3516 8726 3528
rect 9122 3516 9128 3528
rect 8720 3488 9128 3516
rect 8720 3476 8726 3488
rect 9122 3476 9128 3488
rect 9180 3476 9186 3528
rect 9232 3516 9260 3556
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 9508 3516 9536 3547
rect 9582 3544 9588 3596
rect 9640 3584 9646 3596
rect 12069 3587 12127 3593
rect 9640 3556 10824 3584
rect 9640 3544 9646 3556
rect 9232 3488 9536 3516
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 2225 3411 2283 3417
rect 3436 3420 7052 3448
rect 3436 3389 3464 3420
rect 8018 3408 8024 3460
rect 8076 3448 8082 3460
rect 10152 3448 10180 3479
rect 8076 3420 10180 3448
rect 8076 3408 8082 3420
rect 3421 3383 3479 3389
rect 3421 3349 3433 3383
rect 3467 3349 3479 3383
rect 3421 3343 3479 3349
rect 3878 3340 3884 3392
rect 3936 3380 3942 3392
rect 4430 3380 4436 3392
rect 3936 3352 4436 3380
rect 3936 3340 3942 3352
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 5258 3380 5264 3392
rect 5219 3352 5264 3380
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 5408 3352 5453 3380
rect 5408 3340 5414 3352
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 5902 3380 5908 3392
rect 5684 3352 5908 3380
rect 5684 3340 5690 3352
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6273 3383 6331 3389
rect 6273 3380 6285 3383
rect 6052 3352 6285 3380
rect 6052 3340 6058 3352
rect 6273 3349 6285 3352
rect 6319 3349 6331 3383
rect 6730 3380 6736 3392
rect 6691 3352 6736 3380
rect 6273 3343 6331 3349
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7193 3383 7251 3389
rect 7193 3349 7205 3383
rect 7239 3380 7251 3383
rect 7282 3380 7288 3392
rect 7239 3352 7288 3380
rect 7239 3349 7251 3352
rect 7193 3343 7251 3349
rect 7282 3340 7288 3352
rect 7340 3340 7346 3392
rect 7650 3380 7656 3392
rect 7611 3352 7656 3380
rect 7650 3340 7656 3352
rect 7708 3340 7714 3392
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8478 3380 8484 3392
rect 8435 3352 8484 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8938 3380 8944 3392
rect 8899 3352 8944 3380
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10502 3380 10508 3392
rect 10367 3352 10508 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10796 3380 10824 3556
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12434 3584 12440 3596
rect 12115 3556 12440 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 12434 3544 12440 3556
rect 12492 3544 12498 3596
rect 12544 3584 12572 3615
rect 12986 3612 12992 3664
rect 13044 3652 13050 3664
rect 16761 3655 16819 3661
rect 13044 3624 16160 3652
rect 13044 3612 13050 3624
rect 13814 3584 13820 3596
rect 12544 3556 13820 3584
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 15010 3584 15016 3596
rect 14971 3556 15016 3584
rect 15010 3544 15016 3556
rect 15068 3544 15074 3596
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 12345 3519 12403 3525
rect 12345 3516 12357 3519
rect 11020 3488 12357 3516
rect 11020 3476 11026 3488
rect 12345 3485 12357 3488
rect 12391 3485 12403 3519
rect 12345 3479 12403 3485
rect 12894 3476 12900 3528
rect 12952 3516 12958 3528
rect 12989 3519 13047 3525
rect 12989 3516 13001 3519
rect 12952 3488 13001 3516
rect 12952 3476 12958 3488
rect 12989 3485 13001 3488
rect 13035 3485 13047 3519
rect 12989 3479 13047 3485
rect 13446 3476 13452 3528
rect 13504 3516 13510 3528
rect 13541 3519 13599 3525
rect 13541 3516 13553 3519
rect 13504 3488 13553 3516
rect 13504 3476 13510 3488
rect 13541 3485 13553 3488
rect 13587 3485 13599 3519
rect 14734 3516 14740 3528
rect 14695 3488 14740 3516
rect 13541 3479 13599 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 15378 3516 15384 3528
rect 15339 3488 15384 3516
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15470 3476 15476 3528
rect 15528 3516 15534 3528
rect 16025 3519 16083 3525
rect 16025 3516 16037 3519
rect 15528 3488 16037 3516
rect 15528 3476 15534 3488
rect 16025 3485 16037 3488
rect 16071 3485 16083 3519
rect 16132 3516 16160 3624
rect 16761 3621 16773 3655
rect 16807 3652 16819 3655
rect 16807 3624 19012 3652
rect 16807 3621 16819 3624
rect 16761 3615 16819 3621
rect 16390 3544 16396 3596
rect 16448 3584 16454 3596
rect 16448 3556 16712 3584
rect 16448 3544 16454 3556
rect 16577 3519 16635 3525
rect 16577 3516 16589 3519
rect 16132 3488 16589 3516
rect 16025 3479 16083 3485
rect 16577 3485 16589 3488
rect 16623 3485 16635 3519
rect 16684 3516 16712 3556
rect 17126 3544 17132 3596
rect 17184 3584 17190 3596
rect 17221 3587 17279 3593
rect 17221 3584 17233 3587
rect 17184 3556 17233 3584
rect 17184 3544 17190 3556
rect 17221 3553 17233 3556
rect 17267 3553 17279 3587
rect 17221 3547 17279 3553
rect 17405 3587 17463 3593
rect 17405 3553 17417 3587
rect 17451 3584 17463 3587
rect 18598 3584 18604 3596
rect 17451 3556 18604 3584
rect 17451 3553 17463 3556
rect 17405 3547 17463 3553
rect 18598 3544 18604 3556
rect 18656 3544 18662 3596
rect 18785 3587 18843 3593
rect 18785 3553 18797 3587
rect 18831 3584 18843 3587
rect 18874 3584 18880 3596
rect 18831 3556 18880 3584
rect 18831 3553 18843 3556
rect 18785 3547 18843 3553
rect 18874 3544 18880 3556
rect 18932 3544 18938 3596
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 16684 3488 17509 3516
rect 16577 3479 16635 3485
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 18984 3516 19012 3624
rect 19058 3516 19064 3528
rect 18984 3488 19064 3516
rect 17497 3479 17555 3485
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 19168 3516 19196 3692
rect 19610 3680 19616 3692
rect 19668 3680 19674 3732
rect 20622 3720 20628 3732
rect 20583 3692 20628 3720
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 19337 3655 19395 3661
rect 19337 3621 19349 3655
rect 19383 3652 19395 3655
rect 19702 3652 19708 3664
rect 19383 3624 19708 3652
rect 19383 3621 19395 3624
rect 19337 3615 19395 3621
rect 19702 3612 19708 3624
rect 19760 3612 19766 3664
rect 19242 3544 19248 3596
rect 19300 3584 19306 3596
rect 20257 3587 20315 3593
rect 19300 3556 19932 3584
rect 19300 3544 19306 3556
rect 19794 3516 19800 3528
rect 19168 3488 19800 3516
rect 19794 3476 19800 3488
rect 19852 3476 19858 3528
rect 19904 3516 19932 3556
rect 20257 3553 20269 3587
rect 20303 3584 20315 3587
rect 20530 3584 20536 3596
rect 20303 3556 20536 3584
rect 20303 3553 20315 3556
rect 20257 3547 20315 3553
rect 20530 3544 20536 3556
rect 20588 3584 20594 3596
rect 21177 3587 21235 3593
rect 21177 3584 21189 3587
rect 20588 3556 21189 3584
rect 20588 3544 20594 3556
rect 21177 3553 21189 3556
rect 21223 3553 21235 3587
rect 21177 3547 21235 3553
rect 20993 3519 21051 3525
rect 20993 3516 21005 3519
rect 19904 3488 21005 3516
rect 20993 3485 21005 3488
rect 21039 3485 21051 3519
rect 20993 3479 21051 3485
rect 21085 3519 21143 3525
rect 21085 3485 21097 3519
rect 21131 3516 21143 3519
rect 21450 3516 21456 3528
rect 21131 3488 21456 3516
rect 21131 3485 21143 3488
rect 21085 3479 21143 3485
rect 21450 3476 21456 3488
rect 21508 3476 21514 3528
rect 11824 3451 11882 3457
rect 11824 3417 11836 3451
rect 11870 3448 11882 3451
rect 11974 3448 11980 3460
rect 11870 3420 11980 3448
rect 11870 3417 11882 3420
rect 11824 3411 11882 3417
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 12158 3408 12164 3460
rect 12216 3448 12222 3460
rect 12912 3448 12940 3476
rect 12216 3420 12940 3448
rect 14829 3451 14887 3457
rect 12216 3408 12222 3420
rect 14829 3417 14841 3451
rect 14875 3448 14887 3451
rect 14875 3420 18184 3448
rect 14875 3417 14887 3420
rect 14829 3411 14887 3417
rect 12805 3383 12863 3389
rect 12805 3380 12817 3383
rect 10796 3352 12817 3380
rect 12805 3349 12817 3352
rect 12851 3349 12863 3383
rect 12805 3343 12863 3349
rect 16209 3383 16267 3389
rect 16209 3349 16221 3383
rect 16255 3380 16267 3383
rect 17770 3380 17776 3392
rect 16255 3352 17776 3380
rect 16255 3349 16267 3352
rect 16209 3343 16267 3349
rect 17770 3340 17776 3352
rect 17828 3340 17834 3392
rect 18156 3389 18184 3420
rect 18322 3408 18328 3460
rect 18380 3448 18386 3460
rect 18509 3451 18567 3457
rect 18509 3448 18521 3451
rect 18380 3420 18521 3448
rect 18380 3408 18386 3420
rect 18509 3417 18521 3420
rect 18555 3417 18567 3451
rect 18509 3411 18567 3417
rect 18601 3451 18659 3457
rect 18601 3417 18613 3451
rect 18647 3448 18659 3451
rect 18966 3448 18972 3460
rect 18647 3420 18972 3448
rect 18647 3417 18659 3420
rect 18601 3411 18659 3417
rect 18966 3408 18972 3420
rect 19024 3448 19030 3460
rect 20073 3451 20131 3457
rect 20073 3448 20085 3451
rect 19024 3420 20085 3448
rect 19024 3408 19030 3420
rect 20073 3417 20085 3420
rect 20119 3417 20131 3451
rect 20073 3411 20131 3417
rect 18141 3383 18199 3389
rect 18141 3349 18153 3383
rect 18187 3349 18199 3383
rect 19978 3380 19984 3392
rect 19939 3352 19984 3380
rect 18141 3343 18199 3349
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1118 3136 1124 3188
rect 1176 3176 1182 3188
rect 2590 3176 2596 3188
rect 1176 3148 2596 3176
rect 1176 3136 1182 3148
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 3237 3179 3295 3185
rect 2832 3148 2877 3176
rect 2832 3136 2838 3148
rect 3237 3145 3249 3179
rect 3283 3145 3295 3179
rect 3237 3139 3295 3145
rect 3789 3179 3847 3185
rect 3789 3145 3801 3179
rect 3835 3176 3847 3179
rect 3878 3176 3884 3188
rect 3835 3148 3884 3176
rect 3835 3145 3847 3148
rect 3789 3139 3847 3145
rect 934 3068 940 3120
rect 992 3108 998 3120
rect 3252 3108 3280 3139
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4246 3176 4252 3188
rect 4207 3148 4252 3176
rect 4246 3136 4252 3148
rect 4304 3136 4310 3188
rect 8662 3136 8668 3188
rect 8720 3176 8726 3188
rect 13541 3179 13599 3185
rect 13541 3176 13553 3179
rect 8720 3148 13553 3176
rect 8720 3136 8726 3148
rect 13541 3145 13553 3148
rect 13587 3145 13599 3179
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 13541 3139 13599 3145
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 16669 3179 16727 3185
rect 16669 3145 16681 3179
rect 16715 3176 16727 3179
rect 16942 3176 16948 3188
rect 16715 3148 16948 3176
rect 16715 3145 16727 3148
rect 16669 3139 16727 3145
rect 16942 3136 16948 3148
rect 17000 3136 17006 3188
rect 17037 3179 17095 3185
rect 17037 3145 17049 3179
rect 17083 3176 17095 3179
rect 17681 3179 17739 3185
rect 17681 3176 17693 3179
rect 17083 3148 17693 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17681 3145 17693 3148
rect 17727 3145 17739 3179
rect 17681 3139 17739 3145
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 19518 3176 19524 3188
rect 17828 3148 19524 3176
rect 17828 3136 17834 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 5994 3108 6000 3120
rect 992 3080 2774 3108
rect 3252 3080 6000 3108
rect 992 3068 998 3080
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2130 3040 2136 3052
rect 1995 3012 2136 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2590 3040 2596 3052
rect 2551 3012 2596 3040
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 2746 3040 2774 3080
rect 5994 3068 6000 3080
rect 6052 3108 6058 3120
rect 6825 3111 6883 3117
rect 6825 3108 6837 3111
rect 6052 3080 6837 3108
rect 6052 3068 6058 3080
rect 6825 3077 6837 3080
rect 6871 3077 6883 3111
rect 9490 3108 9496 3120
rect 6825 3071 6883 3077
rect 8864 3080 9496 3108
rect 3053 3043 3111 3049
rect 3053 3040 3065 3043
rect 2746 3012 3065 3040
rect 3053 3009 3065 3012
rect 3099 3040 3111 3043
rect 3881 3043 3939 3049
rect 3099 3012 3740 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 14 2932 20 2984
rect 72 2972 78 2984
rect 934 2972 940 2984
rect 72 2944 940 2972
rect 72 2932 78 2944
rect 934 2932 940 2944
rect 992 2972 998 2984
rect 2225 2975 2283 2981
rect 2225 2972 2237 2975
rect 992 2944 2237 2972
rect 992 2932 998 2944
rect 2225 2941 2237 2944
rect 2271 2941 2283 2975
rect 3605 2975 3663 2981
rect 3605 2972 3617 2975
rect 2225 2935 2283 2941
rect 2746 2944 3617 2972
rect 2314 2864 2320 2916
rect 2372 2904 2378 2916
rect 2746 2904 2774 2944
rect 3605 2941 3617 2944
rect 3651 2941 3663 2975
rect 3712 2972 3740 3012
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 4246 3040 4252 3052
rect 3927 3012 4252 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4430 3000 4436 3052
rect 4488 3040 4494 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 4488 3012 5365 3040
rect 4488 3000 4494 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 6638 3040 6644 3052
rect 5859 3012 6644 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3009 6791 3043
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 6733 3003 6791 3009
rect 5077 2975 5135 2981
rect 3712 2944 4660 2972
rect 3605 2935 3663 2941
rect 2372 2876 2774 2904
rect 4632 2904 4660 2944
rect 5077 2941 5089 2975
rect 5123 2972 5135 2975
rect 5442 2972 5448 2984
rect 5123 2944 5448 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 6546 2932 6552 2984
rect 6604 2972 6610 2984
rect 6748 2972 6776 3003
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8202 3040 8208 3052
rect 7883 3012 8208 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 8864 3040 8892 3080
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9766 3068 9772 3120
rect 9824 3108 9830 3120
rect 10882 3111 10940 3117
rect 10882 3108 10894 3111
rect 9824 3080 10894 3108
rect 9824 3068 9830 3080
rect 10882 3077 10894 3080
rect 10928 3077 10940 3111
rect 10882 3071 10940 3077
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 12342 3108 12348 3120
rect 11388 3080 12348 3108
rect 11388 3068 11394 3080
rect 12342 3068 12348 3080
rect 12400 3108 12406 3120
rect 12400 3080 12940 3108
rect 12400 3068 12406 3080
rect 8481 3027 8539 3033
rect 8481 2993 8493 3027
rect 8527 3024 8539 3027
rect 8680 3024 8892 3040
rect 8527 3012 8892 3024
rect 8941 3043 8999 3049
rect 8527 2996 8708 3012
rect 8941 3009 8953 3043
rect 8987 3009 8999 3043
rect 9214 3040 9220 3052
rect 9175 3012 9220 3040
rect 8941 3003 8999 3009
rect 8527 2993 8539 2996
rect 8481 2987 8539 2993
rect 6604 2944 6776 2972
rect 7009 2975 7067 2981
rect 6604 2932 6610 2944
rect 7009 2941 7021 2975
rect 7055 2972 7067 2975
rect 7098 2972 7104 2984
rect 7055 2944 7104 2972
rect 7055 2941 7067 2944
rect 7009 2935 7067 2941
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 8294 2972 8300 2984
rect 8220 2944 8300 2972
rect 5534 2904 5540 2916
rect 4632 2876 5540 2904
rect 2372 2864 2378 2876
rect 5534 2864 5540 2876
rect 5592 2864 5598 2916
rect 5997 2907 6055 2913
rect 5997 2873 6009 2907
rect 6043 2904 6055 2907
rect 8220 2904 8248 2944
rect 8294 2932 8300 2944
rect 8352 2932 8358 2984
rect 8386 2932 8392 2984
rect 8444 2932 8450 2984
rect 8956 2972 8984 3003
rect 9214 3000 9220 3012
rect 9272 3000 9278 3052
rect 10594 3000 10600 3052
rect 10652 3040 10658 3052
rect 11149 3043 11207 3049
rect 10652 3012 11100 3040
rect 10652 3000 10658 3012
rect 9950 2972 9956 2984
rect 8956 2944 9956 2972
rect 9950 2932 9956 2944
rect 10008 2932 10014 2984
rect 11072 2972 11100 3012
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11348 3040 11376 3068
rect 11195 3012 11376 3040
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 12618 3000 12624 3052
rect 12676 3049 12682 3052
rect 12912 3049 12940 3080
rect 14090 3068 14096 3120
rect 14148 3108 14154 3120
rect 18046 3108 18052 3120
rect 14148 3080 15884 3108
rect 18007 3080 18052 3108
rect 14148 3068 14154 3080
rect 12676 3040 12688 3049
rect 12897 3043 12955 3049
rect 12676 3012 12721 3040
rect 12676 3003 12688 3012
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 12897 3003 12955 3009
rect 13188 3012 14197 3040
rect 12676 3000 12682 3003
rect 11072 2944 11560 2972
rect 6043 2876 8248 2904
rect 8404 2904 8432 2932
rect 11532 2913 11560 2944
rect 11517 2907 11575 2913
rect 8404 2876 9904 2904
rect 6043 2873 6055 2876
rect 5997 2867 6055 2873
rect 1026 2796 1032 2848
rect 1084 2836 1090 2848
rect 4062 2836 4068 2848
rect 1084 2808 4068 2836
rect 1084 2796 1090 2808
rect 4062 2796 4068 2808
rect 4120 2836 4126 2848
rect 4522 2836 4528 2848
rect 4120 2808 4528 2836
rect 4120 2796 4126 2808
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 4982 2796 4988 2848
rect 5040 2836 5046 2848
rect 5902 2836 5908 2848
rect 5040 2808 5908 2836
rect 5040 2796 5046 2808
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6362 2836 6368 2848
rect 6323 2808 6368 2836
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6914 2796 6920 2848
rect 6972 2836 6978 2848
rect 7374 2836 7380 2848
rect 6972 2808 7380 2836
rect 6972 2796 6978 2808
rect 7374 2796 7380 2808
rect 7432 2796 7438 2848
rect 7558 2836 7564 2848
rect 7519 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 8018 2836 8024 2848
rect 7979 2808 8024 2836
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8352 2808 8397 2836
rect 8352 2796 8358 2808
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8628 2808 8769 2836
rect 8628 2796 8634 2808
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8757 2799 8815 2805
rect 9401 2839 9459 2845
rect 9401 2805 9413 2839
rect 9447 2836 9459 2839
rect 9582 2836 9588 2848
rect 9447 2808 9588 2836
rect 9447 2805 9459 2808
rect 9401 2799 9459 2805
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 9766 2836 9772 2848
rect 9727 2808 9772 2836
rect 9766 2796 9772 2808
rect 9824 2796 9830 2848
rect 9876 2836 9904 2876
rect 11517 2873 11529 2907
rect 11563 2873 11575 2907
rect 11517 2867 11575 2873
rect 13188 2836 13216 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 15856 3049 15884 3080
rect 18046 3068 18052 3080
rect 18104 3068 18110 3120
rect 18138 3068 18144 3120
rect 18196 3108 18202 3120
rect 19242 3108 19248 3120
rect 18196 3080 19248 3108
rect 18196 3068 18202 3080
rect 19242 3068 19248 3080
rect 19300 3068 19306 3120
rect 19334 3068 19340 3120
rect 19392 3108 19398 3120
rect 20070 3108 20076 3120
rect 19392 3080 20076 3108
rect 19392 3068 19398 3080
rect 20070 3068 20076 3080
rect 20128 3068 20134 3120
rect 14737 3043 14795 3049
rect 14737 3040 14749 3043
rect 14700 3012 14749 3040
rect 14700 3000 14706 3012
rect 14737 3009 14749 3012
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 15289 3043 15347 3049
rect 15289 3009 15301 3043
rect 15335 3009 15347 3043
rect 15289 3003 15347 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 15841 3003 15899 3009
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13446 2972 13452 2984
rect 13320 2944 13365 2972
rect 13407 2944 13452 2972
rect 13320 2932 13326 2944
rect 13446 2932 13452 2944
rect 13504 2932 13510 2984
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 15304 2972 15332 3003
rect 17494 3000 17500 3052
rect 17552 3040 17558 3052
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 17552 3012 19073 3040
rect 17552 3000 17558 3012
rect 19061 3009 19073 3012
rect 19107 3040 19119 3043
rect 19978 3040 19984 3052
rect 19107 3012 19984 3040
rect 19107 3009 19119 3012
rect 19061 3003 19119 3009
rect 19978 3000 19984 3012
rect 20036 3000 20042 3052
rect 20162 3040 20168 3052
rect 20123 3012 20168 3040
rect 20162 3000 20168 3012
rect 20220 3040 20226 3052
rect 20622 3040 20628 3052
rect 20220 3012 20628 3040
rect 20220 3000 20226 3012
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 13688 2944 15332 2972
rect 17129 2975 17187 2981
rect 13688 2932 13694 2944
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17310 2972 17316 2984
rect 17271 2944 17316 2972
rect 17129 2935 17187 2941
rect 13280 2876 14044 2904
rect 13280 2848 13308 2876
rect 9876 2808 13216 2836
rect 13262 2796 13268 2848
rect 13320 2796 13326 2848
rect 14016 2836 14044 2876
rect 14274 2864 14280 2916
rect 14332 2904 14338 2916
rect 14332 2876 14504 2904
rect 14332 2864 14338 2876
rect 14369 2839 14427 2845
rect 14369 2836 14381 2839
rect 14016 2808 14381 2836
rect 14369 2805 14381 2808
rect 14415 2805 14427 2839
rect 14476 2836 14504 2876
rect 14734 2864 14740 2916
rect 14792 2904 14798 2916
rect 14792 2876 15056 2904
rect 14792 2864 14798 2876
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 14476 2808 14933 2836
rect 14369 2799 14427 2805
rect 14921 2805 14933 2808
rect 14967 2805 14979 2839
rect 15028 2836 15056 2876
rect 15102 2864 15108 2916
rect 15160 2904 15166 2916
rect 16025 2907 16083 2913
rect 16025 2904 16037 2907
rect 15160 2876 16037 2904
rect 15160 2864 15166 2876
rect 16025 2873 16037 2876
rect 16071 2873 16083 2907
rect 17144 2904 17172 2935
rect 17310 2932 17316 2944
rect 17368 2932 17374 2984
rect 18230 2972 18236 2984
rect 18191 2944 18236 2972
rect 18230 2932 18236 2944
rect 18288 2972 18294 2984
rect 19153 2975 19211 2981
rect 18288 2944 19104 2972
rect 18288 2932 18294 2944
rect 18693 2907 18751 2913
rect 18693 2904 18705 2907
rect 17144 2876 18705 2904
rect 16025 2867 16083 2873
rect 18693 2873 18705 2876
rect 18739 2873 18751 2907
rect 19076 2904 19104 2944
rect 19153 2941 19165 2975
rect 19199 2972 19211 2975
rect 19242 2972 19248 2984
rect 19199 2944 19248 2972
rect 19199 2941 19211 2944
rect 19153 2935 19211 2941
rect 19242 2932 19248 2944
rect 19300 2932 19306 2984
rect 19337 2975 19395 2981
rect 19337 2941 19349 2975
rect 19383 2941 19395 2975
rect 19337 2935 19395 2941
rect 19352 2904 19380 2935
rect 19886 2932 19892 2984
rect 19944 2972 19950 2984
rect 20349 2975 20407 2981
rect 20349 2972 20361 2975
rect 19944 2944 20361 2972
rect 19944 2932 19950 2944
rect 20349 2941 20361 2944
rect 20395 2941 20407 2975
rect 20349 2935 20407 2941
rect 19076 2876 19380 2904
rect 18693 2867 18751 2873
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 15028 2808 15485 2836
rect 14921 2799 14979 2805
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 17954 2796 17960 2848
rect 18012 2836 18018 2848
rect 21269 2839 21327 2845
rect 21269 2836 21281 2839
rect 18012 2808 21281 2836
rect 18012 2796 18018 2808
rect 21269 2805 21281 2808
rect 21315 2805 21327 2839
rect 21269 2799 21327 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 3418 2632 3424 2644
rect 1903 2604 3424 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 3418 2592 3424 2604
rect 3476 2632 3482 2644
rect 4246 2632 4252 2644
rect 3476 2604 4252 2632
rect 3476 2592 3482 2604
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4614 2592 4620 2644
rect 4672 2592 4678 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 8938 2632 8944 2644
rect 5408 2604 8944 2632
rect 5408 2592 5414 2604
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 11054 2632 11060 2644
rect 9079 2604 11060 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 11054 2592 11060 2604
rect 11112 2632 11118 2644
rect 11330 2632 11336 2644
rect 11112 2604 11336 2632
rect 11112 2592 11118 2604
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 13446 2592 13452 2644
rect 13504 2632 13510 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 13504 2604 13645 2632
rect 13504 2592 13510 2604
rect 13633 2601 13645 2604
rect 13679 2601 13691 2635
rect 13633 2595 13691 2601
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 15933 2635 15991 2641
rect 15933 2632 15945 2635
rect 14424 2604 15945 2632
rect 14424 2592 14430 2604
rect 15933 2601 15945 2604
rect 15979 2601 15991 2635
rect 15933 2595 15991 2601
rect 16022 2592 16028 2644
rect 16080 2632 16086 2644
rect 16080 2604 17908 2632
rect 16080 2592 16086 2604
rect 2409 2567 2467 2573
rect 2409 2533 2421 2567
rect 2455 2564 2467 2567
rect 2590 2564 2596 2576
rect 2455 2536 2596 2564
rect 2455 2533 2467 2536
rect 2409 2527 2467 2533
rect 2590 2524 2596 2536
rect 2648 2524 2654 2576
rect 2961 2567 3019 2573
rect 2961 2533 2973 2567
rect 3007 2564 3019 2567
rect 4632 2564 4660 2592
rect 3007 2536 4660 2564
rect 6825 2567 6883 2573
rect 3007 2533 3019 2536
rect 2961 2527 3019 2533
rect 6825 2533 6837 2567
rect 6871 2564 6883 2567
rect 9306 2564 9312 2576
rect 6871 2536 9312 2564
rect 6871 2533 6883 2536
rect 6825 2527 6883 2533
rect 9306 2524 9312 2536
rect 9364 2524 9370 2576
rect 9766 2564 9772 2576
rect 9727 2536 9772 2564
rect 9766 2524 9772 2536
rect 9824 2524 9830 2576
rect 15381 2567 15439 2573
rect 15381 2564 15393 2567
rect 9876 2536 12434 2564
rect 4522 2456 4528 2508
rect 4580 2496 4586 2508
rect 4617 2499 4675 2505
rect 4617 2496 4629 2499
rect 4580 2468 4629 2496
rect 4580 2456 4586 2468
rect 4617 2465 4629 2468
rect 4663 2465 4675 2499
rect 5442 2496 5448 2508
rect 5403 2468 5448 2496
rect 4617 2459 4675 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 7098 2456 7104 2508
rect 7156 2496 7162 2508
rect 7929 2499 7987 2505
rect 7929 2496 7941 2499
rect 7156 2468 7941 2496
rect 7156 2456 7162 2468
rect 7929 2465 7941 2468
rect 7975 2496 7987 2499
rect 8202 2496 8208 2508
rect 7975 2468 8208 2496
rect 7975 2465 7987 2468
rect 7929 2459 7987 2465
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 9582 2456 9588 2508
rect 9640 2496 9646 2508
rect 9876 2496 9904 2536
rect 11974 2496 11980 2508
rect 9640 2468 9904 2496
rect 11935 2468 11980 2496
rect 9640 2456 9646 2468
rect 11974 2456 11980 2468
rect 12032 2456 12038 2508
rect 1302 2388 1308 2440
rect 1360 2428 1366 2440
rect 1673 2431 1731 2437
rect 1673 2428 1685 2431
rect 1360 2400 1685 2428
rect 1360 2388 1366 2400
rect 1673 2397 1685 2400
rect 1719 2428 1731 2431
rect 1719 2400 2636 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 750 2320 756 2372
rect 808 2360 814 2372
rect 2222 2360 2228 2372
rect 808 2332 2228 2360
rect 808 2320 814 2332
rect 2222 2320 2228 2332
rect 2280 2320 2286 2372
rect 2608 2292 2636 2400
rect 2774 2388 2780 2440
rect 2832 2428 2838 2440
rect 3237 2431 3295 2437
rect 2832 2400 2877 2428
rect 2832 2388 2838 2400
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 4341 2431 4399 2437
rect 3283 2400 4292 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3694 2360 3700 2372
rect 2746 2332 3700 2360
rect 2746 2292 2774 2332
rect 3694 2320 3700 2332
rect 3752 2320 3758 2372
rect 2608 2264 2774 2292
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 4154 2292 4160 2304
rect 3467 2264 4160 2292
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4264 2292 4292 2400
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 5718 2428 5724 2440
rect 5679 2400 5724 2428
rect 4341 2391 4399 2397
rect 4356 2360 4384 2391
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6641 2431 6699 2437
rect 6641 2397 6653 2431
rect 6687 2428 6699 2431
rect 7650 2428 7656 2440
rect 6687 2400 7512 2428
rect 7611 2400 7656 2428
rect 6687 2397 6699 2400
rect 6641 2391 6699 2397
rect 7006 2360 7012 2372
rect 4356 2332 7012 2360
rect 7006 2320 7012 2332
rect 7064 2320 7070 2372
rect 7484 2360 7512 2400
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8570 2428 8576 2440
rect 8531 2400 8576 2428
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9674 2428 9680 2440
rect 9539 2400 9680 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10318 2428 10324 2440
rect 10279 2400 10324 2428
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10594 2428 10600 2440
rect 10555 2400 10600 2428
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12250 2428 12256 2440
rect 11848 2400 12256 2428
rect 11848 2388 11854 2400
rect 12250 2388 12256 2400
rect 12308 2388 12314 2440
rect 7484 2332 8524 2360
rect 6638 2292 6644 2304
rect 4264 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 8386 2292 8392 2304
rect 8347 2264 8392 2292
rect 8386 2252 8392 2264
rect 8444 2252 8450 2304
rect 8496 2292 8524 2332
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 9858 2360 9864 2372
rect 8720 2332 9864 2360
rect 8720 2320 8726 2332
rect 9858 2320 9864 2332
rect 9916 2360 9922 2372
rect 9953 2363 10011 2369
rect 9953 2360 9965 2363
rect 9916 2332 9965 2360
rect 9916 2320 9922 2332
rect 9953 2329 9965 2332
rect 9999 2329 10011 2363
rect 12406 2360 12434 2536
rect 13648 2536 15393 2564
rect 13648 2508 13676 2536
rect 15381 2533 15393 2536
rect 15427 2533 15439 2567
rect 15381 2527 15439 2533
rect 15470 2524 15476 2576
rect 15528 2564 15534 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 15528 2536 16865 2564
rect 15528 2524 15534 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 13078 2496 13084 2508
rect 13039 2468 13084 2496
rect 13078 2456 13084 2468
rect 13136 2456 13142 2508
rect 13173 2499 13231 2505
rect 13173 2465 13185 2499
rect 13219 2496 13231 2499
rect 13354 2496 13360 2508
rect 13219 2468 13360 2496
rect 13219 2465 13231 2468
rect 13173 2459 13231 2465
rect 13354 2456 13360 2468
rect 13412 2456 13418 2508
rect 13630 2456 13636 2508
rect 13688 2456 13694 2508
rect 15010 2496 15016 2508
rect 13924 2468 15016 2496
rect 13265 2431 13323 2437
rect 13265 2397 13277 2431
rect 13311 2428 13323 2431
rect 13924 2428 13952 2468
rect 15010 2456 15016 2468
rect 15068 2456 15074 2508
rect 15120 2468 15884 2496
rect 14090 2428 14096 2440
rect 13311 2400 13952 2428
rect 14051 2400 14096 2428
rect 13311 2397 13323 2400
rect 13265 2391 13323 2397
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 14642 2428 14648 2440
rect 14603 2400 14648 2428
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15120 2428 15148 2468
rect 14976 2400 15148 2428
rect 14976 2388 14982 2400
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15749 2431 15807 2437
rect 15252 2400 15297 2428
rect 15252 2388 15258 2400
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 15856 2428 15884 2468
rect 16298 2456 16304 2508
rect 16356 2496 16362 2508
rect 16356 2468 17816 2496
rect 16356 2456 16362 2468
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 15856 2400 16681 2428
rect 15749 2391 15807 2397
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 17218 2428 17224 2440
rect 17179 2400 17224 2428
rect 16669 2391 16727 2397
rect 15764 2360 15792 2391
rect 17218 2388 17224 2400
rect 17276 2388 17282 2440
rect 17788 2437 17816 2468
rect 17773 2431 17831 2437
rect 17773 2397 17785 2431
rect 17819 2397 17831 2431
rect 17880 2428 17908 2604
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 18012 2604 20545 2632
rect 18012 2592 18018 2604
rect 20533 2601 20545 2604
rect 20579 2601 20591 2635
rect 20533 2595 20591 2601
rect 18138 2456 18144 2508
rect 18196 2496 18202 2508
rect 18196 2468 19288 2496
rect 18196 2456 18202 2468
rect 19260 2437 19288 2468
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 17880 2400 18337 2428
rect 17773 2391 17831 2397
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19794 2428 19800 2440
rect 19755 2400 19800 2428
rect 19245 2391 19303 2397
rect 19794 2388 19800 2400
rect 19852 2388 19858 2440
rect 20346 2428 20352 2440
rect 20307 2400 20352 2428
rect 20346 2388 20352 2400
rect 20404 2388 20410 2440
rect 20898 2428 20904 2440
rect 20859 2400 20904 2428
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 9953 2323 10011 2329
rect 10152 2332 12296 2360
rect 12406 2332 15792 2360
rect 8846 2292 8852 2304
rect 8496 2264 8852 2292
rect 8846 2252 8852 2264
rect 8904 2252 8910 2304
rect 8938 2252 8944 2304
rect 8996 2292 9002 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 8996 2264 9321 2292
rect 8996 2252 9002 2264
rect 9309 2261 9321 2264
rect 9355 2292 9367 2295
rect 10152 2292 10180 2332
rect 9355 2264 10180 2292
rect 11609 2295 11667 2301
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 11609 2261 11621 2295
rect 11655 2292 11667 2295
rect 11790 2292 11796 2304
rect 11655 2264 11796 2292
rect 11655 2261 11667 2264
rect 11609 2255 11667 2261
rect 11790 2252 11796 2264
rect 11848 2252 11854 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 12268 2301 12296 2332
rect 16206 2320 16212 2372
rect 16264 2360 16270 2372
rect 16264 2332 18000 2360
rect 16264 2320 16270 2332
rect 12161 2295 12219 2301
rect 12161 2292 12173 2295
rect 11940 2264 12173 2292
rect 11940 2252 11946 2264
rect 12161 2261 12173 2264
rect 12207 2261 12219 2295
rect 12161 2255 12219 2261
rect 12253 2295 12311 2301
rect 12253 2261 12265 2295
rect 12299 2261 12311 2295
rect 12618 2292 12624 2304
rect 12579 2264 12624 2292
rect 12253 2255 12311 2261
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 13906 2252 13912 2304
rect 13964 2292 13970 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13964 2264 14289 2292
rect 13964 2252 13970 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14826 2292 14832 2304
rect 14787 2264 14832 2292
rect 14277 2255 14335 2261
rect 14826 2252 14832 2264
rect 14884 2252 14890 2304
rect 15838 2252 15844 2304
rect 15896 2292 15902 2304
rect 17972 2301 18000 2332
rect 18046 2320 18052 2372
rect 18104 2360 18110 2372
rect 18104 2332 21128 2360
rect 18104 2320 18110 2332
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 15896 2264 17417 2292
rect 15896 2252 15902 2264
rect 17405 2261 17417 2264
rect 17451 2261 17463 2295
rect 17405 2255 17463 2261
rect 17957 2295 18015 2301
rect 17957 2261 17969 2295
rect 18003 2261 18015 2295
rect 18506 2292 18512 2304
rect 18467 2264 18512 2292
rect 17957 2255 18015 2261
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 19426 2292 19432 2304
rect 19387 2264 19432 2292
rect 19426 2252 19432 2264
rect 19484 2252 19490 2304
rect 19978 2292 19984 2304
rect 19939 2264 19984 2292
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 21100 2301 21128 2332
rect 21085 2295 21143 2301
rect 21085 2261 21097 2295
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 7190 2088 7196 2100
rect 4028 2060 7196 2088
rect 4028 2048 4034 2060
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 11054 2088 11060 2100
rect 8628 2060 11060 2088
rect 8628 2048 8634 2060
rect 11054 2048 11060 2060
rect 11112 2088 11118 2100
rect 12066 2088 12072 2100
rect 11112 2060 12072 2088
rect 11112 2048 11118 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 14642 2088 14648 2100
rect 12176 2060 14648 2088
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 7616 1992 8524 2020
rect 7616 1980 7622 1992
rect 842 1912 848 1964
rect 900 1952 906 1964
rect 8386 1952 8392 1964
rect 900 1924 8392 1952
rect 900 1912 906 1924
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 8496 1952 8524 1992
rect 9306 1980 9312 2032
rect 9364 2020 9370 2032
rect 11882 2020 11888 2032
rect 9364 1992 11888 2020
rect 9364 1980 9370 1992
rect 11882 1980 11888 1992
rect 11940 1980 11946 2032
rect 12176 1952 12204 2060
rect 14642 2048 14648 2060
rect 14700 2048 14706 2100
rect 17034 2048 17040 2100
rect 17092 2088 17098 2100
rect 19426 2088 19432 2100
rect 17092 2060 19432 2088
rect 17092 2048 17098 2060
rect 19426 2048 19432 2060
rect 19484 2048 19490 2100
rect 14090 2020 14096 2032
rect 8496 1924 12204 1952
rect 12406 1992 14096 2020
rect 2958 1844 2964 1896
rect 3016 1884 3022 1896
rect 6546 1884 6552 1896
rect 3016 1856 6552 1884
rect 3016 1844 3022 1856
rect 6546 1844 6552 1856
rect 6604 1844 6610 1896
rect 7282 1844 7288 1896
rect 7340 1884 7346 1896
rect 12406 1884 12434 1992
rect 14090 1980 14096 1992
rect 14148 1980 14154 2032
rect 17310 1980 17316 2032
rect 17368 2020 17374 2032
rect 19978 2020 19984 2032
rect 17368 1992 19984 2020
rect 17368 1980 17374 1992
rect 19978 1980 19984 1992
rect 20036 1980 20042 2032
rect 12894 1912 12900 1964
rect 12952 1952 12958 1964
rect 14826 1952 14832 1964
rect 12952 1924 14832 1952
rect 12952 1912 12958 1924
rect 14826 1912 14832 1924
rect 14884 1912 14890 1964
rect 17402 1912 17408 1964
rect 17460 1952 17466 1964
rect 19794 1952 19800 1964
rect 17460 1924 19800 1952
rect 17460 1912 17466 1924
rect 19794 1912 19800 1924
rect 19852 1912 19858 1964
rect 7340 1856 12434 1884
rect 7340 1844 7346 1856
rect 13814 1844 13820 1896
rect 13872 1884 13878 1896
rect 14918 1884 14924 1896
rect 13872 1856 14924 1884
rect 13872 1844 13878 1856
rect 14918 1844 14924 1856
rect 14976 1844 14982 1896
rect 17586 1844 17592 1896
rect 17644 1884 17650 1896
rect 20346 1884 20352 1896
rect 17644 1856 20352 1884
rect 17644 1844 17650 1856
rect 20346 1844 20352 1856
rect 20404 1844 20410 1896
rect 10502 1776 10508 1828
rect 10560 1816 10566 1828
rect 17218 1816 17224 1828
rect 10560 1788 17224 1816
rect 10560 1776 10566 1788
rect 17218 1776 17224 1788
rect 17276 1776 17282 1828
rect 7834 1708 7840 1760
rect 7892 1748 7898 1760
rect 15194 1748 15200 1760
rect 7892 1720 15200 1748
rect 7892 1708 7898 1720
rect 15194 1708 15200 1720
rect 15252 1708 15258 1760
rect 16574 1708 16580 1760
rect 16632 1748 16638 1760
rect 18506 1748 18512 1760
rect 16632 1720 18512 1748
rect 16632 1708 16638 1720
rect 18506 1708 18512 1720
rect 18564 1708 18570 1760
rect 8846 1640 8852 1692
rect 8904 1680 8910 1692
rect 11146 1680 11152 1692
rect 8904 1652 11152 1680
rect 8904 1640 8910 1652
rect 11146 1640 11152 1652
rect 11204 1640 11210 1692
rect 14550 1640 14556 1692
rect 14608 1680 14614 1692
rect 18230 1680 18236 1692
rect 14608 1652 18236 1680
rect 14608 1640 14614 1652
rect 18230 1640 18236 1652
rect 18288 1640 18294 1692
rect 9674 1572 9680 1624
rect 9732 1612 9738 1624
rect 11238 1612 11244 1624
rect 9732 1584 11244 1612
rect 9732 1572 9738 1584
rect 11238 1572 11244 1584
rect 11296 1572 11302 1624
rect 12618 1572 12624 1624
rect 12676 1612 12682 1624
rect 16390 1612 16396 1624
rect 12676 1584 16396 1612
rect 12676 1572 12682 1584
rect 16390 1572 16396 1584
rect 16448 1572 16454 1624
rect 9858 1504 9864 1556
rect 9916 1544 9922 1556
rect 10686 1544 10692 1556
rect 9916 1516 10692 1544
rect 9916 1504 9922 1516
rect 10686 1504 10692 1516
rect 10744 1504 10750 1556
rect 14458 1504 14464 1556
rect 14516 1544 14522 1556
rect 17954 1544 17960 1556
rect 14516 1516 17960 1544
rect 14516 1504 14522 1516
rect 17954 1504 17960 1516
rect 18012 1504 18018 1556
rect 12526 1368 12532 1420
rect 12584 1408 12590 1420
rect 13906 1408 13912 1420
rect 12584 1380 13912 1408
rect 12584 1368 12590 1380
rect 13906 1368 13912 1380
rect 13964 1368 13970 1420
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 2044 20587 2096 20596
rect 2044 20553 2053 20587
rect 2053 20553 2087 20587
rect 2087 20553 2096 20587
rect 2044 20544 2096 20553
rect 17224 20544 17276 20596
rect 20168 20587 20220 20596
rect 20168 20553 20177 20587
rect 20177 20553 20211 20587
rect 20211 20553 20220 20587
rect 20168 20544 20220 20553
rect 21180 20476 21232 20528
rect 2136 20408 2188 20460
rect 2964 20451 3016 20460
rect 2964 20417 2973 20451
rect 2973 20417 3007 20451
rect 3007 20417 3016 20451
rect 2964 20408 3016 20417
rect 5724 20408 5776 20460
rect 16856 20451 16908 20460
rect 16856 20417 16865 20451
rect 16865 20417 16899 20451
rect 16899 20417 16908 20451
rect 16856 20408 16908 20417
rect 17776 20451 17828 20460
rect 17776 20417 17785 20451
rect 17785 20417 17819 20451
rect 17819 20417 17828 20451
rect 17776 20408 17828 20417
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 19524 20451 19576 20460
rect 19524 20417 19533 20451
rect 19533 20417 19567 20451
rect 19567 20417 19576 20451
rect 19524 20408 19576 20417
rect 20536 20451 20588 20460
rect 4068 20340 4120 20392
rect 4528 20383 4580 20392
rect 4528 20349 4537 20383
rect 4537 20349 4571 20383
rect 4571 20349 4580 20383
rect 4528 20340 4580 20349
rect 7840 20383 7892 20392
rect 7840 20349 7849 20383
rect 7849 20349 7883 20383
rect 7883 20349 7892 20383
rect 7840 20340 7892 20349
rect 14648 20272 14700 20324
rect 1492 20247 1544 20256
rect 1492 20213 1501 20247
rect 1501 20213 1535 20247
rect 1535 20213 1544 20247
rect 1492 20204 1544 20213
rect 3148 20247 3200 20256
rect 3148 20213 3157 20247
rect 3157 20213 3191 20247
rect 3191 20213 3200 20247
rect 3148 20204 3200 20213
rect 12532 20204 12584 20256
rect 12992 20204 13044 20256
rect 16396 20272 16448 20324
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 16488 20204 16540 20256
rect 17684 20204 17736 20256
rect 20444 20204 20496 20256
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 21272 20247 21324 20256
rect 21272 20213 21281 20247
rect 21281 20213 21315 20247
rect 21315 20213 21324 20247
rect 21272 20204 21324 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1952 20000 2004 20052
rect 12900 19932 12952 19984
rect 15016 19932 15068 19984
rect 8484 19864 8536 19916
rect 10508 19907 10560 19916
rect 10508 19873 10517 19907
rect 10517 19873 10551 19907
rect 10551 19873 10560 19907
rect 10508 19864 10560 19873
rect 11244 19864 11296 19916
rect 11796 19907 11848 19916
rect 11796 19873 11805 19907
rect 11805 19873 11839 19907
rect 11839 19873 11848 19907
rect 11796 19864 11848 19873
rect 14740 19907 14792 19916
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 4712 19796 4764 19848
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 9864 19796 9916 19848
rect 14740 19873 14749 19907
rect 14749 19873 14783 19907
rect 14783 19873 14792 19907
rect 14740 19864 14792 19873
rect 19524 20000 19576 20052
rect 21088 20000 21140 20052
rect 15200 19932 15252 19984
rect 16212 19932 16264 19984
rect 20536 19932 20588 19984
rect 20628 19932 20680 19984
rect 12532 19839 12584 19848
rect 12532 19805 12541 19839
rect 12541 19805 12575 19839
rect 12575 19805 12584 19839
rect 12532 19796 12584 19805
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 4528 19771 4580 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 4528 19737 4537 19771
rect 4537 19737 4571 19771
rect 4571 19737 4580 19771
rect 4528 19728 4580 19737
rect 3884 19703 3936 19712
rect 3884 19669 3893 19703
rect 3893 19669 3927 19703
rect 3927 19669 3936 19703
rect 3884 19660 3936 19669
rect 4252 19703 4304 19712
rect 4252 19669 4261 19703
rect 4261 19669 4295 19703
rect 4295 19669 4304 19703
rect 4252 19660 4304 19669
rect 4896 19703 4948 19712
rect 4896 19669 4905 19703
rect 4905 19669 4939 19703
rect 4939 19669 4948 19703
rect 4896 19660 4948 19669
rect 5448 19660 5500 19712
rect 7932 19660 7984 19712
rect 10416 19703 10468 19712
rect 10416 19669 10425 19703
rect 10425 19669 10459 19703
rect 10459 19669 10468 19703
rect 10416 19660 10468 19669
rect 11244 19660 11296 19712
rect 11704 19703 11756 19712
rect 11704 19669 11713 19703
rect 11713 19669 11747 19703
rect 11747 19669 11756 19703
rect 11704 19660 11756 19669
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 13176 19660 13228 19669
rect 14832 19796 14884 19848
rect 15936 19796 15988 19848
rect 17316 19907 17368 19916
rect 17316 19873 17325 19907
rect 17325 19873 17359 19907
rect 17359 19873 17368 19907
rect 17316 19864 17368 19873
rect 17776 19864 17828 19916
rect 18880 19864 18932 19916
rect 14556 19703 14608 19712
rect 14556 19669 14565 19703
rect 14565 19669 14599 19703
rect 14599 19669 14608 19703
rect 14556 19660 14608 19669
rect 15936 19660 15988 19712
rect 16212 19728 16264 19780
rect 17868 19728 17920 19780
rect 16488 19703 16540 19712
rect 16488 19669 16497 19703
rect 16497 19669 16531 19703
rect 16531 19669 16540 19703
rect 16488 19660 16540 19669
rect 16948 19660 17000 19712
rect 17500 19703 17552 19712
rect 17500 19669 17509 19703
rect 17509 19669 17543 19703
rect 17543 19669 17552 19703
rect 17500 19660 17552 19669
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18236 19703 18288 19712
rect 18236 19669 18245 19703
rect 18245 19669 18279 19703
rect 18279 19669 18288 19703
rect 18236 19660 18288 19669
rect 20536 19839 20588 19848
rect 20536 19805 20545 19839
rect 20545 19805 20579 19839
rect 20579 19805 20588 19839
rect 20536 19796 20588 19805
rect 21364 19660 21416 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2228 19456 2280 19508
rect 3700 19456 3752 19508
rect 4712 19499 4764 19508
rect 2136 19388 2188 19440
rect 1952 19320 2004 19372
rect 2228 19363 2280 19372
rect 2228 19329 2237 19363
rect 2237 19329 2271 19363
rect 2271 19329 2280 19363
rect 2228 19320 2280 19329
rect 1216 19184 1268 19236
rect 2044 19227 2096 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 2044 19193 2053 19227
rect 2053 19193 2087 19227
rect 2087 19193 2096 19227
rect 2044 19184 2096 19193
rect 2688 19363 2740 19372
rect 2688 19329 2697 19363
rect 2697 19329 2731 19363
rect 2731 19329 2740 19363
rect 2688 19320 2740 19329
rect 3516 19320 3568 19372
rect 4712 19465 4721 19499
rect 4721 19465 4755 19499
rect 4755 19465 4764 19499
rect 4712 19456 4764 19465
rect 5172 19499 5224 19508
rect 5172 19465 5181 19499
rect 5181 19465 5215 19499
rect 5215 19465 5224 19499
rect 5172 19456 5224 19465
rect 7564 19499 7616 19508
rect 7564 19465 7573 19499
rect 7573 19465 7607 19499
rect 7607 19465 7616 19499
rect 7564 19456 7616 19465
rect 7932 19499 7984 19508
rect 7932 19465 7941 19499
rect 7941 19465 7975 19499
rect 7975 19465 7984 19499
rect 7932 19456 7984 19465
rect 10416 19499 10468 19508
rect 10416 19465 10425 19499
rect 10425 19465 10459 19499
rect 10459 19465 10468 19499
rect 10416 19456 10468 19465
rect 11704 19456 11756 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 14832 19499 14884 19508
rect 14832 19465 14841 19499
rect 14841 19465 14875 19499
rect 14875 19465 14884 19499
rect 14832 19456 14884 19465
rect 17592 19456 17644 19508
rect 18236 19456 18288 19508
rect 5264 19388 5316 19440
rect 13176 19388 13228 19440
rect 17684 19388 17736 19440
rect 17868 19388 17920 19440
rect 19708 19456 19760 19508
rect 20536 19456 20588 19508
rect 20628 19456 20680 19508
rect 5080 19363 5132 19372
rect 4160 19252 4212 19304
rect 5080 19329 5089 19363
rect 5089 19329 5123 19363
rect 5123 19329 5132 19363
rect 5080 19320 5132 19329
rect 4988 19252 5040 19304
rect 8576 19320 8628 19372
rect 14464 19363 14516 19372
rect 14464 19329 14473 19363
rect 14473 19329 14507 19363
rect 14507 19329 14516 19363
rect 14464 19320 14516 19329
rect 18696 19363 18748 19372
rect 5356 19252 5408 19304
rect 8024 19295 8076 19304
rect 6368 19184 6420 19236
rect 8024 19261 8033 19295
rect 8033 19261 8067 19295
rect 8067 19261 8076 19295
rect 8024 19252 8076 19261
rect 9496 19252 9548 19304
rect 9864 19295 9916 19304
rect 9864 19261 9873 19295
rect 9873 19261 9907 19295
rect 9907 19261 9916 19295
rect 9864 19252 9916 19261
rect 12348 19295 12400 19304
rect 12348 19261 12357 19295
rect 12357 19261 12391 19295
rect 12391 19261 12400 19295
rect 12348 19252 12400 19261
rect 15476 19252 15528 19304
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18696 19329 18705 19363
rect 18705 19329 18739 19363
rect 18739 19329 18748 19363
rect 18696 19320 18748 19329
rect 20076 19363 20128 19372
rect 15844 19184 15896 19236
rect 16396 19184 16448 19236
rect 17224 19184 17276 19236
rect 17776 19184 17828 19236
rect 18236 19252 18288 19304
rect 20076 19329 20085 19363
rect 20085 19329 20119 19363
rect 20119 19329 20128 19363
rect 20076 19320 20128 19329
rect 20904 19320 20956 19372
rect 3516 19159 3568 19168
rect 3516 19125 3525 19159
rect 3525 19125 3559 19159
rect 3559 19125 3568 19159
rect 3516 19116 3568 19125
rect 4068 19116 4120 19168
rect 4160 19116 4212 19168
rect 4712 19116 4764 19168
rect 5356 19116 5408 19168
rect 5724 19159 5776 19168
rect 5724 19125 5733 19159
rect 5733 19125 5767 19159
rect 5767 19125 5776 19159
rect 5724 19116 5776 19125
rect 6552 19116 6604 19168
rect 11888 19116 11940 19168
rect 12992 19116 13044 19168
rect 13084 19116 13136 19168
rect 15660 19116 15712 19168
rect 17040 19159 17092 19168
rect 17040 19125 17049 19159
rect 17049 19125 17083 19159
rect 17083 19125 17092 19159
rect 17040 19116 17092 19125
rect 17868 19116 17920 19168
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 21272 19159 21324 19168
rect 21272 19125 21281 19159
rect 21281 19125 21315 19159
rect 21315 19125 21324 19159
rect 21272 19116 21324 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 2228 18912 2280 18964
rect 2504 18912 2556 18964
rect 2044 18708 2096 18760
rect 4160 18776 4212 18828
rect 5080 18912 5132 18964
rect 7196 18912 7248 18964
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1676 18572 1728 18624
rect 6000 18844 6052 18896
rect 6368 18844 6420 18896
rect 11888 18912 11940 18964
rect 14464 18912 14516 18964
rect 14648 18912 14700 18964
rect 16304 18912 16356 18964
rect 16948 18912 17000 18964
rect 17960 18912 18012 18964
rect 18144 18912 18196 18964
rect 18696 18912 18748 18964
rect 6552 18776 6604 18828
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 10048 18776 10100 18828
rect 12072 18844 12124 18896
rect 18880 18844 18932 18896
rect 20812 18844 20864 18896
rect 11980 18819 12032 18828
rect 11980 18785 11989 18819
rect 11989 18785 12023 18819
rect 12023 18785 12032 18819
rect 11980 18776 12032 18785
rect 8116 18708 8168 18760
rect 12348 18708 12400 18760
rect 14372 18776 14424 18828
rect 16120 18819 16172 18828
rect 16120 18785 16129 18819
rect 16129 18785 16163 18819
rect 16163 18785 16172 18819
rect 16120 18776 16172 18785
rect 17224 18819 17276 18828
rect 16304 18708 16356 18760
rect 16948 18708 17000 18760
rect 17224 18785 17233 18819
rect 17233 18785 17267 18819
rect 17267 18785 17276 18819
rect 17224 18776 17276 18785
rect 18696 18776 18748 18828
rect 20260 18776 20312 18828
rect 19984 18708 20036 18760
rect 3884 18572 3936 18624
rect 4528 18572 4580 18624
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 7656 18572 7708 18624
rect 8300 18640 8352 18692
rect 14648 18640 14700 18692
rect 15752 18640 15804 18692
rect 16212 18640 16264 18692
rect 17224 18640 17276 18692
rect 19432 18640 19484 18692
rect 9220 18572 9272 18624
rect 9772 18572 9824 18624
rect 11704 18572 11756 18624
rect 12716 18615 12768 18624
rect 12716 18581 12725 18615
rect 12725 18581 12759 18615
rect 12759 18581 12768 18615
rect 12716 18572 12768 18581
rect 12808 18615 12860 18624
rect 12808 18581 12817 18615
rect 12817 18581 12851 18615
rect 12851 18581 12860 18615
rect 13176 18615 13228 18624
rect 12808 18572 12860 18581
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 15016 18615 15068 18624
rect 15016 18581 15025 18615
rect 15025 18581 15059 18615
rect 15059 18581 15068 18615
rect 15016 18572 15068 18581
rect 15200 18572 15252 18624
rect 15660 18572 15712 18624
rect 16028 18615 16080 18624
rect 16028 18581 16037 18615
rect 16037 18581 16071 18615
rect 16071 18581 16080 18615
rect 16948 18615 17000 18624
rect 16028 18572 16080 18581
rect 16948 18581 16957 18615
rect 16957 18581 16991 18615
rect 16991 18581 17000 18615
rect 16948 18572 17000 18581
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 19616 18615 19668 18624
rect 19616 18581 19625 18615
rect 19625 18581 19659 18615
rect 19659 18581 19668 18615
rect 20260 18615 20312 18624
rect 19616 18572 19668 18581
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 20628 18572 20680 18624
rect 21088 18572 21140 18624
rect 21364 18572 21416 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 1952 18411 2004 18420
rect 1952 18377 1961 18411
rect 1961 18377 1995 18411
rect 1995 18377 2004 18411
rect 1952 18368 2004 18377
rect 5264 18411 5316 18420
rect 5264 18377 5273 18411
rect 5273 18377 5307 18411
rect 5307 18377 5316 18411
rect 5264 18368 5316 18377
rect 5448 18368 5500 18420
rect 1032 18300 1084 18352
rect 4804 18300 4856 18352
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 2504 18232 2556 18284
rect 3056 18232 3108 18284
rect 3240 18275 3292 18284
rect 3240 18241 3249 18275
rect 3249 18241 3283 18275
rect 3283 18241 3292 18275
rect 3240 18232 3292 18241
rect 4068 18232 4120 18284
rect 2872 18164 2924 18216
rect 3976 18207 4028 18216
rect 1584 18096 1636 18148
rect 3976 18173 3985 18207
rect 3985 18173 4019 18207
rect 4019 18173 4028 18207
rect 3976 18164 4028 18173
rect 4160 18207 4212 18216
rect 4160 18173 4169 18207
rect 4169 18173 4203 18207
rect 4203 18173 4212 18207
rect 4160 18164 4212 18173
rect 6828 18232 6880 18284
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2136 18028 2188 18080
rect 3424 18096 3476 18148
rect 4068 18096 4120 18148
rect 7012 18207 7064 18216
rect 4620 18071 4672 18080
rect 4620 18037 4629 18071
rect 4629 18037 4663 18071
rect 4663 18037 4672 18071
rect 4620 18028 4672 18037
rect 7012 18173 7021 18207
rect 7021 18173 7055 18207
rect 7055 18173 7064 18207
rect 7012 18164 7064 18173
rect 8024 18368 8076 18420
rect 8116 18368 8168 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 12072 18368 12124 18420
rect 12808 18368 12860 18420
rect 13636 18368 13688 18420
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15660 18411 15712 18420
rect 15292 18368 15344 18377
rect 15660 18377 15669 18411
rect 15669 18377 15703 18411
rect 15703 18377 15712 18411
rect 15660 18368 15712 18377
rect 16856 18368 16908 18420
rect 17684 18368 17736 18420
rect 17868 18368 17920 18420
rect 7656 18300 7708 18352
rect 8300 18275 8352 18284
rect 8300 18241 8309 18275
rect 8309 18241 8343 18275
rect 8343 18241 8352 18275
rect 8300 18232 8352 18241
rect 8668 18232 8720 18284
rect 7656 18164 7708 18216
rect 8484 18207 8536 18216
rect 8484 18173 8493 18207
rect 8493 18173 8527 18207
rect 8527 18173 8536 18207
rect 9404 18207 9456 18216
rect 8484 18164 8536 18173
rect 9404 18173 9413 18207
rect 9413 18173 9447 18207
rect 9447 18173 9456 18207
rect 9404 18164 9456 18173
rect 9956 18275 10008 18284
rect 9956 18241 9965 18275
rect 9965 18241 9999 18275
rect 9999 18241 10008 18275
rect 9956 18232 10008 18241
rect 6000 18096 6052 18148
rect 8116 18096 8168 18148
rect 8208 18096 8260 18148
rect 10968 18164 11020 18216
rect 10784 18096 10836 18148
rect 11888 18207 11940 18216
rect 11888 18173 11897 18207
rect 11897 18173 11931 18207
rect 11931 18173 11940 18207
rect 11888 18164 11940 18173
rect 12532 18164 12584 18216
rect 13176 18300 13228 18352
rect 17224 18300 17276 18352
rect 17408 18300 17460 18352
rect 12992 18232 13044 18284
rect 13636 18275 13688 18284
rect 13636 18241 13645 18275
rect 13645 18241 13679 18275
rect 13679 18241 13688 18275
rect 13636 18232 13688 18241
rect 16856 18232 16908 18284
rect 6276 18028 6328 18080
rect 6552 18028 6604 18080
rect 8300 18028 8352 18080
rect 9312 18028 9364 18080
rect 12992 18028 13044 18080
rect 17040 18164 17092 18216
rect 17592 18164 17644 18216
rect 18604 18300 18656 18352
rect 18144 18275 18196 18284
rect 18144 18241 18153 18275
rect 18153 18241 18187 18275
rect 18187 18241 18196 18275
rect 18144 18232 18196 18241
rect 18052 18207 18104 18216
rect 18052 18173 18061 18207
rect 18061 18173 18095 18207
rect 18095 18173 18104 18207
rect 20260 18232 20312 18284
rect 20444 18232 20496 18284
rect 18052 18164 18104 18173
rect 19064 18164 19116 18216
rect 13360 18028 13412 18080
rect 16212 18071 16264 18080
rect 16212 18037 16221 18071
rect 16221 18037 16255 18071
rect 16255 18037 16264 18071
rect 16212 18028 16264 18037
rect 16948 18028 17000 18080
rect 17132 18071 17184 18080
rect 17132 18037 17141 18071
rect 17141 18037 17175 18071
rect 17175 18037 17184 18071
rect 17132 18028 17184 18037
rect 18052 18028 18104 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 18972 18096 19024 18148
rect 20996 18096 21048 18148
rect 20720 18071 20772 18080
rect 20720 18037 20729 18071
rect 20729 18037 20763 18071
rect 20763 18037 20772 18071
rect 20720 18028 20772 18037
rect 21272 18071 21324 18080
rect 21272 18037 21281 18071
rect 21281 18037 21315 18071
rect 21315 18037 21324 18071
rect 21272 18028 21324 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 2044 17824 2096 17876
rect 3056 17824 3108 17876
rect 4068 17824 4120 17876
rect 5172 17824 5224 17876
rect 6276 17824 6328 17876
rect 7472 17799 7524 17808
rect 2136 17620 2188 17672
rect 2228 17663 2280 17672
rect 2228 17629 2237 17663
rect 2237 17629 2271 17663
rect 2271 17629 2280 17663
rect 3240 17688 3292 17740
rect 3976 17688 4028 17740
rect 5448 17688 5500 17740
rect 6276 17731 6328 17740
rect 6276 17697 6285 17731
rect 6285 17697 6319 17731
rect 6319 17697 6328 17731
rect 6276 17688 6328 17697
rect 6828 17688 6880 17740
rect 7472 17765 7481 17799
rect 7481 17765 7515 17799
rect 7515 17765 7524 17799
rect 7472 17756 7524 17765
rect 9404 17824 9456 17876
rect 9680 17824 9732 17876
rect 13084 17824 13136 17876
rect 17868 17824 17920 17876
rect 19064 17824 19116 17876
rect 20076 17824 20128 17876
rect 10876 17756 10928 17808
rect 15752 17756 15804 17808
rect 2228 17620 2280 17629
rect 4804 17620 4856 17672
rect 7656 17688 7708 17740
rect 8208 17688 8260 17740
rect 10232 17731 10284 17740
rect 10232 17697 10241 17731
rect 10241 17697 10275 17731
rect 10275 17697 10284 17731
rect 10232 17688 10284 17697
rect 15568 17731 15620 17740
rect 6736 17552 6788 17604
rect 7380 17620 7432 17672
rect 7748 17620 7800 17672
rect 9956 17620 10008 17672
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2044 17527 2096 17536
rect 2044 17493 2053 17527
rect 2053 17493 2087 17527
rect 2087 17493 2096 17527
rect 2044 17484 2096 17493
rect 4252 17527 4304 17536
rect 4252 17493 4261 17527
rect 4261 17493 4295 17527
rect 4295 17493 4304 17527
rect 4252 17484 4304 17493
rect 4988 17527 5040 17536
rect 4988 17493 4997 17527
rect 4997 17493 5031 17527
rect 5031 17493 5040 17527
rect 4988 17484 5040 17493
rect 5172 17484 5224 17536
rect 5908 17484 5960 17536
rect 6552 17484 6604 17536
rect 6920 17484 6972 17536
rect 7104 17527 7156 17536
rect 7104 17493 7113 17527
rect 7113 17493 7147 17527
rect 7147 17493 7156 17527
rect 9036 17552 9088 17604
rect 7104 17484 7156 17493
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 9772 17484 9824 17536
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10692 17527 10744 17536
rect 10048 17484 10100 17493
rect 10692 17493 10701 17527
rect 10701 17493 10735 17527
rect 10735 17493 10744 17527
rect 10692 17484 10744 17493
rect 11152 17527 11204 17536
rect 11152 17493 11161 17527
rect 11161 17493 11195 17527
rect 11195 17493 11204 17527
rect 11152 17484 11204 17493
rect 11520 17527 11572 17536
rect 11520 17493 11529 17527
rect 11529 17493 11563 17527
rect 11563 17493 11572 17527
rect 11520 17484 11572 17493
rect 12072 17484 12124 17536
rect 15568 17697 15577 17731
rect 15577 17697 15611 17731
rect 15611 17697 15620 17731
rect 15568 17688 15620 17697
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 20904 17756 20956 17808
rect 17868 17688 17920 17740
rect 19892 17731 19944 17740
rect 19892 17697 19901 17731
rect 19901 17697 19935 17731
rect 19935 17697 19944 17731
rect 19892 17688 19944 17697
rect 17960 17663 18012 17672
rect 13452 17484 13504 17536
rect 15108 17527 15160 17536
rect 15108 17493 15117 17527
rect 15117 17493 15151 17527
rect 15151 17493 15160 17527
rect 15108 17484 15160 17493
rect 15752 17527 15804 17536
rect 15752 17493 15761 17527
rect 15761 17493 15795 17527
rect 15795 17493 15804 17527
rect 15752 17484 15804 17493
rect 17960 17629 17969 17663
rect 17969 17629 18003 17663
rect 18003 17629 18012 17663
rect 17960 17620 18012 17629
rect 18052 17620 18104 17672
rect 20260 17620 20312 17672
rect 20904 17620 20956 17672
rect 21180 17620 21232 17672
rect 17592 17484 17644 17536
rect 17868 17484 17920 17536
rect 18236 17552 18288 17604
rect 20076 17552 20128 17604
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 19708 17527 19760 17536
rect 19708 17493 19717 17527
rect 19717 17493 19751 17527
rect 19751 17493 19760 17527
rect 19708 17484 19760 17493
rect 20444 17484 20496 17536
rect 20628 17527 20680 17536
rect 20628 17493 20637 17527
rect 20637 17493 20671 17527
rect 20671 17493 20680 17527
rect 20628 17484 20680 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 2228 17280 2280 17332
rect 3148 17280 3200 17332
rect 3976 17323 4028 17332
rect 3976 17289 3985 17323
rect 3985 17289 4019 17323
rect 4019 17289 4028 17323
rect 3976 17280 4028 17289
rect 4160 17280 4212 17332
rect 5172 17323 5224 17332
rect 5172 17289 5181 17323
rect 5181 17289 5215 17323
rect 5215 17289 5224 17323
rect 5172 17280 5224 17289
rect 7012 17280 7064 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 8484 17280 8536 17332
rect 8668 17280 8720 17332
rect 9404 17280 9456 17332
rect 10692 17323 10744 17332
rect 10692 17289 10701 17323
rect 10701 17289 10735 17323
rect 10735 17289 10744 17323
rect 10692 17280 10744 17289
rect 11152 17280 11204 17332
rect 15292 17280 15344 17332
rect 15568 17280 15620 17332
rect 17868 17280 17920 17332
rect 19984 17280 20036 17332
rect 20812 17323 20864 17332
rect 20812 17289 20821 17323
rect 20821 17289 20855 17323
rect 20855 17289 20864 17323
rect 20812 17280 20864 17289
rect 2964 17212 3016 17264
rect 4620 17212 4672 17264
rect 8760 17212 8812 17264
rect 18236 17212 18288 17264
rect 19616 17212 19668 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 2320 17144 2372 17196
rect 7012 17144 7064 17196
rect 9128 17144 9180 17196
rect 9680 17144 9732 17196
rect 11060 17144 11112 17196
rect 16948 17144 17000 17196
rect 18880 17187 18932 17196
rect 18880 17153 18889 17187
rect 18889 17153 18923 17187
rect 18923 17153 18932 17187
rect 18880 17144 18932 17153
rect 19524 17144 19576 17196
rect 2872 17076 2924 17128
rect 4068 17076 4120 17128
rect 6092 17076 6144 17128
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 2412 16983 2464 16992
rect 2412 16949 2421 16983
rect 2421 16949 2455 16983
rect 2455 16949 2464 16983
rect 2412 16940 2464 16949
rect 7104 17076 7156 17128
rect 7748 17076 7800 17128
rect 8300 17076 8352 17128
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 10416 17076 10468 17128
rect 11796 17119 11848 17128
rect 11796 17085 11805 17119
rect 11805 17085 11839 17119
rect 11839 17085 11848 17119
rect 11796 17076 11848 17085
rect 11888 17119 11940 17128
rect 11888 17085 11897 17119
rect 11897 17085 11931 17119
rect 11931 17085 11940 17119
rect 11888 17076 11940 17085
rect 12532 17076 12584 17128
rect 15200 17076 15252 17128
rect 16120 17076 16172 17128
rect 7840 17008 7892 17060
rect 3056 16940 3108 16992
rect 5816 16983 5868 16992
rect 5816 16949 5825 16983
rect 5825 16949 5859 16983
rect 5859 16949 5868 16983
rect 5816 16940 5868 16949
rect 7288 16983 7340 16992
rect 7288 16949 7297 16983
rect 7297 16949 7331 16983
rect 7331 16949 7340 16983
rect 7288 16940 7340 16949
rect 7380 16940 7432 16992
rect 8576 16940 8628 16992
rect 8944 17008 8996 17060
rect 10140 17008 10192 17060
rect 21180 17076 21232 17128
rect 20904 17008 20956 17060
rect 10784 16940 10836 16992
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 12992 16940 13044 16992
rect 17500 16983 17552 16992
rect 17500 16949 17509 16983
rect 17509 16949 17543 16983
rect 17543 16949 17552 16983
rect 17500 16940 17552 16949
rect 18604 16983 18656 16992
rect 18604 16949 18613 16983
rect 18613 16949 18647 16983
rect 18647 16949 18656 16983
rect 18604 16940 18656 16949
rect 20168 16940 20220 16992
rect 20352 16983 20404 16992
rect 20352 16949 20361 16983
rect 20361 16949 20395 16983
rect 20395 16949 20404 16983
rect 20352 16940 20404 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 2136 16736 2188 16788
rect 8484 16736 8536 16788
rect 4344 16668 4396 16720
rect 4436 16668 4488 16720
rect 6092 16668 6144 16720
rect 9956 16736 10008 16788
rect 8668 16668 8720 16720
rect 5264 16600 5316 16652
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5724 16600 5776 16652
rect 7380 16600 7432 16652
rect 9404 16600 9456 16652
rect 11980 16736 12032 16788
rect 15568 16736 15620 16788
rect 15752 16736 15804 16788
rect 19524 16779 19576 16788
rect 19524 16745 19533 16779
rect 19533 16745 19567 16779
rect 19567 16745 19576 16779
rect 19524 16736 19576 16745
rect 11152 16668 11204 16720
rect 2412 16532 2464 16584
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 3056 16532 3108 16584
rect 6644 16532 6696 16584
rect 9036 16532 9088 16584
rect 11704 16600 11756 16652
rect 12808 16643 12860 16652
rect 12808 16609 12817 16643
rect 12817 16609 12851 16643
rect 12851 16609 12860 16643
rect 12808 16600 12860 16609
rect 15108 16600 15160 16652
rect 16396 16600 16448 16652
rect 17500 16668 17552 16720
rect 17684 16668 17736 16720
rect 10692 16532 10744 16584
rect 12164 16532 12216 16584
rect 12992 16575 13044 16584
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 16948 16600 17000 16652
rect 21456 16668 21508 16720
rect 20444 16643 20496 16652
rect 20444 16609 20453 16643
rect 20453 16609 20487 16643
rect 20487 16609 20496 16643
rect 20444 16600 20496 16609
rect 20536 16643 20588 16652
rect 20536 16609 20545 16643
rect 20545 16609 20579 16643
rect 20579 16609 20588 16643
rect 20536 16600 20588 16609
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 18788 16532 18840 16584
rect 20352 16532 20404 16584
rect 20996 16532 21048 16584
rect 4160 16507 4212 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2044 16396 2096 16448
rect 2228 16396 2280 16448
rect 4160 16473 4169 16507
rect 4169 16473 4203 16507
rect 4203 16473 4212 16507
rect 4160 16464 4212 16473
rect 6460 16464 6512 16516
rect 4528 16439 4580 16448
rect 4528 16405 4537 16439
rect 4537 16405 4571 16439
rect 4571 16405 4580 16439
rect 4528 16396 4580 16405
rect 4896 16439 4948 16448
rect 4896 16405 4905 16439
rect 4905 16405 4939 16439
rect 4939 16405 4948 16439
rect 4896 16396 4948 16405
rect 5080 16396 5132 16448
rect 6644 16396 6696 16448
rect 7932 16396 7984 16448
rect 8116 16439 8168 16448
rect 8116 16405 8125 16439
rect 8125 16405 8159 16439
rect 8159 16405 8168 16439
rect 8116 16396 8168 16405
rect 8668 16396 8720 16448
rect 10416 16396 10468 16448
rect 11520 16396 11572 16448
rect 15292 16464 15344 16516
rect 16028 16464 16080 16516
rect 12532 16396 12584 16448
rect 13452 16396 13504 16448
rect 16396 16396 16448 16448
rect 18696 16396 18748 16448
rect 18880 16396 18932 16448
rect 20076 16396 20128 16448
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1676 16192 1728 16244
rect 2872 16192 2924 16244
rect 4712 16192 4764 16244
rect 4988 16192 5040 16244
rect 6552 16235 6604 16244
rect 6552 16201 6561 16235
rect 6561 16201 6595 16235
rect 6595 16201 6604 16235
rect 6552 16192 6604 16201
rect 6736 16192 6788 16244
rect 7932 16235 7984 16244
rect 7932 16201 7941 16235
rect 7941 16201 7975 16235
rect 7975 16201 7984 16235
rect 7932 16192 7984 16201
rect 8484 16192 8536 16244
rect 10692 16192 10744 16244
rect 15016 16192 15068 16244
rect 16396 16192 16448 16244
rect 17316 16192 17368 16244
rect 17592 16192 17644 16244
rect 18512 16192 18564 16244
rect 20720 16192 20772 16244
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2228 16099 2280 16108
rect 2228 16065 2237 16099
rect 2237 16065 2271 16099
rect 2271 16065 2280 16099
rect 2228 16056 2280 16065
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 5448 16099 5500 16108
rect 5448 16065 5457 16099
rect 5457 16065 5491 16099
rect 5491 16065 5500 16099
rect 5448 16056 5500 16065
rect 7748 16124 7800 16176
rect 10140 16124 10192 16176
rect 10416 16124 10468 16176
rect 7380 16056 7432 16108
rect 7472 16056 7524 16108
rect 4068 15988 4120 16040
rect 4528 16031 4580 16040
rect 4528 15997 4537 16031
rect 4537 15997 4571 16031
rect 4571 15997 4580 16031
rect 4528 15988 4580 15997
rect 4896 15988 4948 16040
rect 5356 15988 5408 16040
rect 7012 16031 7064 16040
rect 1400 15920 1452 15972
rect 2780 15920 2832 15972
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7564 15988 7616 16040
rect 8024 16031 8076 16040
rect 8024 15997 8033 16031
rect 8033 15997 8067 16031
rect 8067 15997 8076 16031
rect 8024 15988 8076 15997
rect 9680 16056 9732 16108
rect 11244 16056 11296 16108
rect 6736 15920 6788 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4068 15895 4120 15904
rect 4068 15861 4077 15895
rect 4077 15861 4111 15895
rect 4111 15861 4120 15895
rect 4068 15852 4120 15861
rect 4160 15852 4212 15904
rect 6920 15852 6972 15904
rect 7012 15852 7064 15904
rect 7748 15852 7800 15904
rect 8116 15852 8168 15904
rect 8484 15852 8536 15904
rect 9128 15895 9180 15904
rect 9128 15861 9137 15895
rect 9137 15861 9171 15895
rect 9171 15861 9180 15895
rect 9128 15852 9180 15861
rect 13176 15920 13228 15972
rect 10600 15852 10652 15904
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 10876 15852 10928 15904
rect 12072 15852 12124 15904
rect 12624 15852 12676 15904
rect 13636 16056 13688 16108
rect 17040 16124 17092 16176
rect 17316 16056 17368 16108
rect 18052 16056 18104 16108
rect 19984 16099 20036 16108
rect 19984 16065 19993 16099
rect 19993 16065 20027 16099
rect 20027 16065 20036 16099
rect 19984 16056 20036 16065
rect 20536 16099 20588 16108
rect 20536 16065 20545 16099
rect 20545 16065 20579 16099
rect 20579 16065 20588 16099
rect 20536 16056 20588 16065
rect 20904 16056 20956 16108
rect 15384 15988 15436 16040
rect 18880 16031 18932 16040
rect 18880 15997 18889 16031
rect 18889 15997 18923 16031
rect 18923 15997 18932 16031
rect 18880 15988 18932 15997
rect 13360 15920 13412 15972
rect 17684 15920 17736 15972
rect 20352 15920 20404 15972
rect 20720 15963 20772 15972
rect 20720 15929 20729 15963
rect 20729 15929 20763 15963
rect 20763 15929 20772 15963
rect 20720 15920 20772 15929
rect 15384 15852 15436 15904
rect 21364 15852 21416 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 4436 15691 4488 15700
rect 4436 15657 4445 15691
rect 4445 15657 4479 15691
rect 4479 15657 4488 15691
rect 4436 15648 4488 15657
rect 4712 15648 4764 15700
rect 848 15580 900 15632
rect 5448 15580 5500 15632
rect 3424 15512 3476 15564
rect 5080 15555 5132 15564
rect 5080 15521 5089 15555
rect 5089 15521 5123 15555
rect 5123 15521 5132 15555
rect 5080 15512 5132 15521
rect 1400 15444 1452 15496
rect 2596 15487 2648 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 1952 15351 2004 15360
rect 1952 15317 1961 15351
rect 1961 15317 1995 15351
rect 1995 15317 2004 15351
rect 1952 15308 2004 15317
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 5172 15444 5224 15496
rect 6828 15444 6880 15496
rect 7012 15444 7064 15496
rect 7472 15444 7524 15496
rect 8024 15648 8076 15700
rect 9128 15648 9180 15700
rect 10232 15648 10284 15700
rect 8116 15580 8168 15632
rect 10416 15580 10468 15632
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 11980 15623 12032 15632
rect 11980 15589 11989 15623
rect 11989 15589 12023 15623
rect 12023 15589 12032 15623
rect 11980 15580 12032 15589
rect 12072 15580 12124 15632
rect 17224 15648 17276 15700
rect 17684 15648 17736 15700
rect 19708 15648 19760 15700
rect 20536 15648 20588 15700
rect 9128 15512 9180 15564
rect 12440 15512 12492 15564
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 10784 15444 10836 15496
rect 2688 15308 2740 15360
rect 3056 15308 3108 15360
rect 3792 15308 3844 15360
rect 6552 15351 6604 15360
rect 6552 15317 6561 15351
rect 6561 15317 6595 15351
rect 6595 15317 6604 15351
rect 6552 15308 6604 15317
rect 8484 15308 8536 15360
rect 9496 15419 9548 15428
rect 9496 15385 9530 15419
rect 9530 15385 9548 15419
rect 9496 15376 9548 15385
rect 10692 15376 10744 15428
rect 12716 15444 12768 15496
rect 12992 15444 13044 15496
rect 11244 15376 11296 15428
rect 13820 15376 13872 15428
rect 16580 15487 16632 15496
rect 16580 15453 16589 15487
rect 16589 15453 16623 15487
rect 16623 15453 16632 15487
rect 16580 15444 16632 15453
rect 17684 15487 17736 15496
rect 17684 15453 17693 15487
rect 17693 15453 17727 15487
rect 17727 15453 17736 15487
rect 17684 15444 17736 15453
rect 19524 15444 19576 15496
rect 11888 15308 11940 15360
rect 15200 15351 15252 15360
rect 15200 15317 15209 15351
rect 15209 15317 15243 15351
rect 15243 15317 15252 15351
rect 15200 15308 15252 15317
rect 16120 15308 16172 15360
rect 16764 15308 16816 15360
rect 19524 15308 19576 15360
rect 20352 15376 20404 15428
rect 20812 15308 20864 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 4252 15104 4304 15156
rect 5540 15104 5592 15156
rect 5908 15104 5960 15156
rect 6828 15104 6880 15156
rect 6920 15104 6972 15156
rect 9680 15104 9732 15156
rect 7196 15036 7248 15088
rect 7932 15036 7984 15088
rect 8668 15036 8720 15088
rect 10784 15104 10836 15156
rect 12808 15104 12860 15156
rect 13728 15104 13780 15156
rect 16948 15104 17000 15156
rect 19708 15104 19760 15156
rect 20536 15104 20588 15156
rect 11244 15036 11296 15088
rect 17684 15036 17736 15088
rect 2044 14968 2096 15020
rect 2688 15011 2740 15020
rect 2688 14977 2697 15011
rect 2697 14977 2731 15011
rect 2731 14977 2740 15011
rect 2688 14968 2740 14977
rect 4988 15011 5040 15020
rect 1676 14832 1728 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 2136 14807 2188 14816
rect 2136 14773 2145 14807
rect 2145 14773 2179 14807
rect 2179 14773 2188 14807
rect 2136 14764 2188 14773
rect 4988 14977 4997 15011
rect 4997 14977 5031 15011
rect 5031 14977 5040 15011
rect 4988 14968 5040 14977
rect 5908 14968 5960 15020
rect 7012 14968 7064 15020
rect 9220 14968 9272 15020
rect 9680 15011 9732 15020
rect 9680 14977 9689 15011
rect 9689 14977 9723 15011
rect 9723 14977 9732 15011
rect 9680 14968 9732 14977
rect 9772 14968 9824 15020
rect 10324 14968 10376 15020
rect 4896 14900 4948 14952
rect 5356 14900 5408 14952
rect 7840 14900 7892 14952
rect 3332 14832 3384 14884
rect 4436 14764 4488 14816
rect 4896 14764 4948 14816
rect 6552 14764 6604 14816
rect 7196 14764 7248 14816
rect 8668 14900 8720 14952
rect 11612 14900 11664 14952
rect 12992 14900 13044 14952
rect 10784 14832 10836 14884
rect 15936 14968 15988 15020
rect 17224 14968 17276 15020
rect 18696 14968 18748 15020
rect 20720 15036 20772 15088
rect 10048 14764 10100 14816
rect 11428 14764 11480 14816
rect 11980 14807 12032 14816
rect 11980 14773 11989 14807
rect 11989 14773 12023 14807
rect 12023 14773 12032 14807
rect 11980 14764 12032 14773
rect 12716 14807 12768 14816
rect 12716 14773 12725 14807
rect 12725 14773 12759 14807
rect 12759 14773 12768 14807
rect 12716 14764 12768 14773
rect 12992 14807 13044 14816
rect 12992 14773 13001 14807
rect 13001 14773 13035 14807
rect 13035 14773 13044 14807
rect 12992 14764 13044 14773
rect 13084 14764 13136 14816
rect 14740 14832 14792 14884
rect 15016 14832 15068 14884
rect 14924 14764 14976 14816
rect 16396 14832 16448 14884
rect 16028 14807 16080 14816
rect 16028 14773 16037 14807
rect 16037 14773 16071 14807
rect 16071 14773 16080 14807
rect 16028 14764 16080 14773
rect 19800 14900 19852 14952
rect 18696 14764 18748 14816
rect 19892 14764 19944 14816
rect 20996 14764 21048 14816
rect 21180 14764 21232 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 4988 14560 5040 14612
rect 6644 14603 6696 14612
rect 6644 14569 6653 14603
rect 6653 14569 6687 14603
rect 6687 14569 6696 14603
rect 6644 14560 6696 14569
rect 20 14492 72 14544
rect 1676 14492 1728 14544
rect 3240 14492 3292 14544
rect 3976 14492 4028 14544
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 3976 14356 4028 14408
rect 3148 14288 3200 14340
rect 5172 14492 5224 14544
rect 8392 14560 8444 14612
rect 8852 14560 8904 14612
rect 11520 14560 11572 14612
rect 11704 14560 11756 14612
rect 4160 14424 4212 14476
rect 5080 14424 5132 14476
rect 6644 14424 6696 14476
rect 9312 14492 9364 14544
rect 11796 14492 11848 14544
rect 12256 14492 12308 14544
rect 13820 14560 13872 14612
rect 16396 14560 16448 14612
rect 19708 14560 19760 14612
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 9680 14424 9732 14476
rect 10232 14467 10284 14476
rect 10232 14433 10241 14467
rect 10241 14433 10275 14467
rect 10275 14433 10284 14467
rect 10232 14424 10284 14433
rect 4252 14399 4304 14408
rect 4252 14365 4261 14399
rect 4261 14365 4295 14399
rect 4295 14365 4304 14399
rect 4252 14356 4304 14365
rect 5540 14356 5592 14408
rect 7288 14399 7340 14408
rect 7288 14365 7297 14399
rect 7297 14365 7331 14399
rect 7331 14365 7340 14399
rect 7288 14356 7340 14365
rect 10508 14399 10560 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2136 14263 2188 14272
rect 2136 14229 2145 14263
rect 2145 14229 2179 14263
rect 2179 14229 2188 14263
rect 2136 14220 2188 14229
rect 2504 14220 2556 14272
rect 3424 14220 3476 14272
rect 5080 14288 5132 14340
rect 6644 14220 6696 14272
rect 6736 14220 6788 14272
rect 10048 14288 10100 14340
rect 10508 14365 10542 14399
rect 10542 14365 10560 14399
rect 10508 14356 10560 14365
rect 14464 14424 14516 14476
rect 10968 14288 11020 14340
rect 7656 14263 7708 14272
rect 7656 14229 7665 14263
rect 7665 14229 7699 14263
rect 7699 14229 7708 14263
rect 7656 14220 7708 14229
rect 8300 14263 8352 14272
rect 8300 14229 8309 14263
rect 8309 14229 8343 14263
rect 8343 14229 8352 14263
rect 8300 14220 8352 14229
rect 9680 14263 9732 14272
rect 9680 14229 9689 14263
rect 9689 14229 9723 14263
rect 9723 14229 9732 14263
rect 9680 14220 9732 14229
rect 10692 14220 10744 14272
rect 12072 14220 12124 14272
rect 13084 14220 13136 14272
rect 14924 14356 14976 14408
rect 20720 14356 20772 14408
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 15108 14288 15160 14340
rect 15568 14288 15620 14340
rect 15936 14288 15988 14340
rect 16120 14288 16172 14340
rect 19432 14288 19484 14340
rect 20536 14288 20588 14340
rect 13820 14220 13872 14272
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 3148 14059 3200 14068
rect 2320 13948 2372 14000
rect 2412 13880 2464 13932
rect 2688 13923 2740 13932
rect 2688 13889 2697 13923
rect 2697 13889 2731 13923
rect 2731 13889 2740 13923
rect 2688 13880 2740 13889
rect 3148 14025 3157 14059
rect 3157 14025 3191 14059
rect 3191 14025 3200 14059
rect 3148 14016 3200 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 5080 14059 5132 14068
rect 5080 14025 5089 14059
rect 5089 14025 5123 14059
rect 5123 14025 5132 14059
rect 5080 14016 5132 14025
rect 7012 14016 7064 14068
rect 4068 13948 4120 14000
rect 8852 13991 8904 14000
rect 8852 13957 8861 13991
rect 8861 13957 8895 13991
rect 8895 13957 8904 13991
rect 8852 13948 8904 13957
rect 9588 13948 9640 14000
rect 10232 14016 10284 14068
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 14464 14016 14516 14068
rect 15752 14016 15804 14068
rect 15936 14059 15988 14068
rect 15936 14025 15945 14059
rect 15945 14025 15979 14059
rect 15979 14025 15988 14059
rect 15936 14016 15988 14025
rect 18972 14059 19024 14068
rect 18972 14025 18981 14059
rect 18981 14025 19015 14059
rect 19015 14025 19024 14059
rect 18972 14016 19024 14025
rect 20352 14016 20404 14068
rect 11888 13948 11940 14000
rect 13820 13948 13872 14000
rect 17868 13991 17920 14000
rect 5356 13880 5408 13932
rect 2136 13812 2188 13864
rect 5080 13812 5132 13864
rect 5816 13855 5868 13864
rect 5816 13821 5825 13855
rect 5825 13821 5859 13855
rect 5859 13821 5868 13855
rect 5816 13812 5868 13821
rect 6552 13812 6604 13864
rect 6736 13812 6788 13864
rect 5448 13744 5500 13796
rect 6644 13744 6696 13796
rect 1676 13719 1728 13728
rect 1676 13685 1685 13719
rect 1685 13685 1719 13719
rect 1719 13685 1728 13719
rect 1676 13676 1728 13685
rect 3148 13676 3200 13728
rect 5724 13676 5776 13728
rect 9220 13923 9272 13932
rect 9220 13889 9229 13923
rect 9229 13889 9263 13923
rect 9263 13889 9272 13923
rect 9220 13880 9272 13889
rect 7472 13812 7524 13864
rect 10784 13880 10836 13932
rect 12256 13880 12308 13932
rect 12348 13880 12400 13932
rect 13728 13880 13780 13932
rect 7380 13744 7432 13796
rect 10968 13812 11020 13864
rect 7472 13676 7524 13728
rect 10876 13744 10928 13796
rect 17868 13957 17902 13991
rect 17902 13957 17920 13991
rect 17868 13948 17920 13957
rect 17592 13855 17644 13864
rect 12072 13676 12124 13728
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 16028 13676 16080 13728
rect 17592 13821 17601 13855
rect 17601 13821 17635 13855
rect 17635 13821 17644 13855
rect 17592 13812 17644 13821
rect 19984 13948 20036 14000
rect 20720 13948 20772 14000
rect 19984 13812 20036 13864
rect 18512 13676 18564 13728
rect 20168 13676 20220 13728
rect 20352 13676 20404 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2596 13472 2648 13524
rect 4804 13472 4856 13524
rect 5908 13472 5960 13524
rect 6644 13472 6696 13524
rect 2228 13404 2280 13456
rect 7012 13404 7064 13456
rect 1860 13379 1912 13388
rect 1860 13345 1869 13379
rect 1869 13345 1903 13379
rect 1903 13345 1912 13379
rect 1860 13336 1912 13345
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 7748 13404 7800 13456
rect 10508 13472 10560 13524
rect 10876 13472 10928 13524
rect 11888 13472 11940 13524
rect 12808 13472 12860 13524
rect 13176 13472 13228 13524
rect 16948 13472 17000 13524
rect 17040 13472 17092 13524
rect 17500 13472 17552 13524
rect 19984 13472 20036 13524
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 15200 13404 15252 13456
rect 1676 13268 1728 13320
rect 2688 13311 2740 13320
rect 2688 13277 2697 13311
rect 2697 13277 2731 13311
rect 2731 13277 2740 13311
rect 2688 13268 2740 13277
rect 3148 13268 3200 13320
rect 5816 13311 5868 13320
rect 5816 13277 5825 13311
rect 5825 13277 5859 13311
rect 5859 13277 5868 13311
rect 5816 13268 5868 13277
rect 6828 13268 6880 13320
rect 7748 13268 7800 13320
rect 8024 13268 8076 13320
rect 9220 13336 9272 13388
rect 15660 13336 15712 13388
rect 16028 13311 16080 13320
rect 8760 13200 8812 13252
rect 1676 13132 1728 13184
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 2872 13175 2924 13184
rect 2872 13141 2881 13175
rect 2881 13141 2915 13175
rect 2915 13141 2924 13175
rect 2872 13132 2924 13141
rect 4160 13175 4212 13184
rect 4160 13141 4169 13175
rect 4169 13141 4203 13175
rect 4203 13141 4212 13175
rect 4160 13132 4212 13141
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 5816 13132 5868 13184
rect 6736 13132 6788 13184
rect 7012 13132 7064 13184
rect 7472 13175 7524 13184
rect 7472 13141 7481 13175
rect 7481 13141 7515 13175
rect 7515 13141 7524 13175
rect 7472 13132 7524 13141
rect 7748 13132 7800 13184
rect 10232 13200 10284 13252
rect 12440 13200 12492 13252
rect 13084 13200 13136 13252
rect 9772 13132 9824 13184
rect 10968 13132 11020 13184
rect 11612 13132 11664 13184
rect 11796 13175 11848 13184
rect 11796 13141 11805 13175
rect 11805 13141 11839 13175
rect 11839 13141 11848 13175
rect 11796 13132 11848 13141
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16396 13200 16448 13252
rect 13728 13132 13780 13141
rect 17592 13268 17644 13320
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 20720 13268 20772 13277
rect 18420 13243 18472 13252
rect 18420 13209 18429 13243
rect 18429 13209 18463 13243
rect 18463 13209 18472 13243
rect 18420 13200 18472 13209
rect 20996 13200 21048 13252
rect 18328 13132 18380 13184
rect 19340 13175 19392 13184
rect 19340 13141 19349 13175
rect 19349 13141 19383 13175
rect 19383 13141 19392 13175
rect 19340 13132 19392 13141
rect 19708 13132 19760 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 2688 12971 2740 12980
rect 2688 12937 2697 12971
rect 2697 12937 2731 12971
rect 2731 12937 2740 12971
rect 2688 12928 2740 12937
rect 4252 12928 4304 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 7196 12928 7248 12980
rect 8484 12928 8536 12980
rect 2044 12792 2096 12844
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 4068 12860 4120 12912
rect 8208 12860 8260 12912
rect 10876 12971 10928 12980
rect 9864 12860 9916 12912
rect 10232 12860 10284 12912
rect 10324 12903 10376 12912
rect 10324 12869 10342 12903
rect 10342 12869 10376 12903
rect 10324 12860 10376 12869
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 4620 12792 4672 12844
rect 6644 12792 6696 12844
rect 8484 12792 8536 12844
rect 9496 12792 9548 12844
rect 2228 12724 2280 12733
rect 3976 12724 4028 12776
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 6552 12724 6604 12776
rect 7748 12767 7800 12776
rect 6000 12656 6052 12708
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 10876 12937 10885 12971
rect 10885 12937 10919 12971
rect 10919 12937 10928 12971
rect 10876 12928 10928 12937
rect 11060 12860 11112 12912
rect 11704 12860 11756 12912
rect 15108 12928 15160 12980
rect 16212 12971 16264 12980
rect 16212 12937 16221 12971
rect 16221 12937 16255 12971
rect 16255 12937 16264 12971
rect 16212 12928 16264 12937
rect 13176 12860 13228 12912
rect 14464 12792 14516 12844
rect 14924 12792 14976 12844
rect 15844 12860 15896 12912
rect 19340 12860 19392 12912
rect 20536 12928 20588 12980
rect 15660 12792 15712 12844
rect 16396 12792 16448 12844
rect 17500 12792 17552 12844
rect 18880 12792 18932 12844
rect 19800 12792 19852 12844
rect 19892 12792 19944 12844
rect 21456 12792 21508 12844
rect 13728 12767 13780 12776
rect 13728 12733 13737 12767
rect 13737 12733 13771 12767
rect 13771 12733 13780 12767
rect 13728 12724 13780 12733
rect 10600 12656 10652 12708
rect 4252 12588 4304 12640
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 4896 12588 4948 12640
rect 8300 12631 8352 12640
rect 8300 12597 8309 12631
rect 8309 12597 8343 12631
rect 8343 12597 8352 12631
rect 8300 12588 8352 12597
rect 8760 12588 8812 12640
rect 13820 12588 13872 12640
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 20076 12656 20128 12708
rect 14832 12588 14884 12640
rect 15660 12588 15712 12640
rect 18052 12588 18104 12640
rect 18144 12588 18196 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 3884 12427 3936 12436
rect 3884 12393 3893 12427
rect 3893 12393 3927 12427
rect 3927 12393 3936 12427
rect 3884 12384 3936 12393
rect 5540 12384 5592 12436
rect 5816 12384 5868 12436
rect 6092 12427 6144 12436
rect 6092 12393 6101 12427
rect 6101 12393 6135 12427
rect 6135 12393 6144 12427
rect 6092 12384 6144 12393
rect 6828 12384 6880 12436
rect 8024 12384 8076 12436
rect 8944 12384 8996 12436
rect 9220 12427 9272 12436
rect 9220 12393 9229 12427
rect 9229 12393 9263 12427
rect 9263 12393 9272 12427
rect 9220 12384 9272 12393
rect 11520 12384 11572 12436
rect 12624 12384 12676 12436
rect 13636 12384 13688 12436
rect 2964 12316 3016 12368
rect 5632 12316 5684 12368
rect 5724 12316 5776 12368
rect 6552 12316 6604 12368
rect 12808 12316 12860 12368
rect 13820 12316 13872 12368
rect 14280 12316 14332 12368
rect 18604 12384 18656 12436
rect 19708 12427 19760 12436
rect 19708 12393 19717 12427
rect 19717 12393 19751 12427
rect 19751 12393 19760 12427
rect 19708 12384 19760 12393
rect 20628 12384 20680 12436
rect 16948 12316 17000 12368
rect 1216 12248 1268 12300
rect 2504 12248 2556 12300
rect 4436 12291 4488 12300
rect 4436 12257 4445 12291
rect 4445 12257 4479 12291
rect 4479 12257 4488 12291
rect 4436 12248 4488 12257
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 7748 12248 7800 12300
rect 2228 12223 2280 12232
rect 2228 12189 2237 12223
rect 2237 12189 2271 12223
rect 2271 12189 2280 12223
rect 2228 12180 2280 12189
rect 3240 12180 3292 12232
rect 4068 12180 4120 12232
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 14004 12180 14056 12232
rect 15660 12223 15712 12232
rect 10324 12155 10376 12164
rect 2044 12044 2096 12096
rect 2872 12087 2924 12096
rect 2872 12053 2881 12087
rect 2881 12053 2915 12087
rect 2915 12053 2924 12087
rect 2872 12044 2924 12053
rect 3148 12044 3200 12096
rect 3424 12044 3476 12096
rect 3516 12044 3568 12096
rect 4344 12087 4396 12096
rect 4344 12053 4353 12087
rect 4353 12053 4387 12087
rect 4387 12053 4396 12087
rect 4344 12044 4396 12053
rect 4620 12044 4672 12096
rect 10324 12121 10342 12155
rect 10342 12121 10376 12155
rect 10324 12112 10376 12121
rect 8024 12044 8076 12096
rect 9220 12044 9272 12096
rect 13544 12112 13596 12164
rect 13728 12112 13780 12164
rect 15660 12189 15669 12223
rect 15669 12189 15703 12223
rect 15703 12189 15712 12223
rect 15660 12180 15712 12189
rect 16856 12248 16908 12300
rect 19524 12316 19576 12368
rect 15200 12112 15252 12164
rect 16856 12112 16908 12164
rect 21180 12180 21232 12232
rect 19984 12112 20036 12164
rect 14280 12044 14332 12096
rect 14464 12087 14516 12096
rect 14464 12053 14473 12087
rect 14473 12053 14507 12087
rect 14507 12053 14516 12087
rect 14464 12044 14516 12053
rect 15384 12087 15436 12096
rect 15384 12053 15393 12087
rect 15393 12053 15427 12087
rect 15427 12053 15436 12087
rect 15384 12044 15436 12053
rect 17040 12087 17092 12096
rect 17040 12053 17049 12087
rect 17049 12053 17083 12087
rect 17083 12053 17092 12087
rect 17040 12044 17092 12053
rect 17316 12087 17368 12096
rect 17316 12053 17325 12087
rect 17325 12053 17359 12087
rect 17359 12053 17368 12087
rect 17316 12044 17368 12053
rect 18144 12044 18196 12096
rect 20536 12112 20588 12164
rect 21548 12112 21600 12164
rect 21272 12044 21324 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 3516 11883 3568 11892
rect 3516 11849 3525 11883
rect 3525 11849 3559 11883
rect 3559 11849 3568 11883
rect 3516 11840 3568 11849
rect 4252 11883 4304 11892
rect 4252 11849 4261 11883
rect 4261 11849 4295 11883
rect 4295 11849 4304 11883
rect 4252 11840 4304 11849
rect 4344 11840 4396 11892
rect 7288 11883 7340 11892
rect 7288 11849 7297 11883
rect 7297 11849 7331 11883
rect 7331 11849 7340 11883
rect 7288 11840 7340 11849
rect 9128 11840 9180 11892
rect 13176 11883 13228 11892
rect 13176 11849 13185 11883
rect 13185 11849 13219 11883
rect 13219 11849 13228 11883
rect 13176 11840 13228 11849
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 15660 11840 15712 11892
rect 3976 11772 4028 11824
rect 6460 11772 6512 11824
rect 7472 11772 7524 11824
rect 10600 11815 10652 11824
rect 10600 11781 10618 11815
rect 10618 11781 10652 11815
rect 10600 11772 10652 11781
rect 11060 11772 11112 11824
rect 12164 11772 12216 11824
rect 13268 11772 13320 11824
rect 1952 11747 2004 11756
rect 1952 11713 1961 11747
rect 1961 11713 1995 11747
rect 1995 11713 2004 11747
rect 1952 11704 2004 11713
rect 2136 11704 2188 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 4068 11704 4120 11756
rect 5632 11747 5684 11756
rect 5632 11713 5641 11747
rect 5641 11713 5675 11747
rect 5675 11713 5684 11747
rect 5632 11704 5684 11713
rect 8116 11704 8168 11756
rect 8944 11704 8996 11756
rect 2228 11636 2280 11645
rect 1952 11568 2004 11620
rect 4344 11636 4396 11688
rect 4620 11636 4672 11688
rect 5816 11679 5868 11688
rect 3240 11568 3292 11620
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 6644 11679 6696 11688
rect 6644 11645 6653 11679
rect 6653 11645 6687 11679
rect 6687 11645 6696 11679
rect 6644 11636 6696 11645
rect 10876 11679 10928 11688
rect 8392 11568 8444 11620
rect 9404 11568 9456 11620
rect 7380 11500 7432 11552
rect 7748 11500 7800 11552
rect 8208 11500 8260 11552
rect 9496 11500 9548 11552
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 14372 11747 14424 11756
rect 14372 11713 14406 11747
rect 14406 11713 14424 11747
rect 14372 11704 14424 11713
rect 14832 11704 14884 11756
rect 18052 11704 18104 11756
rect 18236 11747 18288 11756
rect 18236 11713 18270 11747
rect 18270 11713 18288 11747
rect 18236 11704 18288 11713
rect 17316 11636 17368 11688
rect 19800 11840 19852 11892
rect 19984 11840 20036 11892
rect 20904 11840 20956 11892
rect 21272 11883 21324 11892
rect 21272 11849 21281 11883
rect 21281 11849 21315 11883
rect 21315 11849 21324 11883
rect 21272 11840 21324 11849
rect 20168 11747 20220 11756
rect 20168 11713 20177 11747
rect 20177 11713 20211 11747
rect 20211 11713 20220 11747
rect 20168 11704 20220 11713
rect 21456 11704 21508 11756
rect 15200 11568 15252 11620
rect 15384 11568 15436 11620
rect 16488 11568 16540 11620
rect 11060 11500 11112 11552
rect 15476 11543 15528 11552
rect 15476 11509 15485 11543
rect 15485 11509 15519 11543
rect 15519 11509 15528 11543
rect 15476 11500 15528 11509
rect 17316 11500 17368 11552
rect 19800 11568 19852 11620
rect 20444 11568 20496 11620
rect 19524 11500 19576 11552
rect 20904 11568 20956 11620
rect 21088 11500 21140 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1860 11296 1912 11348
rect 5172 11296 5224 11348
rect 1952 11228 2004 11280
rect 6920 11296 6972 11348
rect 9680 11296 9732 11348
rect 10232 11296 10284 11348
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 2504 11160 2556 11212
rect 4620 11160 4672 11212
rect 5172 11160 5224 11212
rect 5724 11160 5776 11212
rect 2044 11135 2096 11144
rect 2044 11101 2053 11135
rect 2053 11101 2087 11135
rect 2087 11101 2096 11135
rect 2044 11092 2096 11101
rect 2964 11092 3016 11144
rect 3240 11092 3292 11144
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 4436 11092 4488 11144
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 6000 11135 6052 11144
rect 6000 11101 6009 11135
rect 6009 11101 6043 11135
rect 6043 11101 6052 11135
rect 6000 11092 6052 11101
rect 4712 11024 4764 11076
rect 5356 11024 5408 11076
rect 5724 11024 5776 11076
rect 8024 11160 8076 11212
rect 12624 11228 12676 11280
rect 6644 11092 6696 11144
rect 7472 11092 7524 11144
rect 8208 11135 8260 11144
rect 8208 11101 8217 11135
rect 8217 11101 8251 11135
rect 8251 11101 8260 11135
rect 8208 11092 8260 11101
rect 8300 11092 8352 11144
rect 8576 11092 8628 11144
rect 8760 11092 8812 11144
rect 8668 11024 8720 11076
rect 9128 11092 9180 11144
rect 11060 11160 11112 11212
rect 12532 11203 12584 11212
rect 10784 11092 10836 11144
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 12532 11169 12541 11203
rect 12541 11169 12575 11203
rect 12575 11169 12584 11203
rect 12532 11160 12584 11169
rect 12900 11160 12952 11212
rect 12624 11092 12676 11144
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 5632 10999 5684 11008
rect 5632 10965 5641 10999
rect 5641 10965 5675 10999
rect 5675 10965 5684 10999
rect 5632 10956 5684 10965
rect 6644 10999 6696 11008
rect 6644 10965 6653 10999
rect 6653 10965 6687 10999
rect 6687 10965 6696 10999
rect 6644 10956 6696 10965
rect 6828 10956 6880 11008
rect 7840 10999 7892 11008
rect 7840 10965 7849 10999
rect 7849 10965 7883 10999
rect 7883 10965 7892 10999
rect 7840 10956 7892 10965
rect 8116 10956 8168 11008
rect 11888 11024 11940 11076
rect 10784 10956 10836 11008
rect 11244 10956 11296 11008
rect 13544 11296 13596 11348
rect 14924 11296 14976 11348
rect 18972 11296 19024 11348
rect 15384 11228 15436 11280
rect 16580 11228 16632 11280
rect 18604 11228 18656 11280
rect 19524 11228 19576 11280
rect 14924 11160 14976 11212
rect 15016 11092 15068 11144
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 17408 11092 17460 11144
rect 18052 11092 18104 11144
rect 21272 11296 21324 11348
rect 20996 11092 21048 11144
rect 13268 11024 13320 11076
rect 13360 10999 13412 11008
rect 13360 10965 13369 10999
rect 13369 10965 13403 10999
rect 13403 10965 13412 10999
rect 13360 10956 13412 10965
rect 20904 11024 20956 11076
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 2412 10752 2464 10804
rect 2136 10684 2188 10736
rect 2688 10752 2740 10804
rect 3884 10795 3936 10804
rect 3884 10761 3893 10795
rect 3893 10761 3927 10795
rect 3927 10761 3936 10795
rect 3884 10752 3936 10761
rect 4436 10752 4488 10804
rect 1768 10616 1820 10668
rect 2780 10616 2832 10668
rect 3424 10616 3476 10668
rect 4252 10684 4304 10736
rect 5448 10752 5500 10804
rect 6644 10752 6696 10804
rect 7564 10752 7616 10804
rect 8208 10752 8260 10804
rect 8484 10752 8536 10804
rect 9220 10795 9272 10804
rect 9220 10761 9229 10795
rect 9229 10761 9263 10795
rect 9263 10761 9272 10795
rect 9220 10752 9272 10761
rect 10324 10752 10376 10804
rect 14924 10795 14976 10804
rect 14924 10761 14933 10795
rect 14933 10761 14967 10795
rect 14967 10761 14976 10795
rect 14924 10752 14976 10761
rect 17316 10752 17368 10804
rect 5816 10684 5868 10736
rect 8116 10684 8168 10736
rect 4896 10616 4948 10668
rect 5448 10659 5500 10668
rect 5448 10625 5457 10659
rect 5457 10625 5491 10659
rect 5491 10625 5500 10659
rect 5448 10616 5500 10625
rect 2412 10548 2464 10600
rect 3976 10591 4028 10600
rect 2504 10480 2556 10532
rect 2688 10480 2740 10532
rect 3976 10557 3985 10591
rect 3985 10557 4019 10591
rect 4019 10557 4028 10591
rect 3976 10548 4028 10557
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4620 10548 4672 10600
rect 7288 10548 7340 10600
rect 8576 10684 8628 10736
rect 8760 10727 8812 10736
rect 8760 10693 8769 10727
rect 8769 10693 8803 10727
rect 8803 10693 8812 10727
rect 8760 10684 8812 10693
rect 11244 10684 11296 10736
rect 8116 10591 8168 10600
rect 7564 10480 7616 10532
rect 2964 10412 3016 10464
rect 5264 10455 5316 10464
rect 5264 10421 5273 10455
rect 5273 10421 5307 10455
rect 5307 10421 5316 10455
rect 5264 10412 5316 10421
rect 5356 10412 5408 10464
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 7104 10412 7156 10464
rect 8116 10557 8125 10591
rect 8125 10557 8159 10591
rect 8159 10557 8168 10591
rect 8116 10548 8168 10557
rect 8484 10548 8536 10600
rect 10508 10616 10560 10668
rect 12624 10659 12676 10668
rect 12624 10625 12642 10659
rect 12642 10625 12676 10659
rect 12624 10616 12676 10625
rect 13360 10616 13412 10668
rect 17684 10752 17736 10804
rect 17868 10752 17920 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 21180 10795 21232 10804
rect 21180 10761 21189 10795
rect 21189 10761 21223 10795
rect 21223 10761 21232 10795
rect 21180 10752 21232 10761
rect 17776 10684 17828 10736
rect 19800 10727 19852 10736
rect 19800 10693 19834 10727
rect 19834 10693 19852 10727
rect 19800 10684 19852 10693
rect 17684 10616 17736 10668
rect 20720 10616 20772 10668
rect 20996 10616 21048 10668
rect 21364 10659 21416 10668
rect 21364 10625 21373 10659
rect 21373 10625 21407 10659
rect 21407 10625 21416 10659
rect 21364 10616 21416 10625
rect 10416 10412 10468 10464
rect 10692 10480 10744 10532
rect 11244 10412 11296 10464
rect 17132 10480 17184 10532
rect 14280 10412 14332 10464
rect 17592 10412 17644 10464
rect 19524 10412 19576 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1400 10208 1452 10260
rect 5264 10208 5316 10260
rect 6828 10208 6880 10260
rect 7288 10251 7340 10260
rect 7288 10217 7297 10251
rect 7297 10217 7331 10251
rect 7331 10217 7340 10251
rect 7288 10208 7340 10217
rect 8024 10208 8076 10260
rect 13820 10208 13872 10260
rect 17684 10251 17736 10260
rect 1676 10072 1728 10124
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 3332 10140 3384 10192
rect 3700 10140 3752 10192
rect 4344 10140 4396 10192
rect 4804 10140 4856 10192
rect 6920 10140 6972 10192
rect 8116 10140 8168 10192
rect 10692 10140 10744 10192
rect 15660 10183 15712 10192
rect 2228 10004 2280 10013
rect 3056 10004 3108 10056
rect 3424 10072 3476 10124
rect 5264 10072 5316 10124
rect 8208 10072 8260 10124
rect 9312 10072 9364 10124
rect 10416 10072 10468 10124
rect 11796 10072 11848 10124
rect 15660 10149 15669 10183
rect 15669 10149 15703 10183
rect 15703 10149 15712 10183
rect 15660 10140 15712 10149
rect 17684 10217 17693 10251
rect 17693 10217 17727 10251
rect 17727 10217 17736 10251
rect 17684 10208 17736 10217
rect 19616 10208 19668 10260
rect 3516 10004 3568 10056
rect 8116 10004 8168 10056
rect 3240 9936 3292 9988
rect 4712 9936 4764 9988
rect 7748 9979 7800 9988
rect 7748 9945 7757 9979
rect 7757 9945 7791 9979
rect 7791 9945 7800 9979
rect 7748 9936 7800 9945
rect 2504 9911 2556 9920
rect 2504 9877 2513 9911
rect 2513 9877 2547 9911
rect 2547 9877 2556 9911
rect 2504 9868 2556 9877
rect 2780 9868 2832 9920
rect 3056 9868 3108 9920
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 4804 9911 4856 9920
rect 4804 9877 4813 9911
rect 4813 9877 4847 9911
rect 4847 9877 4856 9911
rect 4804 9868 4856 9877
rect 5356 9868 5408 9920
rect 6000 9868 6052 9920
rect 6644 9868 6696 9920
rect 6920 9911 6972 9920
rect 6920 9877 6929 9911
rect 6929 9877 6963 9911
rect 6963 9877 6972 9911
rect 6920 9868 6972 9877
rect 7104 9868 7156 9920
rect 7932 9868 7984 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 9496 10004 9548 10056
rect 11244 10004 11296 10056
rect 9220 9936 9272 9988
rect 15936 10004 15988 10056
rect 17960 10072 18012 10124
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 19524 10072 19576 10124
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 21088 10072 21140 10124
rect 18788 10004 18840 10056
rect 20628 10004 20680 10056
rect 11244 9911 11296 9920
rect 11244 9877 11253 9911
rect 11253 9877 11287 9911
rect 11287 9877 11296 9911
rect 11244 9868 11296 9877
rect 14096 9936 14148 9988
rect 14464 9936 14516 9988
rect 20168 9936 20220 9988
rect 13820 9868 13872 9920
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 17592 9868 17644 9920
rect 19800 9868 19852 9920
rect 19984 9911 20036 9920
rect 19984 9877 19993 9911
rect 19993 9877 20027 9911
rect 20027 9877 20036 9911
rect 19984 9868 20036 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 2412 9707 2464 9716
rect 2412 9673 2421 9707
rect 2421 9673 2455 9707
rect 2455 9673 2464 9707
rect 2412 9664 2464 9673
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 2228 9528 2280 9580
rect 2412 9528 2464 9580
rect 3884 9664 3936 9716
rect 3056 9596 3108 9648
rect 3700 9596 3752 9648
rect 6920 9664 6972 9716
rect 7564 9664 7616 9716
rect 8116 9707 8168 9716
rect 8116 9673 8125 9707
rect 8125 9673 8159 9707
rect 8159 9673 8168 9707
rect 8116 9664 8168 9673
rect 9036 9664 9088 9716
rect 4160 9528 4212 9580
rect 4896 9596 4948 9648
rect 5908 9596 5960 9648
rect 6644 9596 6696 9648
rect 8300 9596 8352 9648
rect 9312 9596 9364 9648
rect 9864 9596 9916 9648
rect 10784 9596 10836 9648
rect 11244 9596 11296 9648
rect 11520 9596 11572 9648
rect 4620 9528 4672 9580
rect 8668 9528 8720 9580
rect 12440 9596 12492 9648
rect 13728 9596 13780 9648
rect 13820 9596 13872 9648
rect 17408 9664 17460 9716
rect 20996 9664 21048 9716
rect 3056 9503 3108 9512
rect 3056 9469 3065 9503
rect 3065 9469 3099 9503
rect 3099 9469 3108 9503
rect 3056 9460 3108 9469
rect 3332 9460 3384 9512
rect 3976 9460 4028 9512
rect 4252 9503 4304 9512
rect 4252 9469 4261 9503
rect 4261 9469 4295 9503
rect 4295 9469 4304 9503
rect 4252 9460 4304 9469
rect 5172 9460 5224 9512
rect 5448 9503 5500 9512
rect 2780 9392 2832 9444
rect 4068 9392 4120 9444
rect 4528 9392 4580 9444
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 5816 9460 5868 9512
rect 6736 9460 6788 9512
rect 8300 9460 8352 9512
rect 9496 9503 9548 9512
rect 9496 9469 9505 9503
rect 9505 9469 9539 9503
rect 9539 9469 9548 9503
rect 9496 9460 9548 9469
rect 11060 9392 11112 9444
rect 3608 9367 3660 9376
rect 3608 9333 3617 9367
rect 3617 9333 3651 9367
rect 3651 9333 3660 9367
rect 3608 9324 3660 9333
rect 3976 9324 4028 9376
rect 5540 9324 5592 9376
rect 6644 9324 6696 9376
rect 6736 9324 6788 9376
rect 8208 9324 8260 9376
rect 11244 9324 11296 9376
rect 11520 9367 11572 9376
rect 11520 9333 11529 9367
rect 11529 9333 11563 9367
rect 11563 9333 11572 9367
rect 11520 9324 11572 9333
rect 15936 9571 15988 9580
rect 15936 9537 15945 9571
rect 15945 9537 15979 9571
rect 15979 9537 15988 9571
rect 15936 9528 15988 9537
rect 17776 9528 17828 9580
rect 17868 9528 17920 9580
rect 19248 9528 19300 9580
rect 20168 9571 20220 9580
rect 17960 9460 18012 9512
rect 19708 9503 19760 9512
rect 14096 9392 14148 9444
rect 14556 9435 14608 9444
rect 14556 9401 14565 9435
rect 14565 9401 14599 9435
rect 14599 9401 14608 9435
rect 14556 9392 14608 9401
rect 19708 9469 19717 9503
rect 19717 9469 19751 9503
rect 19751 9469 19760 9503
rect 19708 9460 19760 9469
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 14464 9324 14516 9376
rect 14924 9324 14976 9376
rect 17040 9324 17092 9376
rect 17500 9324 17552 9376
rect 17868 9324 17920 9376
rect 20720 9392 20772 9444
rect 21180 9392 21232 9444
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2780 9120 2832 9172
rect 5448 9120 5500 9172
rect 2228 9052 2280 9104
rect 3884 9052 3936 9104
rect 4068 9052 4120 9104
rect 4804 9052 4856 9104
rect 10048 9120 10100 9172
rect 10784 9163 10836 9172
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 10876 9120 10928 9172
rect 13728 9163 13780 9172
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 1584 8984 1636 9036
rect 15108 9052 15160 9104
rect 2136 8916 2188 8968
rect 3148 8959 3200 8968
rect 3148 8925 3157 8959
rect 3157 8925 3191 8959
rect 3191 8925 3200 8959
rect 3148 8916 3200 8925
rect 4252 8916 4304 8968
rect 1768 8848 1820 8900
rect 3056 8848 3108 8900
rect 5632 8984 5684 9036
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 8208 9027 8260 9036
rect 4436 8916 4488 8968
rect 5724 8916 5776 8968
rect 6644 8959 6696 8968
rect 2228 8780 2280 8832
rect 3976 8780 4028 8832
rect 5540 8848 5592 8900
rect 6644 8925 6653 8959
rect 6653 8925 6687 8959
rect 6687 8925 6696 8959
rect 6644 8916 6696 8925
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 11704 8984 11756 9036
rect 13820 8984 13872 9036
rect 15936 9120 15988 9172
rect 16120 9120 16172 9172
rect 17776 9120 17828 9172
rect 19984 9120 20036 9172
rect 21272 9052 21324 9104
rect 8024 8916 8076 8968
rect 9496 8916 9548 8968
rect 4344 8780 4396 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 5724 8780 5776 8832
rect 5908 8780 5960 8832
rect 6828 8848 6880 8900
rect 8116 8848 8168 8900
rect 7104 8780 7156 8832
rect 7748 8780 7800 8832
rect 8668 8780 8720 8832
rect 9036 8780 9088 8832
rect 10968 8848 11020 8900
rect 11520 8916 11572 8968
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 15476 8916 15528 8968
rect 16488 8916 16540 8968
rect 17776 8984 17828 9036
rect 19616 9027 19668 9036
rect 19616 8993 19625 9027
rect 19625 8993 19659 9027
rect 19659 8993 19668 9027
rect 19616 8984 19668 8993
rect 20812 8984 20864 9036
rect 20996 9027 21048 9036
rect 20996 8993 21005 9027
rect 21005 8993 21039 9027
rect 21039 8993 21048 9027
rect 20996 8984 21048 8993
rect 17408 8916 17460 8968
rect 17868 8848 17920 8900
rect 11060 8823 11112 8832
rect 11060 8789 11069 8823
rect 11069 8789 11103 8823
rect 11103 8789 11112 8823
rect 11060 8780 11112 8789
rect 12164 8780 12216 8832
rect 12348 8780 12400 8832
rect 12440 8780 12492 8832
rect 15384 8780 15436 8832
rect 15752 8780 15804 8832
rect 16212 8780 16264 8832
rect 16488 8780 16540 8832
rect 17040 8780 17092 8832
rect 17500 8780 17552 8832
rect 18052 8780 18104 8832
rect 18972 8848 19024 8900
rect 19984 8780 20036 8832
rect 20168 8823 20220 8832
rect 20168 8789 20177 8823
rect 20177 8789 20211 8823
rect 20211 8789 20220 8823
rect 20168 8780 20220 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2320 8576 2372 8628
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 4528 8619 4580 8628
rect 4528 8585 4537 8619
rect 4537 8585 4571 8619
rect 4571 8585 4580 8619
rect 4528 8576 4580 8585
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 5356 8576 5408 8628
rect 7748 8576 7800 8628
rect 7840 8576 7892 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 12624 8576 12676 8628
rect 13820 8619 13872 8628
rect 13820 8585 13829 8619
rect 13829 8585 13863 8619
rect 13863 8585 13872 8619
rect 13820 8576 13872 8585
rect 15200 8576 15252 8628
rect 15476 8576 15528 8628
rect 1584 8508 1636 8560
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2872 8483 2924 8492
rect 2872 8449 2881 8483
rect 2881 8449 2915 8483
rect 2915 8449 2924 8483
rect 2872 8440 2924 8449
rect 6828 8508 6880 8560
rect 9496 8508 9548 8560
rect 9956 8508 10008 8560
rect 10968 8508 11020 8560
rect 11980 8551 12032 8560
rect 6920 8440 6972 8492
rect 8024 8440 8076 8492
rect 9036 8440 9088 8492
rect 11244 8440 11296 8492
rect 11980 8517 11989 8551
rect 11989 8517 12023 8551
rect 12023 8517 12032 8551
rect 11980 8508 12032 8517
rect 12440 8508 12492 8560
rect 15660 8508 15712 8560
rect 14924 8440 14976 8492
rect 15200 8483 15252 8492
rect 15200 8449 15218 8483
rect 15218 8449 15252 8483
rect 15200 8440 15252 8449
rect 15384 8440 15436 8492
rect 15936 8576 15988 8628
rect 18052 8576 18104 8628
rect 18236 8576 18288 8628
rect 18880 8508 18932 8560
rect 17500 8440 17552 8492
rect 17868 8440 17920 8492
rect 18052 8440 18104 8492
rect 21180 8483 21232 8492
rect 21180 8449 21189 8483
rect 21189 8449 21223 8483
rect 21223 8449 21232 8483
rect 21180 8440 21232 8449
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 2688 8372 2740 8424
rect 3148 8372 3200 8424
rect 4988 8415 5040 8424
rect 4988 8381 4997 8415
rect 4997 8381 5031 8415
rect 5031 8381 5040 8415
rect 4988 8372 5040 8381
rect 5172 8415 5224 8424
rect 5172 8381 5181 8415
rect 5181 8381 5215 8415
rect 5215 8381 5224 8415
rect 5172 8372 5224 8381
rect 7564 8372 7616 8424
rect 10876 8372 10928 8424
rect 11336 8372 11388 8424
rect 11980 8372 12032 8424
rect 3884 8304 3936 8356
rect 4068 8304 4120 8356
rect 3516 8236 3568 8288
rect 4620 8236 4672 8288
rect 6552 8304 6604 8356
rect 6920 8304 6972 8356
rect 7656 8304 7708 8356
rect 8668 8304 8720 8356
rect 11060 8304 11112 8356
rect 12440 8304 12492 8356
rect 12624 8304 12676 8356
rect 15476 8304 15528 8356
rect 15844 8304 15896 8356
rect 16120 8347 16172 8356
rect 16120 8313 16129 8347
rect 16129 8313 16163 8347
rect 16163 8313 16172 8347
rect 16120 8304 16172 8313
rect 17408 8372 17460 8424
rect 15568 8236 15620 8288
rect 17408 8236 17460 8288
rect 17776 8304 17828 8356
rect 19064 8236 19116 8288
rect 19616 8236 19668 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2780 8032 2832 8084
rect 4252 8032 4304 8084
rect 6552 8032 6604 8084
rect 6828 8032 6880 8084
rect 8300 8032 8352 8084
rect 8760 8032 8812 8084
rect 9588 8032 9640 8084
rect 10048 8032 10100 8084
rect 14648 8032 14700 8084
rect 15936 8032 15988 8084
rect 16948 8032 17000 8084
rect 1676 7939 1728 7948
rect 1676 7905 1685 7939
rect 1685 7905 1719 7939
rect 1719 7905 1728 7939
rect 1676 7896 1728 7905
rect 4344 7896 4396 7948
rect 4896 7964 4948 8016
rect 5172 7896 5224 7948
rect 3148 7828 3200 7880
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4436 7828 4488 7880
rect 5724 7939 5776 7948
rect 5724 7905 5733 7939
rect 5733 7905 5767 7939
rect 5767 7905 5776 7939
rect 5724 7896 5776 7905
rect 7104 7939 7156 7948
rect 7104 7905 7113 7939
rect 7113 7905 7147 7939
rect 7147 7905 7156 7939
rect 7104 7896 7156 7905
rect 7748 7964 7800 8016
rect 9036 7964 9088 8016
rect 9220 7964 9272 8016
rect 12808 7964 12860 8016
rect 18052 8032 18104 8084
rect 18788 8032 18840 8084
rect 17960 7964 18012 8016
rect 8300 7939 8352 7948
rect 8300 7905 8309 7939
rect 8309 7905 8343 7939
rect 8343 7905 8352 7939
rect 8300 7896 8352 7905
rect 2136 7760 2188 7812
rect 3424 7760 3476 7812
rect 1860 7735 1912 7744
rect 1860 7701 1869 7735
rect 1869 7701 1903 7735
rect 1903 7701 1912 7735
rect 3240 7735 3292 7744
rect 1860 7692 1912 7701
rect 3240 7701 3249 7735
rect 3249 7701 3283 7735
rect 3283 7701 3292 7735
rect 3240 7692 3292 7701
rect 3332 7692 3384 7744
rect 6000 7692 6052 7744
rect 6552 7692 6604 7744
rect 7012 7735 7064 7744
rect 7012 7701 7021 7735
rect 7021 7701 7055 7735
rect 7055 7701 7064 7735
rect 7012 7692 7064 7701
rect 7840 7828 7892 7880
rect 9220 7828 9272 7880
rect 18420 7896 18472 7948
rect 19248 7896 19300 7948
rect 19800 7896 19852 7948
rect 9312 7760 9364 7812
rect 9128 7692 9180 7744
rect 10048 7871 10100 7880
rect 10048 7837 10066 7871
rect 10066 7837 10100 7871
rect 10048 7828 10100 7837
rect 12348 7828 12400 7880
rect 15108 7828 15160 7880
rect 16948 7828 17000 7880
rect 17408 7828 17460 7880
rect 18052 7828 18104 7880
rect 18512 7828 18564 7880
rect 18696 7828 18748 7880
rect 19892 7828 19944 7880
rect 21272 7871 21324 7880
rect 21272 7837 21281 7871
rect 21281 7837 21315 7871
rect 21315 7837 21324 7871
rect 21272 7828 21324 7837
rect 9588 7760 9640 7812
rect 15292 7760 15344 7812
rect 15660 7760 15712 7812
rect 10692 7692 10744 7744
rect 12164 7692 12216 7744
rect 13728 7692 13780 7744
rect 14280 7735 14332 7744
rect 14280 7701 14289 7735
rect 14289 7701 14323 7735
rect 14323 7701 14332 7735
rect 14280 7692 14332 7701
rect 14648 7735 14700 7744
rect 14648 7701 14657 7735
rect 14657 7701 14691 7735
rect 14691 7701 14700 7735
rect 14648 7692 14700 7701
rect 15476 7735 15528 7744
rect 15476 7701 15485 7735
rect 15485 7701 15519 7735
rect 15519 7701 15528 7735
rect 15476 7692 15528 7701
rect 16212 7735 16264 7744
rect 16212 7701 16221 7735
rect 16221 7701 16255 7735
rect 16255 7701 16264 7735
rect 16212 7692 16264 7701
rect 18788 7803 18840 7812
rect 18788 7769 18797 7803
rect 18797 7769 18831 7803
rect 18831 7769 18840 7803
rect 18788 7760 18840 7769
rect 19616 7803 19668 7812
rect 19616 7769 19625 7803
rect 19625 7769 19659 7803
rect 19659 7769 19668 7803
rect 19616 7760 19668 7769
rect 20076 7760 20128 7812
rect 20444 7760 20496 7812
rect 21088 7803 21140 7812
rect 21088 7769 21097 7803
rect 21097 7769 21131 7803
rect 21131 7769 21140 7803
rect 21088 7760 21140 7769
rect 18696 7692 18748 7744
rect 20720 7692 20772 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1584 7531 1636 7540
rect 1584 7497 1593 7531
rect 1593 7497 1627 7531
rect 1627 7497 1636 7531
rect 1584 7488 1636 7497
rect 2504 7488 2556 7540
rect 4344 7531 4396 7540
rect 4344 7497 4353 7531
rect 4353 7497 4387 7531
rect 4387 7497 4396 7531
rect 4344 7488 4396 7497
rect 5448 7488 5500 7540
rect 6000 7531 6052 7540
rect 6000 7497 6009 7531
rect 6009 7497 6043 7531
rect 6043 7497 6052 7531
rect 6000 7488 6052 7497
rect 3056 7420 3108 7472
rect 3240 7420 3292 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 3424 7395 3476 7404
rect 3424 7361 3433 7395
rect 3433 7361 3467 7395
rect 3467 7361 3476 7395
rect 3424 7352 3476 7361
rect 10876 7488 10928 7540
rect 15936 7488 15988 7540
rect 7380 7463 7432 7472
rect 7380 7429 7389 7463
rect 7389 7429 7423 7463
rect 7423 7429 7432 7463
rect 7380 7420 7432 7429
rect 12256 7420 12308 7472
rect 12348 7420 12400 7472
rect 12440 7420 12492 7472
rect 7932 7395 7984 7404
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 7932 7361 7941 7395
rect 7941 7361 7975 7395
rect 7975 7361 7984 7395
rect 7932 7352 7984 7361
rect 8300 7352 8352 7404
rect 9220 7352 9272 7404
rect 12624 7395 12676 7404
rect 16948 7463 17000 7472
rect 12624 7361 12642 7395
rect 12642 7361 12676 7395
rect 12624 7352 12676 7361
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 4068 7284 4120 7336
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 2688 7191 2740 7200
rect 2688 7157 2697 7191
rect 2697 7157 2731 7191
rect 2731 7157 2740 7191
rect 2688 7148 2740 7157
rect 2964 7191 3016 7200
rect 2964 7157 2973 7191
rect 2973 7157 3007 7191
rect 3007 7157 3016 7191
rect 2964 7148 3016 7157
rect 3240 7148 3292 7200
rect 3976 7148 4028 7200
rect 5540 7327 5592 7336
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 9772 7284 9824 7336
rect 15200 7352 15252 7404
rect 16212 7352 16264 7404
rect 16948 7429 16982 7463
rect 16982 7429 17000 7463
rect 16948 7420 17000 7429
rect 17132 7420 17184 7472
rect 18144 7488 18196 7540
rect 18880 7488 18932 7540
rect 19064 7488 19116 7540
rect 21364 7488 21416 7540
rect 19156 7463 19208 7472
rect 17500 7352 17552 7404
rect 18696 7352 18748 7404
rect 19156 7429 19165 7463
rect 19165 7429 19199 7463
rect 19199 7429 19208 7463
rect 19156 7420 19208 7429
rect 19800 7420 19852 7472
rect 20076 7463 20128 7472
rect 20076 7429 20085 7463
rect 20085 7429 20119 7463
rect 20119 7429 20128 7463
rect 20076 7420 20128 7429
rect 5632 7216 5684 7268
rect 7840 7216 7892 7268
rect 8300 7216 8352 7268
rect 6000 7148 6052 7200
rect 7196 7148 7248 7200
rect 7932 7148 7984 7200
rect 8760 7148 8812 7200
rect 10048 7148 10100 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 12164 7148 12216 7200
rect 12256 7148 12308 7200
rect 15568 7284 15620 7336
rect 18328 7327 18380 7336
rect 15016 7191 15068 7200
rect 15016 7157 15025 7191
rect 15025 7157 15059 7191
rect 15059 7157 15068 7191
rect 15016 7148 15068 7157
rect 15936 7148 15988 7200
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 18880 7284 18932 7336
rect 19248 7352 19300 7404
rect 20536 7395 20588 7404
rect 20536 7361 20545 7395
rect 20545 7361 20579 7395
rect 20579 7361 20588 7395
rect 20536 7352 20588 7361
rect 21456 7352 21508 7404
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2136 6987 2188 6996
rect 2136 6953 2145 6987
rect 2145 6953 2179 6987
rect 2179 6953 2188 6987
rect 2136 6944 2188 6953
rect 2228 6944 2280 6996
rect 2504 6944 2556 6996
rect 4896 6944 4948 6996
rect 5172 6944 5224 6996
rect 6920 6944 6972 6996
rect 7012 6944 7064 6996
rect 8024 6944 8076 6996
rect 8484 6987 8536 6996
rect 8484 6953 8493 6987
rect 8493 6953 8527 6987
rect 8527 6953 8536 6987
rect 8484 6944 8536 6953
rect 9220 6987 9272 6996
rect 9220 6953 9229 6987
rect 9229 6953 9263 6987
rect 9263 6953 9272 6987
rect 9220 6944 9272 6953
rect 9864 6944 9916 6996
rect 10600 6944 10652 6996
rect 12256 6944 12308 6996
rect 12348 6944 12400 6996
rect 12808 6944 12860 6996
rect 2780 6876 2832 6928
rect 4620 6876 4672 6928
rect 1492 6783 1544 6792
rect 1492 6749 1501 6783
rect 1501 6749 1535 6783
rect 1535 6749 1544 6783
rect 1492 6740 1544 6749
rect 5816 6851 5868 6860
rect 5816 6817 5825 6851
rect 5825 6817 5859 6851
rect 5859 6817 5868 6851
rect 5816 6808 5868 6817
rect 7380 6876 7432 6928
rect 7472 6808 7524 6860
rect 8208 6808 8260 6860
rect 2780 6783 2832 6792
rect 2780 6749 2789 6783
rect 2789 6749 2823 6783
rect 2823 6749 2832 6783
rect 2780 6740 2832 6749
rect 3332 6740 3384 6792
rect 5356 6740 5408 6792
rect 6000 6740 6052 6792
rect 3240 6604 3292 6656
rect 3424 6604 3476 6656
rect 3976 6604 4028 6656
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4620 6604 4672 6656
rect 5172 6647 5224 6656
rect 5172 6613 5181 6647
rect 5181 6613 5215 6647
rect 5215 6613 5224 6647
rect 5172 6604 5224 6613
rect 5264 6604 5316 6656
rect 5724 6672 5776 6724
rect 7840 6740 7892 6792
rect 7472 6672 7524 6724
rect 7748 6672 7800 6724
rect 9772 6740 9824 6792
rect 13636 6808 13688 6860
rect 18052 6808 18104 6860
rect 20352 6944 20404 6996
rect 19432 6808 19484 6860
rect 19616 6851 19668 6860
rect 19616 6817 19625 6851
rect 19625 6817 19659 6851
rect 19659 6817 19668 6851
rect 19616 6808 19668 6817
rect 20168 6808 20220 6860
rect 11060 6740 11112 6792
rect 10140 6672 10192 6724
rect 6184 6604 6236 6656
rect 7012 6604 7064 6656
rect 7104 6604 7156 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 7840 6604 7892 6613
rect 9772 6604 9824 6656
rect 11060 6604 11112 6656
rect 11796 6715 11848 6724
rect 11796 6681 11805 6715
rect 11805 6681 11839 6715
rect 11839 6681 11848 6715
rect 11796 6672 11848 6681
rect 13820 6740 13872 6792
rect 14832 6783 14884 6792
rect 14832 6749 14866 6783
rect 14866 6749 14884 6783
rect 14832 6740 14884 6749
rect 15292 6740 15344 6792
rect 15200 6672 15252 6724
rect 16028 6604 16080 6656
rect 16948 6647 17000 6656
rect 16948 6613 16957 6647
rect 16957 6613 16991 6647
rect 16991 6613 17000 6647
rect 16948 6604 17000 6613
rect 18328 6740 18380 6792
rect 18788 6740 18840 6792
rect 17960 6672 18012 6724
rect 18604 6672 18656 6724
rect 19616 6672 19668 6724
rect 18420 6647 18472 6656
rect 18420 6613 18429 6647
rect 18429 6613 18463 6647
rect 18463 6613 18472 6647
rect 18420 6604 18472 6613
rect 18788 6604 18840 6656
rect 19248 6604 19300 6656
rect 20260 6647 20312 6656
rect 20260 6613 20269 6647
rect 20269 6613 20303 6647
rect 20303 6613 20312 6647
rect 20260 6604 20312 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 2596 6443 2648 6452
rect 2596 6409 2605 6443
rect 2605 6409 2639 6443
rect 2639 6409 2648 6443
rect 2596 6400 2648 6409
rect 2964 6400 3016 6452
rect 3332 6400 3384 6452
rect 2780 6332 2832 6384
rect 5264 6400 5316 6452
rect 1768 6239 1820 6248
rect 1768 6205 1777 6239
rect 1777 6205 1811 6239
rect 1811 6205 1820 6239
rect 1768 6196 1820 6205
rect 2688 6264 2740 6316
rect 3056 6264 3108 6316
rect 3424 6264 3476 6316
rect 2872 6128 2924 6180
rect 12624 6400 12676 6452
rect 13636 6400 13688 6452
rect 14832 6400 14884 6452
rect 15292 6400 15344 6452
rect 15476 6400 15528 6452
rect 16304 6443 16356 6452
rect 16304 6409 16313 6443
rect 16313 6409 16347 6443
rect 16347 6409 16356 6443
rect 16304 6400 16356 6409
rect 16856 6400 16908 6452
rect 18144 6400 18196 6452
rect 18420 6400 18472 6452
rect 20812 6400 20864 6452
rect 21548 6400 21600 6452
rect 7012 6332 7064 6384
rect 7288 6332 7340 6384
rect 8576 6375 8628 6384
rect 5724 6307 5776 6316
rect 5724 6273 5733 6307
rect 5733 6273 5767 6307
rect 5767 6273 5776 6307
rect 5724 6264 5776 6273
rect 6828 6264 6880 6316
rect 7104 6264 7156 6316
rect 5816 6239 5868 6248
rect 5816 6205 5825 6239
rect 5825 6205 5859 6239
rect 5859 6205 5868 6239
rect 5816 6196 5868 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7472 6239 7524 6248
rect 7472 6205 7481 6239
rect 7481 6205 7515 6239
rect 7515 6205 7524 6239
rect 7472 6196 7524 6205
rect 4344 6128 4396 6180
rect 4804 6171 4856 6180
rect 4804 6137 4813 6171
rect 4813 6137 4847 6171
rect 4847 6137 4856 6171
rect 4804 6128 4856 6137
rect 5448 6128 5500 6180
rect 8576 6341 8585 6375
rect 8585 6341 8619 6375
rect 8619 6341 8628 6375
rect 8576 6332 8628 6341
rect 8760 6332 8812 6384
rect 11796 6332 11848 6384
rect 12808 6332 12860 6384
rect 18052 6332 18104 6384
rect 19340 6332 19392 6384
rect 19524 6332 19576 6384
rect 20720 6332 20772 6384
rect 9864 6307 9916 6316
rect 8024 6196 8076 6248
rect 8484 6239 8536 6248
rect 4528 6060 4580 6112
rect 4896 6060 4948 6112
rect 8024 6060 8076 6112
rect 8484 6205 8493 6239
rect 8493 6205 8527 6239
rect 8527 6205 8536 6239
rect 8484 6196 8536 6205
rect 8760 6128 8812 6180
rect 9864 6273 9873 6307
rect 9873 6273 9907 6307
rect 9907 6273 9916 6307
rect 9864 6264 9916 6273
rect 10876 6264 10928 6316
rect 14556 6264 14608 6316
rect 15292 6307 15344 6316
rect 15292 6273 15301 6307
rect 15301 6273 15335 6307
rect 15335 6273 15344 6307
rect 15292 6264 15344 6273
rect 9220 6196 9272 6248
rect 10692 6196 10744 6248
rect 11520 6196 11572 6248
rect 15660 6239 15712 6248
rect 15660 6205 15669 6239
rect 15669 6205 15703 6239
rect 15703 6205 15712 6239
rect 15660 6196 15712 6205
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 17132 6264 17184 6316
rect 20536 6264 20588 6316
rect 21364 6264 21416 6316
rect 9220 6103 9272 6112
rect 9220 6069 9229 6103
rect 9229 6069 9263 6103
rect 9263 6069 9272 6103
rect 9220 6060 9272 6069
rect 10324 6060 10376 6112
rect 10508 6103 10560 6112
rect 10508 6069 10517 6103
rect 10517 6069 10551 6103
rect 10551 6069 10560 6103
rect 10508 6060 10560 6069
rect 11060 6060 11112 6112
rect 11520 6103 11572 6112
rect 11520 6069 11529 6103
rect 11529 6069 11563 6103
rect 11563 6069 11572 6103
rect 11520 6060 11572 6069
rect 16396 6128 16448 6180
rect 14556 6060 14608 6112
rect 17500 6060 17552 6112
rect 17960 6128 18012 6180
rect 20720 6196 20772 6248
rect 21088 6196 21140 6248
rect 18420 6060 18472 6112
rect 18512 6060 18564 6112
rect 19984 6060 20036 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1584 5856 1636 5908
rect 3332 5856 3384 5908
rect 3792 5899 3844 5908
rect 3792 5865 3801 5899
rect 3801 5865 3835 5899
rect 3835 5865 3844 5899
rect 3792 5856 3844 5865
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4712 5899 4764 5908
rect 4712 5865 4721 5899
rect 4721 5865 4755 5899
rect 4755 5865 4764 5899
rect 4712 5856 4764 5865
rect 5540 5856 5592 5908
rect 7380 5856 7432 5908
rect 3240 5788 3292 5840
rect 7288 5788 7340 5840
rect 8116 5788 8168 5840
rect 9128 5788 9180 5840
rect 9588 5831 9640 5840
rect 9588 5797 9597 5831
rect 9597 5797 9631 5831
rect 9631 5797 9640 5831
rect 9588 5788 9640 5797
rect 10968 5788 11020 5840
rect 13084 5788 13136 5840
rect 13820 5788 13872 5840
rect 2780 5720 2832 5772
rect 3332 5763 3384 5772
rect 3332 5729 3341 5763
rect 3341 5729 3375 5763
rect 3375 5729 3384 5763
rect 3332 5720 3384 5729
rect 3516 5720 3568 5772
rect 2596 5652 2648 5704
rect 3148 5652 3200 5704
rect 4068 5652 4120 5704
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 6920 5720 6972 5772
rect 5080 5652 5132 5704
rect 5724 5652 5776 5704
rect 6736 5652 6788 5704
rect 9772 5720 9824 5772
rect 12164 5763 12216 5772
rect 12164 5729 12173 5763
rect 12173 5729 12207 5763
rect 12207 5729 12216 5763
rect 12164 5720 12216 5729
rect 8392 5695 8444 5704
rect 8392 5661 8401 5695
rect 8401 5661 8435 5695
rect 8435 5661 8444 5695
rect 8392 5652 8444 5661
rect 9404 5652 9456 5704
rect 11060 5652 11112 5704
rect 14464 5652 14516 5704
rect 15292 5856 15344 5908
rect 15660 5856 15712 5908
rect 17684 5856 17736 5908
rect 20904 5856 20956 5908
rect 16212 5788 16264 5840
rect 19708 5788 19760 5840
rect 20996 5788 21048 5840
rect 15568 5695 15620 5704
rect 3792 5584 3844 5636
rect 6184 5627 6236 5636
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2412 5559 2464 5568
rect 2044 5516 2096 5525
rect 2412 5525 2421 5559
rect 2421 5525 2455 5559
rect 2455 5525 2464 5559
rect 2412 5516 2464 5525
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 6184 5593 6193 5627
rect 6193 5593 6227 5627
rect 6227 5593 6236 5627
rect 6184 5584 6236 5593
rect 8944 5584 8996 5636
rect 10048 5584 10100 5636
rect 14372 5584 14424 5636
rect 15568 5661 15577 5695
rect 15577 5661 15611 5695
rect 15611 5661 15620 5695
rect 15568 5652 15620 5661
rect 17408 5652 17460 5704
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 18880 5695 18932 5704
rect 17132 5584 17184 5636
rect 17684 5584 17736 5636
rect 4436 5516 4488 5568
rect 4712 5516 4764 5568
rect 5356 5559 5408 5568
rect 5356 5525 5365 5559
rect 5365 5525 5399 5559
rect 5399 5525 5408 5559
rect 5356 5516 5408 5525
rect 5448 5516 5500 5568
rect 7380 5516 7432 5568
rect 8208 5559 8260 5568
rect 8208 5525 8217 5559
rect 8217 5525 8251 5559
rect 8251 5525 8260 5559
rect 8208 5516 8260 5525
rect 8760 5516 8812 5568
rect 10232 5516 10284 5568
rect 11704 5516 11756 5568
rect 12900 5516 12952 5568
rect 13636 5516 13688 5568
rect 14188 5559 14240 5568
rect 14188 5525 14197 5559
rect 14197 5525 14231 5559
rect 14231 5525 14240 5559
rect 14188 5516 14240 5525
rect 16856 5516 16908 5568
rect 17040 5516 17092 5568
rect 18512 5516 18564 5568
rect 18880 5661 18881 5695
rect 18881 5661 18915 5695
rect 18915 5661 18932 5695
rect 18880 5652 18932 5661
rect 20168 5652 20220 5704
rect 20720 5695 20772 5704
rect 20444 5627 20496 5636
rect 20444 5593 20462 5627
rect 20462 5593 20496 5627
rect 20444 5584 20496 5593
rect 20720 5661 20729 5695
rect 20729 5661 20763 5695
rect 20763 5661 20772 5695
rect 20720 5652 20772 5661
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 2044 5312 2096 5364
rect 4160 5312 4212 5364
rect 4896 5312 4948 5364
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 1492 5287 1544 5296
rect 1492 5253 1501 5287
rect 1501 5253 1535 5287
rect 1535 5253 1544 5287
rect 1492 5244 1544 5253
rect 2504 5244 2556 5296
rect 2780 5244 2832 5296
rect 3792 5244 3844 5296
rect 4528 5244 4580 5296
rect 6920 5312 6972 5364
rect 10968 5312 11020 5364
rect 11060 5312 11112 5364
rect 11796 5312 11848 5364
rect 14648 5312 14700 5364
rect 16764 5312 16816 5364
rect 2320 5151 2372 5160
rect 2320 5117 2329 5151
rect 2329 5117 2363 5151
rect 2363 5117 2372 5151
rect 2320 5108 2372 5117
rect 2228 5040 2280 5092
rect 4988 5176 5040 5228
rect 4620 5108 4672 5160
rect 5816 5244 5868 5296
rect 12348 5244 12400 5296
rect 6736 5176 6788 5228
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 7196 5176 7248 5228
rect 8116 5219 8168 5228
rect 8116 5185 8125 5219
rect 8125 5185 8159 5219
rect 8159 5185 8168 5219
rect 8116 5176 8168 5185
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8944 5176 8996 5228
rect 9404 5219 9456 5228
rect 9404 5185 9413 5219
rect 9413 5185 9447 5219
rect 9447 5185 9456 5219
rect 9404 5176 9456 5185
rect 10048 5176 10100 5228
rect 14188 5244 14240 5296
rect 14280 5244 14332 5296
rect 14648 5176 14700 5228
rect 3792 5040 3844 5092
rect 7748 5040 7800 5092
rect 8116 5040 8168 5092
rect 8576 5040 8628 5092
rect 9220 5040 9272 5092
rect 2964 5015 3016 5024
rect 2964 4981 2973 5015
rect 2973 4981 3007 5015
rect 3007 4981 3016 5015
rect 2964 4972 3016 4981
rect 4712 5015 4764 5024
rect 4712 4981 4721 5015
rect 4721 4981 4755 5015
rect 4755 4981 4764 5015
rect 4712 4972 4764 4981
rect 4896 4972 4948 5024
rect 7380 4972 7432 5024
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 12348 5108 12400 5160
rect 12624 5108 12676 5160
rect 15384 5176 15436 5228
rect 15752 5219 15804 5228
rect 15752 5185 15761 5219
rect 15761 5185 15795 5219
rect 15795 5185 15804 5219
rect 15752 5176 15804 5185
rect 16948 5176 17000 5228
rect 17132 5312 17184 5364
rect 17316 5312 17368 5364
rect 19708 5312 19760 5364
rect 19984 5355 20036 5364
rect 19984 5321 19993 5355
rect 19993 5321 20027 5355
rect 20027 5321 20036 5355
rect 19984 5312 20036 5321
rect 20352 5355 20404 5364
rect 20352 5321 20361 5355
rect 20361 5321 20395 5355
rect 20395 5321 20404 5355
rect 20352 5312 20404 5321
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 21456 5312 21508 5364
rect 18420 5244 18472 5296
rect 17592 5219 17644 5228
rect 17592 5185 17601 5219
rect 17601 5185 17635 5219
rect 17635 5185 17644 5219
rect 17592 5176 17644 5185
rect 17684 5176 17736 5228
rect 18880 5219 18932 5228
rect 18880 5185 18889 5219
rect 18889 5185 18923 5219
rect 18923 5185 18932 5219
rect 18880 5176 18932 5185
rect 10784 5015 10836 5024
rect 10784 4981 10793 5015
rect 10793 4981 10827 5015
rect 10827 4981 10836 5015
rect 10784 4972 10836 4981
rect 11336 4972 11388 5024
rect 11796 4972 11848 5024
rect 14280 5040 14332 5092
rect 18604 5108 18656 5160
rect 19708 5151 19760 5160
rect 19708 5117 19717 5151
rect 19717 5117 19751 5151
rect 19751 5117 19760 5151
rect 19708 5108 19760 5117
rect 20628 5108 20680 5160
rect 21180 5151 21232 5160
rect 21180 5117 21189 5151
rect 21189 5117 21223 5151
rect 21223 5117 21232 5151
rect 21180 5108 21232 5117
rect 20260 5040 20312 5092
rect 14924 4972 14976 5024
rect 15752 4972 15804 5024
rect 16028 4972 16080 5024
rect 16396 4972 16448 5024
rect 17408 4972 17460 5024
rect 17592 4972 17644 5024
rect 17960 4972 18012 5024
rect 18788 4972 18840 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 3240 4811 3292 4820
rect 3240 4777 3249 4811
rect 3249 4777 3283 4811
rect 3283 4777 3292 4811
rect 3240 4768 3292 4777
rect 5540 4768 5592 4820
rect 7104 4768 7156 4820
rect 7472 4768 7524 4820
rect 8116 4768 8168 4820
rect 8944 4768 8996 4820
rect 9404 4768 9456 4820
rect 10416 4811 10468 4820
rect 10416 4777 10425 4811
rect 10425 4777 10459 4811
rect 10459 4777 10468 4811
rect 10416 4768 10468 4777
rect 1952 4675 2004 4684
rect 1952 4641 1961 4675
rect 1961 4641 1995 4675
rect 1995 4641 2004 4675
rect 1952 4632 2004 4641
rect 3884 4700 3936 4752
rect 4712 4700 4764 4752
rect 3700 4632 3752 4684
rect 4620 4675 4672 4684
rect 4620 4641 4629 4675
rect 4629 4641 4663 4675
rect 4663 4641 4672 4675
rect 4620 4632 4672 4641
rect 5172 4632 5224 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 2412 4564 2464 4616
rect 3240 4564 3292 4616
rect 4896 4607 4948 4616
rect 4896 4573 4905 4607
rect 4905 4573 4939 4607
rect 4939 4573 4948 4607
rect 4896 4564 4948 4573
rect 6552 4632 6604 4684
rect 9588 4700 9640 4752
rect 14740 4768 14792 4820
rect 14924 4768 14976 4820
rect 15108 4811 15160 4820
rect 15108 4777 15117 4811
rect 15117 4777 15151 4811
rect 15151 4777 15160 4811
rect 15108 4768 15160 4777
rect 4804 4496 4856 4548
rect 1768 4428 1820 4480
rect 5172 4428 5224 4480
rect 6552 4496 6604 4548
rect 7564 4564 7616 4616
rect 8024 4564 8076 4616
rect 10600 4632 10652 4684
rect 11796 4675 11848 4684
rect 11796 4641 11805 4675
rect 11805 4641 11839 4675
rect 11839 4641 11848 4675
rect 11796 4632 11848 4641
rect 7840 4496 7892 4548
rect 5356 4428 5408 4480
rect 5632 4428 5684 4480
rect 6644 4471 6696 4480
rect 6644 4437 6653 4471
rect 6653 4437 6687 4471
rect 6687 4437 6696 4471
rect 6644 4428 6696 4437
rect 6736 4428 6788 4480
rect 8944 4428 8996 4480
rect 11704 4564 11756 4616
rect 15384 4632 15436 4684
rect 19708 4768 19760 4820
rect 20168 4768 20220 4820
rect 21088 4743 21140 4752
rect 21088 4709 21097 4743
rect 21097 4709 21131 4743
rect 21131 4709 21140 4743
rect 21088 4700 21140 4709
rect 10140 4496 10192 4548
rect 10692 4496 10744 4548
rect 16396 4564 16448 4616
rect 18512 4607 18564 4616
rect 15568 4496 15620 4548
rect 15936 4496 15988 4548
rect 9772 4428 9824 4480
rect 10876 4428 10928 4480
rect 13728 4428 13780 4480
rect 18144 4496 18196 4548
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 20720 4564 20772 4616
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 19892 4496 19944 4548
rect 21180 4496 21232 4548
rect 17316 4428 17368 4480
rect 18420 4428 18472 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 1584 4267 1636 4276
rect 1584 4233 1593 4267
rect 1593 4233 1627 4267
rect 1627 4233 1636 4267
rect 1584 4224 1636 4233
rect 2964 4224 3016 4276
rect 4620 4224 4672 4276
rect 3056 4156 3108 4208
rect 3516 4156 3568 4208
rect 4252 4156 4304 4208
rect 6552 4224 6604 4276
rect 6920 4224 6972 4276
rect 7564 4224 7616 4276
rect 7840 4267 7892 4276
rect 7840 4233 7849 4267
rect 7849 4233 7883 4267
rect 7883 4233 7892 4267
rect 7840 4224 7892 4233
rect 11244 4224 11296 4276
rect 11336 4224 11388 4276
rect 15752 4224 15804 4276
rect 18052 4224 18104 4276
rect 8944 4199 8996 4208
rect 8944 4165 8953 4199
rect 8953 4165 8987 4199
rect 8987 4165 8996 4199
rect 8944 4156 8996 4165
rect 10600 4156 10652 4208
rect 12164 4156 12216 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 2596 4088 2648 4140
rect 4712 4088 4764 4140
rect 4988 4088 5040 4140
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 5816 4131 5868 4140
rect 5816 4097 5825 4131
rect 5825 4097 5859 4131
rect 5859 4097 5868 4131
rect 5816 4088 5868 4097
rect 5908 4088 5960 4140
rect 2688 4020 2740 4072
rect 6184 4020 6236 4072
rect 4160 3952 4212 4004
rect 5080 3995 5132 4004
rect 5080 3961 5089 3995
rect 5089 3961 5123 3995
rect 5123 3961 5132 3995
rect 5080 3952 5132 3961
rect 5172 3952 5224 4004
rect 7656 4131 7708 4140
rect 7656 4097 7665 4131
rect 7665 4097 7699 4131
rect 7699 4097 7708 4131
rect 7656 4088 7708 4097
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 7104 4020 7156 4072
rect 12256 4131 12308 4140
rect 12256 4097 12265 4131
rect 12265 4097 12299 4131
rect 12299 4097 12308 4131
rect 12256 4088 12308 4097
rect 13728 4131 13780 4140
rect 8852 4063 8904 4072
rect 4344 3884 4396 3936
rect 5540 3927 5592 3936
rect 5540 3893 5549 3927
rect 5549 3893 5583 3927
rect 5583 3893 5592 3927
rect 5540 3884 5592 3893
rect 7288 3952 7340 4004
rect 8852 4029 8861 4063
rect 8861 4029 8895 4063
rect 8895 4029 8904 4063
rect 8852 4020 8904 4029
rect 8944 4020 8996 4072
rect 9312 3995 9364 4004
rect 9312 3961 9321 3995
rect 9321 3961 9355 3995
rect 9355 3961 9364 3995
rect 9312 3952 9364 3961
rect 9772 3995 9824 4004
rect 9772 3961 9781 3995
rect 9781 3961 9815 3995
rect 9815 3961 9824 3995
rect 9772 3952 9824 3961
rect 7104 3884 7156 3936
rect 7748 3884 7800 3936
rect 8116 3927 8168 3936
rect 8116 3893 8125 3927
rect 8125 3893 8159 3927
rect 8159 3893 8168 3927
rect 8116 3884 8168 3893
rect 8852 3884 8904 3936
rect 9404 3884 9456 3936
rect 9588 3884 9640 3936
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 11796 4020 11848 4072
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 15200 4156 15252 4208
rect 15384 4156 15436 4208
rect 15292 4131 15344 4140
rect 15292 4097 15310 4131
rect 15310 4097 15344 4131
rect 15568 4131 15620 4140
rect 15292 4088 15344 4097
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16672 4131 16724 4140
rect 14280 4020 14332 4072
rect 13912 3995 13964 4004
rect 11888 3884 11940 3936
rect 12992 3927 13044 3936
rect 12992 3893 13001 3927
rect 13001 3893 13035 3927
rect 13035 3893 13044 3927
rect 12992 3884 13044 3893
rect 13544 3884 13596 3936
rect 13912 3961 13921 3995
rect 13921 3961 13955 3995
rect 13955 3961 13964 3995
rect 13912 3952 13964 3961
rect 14372 3952 14424 4004
rect 14280 3884 14332 3936
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 17500 4088 17552 4140
rect 18144 4131 18196 4140
rect 18144 4097 18153 4131
rect 18153 4097 18187 4131
rect 18187 4097 18196 4131
rect 18144 4088 18196 4097
rect 17776 4063 17828 4072
rect 17776 4029 17785 4063
rect 17785 4029 17819 4063
rect 17819 4029 17828 4063
rect 17776 4020 17828 4029
rect 15936 3952 15988 4004
rect 16304 3884 16356 3936
rect 17868 3952 17920 4004
rect 19340 4088 19392 4140
rect 19800 4156 19852 4208
rect 20720 4199 20772 4208
rect 20720 4165 20729 4199
rect 20729 4165 20763 4199
rect 20763 4165 20772 4199
rect 20720 4156 20772 4165
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 20812 4131 20864 4140
rect 20812 4097 20821 4131
rect 20821 4097 20855 4131
rect 20855 4097 20864 4131
rect 20812 4088 20864 4097
rect 20536 4020 20588 4072
rect 18604 3884 18656 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2504 3680 2556 3732
rect 4804 3680 4856 3732
rect 13636 3680 13688 3732
rect 14280 3680 14332 3732
rect 14372 3723 14424 3732
rect 14372 3689 14381 3723
rect 14381 3689 14415 3723
rect 14415 3689 14424 3723
rect 14372 3680 14424 3689
rect 16672 3680 16724 3732
rect 17224 3680 17276 3732
rect 18144 3680 18196 3732
rect 19616 3723 19668 3732
rect 2320 3544 2372 3596
rect 3056 3476 3108 3528
rect 5080 3612 5132 3664
rect 5540 3612 5592 3664
rect 10692 3655 10744 3664
rect 10692 3621 10701 3655
rect 10701 3621 10735 3655
rect 10735 3621 10744 3655
rect 10692 3612 10744 3621
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 4528 3587 4580 3596
rect 4528 3553 4537 3587
rect 4537 3553 4571 3587
rect 4571 3553 4580 3587
rect 4528 3544 4580 3553
rect 4712 3544 4764 3596
rect 5816 3544 5868 3596
rect 6000 3544 6052 3596
rect 4160 3476 4212 3528
rect 6552 3476 6604 3528
rect 6736 3476 6788 3528
rect 8208 3544 8260 3596
rect 8760 3544 8812 3596
rect 9404 3587 9456 3596
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8668 3476 8720 3528
rect 9128 3476 9180 3528
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 9588 3544 9640 3596
rect 8024 3408 8076 3460
rect 3884 3340 3936 3392
rect 4436 3340 4488 3392
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5356 3383 5408 3392
rect 5356 3349 5365 3383
rect 5365 3349 5399 3383
rect 5399 3349 5408 3383
rect 5356 3340 5408 3349
rect 5632 3340 5684 3392
rect 5908 3340 5960 3392
rect 6000 3340 6052 3392
rect 6736 3383 6788 3392
rect 6736 3349 6745 3383
rect 6745 3349 6779 3383
rect 6779 3349 6788 3383
rect 6736 3340 6788 3349
rect 7288 3340 7340 3392
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 8484 3340 8536 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 10508 3340 10560 3392
rect 12440 3544 12492 3596
rect 12992 3612 13044 3664
rect 13820 3544 13872 3596
rect 15016 3587 15068 3596
rect 15016 3553 15025 3587
rect 15025 3553 15059 3587
rect 15059 3553 15068 3587
rect 15016 3544 15068 3553
rect 10968 3476 11020 3528
rect 12900 3476 12952 3528
rect 13452 3476 13504 3528
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 15384 3519 15436 3528
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15476 3476 15528 3528
rect 16396 3544 16448 3596
rect 17132 3544 17184 3596
rect 18604 3544 18656 3596
rect 18880 3544 18932 3596
rect 19064 3476 19116 3528
rect 19616 3689 19625 3723
rect 19625 3689 19659 3723
rect 19659 3689 19668 3723
rect 19616 3680 19668 3689
rect 20628 3723 20680 3732
rect 20628 3689 20637 3723
rect 20637 3689 20671 3723
rect 20671 3689 20680 3723
rect 20628 3680 20680 3689
rect 19708 3612 19760 3664
rect 19248 3544 19300 3596
rect 19800 3476 19852 3528
rect 20536 3544 20588 3596
rect 21456 3476 21508 3528
rect 11980 3408 12032 3460
rect 12164 3408 12216 3460
rect 17776 3340 17828 3392
rect 18328 3408 18380 3460
rect 18972 3408 19024 3460
rect 19984 3383 20036 3392
rect 19984 3349 19993 3383
rect 19993 3349 20027 3383
rect 20027 3349 20036 3383
rect 19984 3340 20036 3349
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 1124 3136 1176 3188
rect 2596 3136 2648 3188
rect 2780 3179 2832 3188
rect 2780 3145 2789 3179
rect 2789 3145 2823 3179
rect 2823 3145 2832 3179
rect 2780 3136 2832 3145
rect 940 3068 992 3120
rect 3884 3136 3936 3188
rect 4252 3179 4304 3188
rect 4252 3145 4261 3179
rect 4261 3145 4295 3179
rect 4295 3145 4304 3179
rect 4252 3136 4304 3145
rect 8668 3136 8720 3188
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 16948 3136 17000 3188
rect 17776 3136 17828 3188
rect 19524 3136 19576 3188
rect 2136 3000 2188 3052
rect 2596 3043 2648 3052
rect 2596 3009 2605 3043
rect 2605 3009 2639 3043
rect 2639 3009 2648 3043
rect 2596 3000 2648 3009
rect 6000 3068 6052 3120
rect 20 2932 72 2984
rect 940 2932 992 2984
rect 2320 2864 2372 2916
rect 4252 3000 4304 3052
rect 4436 3000 4488 3052
rect 6644 3000 6696 3052
rect 7380 3043 7432 3052
rect 5448 2932 5500 2984
rect 6552 2932 6604 2984
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 8208 3000 8260 3052
rect 9496 3068 9548 3120
rect 9772 3068 9824 3120
rect 11336 3068 11388 3120
rect 12348 3068 12400 3120
rect 9220 3043 9272 3052
rect 7104 2932 7156 2984
rect 5540 2864 5592 2916
rect 8300 2932 8352 2984
rect 8392 2932 8444 2984
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 10600 3000 10652 3052
rect 9956 2932 10008 2984
rect 12624 3043 12676 3052
rect 14096 3068 14148 3120
rect 18052 3111 18104 3120
rect 12624 3009 12642 3043
rect 12642 3009 12676 3043
rect 12624 3000 12676 3009
rect 1032 2796 1084 2848
rect 4068 2796 4120 2848
rect 4528 2796 4580 2848
rect 4988 2796 5040 2848
rect 5908 2796 5960 2848
rect 6368 2839 6420 2848
rect 6368 2805 6377 2839
rect 6377 2805 6411 2839
rect 6411 2805 6420 2839
rect 6368 2796 6420 2805
rect 6920 2796 6972 2848
rect 7380 2796 7432 2848
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 8024 2839 8076 2848
rect 8024 2805 8033 2839
rect 8033 2805 8067 2839
rect 8067 2805 8076 2839
rect 8024 2796 8076 2805
rect 8300 2839 8352 2848
rect 8300 2805 8309 2839
rect 8309 2805 8343 2839
rect 8343 2805 8352 2839
rect 8300 2796 8352 2805
rect 8576 2796 8628 2848
rect 9588 2796 9640 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 14648 3000 14700 3052
rect 18052 3077 18061 3111
rect 18061 3077 18095 3111
rect 18095 3077 18104 3111
rect 18052 3068 18104 3077
rect 18144 3111 18196 3120
rect 18144 3077 18153 3111
rect 18153 3077 18187 3111
rect 18187 3077 18196 3111
rect 18144 3068 18196 3077
rect 19248 3068 19300 3120
rect 19340 3068 19392 3120
rect 20076 3068 20128 3120
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13452 2975 13504 2984
rect 13268 2932 13320 2941
rect 13452 2941 13461 2975
rect 13461 2941 13495 2975
rect 13495 2941 13504 2975
rect 13452 2932 13504 2941
rect 13636 2932 13688 2984
rect 17500 3000 17552 3052
rect 19984 3000 20036 3052
rect 20168 3043 20220 3052
rect 20168 3009 20177 3043
rect 20177 3009 20211 3043
rect 20211 3009 20220 3043
rect 20168 3000 20220 3009
rect 20628 3000 20680 3052
rect 17316 2975 17368 2984
rect 13268 2796 13320 2848
rect 14280 2864 14332 2916
rect 14740 2864 14792 2916
rect 15108 2864 15160 2916
rect 17316 2941 17325 2975
rect 17325 2941 17359 2975
rect 17359 2941 17368 2975
rect 17316 2932 17368 2941
rect 18236 2975 18288 2984
rect 18236 2941 18245 2975
rect 18245 2941 18279 2975
rect 18279 2941 18288 2975
rect 18236 2932 18288 2941
rect 19248 2932 19300 2984
rect 19892 2932 19944 2984
rect 17960 2796 18012 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3424 2592 3476 2644
rect 4252 2592 4304 2644
rect 4620 2592 4672 2644
rect 5356 2592 5408 2644
rect 8944 2592 8996 2644
rect 11060 2592 11112 2644
rect 11336 2592 11388 2644
rect 13452 2592 13504 2644
rect 14372 2592 14424 2644
rect 16028 2592 16080 2644
rect 2596 2524 2648 2576
rect 9312 2524 9364 2576
rect 9772 2567 9824 2576
rect 9772 2533 9781 2567
rect 9781 2533 9815 2567
rect 9815 2533 9824 2567
rect 9772 2524 9824 2533
rect 4528 2456 4580 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 5448 2456 5500 2465
rect 7104 2456 7156 2508
rect 8208 2456 8260 2508
rect 9588 2456 9640 2508
rect 11980 2499 12032 2508
rect 11980 2465 11989 2499
rect 11989 2465 12023 2499
rect 12023 2465 12032 2499
rect 11980 2456 12032 2465
rect 1308 2388 1360 2440
rect 756 2320 808 2372
rect 2228 2363 2280 2372
rect 2228 2329 2237 2363
rect 2237 2329 2271 2363
rect 2271 2329 2280 2363
rect 2228 2320 2280 2329
rect 2780 2431 2832 2440
rect 2780 2397 2789 2431
rect 2789 2397 2823 2431
rect 2823 2397 2832 2431
rect 2780 2388 2832 2397
rect 3700 2320 3752 2372
rect 4160 2252 4212 2304
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 7656 2431 7708 2440
rect 7012 2320 7064 2372
rect 7656 2397 7665 2431
rect 7665 2397 7699 2431
rect 7699 2397 7708 2431
rect 7656 2388 7708 2397
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9680 2388 9732 2440
rect 10324 2431 10376 2440
rect 10324 2397 10333 2431
rect 10333 2397 10367 2431
rect 10367 2397 10376 2431
rect 10324 2388 10376 2397
rect 10600 2431 10652 2440
rect 10600 2397 10609 2431
rect 10609 2397 10643 2431
rect 10643 2397 10652 2431
rect 10600 2388 10652 2397
rect 11796 2388 11848 2440
rect 12256 2388 12308 2440
rect 6644 2252 6696 2304
rect 8392 2295 8444 2304
rect 8392 2261 8401 2295
rect 8401 2261 8435 2295
rect 8435 2261 8444 2295
rect 8392 2252 8444 2261
rect 8668 2320 8720 2372
rect 9864 2320 9916 2372
rect 15476 2524 15528 2576
rect 13084 2499 13136 2508
rect 13084 2465 13093 2499
rect 13093 2465 13127 2499
rect 13127 2465 13136 2499
rect 13084 2456 13136 2465
rect 13360 2456 13412 2508
rect 13636 2456 13688 2508
rect 15016 2456 15068 2508
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 14924 2388 14976 2440
rect 15200 2431 15252 2440
rect 15200 2397 15209 2431
rect 15209 2397 15243 2431
rect 15243 2397 15252 2431
rect 15200 2388 15252 2397
rect 16304 2456 16356 2508
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 17960 2592 18012 2644
rect 18144 2456 18196 2508
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 20352 2431 20404 2440
rect 20352 2397 20361 2431
rect 20361 2397 20395 2431
rect 20395 2397 20404 2431
rect 20352 2388 20404 2397
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 8852 2252 8904 2304
rect 8944 2252 8996 2304
rect 11796 2252 11848 2304
rect 11888 2252 11940 2304
rect 16212 2320 16264 2372
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 13912 2252 13964 2304
rect 14832 2295 14884 2304
rect 14832 2261 14841 2295
rect 14841 2261 14875 2295
rect 14875 2261 14884 2295
rect 14832 2252 14884 2261
rect 15844 2252 15896 2304
rect 18052 2320 18104 2372
rect 18512 2295 18564 2304
rect 18512 2261 18521 2295
rect 18521 2261 18555 2295
rect 18555 2261 18564 2295
rect 18512 2252 18564 2261
rect 19432 2295 19484 2304
rect 19432 2261 19441 2295
rect 19441 2261 19475 2295
rect 19475 2261 19484 2295
rect 19432 2252 19484 2261
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 3976 2048 4028 2100
rect 7196 2048 7248 2100
rect 8576 2048 8628 2100
rect 11060 2048 11112 2100
rect 12072 2048 12124 2100
rect 7564 1980 7616 2032
rect 848 1912 900 1964
rect 8392 1912 8444 1964
rect 9312 1980 9364 2032
rect 11888 1980 11940 2032
rect 14648 2048 14700 2100
rect 17040 2048 17092 2100
rect 19432 2048 19484 2100
rect 2964 1844 3016 1896
rect 6552 1844 6604 1896
rect 7288 1844 7340 1896
rect 14096 1980 14148 2032
rect 17316 1980 17368 2032
rect 19984 1980 20036 2032
rect 12900 1912 12952 1964
rect 14832 1912 14884 1964
rect 17408 1912 17460 1964
rect 19800 1912 19852 1964
rect 13820 1844 13872 1896
rect 14924 1844 14976 1896
rect 17592 1844 17644 1896
rect 20352 1844 20404 1896
rect 10508 1776 10560 1828
rect 17224 1776 17276 1828
rect 7840 1708 7892 1760
rect 15200 1708 15252 1760
rect 16580 1708 16632 1760
rect 18512 1708 18564 1760
rect 8852 1640 8904 1692
rect 11152 1640 11204 1692
rect 14556 1640 14608 1692
rect 18236 1640 18288 1692
rect 9680 1572 9732 1624
rect 11244 1572 11296 1624
rect 12624 1572 12676 1624
rect 16396 1572 16448 1624
rect 9864 1504 9916 1556
rect 10692 1504 10744 1556
rect 14464 1504 14516 1556
rect 17960 1504 18012 1556
rect 12532 1368 12584 1420
rect 13912 1368 13964 1420
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 2962 21312 3018 21321
rect 2962 21247 3018 21256
rect 1950 20904 2006 20913
rect 1950 20839 2006 20848
rect 1306 20360 1362 20369
rect 1306 20295 1362 20304
rect 1122 19816 1178 19825
rect 1122 19751 1178 19760
rect 938 19544 994 19553
rect 768 19502 938 19530
rect 20 14544 72 14550
rect 20 14486 72 14492
rect 32 2990 60 14486
rect 20 2984 72 2990
rect 20 2926 72 2932
rect 768 2378 796 19502
rect 938 19479 994 19488
rect 1032 18352 1084 18358
rect 1032 18294 1084 18300
rect 938 17776 994 17785
rect 938 17711 994 17720
rect 848 15632 900 15638
rect 848 15574 900 15580
rect 756 2372 808 2378
rect 756 2314 808 2320
rect 860 1970 888 15574
rect 952 3126 980 17711
rect 940 3120 992 3126
rect 940 3062 992 3068
rect 940 2984 992 2990
rect 938 2952 940 2961
rect 992 2952 994 2961
rect 938 2887 994 2896
rect 1044 2854 1072 18294
rect 1136 3194 1164 19751
rect 1216 19236 1268 19242
rect 1216 19178 1268 19184
rect 1228 12306 1256 19178
rect 1216 12300 1268 12306
rect 1216 12242 1268 12248
rect 1124 3188 1176 3194
rect 1124 3130 1176 3136
rect 1032 2848 1084 2854
rect 1032 2790 1084 2796
rect 1320 2446 1348 20295
rect 1492 20256 1544 20262
rect 1492 20198 1544 20204
rect 1504 20097 1532 20198
rect 1490 20088 1546 20097
rect 1964 20058 1992 20839
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2056 20505 2084 20538
rect 2042 20496 2098 20505
rect 2976 20466 3004 21247
rect 5262 20496 5318 20505
rect 2042 20431 2098 20440
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 2964 20460 3016 20466
rect 5736 20466 5764 22200
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 17236 20602 17264 22200
rect 18694 21312 18750 21321
rect 18694 21247 18750 21256
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 16854 20496 16910 20505
rect 5262 20431 5318 20440
rect 5724 20460 5776 20466
rect 2964 20402 3016 20408
rect 1490 20023 1546 20032
rect 1952 20052 2004 20058
rect 1952 19994 2004 20000
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 2148 19446 2176 20402
rect 4068 20392 4120 20398
rect 4528 20392 4580 20398
rect 4068 20334 4120 20340
rect 4526 20360 4528 20369
rect 4580 20360 4582 20369
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2240 19514 2268 19790
rect 2686 19544 2742 19553
rect 2228 19508 2280 19514
rect 2686 19479 2742 19488
rect 2228 19450 2280 19456
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2700 19378 2728 19479
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 2228 19372 2280 19378
rect 2228 19314 2280 19320
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1688 18290 1716 18566
rect 1964 18426 1992 19314
rect 2042 19272 2098 19281
rect 2042 19207 2044 19216
rect 2096 19207 2098 19216
rect 2044 19178 2096 19184
rect 2240 18970 2268 19314
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2504 18964 2556 18970
rect 2504 18906 2556 18912
rect 2044 18760 2096 18766
rect 2044 18702 2096 18708
rect 1952 18420 2004 18426
rect 1952 18362 2004 18368
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1584 18148 1636 18154
rect 1584 18090 1636 18096
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1490 16759 1546 16768
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1398 16008 1454 16017
rect 1398 15943 1400 15952
rect 1452 15943 1454 15952
rect 1400 15914 1452 15920
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 10266 1440 15438
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14385 1532 14758
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 13569 1532 14214
rect 1490 13560 1546 13569
rect 1490 13495 1546 13504
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1504 7585 1532 11591
rect 1596 9042 1624 18090
rect 2056 17882 2084 18702
rect 2516 18290 2544 18906
rect 2504 18284 2556 18290
rect 2504 18226 2556 18232
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 2872 18216 2924 18222
rect 2872 18158 2924 18164
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 2148 17678 2176 18022
rect 2136 17672 2188 17678
rect 2042 17640 2098 17649
rect 2136 17614 2188 17620
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2042 17575 2098 17584
rect 2056 17542 2084 17575
rect 2044 17536 2096 17542
rect 2044 17478 2096 17484
rect 2240 17338 2268 17614
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 2320 17196 2372 17202
rect 2320 17138 2372 17144
rect 1688 16250 1716 17138
rect 2136 16788 2188 16794
rect 2136 16730 2188 16736
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 1676 16244 1728 16250
rect 1676 16186 1728 16192
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1688 14890 1716 16050
rect 1952 15360 2004 15366
rect 1952 15302 2004 15308
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1676 14544 1728 14550
rect 1674 14512 1676 14521
rect 1728 14512 1730 14521
rect 1674 14447 1730 14456
rect 1964 14414 1992 15302
rect 2056 15026 2084 16390
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 2148 14906 2176 16730
rect 2228 16448 2280 16454
rect 2228 16390 2280 16396
rect 2240 16114 2268 16390
rect 2228 16108 2280 16114
rect 2228 16050 2280 16056
rect 2056 14878 2176 14906
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13326 1716 13670
rect 1766 13424 1822 13433
rect 1766 13359 1822 13368
rect 1860 13388 1912 13394
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 1688 10130 1716 13126
rect 1780 10674 1808 13359
rect 1860 13330 1912 13336
rect 1872 12209 1900 13330
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1858 12200 1914 12209
rect 1858 12135 1914 12144
rect 1964 11914 1992 13126
rect 2056 12850 2084 14878
rect 2136 14816 2188 14822
rect 2134 14784 2136 14793
rect 2188 14784 2190 14793
rect 2134 14719 2190 14728
rect 2136 14272 2188 14278
rect 2136 14214 2188 14220
rect 2148 13977 2176 14214
rect 2332 14090 2360 17138
rect 2884 17134 2912 18158
rect 3068 17882 3096 18226
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3160 17338 3188 20198
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3896 19553 3924 19654
rect 4080 19553 4108 20334
rect 4526 20295 4582 20304
rect 4712 19848 4764 19854
rect 4526 19816 4582 19825
rect 4712 19790 4764 19796
rect 4526 19751 4528 19760
rect 4580 19751 4582 19760
rect 4528 19722 4580 19728
rect 4252 19712 4304 19718
rect 4252 19654 4304 19660
rect 3698 19544 3754 19553
rect 3698 19479 3700 19488
rect 3752 19479 3754 19488
rect 3882 19544 3938 19553
rect 3882 19479 3938 19488
rect 4066 19544 4122 19553
rect 4066 19479 4122 19488
rect 3700 19450 3752 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 19174 3556 19314
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 4172 19174 4200 19246
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4160 19168 4212 19174
rect 4160 19110 4212 19116
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3240 18284 3292 18290
rect 3240 18226 3292 18232
rect 3252 17746 3280 18226
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3240 17740 3292 17746
rect 3240 17682 3292 17688
rect 3148 17332 3200 17338
rect 3148 17274 3200 17280
rect 2964 17264 3016 17270
rect 2964 17206 3016 17212
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2424 16590 2452 16934
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16250 2912 16526
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 15972 2832 15978
rect 2780 15914 2832 15920
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2240 14062 2360 14090
rect 2134 13968 2190 13977
rect 2134 13903 2190 13912
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 12844 2096 12850
rect 2044 12786 2096 12792
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1872 11886 1992 11914
rect 1872 11354 1900 11886
rect 1950 11792 2006 11801
rect 1950 11727 1952 11736
rect 2004 11727 2006 11736
rect 1952 11698 2004 11704
rect 1952 11620 2004 11626
rect 1952 11562 2004 11568
rect 1860 11348 1912 11354
rect 1860 11290 1912 11296
rect 1964 11286 1992 11562
rect 1952 11280 2004 11286
rect 1952 11222 2004 11228
rect 2056 11150 2084 12038
rect 2148 11762 2176 13806
rect 2240 13462 2268 14062
rect 2320 14000 2372 14006
rect 2320 13942 2372 13948
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12345 2268 12718
rect 2226 12336 2282 12345
rect 2226 12271 2282 12280
rect 2228 12232 2280 12238
rect 2228 12174 2280 12180
rect 2240 11937 2268 12174
rect 2226 11928 2282 11937
rect 2226 11863 2282 11872
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11529 2268 11630
rect 2226 11520 2282 11529
rect 2226 11455 2282 11464
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 2136 10736 2188 10742
rect 2136 10678 2188 10684
rect 1768 10668 1820 10674
rect 1768 10610 1820 10616
rect 1676 10124 1728 10130
rect 1676 10066 1728 10072
rect 1950 9616 2006 9625
rect 1950 9551 2006 9560
rect 2044 9580 2096 9586
rect 1584 9036 1636 9042
rect 1584 8978 1636 8984
rect 1768 8900 1820 8906
rect 1768 8842 1820 8848
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1490 7576 1546 7585
rect 1596 7546 1624 8502
rect 1676 7948 1728 7954
rect 1780 7936 1808 8842
rect 1964 8498 1992 9551
rect 2044 9522 2096 9528
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2056 8378 2084 9522
rect 2148 8974 2176 10678
rect 2240 10577 2268 11154
rect 2226 10568 2282 10577
rect 2226 10503 2282 10512
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2240 9897 2268 9998
rect 2226 9888 2282 9897
rect 2226 9823 2282 9832
rect 2226 9616 2282 9625
rect 2226 9551 2228 9560
rect 2280 9551 2282 9560
rect 2228 9522 2280 9528
rect 2226 9480 2282 9489
rect 2226 9415 2282 9424
rect 2240 9110 2268 9415
rect 2228 9104 2280 9110
rect 2228 9046 2280 9052
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2148 8673 2176 8910
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2134 8664 2190 8673
rect 2134 8599 2190 8608
rect 2240 8430 2268 8774
rect 2332 8634 2360 13942
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2424 10810 2452 13874
rect 2516 12850 2544 14214
rect 2608 13530 2636 15438
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2700 15026 2728 15302
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2700 14929 2728 14962
rect 2686 14920 2742 14929
rect 2686 14855 2742 14864
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2700 13410 2728 13874
rect 2608 13382 2728 13410
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2516 11218 2544 12242
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 9722 2452 10542
rect 2516 10538 2544 11154
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2412 9580 2464 9586
rect 2412 9522 2464 9528
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1728 7908 1808 7936
rect 1676 7890 1728 7896
rect 1490 7511 1546 7520
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1490 7440 1546 7449
rect 1490 7375 1492 7384
rect 1544 7375 1546 7384
rect 1492 7346 1544 7352
rect 1490 7032 1546 7041
rect 1490 6967 1546 6976
rect 1504 6798 1532 6967
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1780 6254 1808 7908
rect 1964 8350 2084 8378
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 1860 7744 1912 7750
rect 1858 7712 1860 7721
rect 1912 7712 1914 7721
rect 1858 7647 1914 7656
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1490 5536 1546 5545
rect 1490 5471 1546 5480
rect 1504 5302 1532 5471
rect 1492 5296 1544 5302
rect 1492 5238 1544 5244
rect 1398 4992 1454 5001
rect 1398 4927 1454 4936
rect 1412 4146 1440 4927
rect 1596 4282 1624 5850
rect 1780 4486 1808 6190
rect 1964 4690 1992 8350
rect 2240 8265 2268 8366
rect 2226 8256 2282 8265
rect 2226 8191 2282 8200
rect 2136 7812 2188 7818
rect 2136 7754 2188 7760
rect 2148 7002 2176 7754
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2240 7002 2268 7278
rect 2136 6996 2188 7002
rect 2136 6938 2188 6944
rect 2228 6996 2280 7002
rect 2228 6938 2280 6944
rect 2424 6882 2452 9522
rect 2516 7546 2544 9862
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2504 6996 2556 7002
rect 2504 6938 2556 6944
rect 2148 6854 2452 6882
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2056 5370 2084 5510
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1584 4276 1636 4282
rect 1584 4218 1636 4224
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 2148 3058 2176 6854
rect 2318 5672 2374 5681
rect 2318 5607 2374 5616
rect 2332 5166 2360 5607
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2320 5160 2372 5166
rect 2226 5128 2282 5137
rect 2320 5102 2372 5108
rect 2226 5063 2228 5072
rect 2280 5063 2282 5072
rect 2228 5034 2280 5040
rect 2228 4616 2280 4622
rect 2226 4584 2228 4593
rect 2280 4584 2282 4593
rect 2226 4519 2282 4528
rect 2332 3602 2360 5102
rect 2424 4622 2452 5510
rect 2516 5302 2544 6938
rect 2608 6458 2636 13382
rect 2688 13320 2740 13326
rect 2688 13262 2740 13268
rect 2700 12986 2728 13262
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2792 12322 2820 15914
rect 2872 13184 2924 13190
rect 2870 13152 2872 13161
rect 2924 13152 2926 13161
rect 2870 13087 2926 13096
rect 2976 12481 3004 17206
rect 3056 16992 3108 16998
rect 3056 16934 3108 16940
rect 3068 16590 3096 16934
rect 3056 16584 3108 16590
rect 3436 16561 3464 18090
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16827 3857 16836
rect 3056 16526 3108 16532
rect 3422 16552 3478 16561
rect 3422 16487 3478 16496
rect 3436 15570 3464 16487
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3424 15564 3476 15570
rect 3424 15506 3476 15512
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 2962 12472 3018 12481
rect 2962 12407 3018 12416
rect 2700 12294 2820 12322
rect 2964 12368 3016 12374
rect 2964 12310 3016 12316
rect 2700 11914 2728 12294
rect 2872 12096 2924 12102
rect 2872 12038 2924 12044
rect 2700 11886 2820 11914
rect 2792 10826 2820 11886
rect 2700 10810 2820 10826
rect 2688 10804 2820 10810
rect 2740 10798 2820 10804
rect 2688 10746 2740 10752
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2688 10532 2740 10538
rect 2688 10474 2740 10480
rect 2700 8430 2728 10474
rect 2792 10305 2820 10610
rect 2778 10296 2834 10305
rect 2778 10231 2834 10240
rect 2778 10160 2834 10169
rect 2778 10095 2834 10104
rect 2792 9926 2820 10095
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2792 9178 2820 9386
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 8616 2912 12038
rect 2976 11150 3004 12310
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2976 10713 3004 11086
rect 2962 10704 3018 10713
rect 2962 10639 3018 10648
rect 2964 10464 3016 10470
rect 2964 10406 3016 10412
rect 2976 8634 3004 10406
rect 3068 10062 3096 15302
rect 3804 15201 3832 15302
rect 3790 15192 3846 15201
rect 3790 15127 3846 15136
rect 3332 14884 3384 14890
rect 3332 14826 3384 14832
rect 3240 14544 3292 14550
rect 3240 14486 3292 14492
rect 3148 14340 3200 14346
rect 3148 14282 3200 14288
rect 3160 14074 3188 14282
rect 3148 14068 3200 14074
rect 3148 14010 3200 14016
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13326 3188 13670
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3160 12753 3188 13262
rect 3146 12744 3202 12753
rect 3146 12679 3202 12688
rect 3252 12238 3280 14486
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3068 9654 3096 9862
rect 3056 9648 3108 9654
rect 3056 9590 3108 9596
rect 3056 9512 3108 9518
rect 3056 9454 3108 9460
rect 3068 8906 3096 9454
rect 3160 9081 3188 12038
rect 3240 11620 3292 11626
rect 3240 11562 3292 11568
rect 3252 11150 3280 11562
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3252 10169 3280 10950
rect 3344 10198 3372 14826
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3424 14272 3476 14278
rect 3424 14214 3476 14220
rect 3436 12102 3464 14214
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3896 12442 3924 18566
rect 4080 18290 4108 19110
rect 4172 18834 4200 19110
rect 4160 18828 4212 18834
rect 4160 18770 4212 18776
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 3976 18216 4028 18222
rect 3976 18158 4028 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 3988 17746 4016 18158
rect 4068 18148 4120 18154
rect 4068 18090 4120 18096
rect 4080 17882 4108 18090
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 4172 17338 4200 18158
rect 4264 17785 4292 19654
rect 4724 19514 4752 19790
rect 4896 19712 4948 19718
rect 4894 19680 4896 19689
rect 4948 19680 4950 19689
rect 4894 19615 4950 19624
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 5172 19508 5224 19514
rect 5172 19450 5224 19456
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4988 19304 5040 19310
rect 4988 19246 5040 19252
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4250 17776 4306 17785
rect 4250 17711 4306 17720
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 3976 17332 4028 17338
rect 3976 17274 4028 17280
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3988 14550 4016 17274
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 4080 16046 4108 17070
rect 4264 16697 4292 17478
rect 4434 17096 4490 17105
rect 4434 17031 4490 17040
rect 4448 16726 4476 17031
rect 4344 16720 4396 16726
rect 4250 16688 4306 16697
rect 4344 16662 4396 16668
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4250 16623 4306 16632
rect 4160 16516 4212 16522
rect 4160 16458 4212 16464
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 4172 15910 4200 16458
rect 4068 15904 4120 15910
rect 4068 15846 4120 15852
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 3976 14544 4028 14550
rect 3976 14486 4028 14492
rect 3976 14408 4028 14414
rect 3976 14350 4028 14356
rect 3988 14074 4016 14350
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4080 14006 4108 15846
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4172 13274 4200 14418
rect 4264 14414 4292 15098
rect 4252 14408 4304 14414
rect 4252 14350 4304 14356
rect 4080 13246 4200 13274
rect 4080 12918 4108 13246
rect 4160 13184 4212 13190
rect 4160 13126 4212 13132
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4068 12912 4120 12918
rect 4172 12889 4200 13126
rect 4264 12986 4292 13126
rect 4252 12980 4304 12986
rect 4252 12922 4304 12928
rect 4068 12854 4120 12860
rect 4158 12880 4214 12889
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3882 12336 3938 12345
rect 3882 12271 3938 12280
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3528 11898 3556 12038
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3792 11144 3844 11150
rect 3790 11112 3792 11121
rect 3844 11112 3846 11121
rect 3790 11047 3846 11056
rect 3896 10810 3924 12271
rect 3988 11830 4016 12718
rect 4080 12322 4108 12854
rect 4158 12815 4214 12824
rect 4252 12640 4304 12646
rect 4252 12582 4304 12588
rect 4080 12294 4200 12322
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4080 11762 4108 12174
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4172 11642 4200 12294
rect 4264 11898 4292 12582
rect 4356 12434 4384 16662
rect 4540 16454 4568 18566
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4632 17270 4660 18022
rect 4620 17264 4672 17270
rect 4620 17206 4672 17212
rect 4528 16448 4580 16454
rect 4724 16402 4752 19110
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 18358 4844 18566
rect 4804 18352 4856 18358
rect 4804 18294 4856 18300
rect 4804 17672 4856 17678
rect 4804 17614 4856 17620
rect 5000 17626 5028 19246
rect 5092 18970 5120 19314
rect 5080 18964 5132 18970
rect 5080 18906 5132 18912
rect 5184 17882 5212 19450
rect 5276 19446 5304 20431
rect 18708 20466 18736 21247
rect 20626 20904 20682 20913
rect 20626 20839 20682 20848
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 20180 20505 20208 20538
rect 20166 20496 20222 20505
rect 16854 20431 16856 20440
rect 5724 20402 5776 20408
rect 16908 20431 16910 20440
rect 17776 20460 17828 20466
rect 16856 20402 16908 20408
rect 17776 20402 17828 20408
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 19524 20460 19576 20466
rect 20166 20431 20222 20440
rect 20536 20460 20588 20466
rect 19524 20402 19576 20408
rect 20536 20402 20588 20408
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7852 19854 7880 20334
rect 14648 20324 14700 20330
rect 14648 20266 14700 20272
rect 16396 20324 16448 20330
rect 16396 20266 16448 20272
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12992 20256 13044 20262
rect 12992 20198 13044 20204
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8484 19916 8536 19922
rect 8484 19858 8536 19864
rect 10508 19916 10560 19922
rect 10508 19858 10560 19864
rect 11244 19916 11296 19922
rect 11244 19858 11296 19864
rect 11796 19916 11848 19922
rect 11796 19858 11848 19864
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 5448 19712 5500 19718
rect 5448 19654 5500 19660
rect 7932 19712 7984 19718
rect 7932 19654 7984 19660
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5356 19304 5408 19310
rect 5356 19246 5408 19252
rect 5368 19174 5396 19246
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5460 18578 5488 19654
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 5814 19544 5870 19553
rect 6148 19547 6456 19556
rect 7944 19514 7972 19654
rect 5814 19479 5870 19488
rect 7564 19508 7616 19514
rect 5724 19168 5776 19174
rect 5724 19110 5776 19116
rect 5736 18737 5764 19110
rect 5722 18728 5778 18737
rect 5722 18663 5778 18672
rect 5368 18550 5488 18578
rect 5264 18420 5316 18426
rect 5264 18362 5316 18368
rect 5172 17876 5224 17882
rect 5172 17818 5224 17824
rect 4528 16390 4580 16396
rect 4632 16374 4752 16402
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 4448 15706 4476 16050
rect 4528 16040 4580 16046
rect 4528 15982 4580 15988
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4448 14074 4476 14758
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4448 13297 4476 13330
rect 4434 13288 4490 13297
rect 4434 13223 4490 13232
rect 4356 12406 4476 12434
rect 4448 12306 4476 12406
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4356 11898 4384 12038
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4080 11614 4200 11642
rect 4344 11688 4396 11694
rect 4448 11665 4476 12242
rect 4344 11630 4396 11636
rect 4434 11656 4490 11665
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10192 3384 10198
rect 3238 10160 3294 10169
rect 3332 10134 3384 10140
rect 3436 10130 3464 10610
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3238 10095 3294 10104
rect 3424 10124 3476 10130
rect 3424 10066 3476 10072
rect 3516 10056 3568 10062
rect 3516 9998 3568 10004
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 3146 9072 3202 9081
rect 3146 9007 3202 9016
rect 3160 8974 3188 9007
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2792 8588 2912 8616
rect 2964 8628 3016 8634
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2792 8090 2820 8588
rect 2964 8570 3016 8576
rect 3252 8514 3280 9930
rect 3332 9512 3384 9518
rect 3332 9454 3384 9460
rect 2872 8492 2924 8498
rect 2872 8434 2924 8440
rect 2976 8486 3280 8514
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2778 7848 2834 7857
rect 2778 7783 2834 7792
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6322 2728 7142
rect 2792 6934 2820 7783
rect 2780 6928 2832 6934
rect 2780 6870 2832 6876
rect 2780 6792 2832 6798
rect 2780 6734 2832 6740
rect 2792 6390 2820 6734
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2792 5778 2820 6326
rect 2884 6186 2912 8434
rect 2976 7290 3004 8486
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3054 7984 3110 7993
rect 3054 7919 3110 7928
rect 3068 7478 3096 7919
rect 3160 7886 3188 8366
rect 3344 8004 3372 9454
rect 3528 9364 3556 9998
rect 3712 9654 3740 10134
rect 3896 9722 3924 10746
rect 4080 10606 4108 11614
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 3976 10600 4028 10606
rect 3976 10542 4028 10548
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3700 9648 3752 9654
rect 3606 9616 3662 9625
rect 3700 9590 3752 9596
rect 3606 9551 3662 9560
rect 3620 9382 3648 9551
rect 3988 9518 4016 10542
rect 3976 9512 4028 9518
rect 3882 9480 3938 9489
rect 3976 9454 4028 9460
rect 4080 9450 4108 10542
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3882 9415 3938 9424
rect 4068 9444 4120 9450
rect 3436 9336 3556 9364
rect 3608 9376 3660 9382
rect 3436 9160 3464 9336
rect 3608 9318 3660 9324
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3436 9132 3556 9160
rect 3528 8294 3556 9132
rect 3896 9110 3924 9415
rect 4068 9386 4120 9392
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3988 8838 4016 9318
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 4080 8362 4108 9046
rect 3884 8356 3936 8362
rect 3884 8298 3936 8304
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 3516 8288 3568 8294
rect 3516 8230 3568 8236
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 3344 7976 3556 8004
rect 3148 7880 3200 7886
rect 3148 7822 3200 7828
rect 3424 7812 3476 7818
rect 3424 7754 3476 7760
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3252 7478 3280 7686
rect 3056 7472 3108 7478
rect 3056 7414 3108 7420
rect 3240 7472 3292 7478
rect 3240 7414 3292 7420
rect 2976 7262 3096 7290
rect 2964 7200 3016 7206
rect 2964 7142 3016 7148
rect 2976 6458 3004 7142
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2962 6352 3018 6361
rect 3068 6322 3096 7262
rect 3240 7200 3292 7206
rect 3240 7142 3292 7148
rect 3146 7032 3202 7041
rect 3146 6967 3202 6976
rect 2962 6287 3018 6296
rect 3056 6316 3108 6322
rect 2872 6180 2924 6186
rect 2872 6122 2924 6128
rect 2780 5772 2832 5778
rect 2780 5714 2832 5720
rect 2596 5704 2648 5710
rect 2596 5646 2648 5652
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 4434 2544 5238
rect 2424 4406 2544 4434
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2332 2922 2360 3538
rect 2320 2916 2372 2922
rect 2320 2858 2372 2864
rect 2424 2774 2452 4406
rect 2608 4146 2636 5646
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2516 3738 2544 4082
rect 2700 4078 2728 5510
rect 2780 5296 2832 5302
rect 2780 5238 2832 5244
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2792 3194 2820 5238
rect 2976 5114 3004 6287
rect 3056 6258 3108 6264
rect 3068 6225 3096 6258
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 3160 5710 3188 6967
rect 3252 6769 3280 7142
rect 3344 6798 3372 7686
rect 3436 7410 3464 7754
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3528 7290 3556 7976
rect 3436 7262 3556 7290
rect 3332 6792 3384 6798
rect 3238 6760 3294 6769
rect 3332 6734 3384 6740
rect 3238 6695 3294 6704
rect 3436 6662 3464 7262
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3252 5846 3280 6598
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3344 5914 3372 6394
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3332 5908 3384 5914
rect 3332 5850 3384 5856
rect 3240 5840 3292 5846
rect 3436 5817 3464 6258
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3240 5782 3292 5788
rect 3422 5808 3478 5817
rect 3332 5772 3384 5778
rect 3422 5743 3478 5752
rect 3516 5772 3568 5778
rect 3332 5714 3384 5720
rect 3516 5714 3568 5720
rect 3148 5704 3200 5710
rect 3344 5681 3372 5714
rect 3148 5646 3200 5652
rect 3330 5672 3386 5681
rect 3160 5409 3188 5646
rect 3330 5607 3386 5616
rect 3146 5400 3202 5409
rect 3528 5386 3556 5714
rect 3804 5642 3832 5850
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3896 5522 3924 8298
rect 3974 8256 4030 8265
rect 3974 8191 4030 8200
rect 3988 7886 4016 8191
rect 4172 7970 4200 9522
rect 4264 9518 4292 10678
rect 4356 10198 4384 11630
rect 4434 11591 4490 11600
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4448 10810 4476 11086
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4448 8974 4476 9862
rect 4540 9450 4568 15982
rect 4632 12850 4660 16374
rect 4712 16244 4764 16250
rect 4712 16186 4764 16192
rect 4724 15706 4752 16186
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4632 12102 4660 12786
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4620 11688 4672 11694
rect 4620 11630 4672 11636
rect 4632 11218 4660 11630
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10606 4660 11154
rect 4724 11082 4752 15642
rect 4816 13530 4844 17614
rect 5000 17598 5120 17626
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 4896 16448 4948 16454
rect 4896 16390 4948 16396
rect 4908 16046 4936 16390
rect 5000 16250 5028 17478
rect 5092 16538 5120 17598
rect 5172 17536 5224 17542
rect 5172 17478 5224 17484
rect 5184 17338 5212 17478
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5276 16658 5304 18362
rect 5264 16652 5316 16658
rect 5264 16594 5316 16600
rect 5092 16510 5212 16538
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4908 14958 4936 15982
rect 5092 15570 5120 16390
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 4988 15020 5040 15026
rect 4988 14962 5040 14968
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 4804 13524 4856 13530
rect 4804 13466 4856 13472
rect 4908 13410 4936 14758
rect 5000 14618 5028 14962
rect 4988 14612 5040 14618
rect 4988 14554 5040 14560
rect 5092 14482 5120 15506
rect 5184 15502 5212 16510
rect 5368 16130 5396 18550
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5460 18193 5488 18362
rect 5446 18184 5502 18193
rect 5630 18184 5686 18193
rect 5446 18119 5502 18128
rect 5552 18142 5630 18170
rect 5448 17740 5500 17746
rect 5448 17682 5500 17688
rect 5460 17649 5488 17682
rect 5446 17640 5502 17649
rect 5446 17575 5502 17584
rect 5276 16102 5396 16130
rect 5448 16108 5500 16114
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 5172 14544 5224 14550
rect 5172 14486 5224 14492
rect 5080 14476 5132 14482
rect 5080 14418 5132 14424
rect 5080 14340 5132 14346
rect 5080 14282 5132 14288
rect 5092 14074 5120 14282
rect 5080 14068 5132 14074
rect 5080 14010 5132 14016
rect 5092 13870 5120 14010
rect 5080 13864 5132 13870
rect 5080 13806 5132 13812
rect 4816 13382 4936 13410
rect 4816 12646 4844 13382
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4896 12640 4948 12646
rect 4896 12582 4948 12588
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10600 4672 10606
rect 4620 10542 4672 10548
rect 4816 10554 4844 12582
rect 4908 10674 4936 12582
rect 5184 12434 5212 14486
rect 5092 12406 5212 12434
rect 4988 11144 5040 11150
rect 4986 11112 4988 11121
rect 5040 11112 5042 11121
rect 4986 11047 5042 11056
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4816 10526 5028 10554
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 4712 9988 4764 9994
rect 4712 9930 4764 9936
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4528 9444 4580 9450
rect 4528 9386 4580 9392
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4264 8090 4292 8910
rect 4344 8832 4396 8838
rect 4528 8832 4580 8838
rect 4396 8792 4476 8820
rect 4344 8774 4396 8780
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4172 7942 4292 7970
rect 3976 7880 4028 7886
rect 3976 7822 4028 7828
rect 3988 7206 4016 7822
rect 4068 7336 4120 7342
rect 4068 7278 4120 7284
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3976 6656 4028 6662
rect 4080 6644 4108 7278
rect 4028 6616 4108 6644
rect 4160 6656 4212 6662
rect 3976 6598 4028 6604
rect 4160 6598 4212 6604
rect 3146 5335 3202 5344
rect 3344 5358 3556 5386
rect 3712 5494 3924 5522
rect 2884 5086 3004 5114
rect 2884 3369 2912 5086
rect 2964 5024 3016 5030
rect 2964 4966 3016 4972
rect 2976 4282 3004 4966
rect 3238 4856 3294 4865
rect 3238 4791 3240 4800
rect 3292 4791 3294 4800
rect 3240 4762 3292 4768
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3068 3534 3096 4150
rect 3056 3528 3108 3534
rect 3252 3505 3280 4558
rect 3056 3470 3108 3476
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2608 3058 2636 3130
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2608 2961 2636 2994
rect 2594 2952 2650 2961
rect 2594 2887 2650 2896
rect 2778 2816 2834 2825
rect 2424 2746 2636 2774
rect 3344 2774 3372 5358
rect 3712 5284 3740 5494
rect 2778 2751 2834 2760
rect 2608 2582 2636 2746
rect 2596 2576 2648 2582
rect 2596 2518 2648 2524
rect 2792 2446 2820 2751
rect 3252 2746 3372 2774
rect 3436 5256 3740 5284
rect 3792 5296 3844 5302
rect 1308 2440 1360 2446
rect 2780 2440 2832 2446
rect 1308 2382 1360 2388
rect 2608 2400 2780 2428
rect 2228 2372 2280 2378
rect 2228 2314 2280 2320
rect 848 1964 900 1970
rect 848 1906 900 1912
rect 2240 800 2268 2314
rect 2608 800 2636 2400
rect 2780 2382 2832 2388
rect 2964 1896 3016 1902
rect 2964 1838 3016 1844
rect 2976 1737 3004 1838
rect 2962 1728 3018 1737
rect 2962 1663 3018 1672
rect 2976 870 3096 898
rect 2976 800 3004 870
rect 2226 0 2282 800
rect 2594 0 2650 800
rect 2962 0 3018 800
rect 3068 762 3096 870
rect 3252 762 3280 2746
rect 3436 2650 3464 5256
rect 3792 5238 3844 5244
rect 3804 5098 3832 5238
rect 3882 5128 3938 5137
rect 3792 5092 3844 5098
rect 3882 5063 3938 5072
rect 3792 5034 3844 5040
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3896 4758 3924 5063
rect 3884 4752 3936 4758
rect 3884 4694 3936 4700
rect 3700 4684 3752 4690
rect 3700 4626 3752 4632
rect 3712 4593 3740 4626
rect 3698 4584 3754 4593
rect 3698 4519 3754 4528
rect 3514 4312 3570 4321
rect 3514 4247 3570 4256
rect 3528 4214 3556 4247
rect 3516 4208 3568 4214
rect 3516 4150 3568 4156
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 3712 2938 3740 3431
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3896 3194 3924 3334
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3712 2910 3924 2938
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3424 2644 3476 2650
rect 3424 2586 3476 2592
rect 3896 2530 3924 2910
rect 3620 2502 3924 2530
rect 3344 870 3464 898
rect 3344 800 3372 870
rect 3068 734 3280 762
rect 3330 0 3386 800
rect 3436 762 3464 870
rect 3620 762 3648 2502
rect 3988 2417 4016 6598
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 4080 4185 4108 5646
rect 4172 5370 4200 6598
rect 4264 5914 4292 7942
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4356 7546 4384 7890
rect 4448 7886 4476 8792
rect 4528 8774 4580 8780
rect 4540 8634 4568 8774
rect 4528 8628 4580 8634
rect 4528 8570 4580 8576
rect 4632 8514 4660 9522
rect 4540 8486 4660 8514
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4342 6216 4398 6225
rect 4342 6151 4344 6160
rect 4396 6151 4398 6160
rect 4344 6122 4396 6128
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4160 5364 4212 5370
rect 4160 5306 4212 5312
rect 4356 4321 4384 6122
rect 4540 6118 4568 8486
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 7342 4660 8230
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4632 6934 4660 7278
rect 4620 6928 4672 6934
rect 4620 6870 4672 6876
rect 4618 6760 4674 6769
rect 4618 6695 4674 6704
rect 4632 6662 4660 6695
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4434 5808 4490 5817
rect 4434 5743 4490 5752
rect 4448 5710 4476 5743
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4436 5568 4488 5574
rect 4436 5510 4488 5516
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4252 4208 4304 4214
rect 4066 4176 4122 4185
rect 4252 4150 4304 4156
rect 4066 4111 4122 4120
rect 4160 4004 4212 4010
rect 4160 3946 4212 3952
rect 4172 3534 4200 3946
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4264 3194 4292 4150
rect 4344 3936 4396 3942
rect 4344 3878 4396 3884
rect 4356 3602 4384 3878
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4448 3398 4476 5510
rect 4540 5302 4568 6054
rect 4632 5386 4660 6598
rect 4724 5914 4752 9930
rect 4816 9926 4844 10134
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9110 4844 9862
rect 4896 9648 4948 9654
rect 4896 9590 4948 9596
rect 4804 9104 4856 9110
rect 4804 9046 4856 9052
rect 4802 8936 4858 8945
rect 4802 8871 4858 8880
rect 4816 6882 4844 8871
rect 4908 8634 4936 9590
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4908 8022 4936 8570
rect 5000 8430 5028 10526
rect 4988 8424 5040 8430
rect 4988 8366 5040 8372
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4908 7002 4936 7958
rect 4896 6996 4948 7002
rect 4896 6938 4948 6944
rect 4816 6854 5028 6882
rect 4802 6352 4858 6361
rect 4802 6287 4858 6296
rect 4816 6186 4844 6287
rect 4804 6180 4856 6186
rect 4804 6122 4856 6128
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4712 5908 4764 5914
rect 4712 5850 4764 5856
rect 4724 5574 4752 5850
rect 4712 5568 4764 5574
rect 4712 5510 4764 5516
rect 4632 5358 4752 5386
rect 4908 5370 4936 6054
rect 4528 5296 4580 5302
rect 4528 5238 4580 5244
rect 4620 5160 4672 5166
rect 4620 5102 4672 5108
rect 4724 5114 4752 5358
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 5000 5234 5028 6854
rect 5092 5710 5120 12406
rect 5276 11370 5304 16102
rect 5448 16050 5500 16056
rect 5356 16040 5408 16046
rect 5354 16008 5356 16017
rect 5408 16008 5410 16017
rect 5354 15943 5410 15952
rect 5460 15638 5488 16050
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5552 15162 5580 18142
rect 5630 18119 5686 18128
rect 5828 17082 5856 19479
rect 7564 19450 7616 19456
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 7576 19417 7604 19450
rect 7562 19408 7618 19417
rect 7562 19343 7618 19352
rect 8024 19304 8076 19310
rect 8024 19246 8076 19252
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6380 18902 6408 19178
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6000 18896 6052 18902
rect 6000 18838 6052 18844
rect 6368 18896 6420 18902
rect 6368 18838 6420 18844
rect 6012 18329 6040 18838
rect 6564 18834 6592 19110
rect 7196 18964 7248 18970
rect 7196 18906 7248 18912
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 5998 18320 6054 18329
rect 5998 18255 6054 18264
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5920 17241 5948 17478
rect 5906 17232 5962 17241
rect 5906 17167 5962 17176
rect 5828 17054 5948 17082
rect 5816 16992 5868 16998
rect 5816 16934 5868 16940
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5724 16652 5776 16658
rect 5724 16594 5776 16600
rect 5540 15156 5592 15162
rect 5540 15098 5592 15104
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5368 13938 5396 14894
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5356 13932 5408 13938
rect 5356 13874 5408 13880
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5184 11354 5304 11370
rect 5172 11348 5304 11354
rect 5224 11342 5304 11348
rect 5172 11290 5224 11296
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5184 9518 5212 11154
rect 5356 11076 5408 11082
rect 5356 11018 5408 11024
rect 5368 10470 5396 11018
rect 5460 10810 5488 13738
rect 5552 12442 5580 14350
rect 5644 12481 5672 16594
rect 5736 13841 5764 16594
rect 5828 14793 5856 16934
rect 5920 15162 5948 17054
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5814 14784 5870 14793
rect 5814 14719 5870 14728
rect 5816 13864 5868 13870
rect 5722 13832 5778 13841
rect 5816 13806 5868 13812
rect 5722 13767 5778 13776
rect 5724 13728 5776 13734
rect 5724 13670 5776 13676
rect 5736 12986 5764 13670
rect 5828 13326 5856 13806
rect 5920 13530 5948 14962
rect 5908 13524 5960 13530
rect 5908 13466 5960 13472
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5828 12628 5856 13126
rect 6012 12832 6040 18090
rect 6564 18086 6592 18770
rect 6840 18290 6868 18770
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 7012 18216 7064 18222
rect 7012 18158 7064 18164
rect 6276 18080 6328 18086
rect 6276 18022 6328 18028
rect 6552 18080 6604 18086
rect 6552 18022 6604 18028
rect 6288 17882 6316 18022
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6288 17746 6316 17818
rect 6276 17740 6328 17746
rect 6276 17682 6328 17688
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6552 17536 6604 17542
rect 6552 17478 6604 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6104 16726 6132 17070
rect 6092 16720 6144 16726
rect 6092 16662 6144 16668
rect 6458 16552 6514 16561
rect 6458 16487 6460 16496
rect 6512 16487 6514 16496
rect 6460 16458 6512 16464
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6564 16250 6592 17478
rect 6644 16584 6696 16590
rect 6644 16526 6696 16532
rect 6656 16454 6684 16526
rect 6644 16448 6696 16454
rect 6644 16390 6696 16396
rect 6552 16244 6604 16250
rect 6552 16186 6604 16192
rect 6552 15360 6604 15366
rect 6552 15302 6604 15308
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 6564 14822 6592 15302
rect 6656 15042 6684 16390
rect 6748 16250 6776 17546
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6748 15881 6776 15914
rect 6734 15872 6790 15881
rect 6734 15807 6790 15816
rect 6840 15502 6868 17682
rect 6920 17536 6972 17542
rect 6920 17478 6972 17484
rect 6932 16153 6960 17478
rect 7024 17338 7052 18158
rect 7104 17536 7156 17542
rect 7102 17504 7104 17513
rect 7156 17504 7158 17513
rect 7102 17439 7158 17448
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6918 16144 6974 16153
rect 6918 16079 6974 16088
rect 7024 16046 7052 17138
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7024 15910 7052 15982
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 7012 15904 7064 15910
rect 7012 15846 7064 15852
rect 6828 15496 6880 15502
rect 6932 15484 6960 15846
rect 7012 15496 7064 15502
rect 6932 15456 7012 15484
rect 6828 15438 6880 15444
rect 7012 15438 7064 15444
rect 6840 15162 6868 15438
rect 6828 15156 6880 15162
rect 6828 15098 6880 15104
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6656 15014 6868 15042
rect 6642 14920 6698 14929
rect 6642 14855 6698 14864
rect 6552 14816 6604 14822
rect 6552 14758 6604 14764
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6564 14113 6592 14758
rect 6656 14618 6684 14855
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6644 14476 6696 14482
rect 6644 14418 6696 14424
rect 6656 14278 6684 14418
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6550 14104 6606 14113
rect 6550 14039 6606 14048
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6564 13002 6592 13806
rect 6656 13802 6684 14214
rect 6748 13870 6776 14214
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6656 13530 6684 13738
rect 6840 13716 6868 15014
rect 6748 13688 6868 13716
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6748 13190 6776 13688
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6736 13184 6788 13190
rect 6736 13126 6788 13132
rect 6564 12974 6776 13002
rect 6644 12844 6696 12850
rect 6012 12804 6132 12832
rect 5908 12776 5960 12782
rect 5906 12744 5908 12753
rect 5960 12744 5962 12753
rect 5906 12679 5962 12688
rect 6000 12708 6052 12714
rect 6000 12650 6052 12656
rect 5828 12600 5948 12628
rect 5630 12472 5686 12481
rect 5540 12436 5592 12442
rect 5630 12407 5686 12416
rect 5816 12436 5868 12442
rect 5540 12378 5592 12384
rect 5816 12378 5868 12384
rect 5632 12368 5684 12374
rect 5538 12336 5594 12345
rect 5632 12310 5684 12316
rect 5724 12368 5776 12374
rect 5724 12310 5776 12316
rect 5538 12271 5594 12280
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5276 10266 5304 10406
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5172 9512 5224 9518
rect 5172 9454 5224 9460
rect 5172 8424 5224 8430
rect 5276 8412 5304 10066
rect 5356 9920 5408 9926
rect 5460 9908 5488 10610
rect 5408 9880 5488 9908
rect 5356 9862 5408 9868
rect 5368 8634 5396 9862
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5552 9382 5580 12271
rect 5644 11762 5672 12310
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5644 11393 5672 11698
rect 5630 11384 5686 11393
rect 5630 11319 5686 11328
rect 5736 11218 5764 12310
rect 5828 11694 5856 12378
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5540 9376 5592 9382
rect 5540 9318 5592 9324
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5644 9042 5672 10950
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5736 8974 5764 11018
rect 5828 10742 5856 11630
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10169 5856 10406
rect 5814 10160 5870 10169
rect 5814 10095 5870 10104
rect 5920 9654 5948 12600
rect 6012 11150 6040 12650
rect 6104 12442 6132 12804
rect 6644 12786 6696 12792
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6092 12436 6144 12442
rect 6092 12378 6144 12384
rect 6564 12374 6592 12718
rect 6656 12481 6684 12786
rect 6642 12472 6698 12481
rect 6642 12407 6698 12416
rect 6552 12368 6604 12374
rect 6552 12310 6604 12316
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6550 11928 6606 11937
rect 6550 11863 6606 11872
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6472 11098 6500 11766
rect 6564 11529 6592 11863
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 6550 11520 6606 11529
rect 6550 11455 6606 11464
rect 6656 11150 6684 11630
rect 6644 11144 6696 11150
rect 6472 11070 6592 11098
rect 6644 11086 6696 11092
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6000 9920 6052 9926
rect 6000 9862 6052 9868
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5724 8968 5776 8974
rect 5724 8910 5776 8916
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5224 8384 5304 8412
rect 5172 8366 5224 8372
rect 5184 7954 5212 8366
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7002 5212 7890
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5368 6798 5396 8570
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4526 4720 4582 4729
rect 4632 4690 4660 5102
rect 4724 5086 5028 5114
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4724 4758 4752 4966
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4526 4655 4582 4664
rect 4620 4684 4672 4690
rect 4540 3602 4568 4655
rect 4620 4626 4672 4632
rect 4632 4282 4660 4626
rect 4908 4622 4936 4966
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4724 3602 4752 4082
rect 4816 3738 4844 4490
rect 5000 4434 5028 5086
rect 5184 4690 5212 6598
rect 5276 6458 5304 6598
rect 5264 6452 5316 6458
rect 5264 6394 5316 6400
rect 5460 6186 5488 7482
rect 5552 7426 5580 8842
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 7954 5764 8774
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5552 7398 5672 7426
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 6066 5488 6122
rect 5276 6038 5488 6066
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 4908 4406 5028 4434
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 4804 3732 4856 3738
rect 4804 3674 4856 3680
rect 4528 3596 4580 3602
rect 4528 3538 4580 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4252 3188 4304 3194
rect 4252 3130 4304 3136
rect 4158 3088 4214 3097
rect 4158 3023 4214 3032
rect 4252 3052 4304 3058
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3974 2408 4030 2417
rect 3700 2372 3752 2378
rect 3974 2343 4030 2352
rect 3700 2314 3752 2320
rect 3712 800 3740 2314
rect 3974 2136 4030 2145
rect 3974 2071 3976 2080
rect 4028 2071 4030 2080
rect 3976 2042 4028 2048
rect 4080 800 4108 2790
rect 4172 2310 4200 3023
rect 4252 2994 4304 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4264 2650 4292 2994
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4448 1601 4476 2994
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4540 2514 4568 2790
rect 4908 2774 4936 4406
rect 4986 4312 5042 4321
rect 4986 4247 5042 4256
rect 5000 4146 5028 4247
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 5000 2854 5028 4082
rect 5078 4040 5134 4049
rect 5184 4010 5212 4422
rect 5078 3975 5080 3984
rect 5132 3975 5134 3984
rect 5172 4004 5224 4010
rect 5080 3946 5132 3952
rect 5172 3946 5224 3952
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 4988 2848 5040 2854
rect 4988 2790 5040 2796
rect 4632 2746 4936 2774
rect 4632 2650 4660 2746
rect 5092 2689 5120 3606
rect 5276 3398 5304 6038
rect 5552 5914 5580 7278
rect 5644 7274 5672 7398
rect 5632 7268 5684 7274
rect 5632 7210 5684 7216
rect 5828 6984 5856 9454
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5644 6956 5856 6984
rect 5540 5908 5592 5914
rect 5540 5850 5592 5856
rect 5538 5808 5594 5817
rect 5538 5743 5594 5752
rect 5356 5568 5408 5574
rect 5356 5510 5408 5516
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5368 5370 5396 5510
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5368 4146 5396 4422
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5170 2952 5226 2961
rect 5170 2887 5226 2896
rect 5078 2680 5134 2689
rect 4620 2644 4672 2650
rect 5078 2615 5134 2624
rect 4620 2586 4672 2592
rect 4528 2508 4580 2514
rect 4528 2450 4580 2456
rect 4802 1728 4858 1737
rect 4802 1663 4858 1672
rect 4434 1592 4490 1601
rect 4434 1527 4490 1536
rect 4448 800 4476 1527
rect 4816 800 4844 1663
rect 5184 800 5212 2887
rect 5368 2650 5396 3334
rect 5460 2990 5488 5510
rect 5552 4826 5580 5743
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5644 4486 5672 6956
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5736 6322 5764 6666
rect 5724 6316 5776 6322
rect 5724 6258 5776 6264
rect 5736 5817 5764 6258
rect 5828 6254 5856 6802
rect 5816 6248 5868 6254
rect 5816 6190 5868 6196
rect 5722 5808 5778 5817
rect 5722 5743 5778 5752
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5552 3670 5580 3878
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5644 3398 5672 4422
rect 5632 3392 5684 3398
rect 5632 3334 5684 3340
rect 5736 3074 5764 5646
rect 5828 5302 5856 6190
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5920 4146 5948 8774
rect 6012 7993 6040 9862
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6564 8480 6592 11070
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10810 6684 10950
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6656 9654 6684 9862
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6748 9518 6776 12974
rect 6840 12442 6868 13262
rect 6828 12436 6880 12442
rect 6828 12378 6880 12384
rect 6932 12186 6960 15098
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 7024 14074 7052 14962
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 7116 13569 7144 17070
rect 7208 15094 7236 18906
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18358 7696 18566
rect 8036 18426 8064 19246
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 8128 18426 8156 18702
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8024 18420 8076 18426
rect 8024 18362 8076 18368
rect 8116 18420 8168 18426
rect 8116 18362 8168 18368
rect 7656 18352 7708 18358
rect 7656 18294 7708 18300
rect 7668 18222 7696 18294
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 8128 18154 8156 18362
rect 8312 18290 8340 18634
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8496 18222 8524 19858
rect 9864 19848 9916 19854
rect 9864 19790 9916 19796
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8484 18216 8536 18222
rect 8484 18158 8536 18164
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 8208 18148 8260 18154
rect 8208 18090 8260 18096
rect 7472 17808 7524 17814
rect 7470 17776 7472 17785
rect 7524 17776 7526 17785
rect 8220 17746 8248 18090
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 7470 17711 7526 17720
rect 7656 17740 7708 17746
rect 7656 17682 7708 17688
rect 8208 17740 8260 17746
rect 8208 17682 8260 17688
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7392 16998 7420 17614
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7196 15088 7248 15094
rect 7196 15030 7248 15036
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 7208 14482 7236 14758
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7300 14414 7328 16934
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7392 16114 7420 16594
rect 7562 16552 7618 16561
rect 7562 16487 7618 16496
rect 7380 16108 7432 16114
rect 7380 16050 7432 16056
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7392 13802 7420 16050
rect 7484 15881 7512 16050
rect 7576 16046 7604 16487
rect 7564 16040 7616 16046
rect 7564 15982 7616 15988
rect 7470 15872 7526 15881
rect 7470 15807 7526 15816
rect 7472 15496 7524 15502
rect 7524 15456 7604 15484
rect 7472 15438 7524 15444
rect 7472 13864 7524 13870
rect 7472 13806 7524 13812
rect 7380 13796 7432 13802
rect 7380 13738 7432 13744
rect 7484 13734 7512 13806
rect 7472 13728 7524 13734
rect 7472 13670 7524 13676
rect 7102 13560 7158 13569
rect 7102 13495 7158 13504
rect 7012 13456 7064 13462
rect 7012 13398 7064 13404
rect 7024 13274 7052 13398
rect 7024 13246 7328 13274
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6840 12158 6960 12186
rect 6840 11234 6868 12158
rect 6918 12064 6974 12073
rect 6918 11999 6974 12008
rect 6932 11354 6960 11999
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6840 11206 6960 11234
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10266 6868 10950
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 9512 6788 9518
rect 6840 9489 6868 10202
rect 6932 10198 6960 11206
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6918 10024 6974 10033
rect 6918 9959 6974 9968
rect 6932 9926 6960 9959
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6932 9722 6960 9862
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6736 9454 6788 9460
rect 6826 9480 6882 9489
rect 6826 9415 6882 9424
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6656 8974 6684 9318
rect 6748 9042 6776 9318
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6840 8566 6868 8842
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6932 8498 6960 9658
rect 6920 8492 6972 8498
rect 6564 8452 6684 8480
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6564 8090 6592 8298
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 5998 7984 6054 7993
rect 5998 7919 6054 7928
rect 6000 7744 6052 7750
rect 6000 7686 6052 7692
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6012 7546 6040 7686
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6012 6798 6040 7142
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6182 6760 6238 6769
rect 6012 6633 6040 6734
rect 6182 6695 6238 6704
rect 6196 6662 6224 6695
rect 6184 6656 6236 6662
rect 5998 6624 6054 6633
rect 6184 6598 6236 6604
rect 5998 6559 6054 6568
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6182 5944 6238 5953
rect 6182 5879 6238 5888
rect 5998 5808 6054 5817
rect 5998 5743 6054 5752
rect 5816 4140 5868 4146
rect 5816 4082 5868 4088
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 5828 3913 5856 4082
rect 5814 3904 5870 3913
rect 5814 3839 5870 3848
rect 5814 3632 5870 3641
rect 6012 3602 6040 5743
rect 6196 5642 6224 5879
rect 6184 5636 6236 5642
rect 6184 5578 6236 5584
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 6564 4690 6592 7686
rect 6656 4865 6684 8452
rect 6920 8434 6972 8440
rect 6920 8356 6972 8362
rect 6748 8316 6920 8344
rect 6748 5710 6776 8316
rect 6920 8298 6972 8304
rect 6828 8084 6880 8090
rect 6828 8026 6880 8032
rect 6840 6322 6868 8026
rect 7024 7834 7052 13126
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7116 9926 7144 10406
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7116 7954 7144 8774
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7024 7806 7144 7834
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7002 7052 7686
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 7012 6996 7064 7002
rect 7012 6938 7064 6944
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6734 5400 6790 5409
rect 6734 5335 6790 5344
rect 6748 5234 6776 5335
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6642 4856 6698 4865
rect 6642 4791 6698 4800
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6564 4282 6592 4490
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6736 4480 6788 4486
rect 6736 4422 6788 4428
rect 6552 4276 6604 4282
rect 6552 4218 6604 4224
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 6196 3913 6224 4014
rect 6182 3904 6238 3913
rect 6182 3839 6238 3848
rect 5814 3567 5816 3576
rect 5868 3567 5870 3576
rect 6000 3596 6052 3602
rect 5816 3538 5868 3544
rect 6000 3538 6052 3544
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 5908 3392 5960 3398
rect 5908 3334 5960 3340
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5644 3046 5764 3074
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5540 2916 5592 2922
rect 5540 2858 5592 2864
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5446 2544 5502 2553
rect 5446 2479 5448 2488
rect 5500 2479 5502 2488
rect 5448 2450 5500 2456
rect 5552 800 5580 2858
rect 5644 2825 5672 3046
rect 5920 2938 5948 3334
rect 6012 3126 6040 3334
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6000 3120 6052 3126
rect 6000 3062 6052 3068
rect 6564 2990 6592 3470
rect 6656 3058 6684 4422
rect 6748 3534 6776 4422
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3233 6776 3334
rect 6734 3224 6790 3233
rect 6734 3159 6790 3168
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6552 2984 6604 2990
rect 6366 2952 6422 2961
rect 5920 2910 6040 2938
rect 5908 2848 5960 2854
rect 5630 2816 5686 2825
rect 5908 2790 5960 2796
rect 5630 2751 5686 2760
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5736 1737 5764 2382
rect 5722 1728 5778 1737
rect 5722 1663 5778 1672
rect 5920 800 5948 2790
rect 3436 734 3648 762
rect 3698 0 3754 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5538 0 5594 800
rect 5906 0 5962 800
rect 6012 762 6040 2910
rect 6552 2926 6604 2932
rect 6366 2887 6422 2896
rect 6380 2854 6408 2887
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6840 2774 6868 6258
rect 6932 5778 6960 6938
rect 7116 6662 7144 7806
rect 7208 7290 7236 12922
rect 7300 11898 7328 13246
rect 7472 13184 7524 13190
rect 7472 13126 7524 13132
rect 7378 12336 7434 12345
rect 7378 12271 7380 12280
rect 7432 12271 7434 12280
rect 7380 12242 7432 12248
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7484 11830 7512 13126
rect 7472 11824 7524 11830
rect 7472 11766 7524 11772
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7300 10266 7328 10542
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7392 7478 7420 11494
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 8945 7512 11086
rect 7576 10810 7604 15456
rect 7668 14362 7696 17682
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7760 17134 7788 17614
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 7840 17060 7892 17066
rect 7840 17002 7892 17008
rect 7746 16416 7802 16425
rect 7746 16351 7802 16360
rect 7760 16182 7788 16351
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7748 15904 7800 15910
rect 7748 15846 7800 15852
rect 7760 14804 7788 15846
rect 7852 14958 7880 17002
rect 7932 16448 7984 16454
rect 7930 16416 7932 16425
rect 8116 16448 8168 16454
rect 7984 16416 7986 16425
rect 8116 16390 8168 16396
rect 7930 16351 7986 16360
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7944 16153 7972 16186
rect 7930 16144 7986 16153
rect 7930 16079 7986 16088
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8036 15706 8064 15982
rect 8128 15910 8156 16390
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8024 15700 8076 15706
rect 8024 15642 8076 15648
rect 8116 15632 8168 15638
rect 8116 15574 8168 15580
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7760 14776 7880 14804
rect 7668 14334 7788 14362
rect 7656 14272 7708 14278
rect 7656 14214 7708 14220
rect 7668 13841 7696 14214
rect 7654 13832 7710 13841
rect 7654 13767 7710 13776
rect 7760 13462 7788 14334
rect 7748 13456 7800 13462
rect 7748 13398 7800 13404
rect 7760 13326 7788 13398
rect 7748 13320 7800 13326
rect 7748 13262 7800 13268
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12782 7788 13126
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 12434 7788 12718
rect 7668 12406 7788 12434
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7576 9722 7604 10474
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7668 8514 7696 12406
rect 7748 12300 7800 12306
rect 7748 12242 7800 12248
rect 7760 11558 7788 12242
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 7852 11098 7880 14776
rect 7760 11070 7880 11098
rect 7760 9994 7788 11070
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8634 7788 8774
rect 7852 8634 7880 10950
rect 7944 10010 7972 15030
rect 8024 13320 8076 13326
rect 8024 13262 8076 13268
rect 8036 12442 8064 13262
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8036 12102 8064 12378
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8128 11880 8156 15574
rect 8220 12918 8248 17682
rect 8312 17338 8340 18022
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 17338 8524 17478
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8588 17184 8616 19314
rect 9876 19310 9904 19790
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 19514 10456 19654
rect 10416 19508 10468 19514
rect 10416 19450 10468 19456
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9864 19304 9916 19310
rect 9864 19246 9916 19252
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 8668 18284 8720 18290
rect 8668 18226 8720 18232
rect 8680 17338 8708 18226
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 9034 17640 9090 17649
rect 9034 17575 9036 17584
rect 9088 17575 9090 17584
rect 9036 17546 9088 17552
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8760 17264 8812 17270
rect 8760 17206 8812 17212
rect 8404 17156 8616 17184
rect 8300 17128 8352 17134
rect 8298 17096 8300 17105
rect 8352 17096 8354 17105
rect 8298 17031 8354 17040
rect 8404 14770 8432 17156
rect 8772 17116 8800 17206
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 8496 17088 8800 17116
rect 8942 17096 8998 17105
rect 8496 16794 8524 17088
rect 8942 17031 8944 17040
rect 8996 17031 8998 17040
rect 8944 17002 8996 17008
rect 8576 16992 8628 16998
rect 8576 16934 8628 16940
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8588 16697 8616 16934
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8668 16720 8720 16726
rect 8574 16688 8630 16697
rect 8668 16662 8720 16668
rect 8574 16623 8630 16632
rect 8680 16572 8708 16662
rect 8588 16544 8708 16572
rect 9036 16584 9088 16590
rect 8484 16244 8536 16250
rect 8484 16186 8536 16192
rect 8496 15910 8524 16186
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 8496 15366 8524 15846
rect 8484 15360 8536 15366
rect 8484 15302 8536 15308
rect 8404 14742 8524 14770
rect 8392 14612 8444 14618
rect 8392 14554 8444 14560
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 13433 8340 14214
rect 8298 13424 8354 13433
rect 8298 13359 8354 13368
rect 8208 12912 8260 12918
rect 8208 12854 8260 12860
rect 8298 12880 8354 12889
rect 8298 12815 8354 12824
rect 8312 12646 8340 12815
rect 8300 12640 8352 12646
rect 8298 12608 8300 12617
rect 8352 12608 8354 12617
rect 8298 12543 8354 12552
rect 8404 12434 8432 14554
rect 8496 12986 8524 14742
rect 8484 12980 8536 12986
rect 8484 12922 8536 12928
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8036 11852 8156 11880
rect 8312 12406 8432 12434
rect 8036 11218 8064 11852
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 8036 10713 8064 11154
rect 8128 11014 8156 11698
rect 8312 11642 8340 12406
rect 8220 11614 8340 11642
rect 8392 11620 8444 11626
rect 8220 11558 8248 11614
rect 8392 11562 8444 11568
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8220 11150 8248 11494
rect 8208 11144 8260 11150
rect 8208 11086 8260 11092
rect 8300 11144 8352 11150
rect 8300 11086 8352 11092
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 8206 10840 8262 10849
rect 8206 10775 8208 10784
rect 8260 10775 8262 10784
rect 8208 10746 8260 10752
rect 8116 10736 8168 10742
rect 8022 10704 8078 10713
rect 8116 10678 8168 10684
rect 8206 10704 8262 10713
rect 8022 10639 8078 10648
rect 8128 10606 8156 10678
rect 8206 10639 8262 10648
rect 8116 10600 8168 10606
rect 8022 10568 8078 10577
rect 8116 10542 8168 10548
rect 8022 10503 8078 10512
rect 8036 10266 8064 10503
rect 8024 10260 8076 10266
rect 8024 10202 8076 10208
rect 8128 10198 8156 10542
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8128 10062 8156 10134
rect 8220 10130 8248 10639
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 10056 8168 10062
rect 7944 9982 8064 10010
rect 8116 9998 8168 10004
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7484 8486 7696 8514
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7208 7262 7328 7290
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7024 6474 7052 6598
rect 7024 6446 7144 6474
rect 7012 6384 7064 6390
rect 7012 6326 7064 6332
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6918 5536 6974 5545
rect 6918 5471 6974 5480
rect 6932 5370 6960 5471
rect 6920 5364 6972 5370
rect 6920 5306 6972 5312
rect 6920 4276 6972 4282
rect 6920 4218 6972 4224
rect 6932 2854 6960 4218
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6564 2746 6868 2774
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 1902 6592 2746
rect 7024 2378 7052 6326
rect 7116 6322 7144 6446
rect 7104 6316 7156 6322
rect 7104 6258 7156 6264
rect 7116 5409 7144 6258
rect 7102 5400 7158 5409
rect 7102 5335 7158 5344
rect 7208 5234 7236 7142
rect 7300 6390 7328 7262
rect 7392 6934 7420 7414
rect 7380 6928 7432 6934
rect 7380 6870 7432 6876
rect 7484 6866 7512 8486
rect 7564 8424 7616 8430
rect 7564 8366 7616 8372
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7472 6724 7524 6730
rect 7472 6666 7524 6672
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7484 6254 7512 6666
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7392 5914 7420 6190
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7288 5840 7340 5846
rect 7288 5782 7340 5788
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7116 4826 7144 5170
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7104 4072 7156 4078
rect 7104 4014 7156 4020
rect 7116 3942 7144 4014
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7116 2990 7144 3878
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7208 2774 7236 5170
rect 7300 4010 7328 5782
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5137 7420 5510
rect 7378 5128 7434 5137
rect 7378 5063 7434 5072
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4004 7340 4010
rect 7288 3946 7340 3952
rect 7288 3392 7340 3398
rect 7288 3334 7340 3340
rect 7116 2746 7236 2774
rect 7116 2666 7144 2746
rect 7116 2638 7236 2666
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7012 2372 7064 2378
rect 7012 2314 7064 2320
rect 6644 2304 6696 2310
rect 7116 2258 7144 2450
rect 6644 2246 6696 2252
rect 6552 1896 6604 1902
rect 6656 1873 6684 2246
rect 7024 2230 7144 2258
rect 6552 1838 6604 1844
rect 6642 1864 6698 1873
rect 6642 1799 6698 1808
rect 6196 870 6316 898
rect 6196 762 6224 870
rect 6288 800 6316 870
rect 6656 800 6684 1799
rect 7024 800 7052 2230
rect 7208 2106 7236 2638
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7300 1902 7328 3334
rect 7392 3058 7420 4966
rect 7484 4826 7512 6190
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7576 4622 7604 8366
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7576 4282 7604 4558
rect 7564 4276 7616 4282
rect 7564 4218 7616 4224
rect 7668 4146 7696 8298
rect 7748 8016 7800 8022
rect 7746 7984 7748 7993
rect 7800 7984 7802 7993
rect 7746 7919 7802 7928
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7274 7880 7822
rect 7944 7410 7972 9862
rect 8036 8974 8064 9982
rect 8116 9716 8168 9722
rect 8116 9658 8168 9664
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8498 8064 8910
rect 8128 8906 8156 9658
rect 8312 9654 8340 11086
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8220 9042 8248 9318
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8114 8664 8170 8673
rect 8114 8599 8116 8608
rect 8168 8599 8170 8608
rect 8116 8570 8168 8576
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 7404 7984 7410
rect 7932 7346 7984 7352
rect 7840 7268 7892 7274
rect 7840 7210 7892 7216
rect 7852 6798 7880 7210
rect 7932 7200 7984 7206
rect 7932 7142 7984 7148
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7760 5098 7788 6666
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7748 5092 7800 5098
rect 7748 5034 7800 5040
rect 7852 4554 7880 6598
rect 7840 4548 7892 4554
rect 7840 4490 7892 4496
rect 7852 4282 7880 4490
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7656 4140 7708 4146
rect 7576 4100 7656 4128
rect 7380 3052 7432 3058
rect 7380 2994 7432 3000
rect 7576 2938 7604 4100
rect 7656 4082 7708 4088
rect 7748 3936 7800 3942
rect 7748 3878 7800 3884
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7760 3346 7788 3878
rect 7944 3534 7972 7142
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 8036 6254 8064 6938
rect 8220 6866 8248 8978
rect 8312 8090 8340 9454
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8312 7410 8340 7890
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 8300 7268 8352 7274
rect 8300 7210 8352 7216
rect 8208 6860 8260 6866
rect 8208 6802 8260 6808
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8114 6216 8170 6225
rect 8114 6151 8170 6160
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 8036 4622 8064 6054
rect 8128 5846 8156 6151
rect 8116 5840 8168 5846
rect 8116 5782 8168 5788
rect 8208 5568 8260 5574
rect 8114 5536 8170 5545
rect 8208 5510 8260 5516
rect 8114 5471 8170 5480
rect 8128 5234 8156 5471
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 8128 4826 8156 5034
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 8036 3754 8064 4558
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8128 3942 8156 3975
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8036 3726 8156 3754
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8024 3460 8076 3466
rect 8024 3402 8076 3408
rect 7668 3097 7696 3334
rect 7760 3318 7880 3346
rect 7654 3088 7710 3097
rect 7654 3023 7710 3032
rect 7576 2910 7788 2938
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7288 1896 7340 1902
rect 7288 1838 7340 1844
rect 7392 800 7420 2790
rect 7576 2038 7604 2790
rect 7656 2440 7708 2446
rect 7654 2408 7656 2417
rect 7708 2408 7710 2417
rect 7654 2343 7710 2352
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7760 800 7788 2910
rect 7852 1766 7880 3318
rect 8036 2854 8064 3402
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 7840 1760 7892 1766
rect 7840 1702 7892 1708
rect 8128 800 8156 3726
rect 8220 3602 8248 5510
rect 8312 4146 8340 7210
rect 8404 5710 8432 11562
rect 8496 10810 8524 12786
rect 8588 11150 8616 16544
rect 9140 16572 9168 17138
rect 9088 16544 9168 16572
rect 9036 16526 9088 16532
rect 9232 16538 9260 18566
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9324 18086 9352 18362
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9416 17882 9444 18158
rect 9404 17876 9456 17882
rect 9404 17818 9456 17824
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9416 16658 9444 17274
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9232 16510 9444 16538
rect 8668 16448 8720 16454
rect 8668 16390 8720 16396
rect 8680 15094 8708 16390
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15706 9168 15846
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9128 15564 9180 15570
rect 9128 15506 9180 15512
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8680 11234 8708 14894
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8864 14006 8892 14554
rect 8852 14000 8904 14006
rect 8852 13942 8904 13948
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 8760 13252 8812 13258
rect 8760 13194 8812 13200
rect 8772 12646 8800 13194
rect 8760 12640 8812 12646
rect 8760 12582 8812 12588
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8944 12436 8996 12442
rect 8944 12378 8996 12384
rect 8956 11762 8984 12378
rect 9140 11898 9168 15506
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 9232 15026 9260 15438
rect 9416 15314 9444 16510
rect 9508 15434 9536 19246
rect 9772 18624 9824 18630
rect 9772 18566 9824 18572
rect 9680 17876 9732 17882
rect 9680 17818 9732 17824
rect 9692 17202 9720 17818
rect 9784 17542 9812 18566
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9588 17128 9640 17134
rect 9588 17070 9640 17076
rect 9496 15428 9548 15434
rect 9496 15370 9548 15376
rect 9416 15286 9536 15314
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 9232 13938 9260 14962
rect 9312 14544 9364 14550
rect 9312 14486 9364 14492
rect 9220 13932 9272 13938
rect 9220 13874 9272 13880
rect 9232 13394 9260 13874
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 9324 13274 9352 14486
rect 9232 13246 9352 13274
rect 9232 12442 9260 13246
rect 9508 12850 9536 15286
rect 9600 14006 9628 17070
rect 9680 16108 9732 16114
rect 9680 16050 9732 16056
rect 9692 15348 9720 16050
rect 9784 15473 9812 17478
rect 9770 15464 9826 15473
rect 9770 15399 9826 15408
rect 9692 15320 9812 15348
rect 9678 15192 9734 15201
rect 9678 15127 9680 15136
rect 9732 15127 9734 15136
rect 9680 15098 9732 15104
rect 9784 15026 9812 15320
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9772 15020 9824 15026
rect 9772 14962 9824 14968
rect 9692 14482 9720 14962
rect 9680 14476 9732 14482
rect 9680 14418 9732 14424
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9588 14000 9640 14006
rect 9692 13977 9720 14214
rect 9588 13942 9640 13948
rect 9678 13968 9734 13977
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9232 12102 9260 12378
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 8944 11756 8996 11762
rect 8944 11698 8996 11704
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 8680 11206 9076 11234
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8484 10804 8536 10810
rect 8484 10746 8536 10752
rect 8576 10736 8628 10742
rect 8680 10713 8708 11018
rect 8772 10742 8800 11086
rect 8760 10736 8812 10742
rect 8576 10678 8628 10684
rect 8666 10704 8722 10713
rect 8484 10600 8536 10606
rect 8484 10542 8536 10548
rect 8496 7002 8524 10542
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8482 6488 8538 6497
rect 8482 6423 8538 6432
rect 8496 6254 8524 6423
rect 8588 6390 8616 10678
rect 8760 10678 8812 10684
rect 8666 10639 8722 10648
rect 9048 10520 9076 11206
rect 9140 11150 9168 11834
rect 9404 11620 9456 11626
rect 9404 11562 9456 11568
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 9220 10804 9272 10810
rect 9220 10746 9272 10752
rect 9048 10492 9168 10520
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9722 9076 9862
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8668 9580 8720 9586
rect 9140 9568 9168 10492
rect 9232 9994 9260 10746
rect 9312 10124 9364 10130
rect 9312 10066 9364 10072
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9324 9654 9352 10066
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9140 9540 9260 9568
rect 8668 9522 8720 9528
rect 8680 8838 8708 9522
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8498 9076 8774
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8484 6248 8536 6254
rect 8484 6190 8536 6196
rect 8392 5704 8444 5710
rect 8588 5658 8616 6326
rect 8392 5646 8444 5652
rect 8496 5630 8616 5658
rect 8390 5400 8446 5409
rect 8390 5335 8446 5344
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8206 3496 8262 3505
rect 8206 3431 8262 3440
rect 8220 3058 8248 3431
rect 8312 3074 8340 4082
rect 8404 3210 8432 5335
rect 8496 3398 8524 5630
rect 8574 5536 8630 5545
rect 8574 5471 8630 5480
rect 8588 5234 8616 5471
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8576 5092 8628 5098
rect 8576 5034 8628 5040
rect 8588 3641 8616 5034
rect 8574 3632 8630 3641
rect 8574 3567 8630 3576
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8588 3346 8616 3567
rect 8680 3534 8708 8298
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8772 7206 8800 8026
rect 9232 8022 9260 9540
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9048 7857 9076 7958
rect 9220 7880 9272 7886
rect 9034 7848 9090 7857
rect 9220 7822 9272 7828
rect 9034 7783 9090 7792
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8760 7200 8812 7206
rect 8760 7142 8812 7148
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8760 6384 8812 6390
rect 8760 6326 8812 6332
rect 8772 6186 8800 6326
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 9140 5953 9168 7686
rect 9232 7410 9260 7822
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9232 7002 9260 7346
rect 9220 6996 9272 7002
rect 9220 6938 9272 6944
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9232 6118 9260 6190
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9126 5944 9182 5953
rect 9126 5879 9182 5888
rect 9128 5840 9180 5846
rect 9324 5794 9352 7754
rect 9128 5782 9180 5788
rect 9140 5681 9168 5782
rect 9232 5766 9352 5794
rect 9416 5794 9444 11562
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9508 10577 9536 11494
rect 9494 10568 9550 10577
rect 9494 10503 9550 10512
rect 9496 10056 9548 10062
rect 9496 9998 9548 10004
rect 9508 9518 9536 9998
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9508 8974 9536 9454
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9508 7970 9536 8502
rect 9600 8090 9628 13942
rect 9678 13903 9734 13912
rect 9784 13512 9812 14962
rect 9683 13484 9812 13512
rect 9683 13138 9711 13484
rect 9772 13184 9824 13190
rect 9683 13110 9720 13138
rect 9876 13172 9904 19246
rect 10048 18828 10100 18834
rect 10048 18770 10100 18776
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9968 17678 9996 18226
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10060 17542 10088 18770
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10140 17060 10192 17066
rect 10140 17002 10192 17008
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9968 13569 9996 16730
rect 10152 16182 10180 17002
rect 10140 16176 10192 16182
rect 10140 16118 10192 16124
rect 10244 15706 10272 17682
rect 10416 17128 10468 17134
rect 10414 17096 10416 17105
rect 10468 17096 10470 17105
rect 10414 17031 10470 17040
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 16182 10456 16390
rect 10416 16176 10468 16182
rect 10416 16118 10468 16124
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10048 14816 10100 14822
rect 10100 14776 10180 14804
rect 10048 14758 10100 14764
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 9954 13560 10010 13569
rect 9954 13495 10010 13504
rect 9824 13144 9904 13172
rect 9772 13126 9824 13132
rect 9692 11354 9720 13110
rect 9784 12617 9812 13126
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9770 12608 9826 12617
rect 9770 12543 9826 12552
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9876 9654 9904 12854
rect 10060 12434 10088 14282
rect 9968 12406 10088 12434
rect 10152 12434 10180 14776
rect 10244 14634 10272 15642
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10322 15192 10378 15201
rect 10322 15127 10378 15136
rect 10336 15026 10364 15127
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10244 14606 10364 14634
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10244 14074 10272 14418
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10244 12918 10272 13194
rect 10336 12918 10364 14606
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10152 12406 10364 12434
rect 9864 9648 9916 9654
rect 9864 9590 9916 9596
rect 9968 8650 9996 12406
rect 10336 12170 10364 12406
rect 10324 12164 10376 12170
rect 10324 12106 10376 12112
rect 10232 11348 10284 11354
rect 10232 11290 10284 11296
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9692 8622 9996 8650
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9508 7942 9628 7970
rect 9600 7818 9628 7942
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 5846 9628 7754
rect 9588 5840 9640 5846
rect 9416 5766 9536 5794
rect 9588 5782 9640 5788
rect 9126 5672 9182 5681
rect 8944 5636 8996 5642
rect 9126 5607 9182 5616
rect 8944 5578 8996 5584
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 5137 8800 5510
rect 8956 5234 8984 5578
rect 9232 5250 9260 5766
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 8944 5228 8996 5234
rect 9232 5222 9352 5250
rect 9416 5234 9444 5646
rect 8944 5170 8996 5176
rect 8758 5128 8814 5137
rect 8758 5063 8814 5072
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8956 4486 8984 4762
rect 8944 4480 8996 4486
rect 8944 4422 8996 4428
rect 8944 4208 8996 4214
rect 8942 4176 8944 4185
rect 9140 4185 9168 4966
rect 8996 4176 8998 4185
rect 8942 4111 8998 4120
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 8852 4072 8904 4078
rect 8944 4072 8996 4078
rect 8852 4014 8904 4020
rect 8942 4040 8944 4049
rect 8996 4040 8998 4049
rect 8864 3942 8892 4014
rect 8942 3975 8998 3984
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8760 3596 8812 3602
rect 8760 3538 8812 3544
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8772 3346 8800 3538
rect 9128 3528 9180 3534
rect 8942 3496 8998 3505
rect 9128 3470 9180 3476
rect 8942 3431 8998 3440
rect 8956 3398 8984 3431
rect 8588 3318 8800 3346
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8666 3224 8722 3233
rect 8404 3182 8616 3210
rect 8208 3052 8260 3058
rect 8312 3046 8524 3074
rect 8208 2994 8260 3000
rect 8300 2984 8352 2990
rect 8206 2952 8262 2961
rect 8392 2984 8444 2990
rect 8352 2944 8392 2972
rect 8300 2926 8352 2932
rect 8392 2926 8444 2932
rect 8206 2887 8262 2896
rect 8220 2514 8248 2887
rect 8300 2848 8352 2854
rect 8300 2790 8352 2796
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8312 2281 8340 2790
rect 8392 2304 8444 2310
rect 8298 2272 8354 2281
rect 8392 2246 8444 2252
rect 8298 2207 8354 2216
rect 8404 1970 8432 2246
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8496 800 8524 3046
rect 8588 2854 8616 3182
rect 8666 3159 8668 3168
rect 8720 3159 8722 3168
rect 8668 3130 8720 3136
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 9140 2774 9168 3470
rect 9232 3058 9260 5034
rect 9324 4162 9352 5222
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 9416 4826 9444 5170
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9324 4134 9444 4162
rect 9310 4040 9366 4049
rect 9310 3975 9312 3984
rect 9364 3975 9366 3984
rect 9312 3946 9364 3952
rect 9416 3942 9444 4134
rect 9404 3936 9456 3942
rect 9404 3878 9456 3884
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9416 3505 9444 3538
rect 9402 3496 9458 3505
rect 9402 3431 9458 3440
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 9140 2746 9260 2774
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8574 2680 8630 2689
rect 8747 2683 9055 2692
rect 8630 2638 8708 2666
rect 8574 2615 8630 2624
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8588 2106 8616 2382
rect 8680 2378 8708 2638
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8956 2310 8984 2586
rect 8852 2304 8904 2310
rect 8852 2246 8904 2252
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8864 1698 8892 2246
rect 8852 1692 8904 1698
rect 8852 1634 8904 1640
rect 8864 800 8892 1634
rect 9232 800 9260 2746
rect 9324 2582 9352 3334
rect 9508 3126 9536 5766
rect 9588 4752 9640 4758
rect 9588 4694 9640 4700
rect 9600 4593 9628 4694
rect 9586 4584 9642 4593
rect 9586 4519 9642 4528
rect 9588 3936 9640 3942
rect 9588 3878 9640 3884
rect 9600 3602 9628 3878
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9324 2038 9352 2518
rect 9508 2394 9536 3062
rect 9692 2961 9720 8622
rect 9956 8560 10008 8566
rect 9956 8502 10008 8508
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9784 6798 9812 7278
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9772 6792 9824 6798
rect 9772 6734 9824 6740
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9784 5778 9812 6598
rect 9876 6322 9904 6938
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9772 5772 9824 5778
rect 9824 5732 9904 5760
rect 9772 5714 9824 5720
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9784 4010 9812 4422
rect 9772 4004 9824 4010
rect 9772 3946 9824 3952
rect 9784 3126 9812 3946
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9678 2952 9734 2961
rect 9678 2887 9734 2896
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9772 2848 9824 2854
rect 9876 2836 9904 5732
rect 9968 2990 9996 8502
rect 10060 8090 10088 9114
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10060 7886 10088 8026
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 10060 5642 10088 7142
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10048 5636 10100 5642
rect 10048 5578 10100 5584
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 10060 4729 10088 5170
rect 10046 4720 10102 4729
rect 10046 4655 10102 4664
rect 10152 4554 10180 6666
rect 10244 5574 10272 11290
rect 10336 10810 10364 12106
rect 10428 11937 10456 15574
rect 10520 14414 10548 19858
rect 11256 19718 11284 19858
rect 11808 19825 11836 19858
rect 12544 19854 12572 20198
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12532 19848 12584 19854
rect 11794 19816 11850 19825
rect 12532 19790 12584 19796
rect 11794 19751 11850 19760
rect 11244 19712 11296 19718
rect 11244 19654 11296 19660
rect 11704 19712 11756 19718
rect 11704 19654 11756 19660
rect 10968 18216 11020 18222
rect 10968 18158 11020 18164
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 10692 17536 10744 17542
rect 10690 17504 10692 17513
rect 10744 17504 10746 17513
rect 10690 17439 10746 17448
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10704 16590 10732 17274
rect 10796 16998 10824 18090
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 16584 10744 16590
rect 10692 16526 10744 16532
rect 10704 16250 10732 16526
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10888 15910 10916 17750
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10876 15904 10928 15910
rect 10876 15846 10928 15852
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10520 13530 10548 14350
rect 10612 14090 10640 15846
rect 10796 15502 10824 15846
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10704 14278 10732 15370
rect 10796 15162 10824 15438
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10796 14890 10824 15098
rect 10784 14884 10836 14890
rect 10784 14826 10836 14832
rect 10980 14346 11008 18158
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17338 11192 17478
rect 11152 17332 11204 17338
rect 11152 17274 11204 17280
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 10968 14340 11020 14346
rect 10968 14282 11020 14288
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10612 14062 10732 14090
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10600 12708 10652 12714
rect 10600 12650 10652 12656
rect 10612 12434 10640 12650
rect 10520 12406 10640 12434
rect 10414 11928 10470 11937
rect 10414 11863 10470 11872
rect 10414 11656 10470 11665
rect 10520 11642 10548 12406
rect 10598 12200 10654 12209
rect 10598 12135 10654 12144
rect 10612 11830 10640 12135
rect 10600 11824 10652 11830
rect 10600 11766 10652 11772
rect 10612 11665 10640 11766
rect 10470 11614 10548 11642
rect 10414 11591 10470 11600
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10520 10674 10548 11614
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10704 10538 10732 14062
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 12209 10824 13874
rect 10888 13802 10916 14010
rect 10980 13870 11008 14282
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13796 10928 13802
rect 10876 13738 10928 13744
rect 10888 13530 10916 13738
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10888 12986 10916 13466
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10876 12980 10928 12986
rect 10876 12922 10928 12928
rect 10888 12238 10916 12922
rect 10980 12730 11008 13126
rect 11072 12918 11100 17138
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16726 11192 16934
rect 11152 16720 11204 16726
rect 11152 16662 11204 16668
rect 11256 16572 11284 19654
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11716 19514 11744 19654
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 12348 19304 12400 19310
rect 12348 19246 12400 19252
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18970 11928 19110
rect 11888 18964 11940 18970
rect 11888 18906 11940 18912
rect 12072 18896 12124 18902
rect 12072 18838 12124 18844
rect 11980 18828 12032 18834
rect 11980 18770 12032 18776
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11518 17640 11574 17649
rect 11518 17575 11574 17584
rect 11532 17542 11560 17575
rect 11520 17536 11572 17542
rect 11520 17478 11572 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17371 11654 17380
rect 11716 16810 11744 18566
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11900 17134 11928 18158
rect 11796 17128 11848 17134
rect 11794 17096 11796 17105
rect 11888 17128 11940 17134
rect 11848 17096 11850 17105
rect 11888 17070 11940 17076
rect 11794 17031 11850 17040
rect 11164 16544 11284 16572
rect 11532 16782 11744 16810
rect 11060 12912 11112 12918
rect 11060 12854 11112 12860
rect 10980 12702 11100 12730
rect 10876 12232 10928 12238
rect 10782 12200 10838 12209
rect 10876 12174 10928 12180
rect 10782 12135 10838 12144
rect 10888 11694 10916 12174
rect 11072 11830 11100 12702
rect 11164 12073 11192 16544
rect 11532 16454 11560 16782
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11520 16448 11572 16454
rect 11520 16390 11572 16396
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11244 16108 11296 16114
rect 11244 16050 11296 16056
rect 11256 15434 11284 16050
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11150 12064 11206 12073
rect 11150 11999 11206 12008
rect 11256 11914 11284 15030
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11440 14498 11468 14758
rect 11624 14634 11652 14894
rect 11532 14618 11652 14634
rect 11716 14618 11744 16594
rect 11520 14612 11652 14618
rect 11572 14606 11652 14612
rect 11704 14612 11756 14618
rect 11520 14554 11572 14560
rect 11704 14554 11756 14560
rect 11808 14550 11836 17031
rect 11992 16794 12020 18770
rect 12084 18426 12112 18838
rect 12360 18766 12388 19246
rect 12348 18760 12400 18766
rect 12348 18702 12400 18708
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12544 18222 12572 19790
rect 12716 18624 12768 18630
rect 12716 18566 12768 18572
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12532 18216 12584 18222
rect 12532 18158 12584 18164
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 12084 16538 12112 17478
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 11900 16510 12112 16538
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 11900 15484 11928 16510
rect 12072 15904 12124 15910
rect 12072 15846 12124 15852
rect 12084 15638 12112 15846
rect 11980 15632 12032 15638
rect 11978 15600 11980 15609
rect 12072 15632 12124 15638
rect 12032 15600 12034 15609
rect 12072 15574 12124 15580
rect 11978 15535 12034 15544
rect 11900 15456 12020 15484
rect 11888 15360 11940 15366
rect 11886 15328 11888 15337
rect 11940 15328 11942 15337
rect 11886 15263 11942 15272
rect 11992 15178 12020 15456
rect 11900 15150 12020 15178
rect 11796 14544 11848 14550
rect 11440 14470 11744 14498
rect 11796 14486 11848 14492
rect 11716 14362 11744 14470
rect 11900 14362 11928 15150
rect 11980 14816 12032 14822
rect 11980 14758 12032 14764
rect 11716 14334 11928 14362
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11612 13184 11664 13190
rect 11716 13172 11744 14334
rect 11888 14000 11940 14006
rect 11888 13942 11940 13948
rect 11900 13530 11928 13942
rect 11992 13841 12020 14758
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 11978 13832 12034 13841
rect 11978 13767 12034 13776
rect 12084 13734 12112 14214
rect 12072 13728 12124 13734
rect 12072 13670 12124 13676
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11664 13144 11744 13172
rect 11796 13184 11848 13190
rect 11612 13126 11664 13132
rect 11796 13126 11848 13132
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11704 12912 11756 12918
rect 11808 12889 11836 13126
rect 11704 12854 11756 12860
rect 11794 12880 11850 12889
rect 11518 12608 11574 12617
rect 11518 12543 11574 12552
rect 11532 12442 11560 12543
rect 11520 12436 11572 12442
rect 11520 12378 11572 12384
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11164 11886 11284 11914
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11144 10836 11150
rect 10888 11132 10916 11630
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 11072 11218 11100 11494
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 10836 11104 10916 11132
rect 10784 11086 10836 11092
rect 10796 11014 10824 11086
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10692 10532 10744 10538
rect 10692 10474 10744 10480
rect 10416 10464 10468 10470
rect 10416 10406 10468 10412
rect 10428 10130 10456 10406
rect 10704 10198 10732 10474
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10324 6112 10376 6118
rect 10324 6054 10376 6060
rect 10232 5568 10284 5574
rect 10232 5510 10284 5516
rect 10140 4548 10192 4554
rect 10140 4490 10192 4496
rect 9956 2984 10008 2990
rect 9956 2926 10008 2932
rect 9824 2808 9904 2836
rect 9772 2790 9824 2796
rect 9600 2514 9628 2790
rect 9770 2680 9826 2689
rect 9770 2615 9826 2624
rect 9784 2582 9812 2615
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 9680 2440 9732 2446
rect 9508 2366 9628 2394
rect 9680 2382 9732 2388
rect 9312 2032 9364 2038
rect 9312 1974 9364 1980
rect 9600 800 9628 2366
rect 9692 1630 9720 2382
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9680 1624 9732 1630
rect 9680 1566 9732 1572
rect 9876 1562 9904 2314
rect 9864 1556 9916 1562
rect 9864 1498 9916 1504
rect 9968 800 9996 2926
rect 10336 2446 10364 6054
rect 10428 4826 10456 10066
rect 10704 7750 10732 10134
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10796 9178 10824 9590
rect 11072 9450 11100 11154
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10782 8936 10838 8945
rect 10782 8871 10838 8880
rect 10692 7744 10744 7750
rect 10692 7686 10744 7692
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6112 10560 6118
rect 10508 6054 10560 6060
rect 10520 5817 10548 6054
rect 10506 5808 10562 5817
rect 10506 5743 10562 5752
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10612 4690 10640 6938
rect 10692 6248 10744 6254
rect 10692 6190 10744 6196
rect 10704 5137 10732 6190
rect 10690 5128 10746 5137
rect 10690 5063 10746 5072
rect 10796 5030 10824 8871
rect 10888 8430 10916 9114
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10980 8566 11008 8842
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11072 8362 11100 8774
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10888 6322 10916 7482
rect 11072 7206 11100 8298
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11072 6798 11100 7142
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11072 6662 11100 6734
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10876 6316 10928 6322
rect 10876 6258 10928 6264
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10600 4684 10652 4690
rect 10600 4626 10652 4632
rect 10692 4548 10744 4554
rect 10692 4490 10744 4496
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10336 800 10364 2382
rect 10520 1834 10548 3334
rect 10612 3058 10640 4150
rect 10704 3670 10732 4490
rect 10796 4457 10824 4966
rect 10888 4486 10916 6258
rect 11072 6118 11100 6598
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 10968 5840 11020 5846
rect 10966 5808 10968 5817
rect 11020 5808 11022 5817
rect 10966 5743 11022 5752
rect 11072 5710 11100 6054
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 11072 5370 11100 5646
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10876 4480 10928 4486
rect 10782 4448 10838 4457
rect 10876 4422 10928 4428
rect 10782 4383 10838 4392
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10980 3534 11008 5306
rect 11164 4162 11192 11886
rect 11716 11354 11744 12854
rect 11794 12815 11850 12824
rect 12176 11830 12204 16526
rect 12544 16454 12572 17070
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12440 15564 12492 15570
rect 12440 15506 12492 15512
rect 12256 14544 12308 14550
rect 12308 14504 12388 14532
rect 12256 14486 12308 14492
rect 12360 13938 12388 14504
rect 12256 13932 12308 13938
rect 12256 13874 12308 13880
rect 12348 13932 12400 13938
rect 12348 13874 12400 13880
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11244 11008 11296 11014
rect 11244 10950 11296 10956
rect 11256 10742 11284 10950
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10470 11284 10678
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11256 10062 11284 10406
rect 11796 10124 11848 10130
rect 11796 10066 11848 10072
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11256 9926 11284 9998
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11256 9654 11284 9862
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11532 9382 11560 9590
rect 11702 9480 11758 9489
rect 11702 9415 11758 9424
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 11520 9376 11572 9382
rect 11520 9318 11572 9324
rect 11256 8616 11284 9318
rect 11532 8974 11560 9318
rect 11716 9042 11744 9415
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11520 8968 11572 8974
rect 11520 8910 11572 8916
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11256 8588 11376 8616
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11256 4282 11284 8434
rect 11348 8430 11376 8588
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11520 6248 11572 6254
rect 11716 6225 11744 8978
rect 11808 8401 11836 10066
rect 11794 8392 11850 8401
rect 11794 8327 11850 8336
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11808 6497 11836 6666
rect 11794 6488 11850 6497
rect 11794 6423 11850 6432
rect 11796 6384 11848 6390
rect 11796 6326 11848 6332
rect 11520 6190 11572 6196
rect 11702 6216 11758 6225
rect 11532 6118 11560 6190
rect 11702 6151 11758 6160
rect 11520 6112 11572 6118
rect 11808 6089 11836 6326
rect 11520 6054 11572 6060
rect 11794 6080 11850 6089
rect 11794 6015 11850 6024
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11336 5024 11388 5030
rect 11334 4992 11336 5001
rect 11388 4992 11390 5001
rect 11334 4927 11390 4936
rect 11716 4622 11744 5510
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11808 5030 11836 5306
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4690 11836 4966
rect 11796 4684 11848 4690
rect 11796 4626 11848 4632
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11336 4276 11388 4282
rect 11336 4218 11388 4224
rect 11164 4134 11284 4162
rect 11152 4072 11204 4078
rect 11072 4032 11152 4060
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 11072 2650 11100 4032
rect 11152 4014 11204 4020
rect 11256 3890 11284 4134
rect 11164 3862 11284 3890
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10598 2544 10654 2553
rect 10598 2479 10654 2488
rect 10612 2446 10640 2479
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 11060 2100 11112 2106
rect 11060 2042 11112 2048
rect 10508 1828 10560 1834
rect 10508 1770 10560 1776
rect 10692 1556 10744 1562
rect 10692 1498 10744 1504
rect 10704 800 10732 1498
rect 11072 800 11100 2042
rect 11164 1698 11192 3862
rect 11348 3754 11376 4218
rect 11808 4078 11836 4626
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11900 3942 11928 11018
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11992 9081 12020 9551
rect 11978 9072 12034 9081
rect 11978 9007 12034 9016
rect 11992 8566 12020 9007
rect 11980 8560 12032 8566
rect 11980 8502 12032 8508
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11256 3726 11376 3754
rect 11256 1714 11284 3726
rect 11992 3466 12020 8366
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 11336 3120 11388 3126
rect 11336 3062 11388 3068
rect 11348 2650 11376 3062
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11980 2508 12032 2514
rect 11980 2450 12032 2456
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11808 2310 11836 2382
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11152 1692 11204 1698
rect 11152 1634 11204 1640
rect 11256 1686 11468 1714
rect 11256 1630 11284 1686
rect 11244 1624 11296 1630
rect 11244 1566 11296 1572
rect 11440 800 11468 1686
rect 11808 800 11836 2246
rect 11900 2038 11928 2246
rect 11888 2032 11940 2038
rect 11992 2009 12020 2450
rect 12084 2106 12112 11086
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12176 7750 12204 8774
rect 12164 7744 12216 7750
rect 12164 7686 12216 7692
rect 12268 7562 12296 13874
rect 12452 13734 12480 15506
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13258 12480 13670
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12346 13152 12402 13161
rect 12346 13087 12402 13096
rect 12360 11506 12388 13087
rect 12544 11801 12572 16390
rect 12624 15904 12676 15910
rect 12624 15846 12676 15852
rect 12636 13682 12664 15846
rect 12728 15502 12756 18566
rect 12820 18426 12848 18566
rect 12808 18420 12860 18426
rect 12808 18362 12860 18368
rect 12808 16652 12860 16658
rect 12808 16594 12860 16600
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12820 15162 12848 16594
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12716 14816 12768 14822
rect 12716 14758 12768 14764
rect 12728 13841 12756 14758
rect 12714 13832 12770 13841
rect 12714 13767 12770 13776
rect 12636 13654 12756 13682
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12530 11792 12586 11801
rect 12530 11727 12586 11736
rect 12360 11478 12480 11506
rect 12452 9654 12480 11478
rect 12636 11286 12664 12378
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12346 8936 12402 8945
rect 12346 8871 12402 8880
rect 12360 8838 12388 8871
rect 12348 8832 12400 8838
rect 12348 8774 12400 8780
rect 12440 8832 12492 8838
rect 12440 8774 12492 8780
rect 12452 8566 12480 8774
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12440 8356 12492 8362
rect 12440 8298 12492 8304
rect 12348 7880 12400 7886
rect 12348 7822 12400 7828
rect 12176 7534 12296 7562
rect 12176 7313 12204 7534
rect 12360 7478 12388 7822
rect 12452 7478 12480 8298
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12162 7304 12218 7313
rect 12268 7290 12296 7414
rect 12268 7262 12388 7290
rect 12162 7239 12218 7248
rect 12164 7200 12216 7206
rect 12164 7142 12216 7148
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12176 5778 12204 7142
rect 12268 7002 12296 7142
rect 12360 7002 12388 7262
rect 12256 6996 12308 7002
rect 12256 6938 12308 6944
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12176 4214 12204 5714
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12360 5166 12388 5238
rect 12348 5160 12400 5166
rect 12348 5102 12400 5108
rect 12544 4706 12572 11154
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12636 10674 12664 11086
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12636 8362 12664 8570
rect 12624 8356 12676 8362
rect 12624 8298 12676 8304
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12636 6458 12664 7346
rect 12624 6452 12676 6458
rect 12624 6394 12676 6400
rect 12624 5160 12676 5166
rect 12624 5102 12676 5108
rect 12360 4678 12572 4706
rect 12164 4208 12216 4214
rect 12164 4150 12216 4156
rect 12256 4140 12308 4146
rect 12256 4082 12308 4088
rect 12164 3460 12216 3466
rect 12164 3402 12216 3408
rect 12072 2100 12124 2106
rect 12072 2042 12124 2048
rect 11888 1974 11940 1980
rect 11978 2000 12034 2009
rect 11978 1935 12034 1944
rect 12176 800 12204 3402
rect 12268 2446 12296 4082
rect 12360 3641 12388 4678
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12452 3482 12480 3538
rect 12360 3454 12480 3482
rect 12360 3126 12388 3454
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12636 3058 12664 5102
rect 12624 3052 12676 3058
rect 12624 2994 12676 3000
rect 12728 2689 12756 13654
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12820 12374 12848 13466
rect 12808 12368 12860 12374
rect 12808 12310 12860 12316
rect 12820 9674 12848 12310
rect 12912 11218 12940 19926
rect 13004 19854 13032 20198
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 12992 19848 13044 19854
rect 12992 19790 13044 19796
rect 13004 19174 13032 19790
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 14556 19712 14608 19718
rect 14556 19654 14608 19660
rect 13188 19446 13216 19654
rect 14370 19544 14426 19553
rect 14370 19479 14372 19488
rect 14424 19479 14426 19488
rect 14372 19450 14424 19456
rect 13176 19440 13228 19446
rect 14568 19417 14596 19654
rect 13176 19382 13228 19388
rect 14554 19408 14610 19417
rect 14464 19372 14516 19378
rect 14554 19343 14610 19352
rect 14464 19314 14516 19320
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 13084 19168 13136 19174
rect 13084 19110 13136 19116
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 18086 13032 18226
rect 12992 18080 13044 18086
rect 12992 18022 13044 18028
rect 13096 17882 13124 19110
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14476 18970 14504 19314
rect 14660 19258 14688 20266
rect 15016 19984 15068 19990
rect 15200 19984 15252 19990
rect 15068 19932 15200 19938
rect 15016 19926 15252 19932
rect 16212 19984 16264 19990
rect 16212 19926 16264 19932
rect 14740 19916 14792 19922
rect 15028 19910 15240 19926
rect 14740 19858 14792 19864
rect 14568 19230 14688 19258
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13188 18358 13216 18566
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13648 18290 13676 18362
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16590 13032 16934
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13372 15978 13400 18022
rect 13452 17536 13504 17542
rect 13452 17478 13504 17484
rect 13464 16574 13492 17478
rect 13464 16546 13584 16574
rect 13452 16448 13504 16454
rect 13452 16390 13504 16396
rect 13176 15972 13228 15978
rect 13176 15914 13228 15920
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13004 14958 13032 15438
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12992 14816 13044 14822
rect 12992 14758 13044 14764
rect 13084 14816 13136 14822
rect 13084 14758 13136 14764
rect 13004 14521 13032 14758
rect 12990 14512 13046 14521
rect 12990 14447 13046 14456
rect 13096 14278 13124 14758
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 13082 13560 13138 13569
rect 13188 13530 13216 15914
rect 13464 13818 13492 16390
rect 13556 13954 13584 16546
rect 13648 16114 13676 18226
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15706 13676 16050
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13728 15156 13780 15162
rect 13728 15098 13780 15104
rect 13556 13926 13676 13954
rect 13740 13938 13768 15098
rect 13832 14618 13860 15370
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13820 14272 13872 14278
rect 13820 14214 13872 14220
rect 13832 14006 13860 14214
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13464 13790 13584 13818
rect 13082 13495 13138 13504
rect 13176 13524 13228 13530
rect 13096 13410 13124 13495
rect 13176 13466 13228 13472
rect 13096 13382 13216 13410
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12481 13032 13126
rect 12990 12472 13046 12481
rect 12990 12407 13046 12416
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12820 9646 12940 9674
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 12820 7002 12848 7958
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12808 6384 12860 6390
rect 12808 6326 12860 6332
rect 12820 6089 12848 6326
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12912 5658 12940 9646
rect 13096 5930 13124 13194
rect 13188 12918 13216 13382
rect 13176 12912 13228 12918
rect 13176 12854 13228 12860
rect 13188 11898 13216 12854
rect 13556 12434 13584 13790
rect 13648 12442 13676 13926
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13740 12782 13768 13126
rect 13728 12776 13780 12782
rect 13728 12718 13780 12724
rect 13464 12406 13584 12434
rect 13636 12436 13688 12442
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13268 11824 13320 11830
rect 13268 11766 13320 11772
rect 13280 11082 13308 11766
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10674 13400 10950
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13004 5902 13124 5930
rect 13004 5681 13032 5902
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 13266 5808 13322 5817
rect 12820 5630 12940 5658
rect 12990 5672 13046 5681
rect 12820 5001 12848 5630
rect 12990 5607 13046 5616
rect 12900 5568 12952 5574
rect 12900 5510 12952 5516
rect 12806 4992 12862 5001
rect 12806 4927 12862 4936
rect 12912 3534 12940 5510
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3670 13032 3878
rect 12992 3664 13044 3670
rect 12992 3606 13044 3612
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12714 2680 12770 2689
rect 12714 2615 12770 2624
rect 13096 2514 13124 5782
rect 13266 5743 13322 5752
rect 13280 2990 13308 5743
rect 13358 5672 13414 5681
rect 13358 5607 13414 5616
rect 13372 3777 13400 5607
rect 13358 3768 13414 3777
rect 13358 3703 13414 3712
rect 13464 3534 13492 12406
rect 13636 12378 13688 12384
rect 13740 12170 13768 12718
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 12374 13860 12582
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12368 13872 12374
rect 13820 12310 13872 12316
rect 14280 12368 14332 12374
rect 14280 12310 14332 12316
rect 14004 12232 14056 12238
rect 14004 12174 14056 12180
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13728 12164 13780 12170
rect 13728 12106 13780 12112
rect 13556 11898 13584 12106
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13556 11354 13584 11834
rect 14016 11642 14044 12174
rect 14292 12102 14320 12310
rect 14280 12096 14332 12102
rect 14280 12038 14332 12044
rect 14384 11762 14412 18770
rect 14568 15337 14596 19230
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14660 18698 14688 18906
rect 14648 18692 14700 18698
rect 14648 18634 14700 18640
rect 14554 15328 14610 15337
rect 14554 15263 14610 15272
rect 14752 14890 14780 19858
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 14844 19514 14872 19790
rect 15948 19718 15976 19790
rect 16224 19786 16252 19926
rect 16212 19780 16264 19786
rect 16212 19722 16264 19728
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 14832 19508 14884 19514
rect 14832 19450 14884 19456
rect 15476 19304 15528 19310
rect 15476 19246 15528 19252
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15028 16250 15056 18566
rect 15212 18426 15240 18566
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 17377 15148 17478
rect 15106 17368 15162 17377
rect 15304 17338 15332 18362
rect 15106 17303 15162 17312
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 16652 15160 16658
rect 15108 16594 15160 16600
rect 15016 16244 15068 16250
rect 15016 16186 15068 16192
rect 15120 15042 15148 16594
rect 15212 15366 15240 17070
rect 15292 16516 15344 16522
rect 15292 16458 15344 16464
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14844 15014 15148 15042
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14464 14476 14516 14482
rect 14464 14418 14516 14424
rect 14476 14074 14504 14418
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14476 12102 14504 12786
rect 14844 12646 14872 15014
rect 15016 14884 15068 14890
rect 15016 14826 15068 14832
rect 14924 14816 14976 14822
rect 14924 14758 14976 14764
rect 14936 14414 14964 14758
rect 14924 14408 14976 14414
rect 14924 14350 14976 14356
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14936 12434 14964 12786
rect 14660 12406 14964 12434
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 11756 14424 11762
rect 14372 11698 14424 11704
rect 14016 11614 14412 11642
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13832 9926 13860 10202
rect 14096 9988 14148 9994
rect 14096 9930 14148 9936
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13832 9654 13860 9862
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13740 9178 13768 9590
rect 14108 9450 14136 9930
rect 14292 9489 14320 10406
rect 14278 9480 14334 9489
rect 14096 9444 14148 9450
rect 14278 9415 14334 9424
rect 14096 9386 14148 9392
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13832 8634 13860 8978
rect 13820 8628 13872 8634
rect 13820 8570 13872 8576
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 14280 7744 14332 7750
rect 14280 7686 14332 7692
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13648 6866 13676 7346
rect 13636 6860 13688 6866
rect 13636 6802 13688 6808
rect 13648 6458 13676 6802
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13740 6225 13768 7686
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 13820 6792 13872 6798
rect 13820 6734 13872 6740
rect 13726 6216 13782 6225
rect 13726 6151 13782 6160
rect 13832 5846 13860 6734
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 13820 5840 13872 5846
rect 13820 5782 13872 5788
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 14188 5568 14240 5574
rect 14188 5510 14240 5516
rect 13542 4720 13598 4729
rect 13542 4655 13598 4664
rect 13556 3942 13584 4655
rect 13648 4026 13676 5510
rect 14200 5302 14228 5510
rect 14292 5302 14320 7686
rect 14384 7313 14412 11614
rect 14476 9994 14504 12038
rect 14554 11656 14610 11665
rect 14554 11591 14610 11600
rect 14464 9988 14516 9994
rect 14464 9930 14516 9936
rect 14568 9450 14596 11591
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14370 7304 14426 7313
rect 14370 7239 14426 7248
rect 14476 7177 14504 9318
rect 14660 8090 14688 12406
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 14660 7834 14688 8026
rect 14660 7806 14780 7834
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14462 7168 14518 7177
rect 14462 7103 14518 7112
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14568 6118 14596 6258
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14372 5636 14424 5642
rect 14372 5578 14424 5584
rect 14188 5296 14240 5302
rect 14188 5238 14240 5244
rect 14280 5296 14332 5302
rect 14280 5238 14332 5244
rect 14280 5092 14332 5098
rect 14280 5034 14332 5040
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 13728 4480 13780 4486
rect 13728 4422 13780 4428
rect 13740 4146 13768 4422
rect 13910 4176 13966 4185
rect 13728 4140 13780 4146
rect 13910 4111 13966 4120
rect 13728 4082 13780 4088
rect 13648 3998 13768 4026
rect 13924 4010 13952 4111
rect 14292 4078 14320 5034
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14384 4010 14412 5578
rect 13544 3936 13596 3942
rect 13544 3878 13596 3884
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13648 2990 13676 3674
rect 13268 2984 13320 2990
rect 13188 2932 13268 2938
rect 13452 2984 13504 2990
rect 13188 2926 13320 2932
rect 13358 2952 13414 2961
rect 13188 2910 13308 2926
rect 13188 2553 13216 2910
rect 13452 2926 13504 2932
rect 13636 2984 13688 2990
rect 13740 2961 13768 3998
rect 13912 4004 13964 4010
rect 13912 3946 13964 3952
rect 14372 4004 14424 4010
rect 14372 3946 14424 3952
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14292 3738 14320 3878
rect 14370 3768 14426 3777
rect 14280 3732 14332 3738
rect 14370 3703 14372 3712
rect 14280 3674 14332 3680
rect 14424 3703 14426 3712
rect 14372 3674 14424 3680
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13636 2926 13688 2932
rect 13726 2952 13782 2961
rect 13358 2887 13414 2896
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13174 2544 13230 2553
rect 13084 2508 13136 2514
rect 13174 2479 13230 2488
rect 13084 2450 13136 2456
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12254 2136 12310 2145
rect 12254 2071 12310 2080
rect 12268 1873 12296 2071
rect 12254 1864 12310 1873
rect 12254 1799 12310 1808
rect 12636 1630 12664 2246
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 12624 1624 12676 1630
rect 12624 1566 12676 1572
rect 12532 1420 12584 1426
rect 12532 1362 12584 1368
rect 12544 800 12572 1362
rect 12912 800 12940 1906
rect 13280 800 13308 2790
rect 13372 2514 13400 2887
rect 13464 2650 13492 2926
rect 13726 2887 13782 2896
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13360 2508 13412 2514
rect 13360 2450 13412 2456
rect 13636 2508 13688 2514
rect 13636 2450 13688 2456
rect 13648 800 13676 2450
rect 13832 1902 13860 3538
rect 13910 3224 13966 3233
rect 13910 3159 13912 3168
rect 13964 3159 13966 3168
rect 13912 3130 13964 3136
rect 14096 3120 14148 3126
rect 14094 3088 14096 3097
rect 14148 3088 14150 3097
rect 14094 3023 14150 3032
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 13912 2304 13964 2310
rect 13912 2246 13964 2252
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 13924 1426 13952 2246
rect 14108 2038 14136 2382
rect 14096 2032 14148 2038
rect 14096 1974 14148 1980
rect 13912 1420 13964 1426
rect 13912 1362 13964 1368
rect 14016 870 14136 898
rect 14016 800 14044 870
rect 6012 734 6224 762
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7378 0 7434 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 9954 0 10010 800
rect 10322 0 10378 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12530 0 12586 800
rect 12898 0 12954 800
rect 13266 0 13322 800
rect 13634 0 13690 800
rect 14002 0 14058 800
rect 14108 762 14136 870
rect 14292 762 14320 2858
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14384 800 14412 2586
rect 14476 1562 14504 5646
rect 14568 1698 14596 6054
rect 14660 5370 14688 7686
rect 14752 6882 14780 7806
rect 14844 7188 14872 11698
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14936 11218 14964 11290
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14936 10810 14964 11154
rect 15028 11150 15056 14826
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15120 12986 15148 14282
rect 15200 13456 15252 13462
rect 15200 13398 15252 13404
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15212 12170 15240 13398
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14936 8498 14964 9318
rect 15108 9104 15160 9110
rect 15108 9046 15160 9052
rect 14924 8492 14976 8498
rect 14924 8434 14976 8440
rect 15120 7886 15148 9046
rect 15212 8786 15240 11562
rect 15304 8974 15332 16458
rect 15384 16040 15436 16046
rect 15384 15982 15436 15988
rect 15396 15910 15424 15982
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 12102 15424 15846
rect 15384 12096 15436 12102
rect 15384 12038 15436 12044
rect 15396 11626 15424 12038
rect 15384 11620 15436 11626
rect 15384 11562 15436 11568
rect 15488 11558 15516 19246
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15672 18630 15700 19110
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15660 18624 15712 18630
rect 15660 18566 15712 18572
rect 15660 18420 15712 18426
rect 15660 18362 15712 18368
rect 15672 18057 15700 18362
rect 15658 18048 15714 18057
rect 15658 17983 15714 17992
rect 15764 17814 15792 18634
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15580 17338 15608 17682
rect 15752 17536 15804 17542
rect 15752 17478 15804 17484
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15764 16794 15792 17478
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15580 14346 15608 16730
rect 15856 14929 15884 19178
rect 15948 15026 15976 19654
rect 16408 19242 16436 20266
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 17684 20256 17736 20262
rect 17684 20198 17736 20204
rect 16500 19718 16528 20198
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 16488 19712 16540 19718
rect 16488 19654 16540 19660
rect 16948 19712 17000 19718
rect 16948 19654 17000 19660
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16960 18970 16988 19654
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17040 19168 17092 19174
rect 17038 19136 17040 19145
rect 17092 19136 17094 19145
rect 17038 19071 17094 19080
rect 16304 18964 16356 18970
rect 16304 18906 16356 18912
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16120 18828 16172 18834
rect 16120 18770 16172 18776
rect 16028 18624 16080 18630
rect 16028 18566 16080 18572
rect 16040 16522 16068 18566
rect 16132 17134 16160 18770
rect 16316 18766 16344 18906
rect 17236 18834 17264 19178
rect 17224 18828 17276 18834
rect 17224 18770 17276 18776
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16948 18760 17000 18766
rect 16948 18702 17000 18708
rect 16212 18692 16264 18698
rect 16212 18634 16264 18640
rect 16224 18193 16252 18634
rect 16960 18630 16988 18702
rect 17224 18692 17276 18698
rect 17224 18634 17276 18640
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16868 18290 16896 18362
rect 16856 18284 16908 18290
rect 16856 18226 16908 18232
rect 16210 18184 16266 18193
rect 16210 18119 16266 18128
rect 16224 18086 16252 18119
rect 16960 18086 16988 18566
rect 17236 18358 17264 18634
rect 17224 18352 17276 18358
rect 17224 18294 17276 18300
rect 17040 18216 17092 18222
rect 17040 18158 17092 18164
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16948 18080 17000 18086
rect 16948 18022 17000 18028
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16408 16658 16436 17614
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16960 17202 16988 18022
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16396 16652 16448 16658
rect 16396 16594 16448 16600
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16408 16250 16436 16390
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16396 16244 16448 16250
rect 16396 16186 16448 16192
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16120 15360 16172 15366
rect 16592 15348 16620 15438
rect 16120 15302 16172 15308
rect 16408 15320 16620 15348
rect 16764 15360 16816 15366
rect 15936 15020 15988 15026
rect 15936 14962 15988 14968
rect 15842 14920 15898 14929
rect 15948 14906 15976 14962
rect 15948 14878 16068 14906
rect 15842 14855 15898 14864
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15752 14068 15804 14074
rect 15752 14010 15804 14016
rect 15660 13388 15712 13394
rect 15660 13330 15712 13336
rect 15672 12850 15700 13330
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15660 12640 15712 12646
rect 15660 12582 15712 12588
rect 15672 12238 15700 12582
rect 15764 12434 15792 14010
rect 15856 12918 15884 14855
rect 16040 14822 16068 14878
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 15936 14340 15988 14346
rect 15936 14282 15988 14288
rect 15948 14074 15976 14282
rect 15936 14068 15988 14074
rect 15936 14010 15988 14016
rect 16040 13818 16068 14758
rect 16132 14346 16160 15302
rect 16408 14890 16436 15320
rect 16960 15348 16988 16594
rect 17052 16182 17080 18158
rect 17132 18080 17184 18086
rect 17132 18022 17184 18028
rect 17040 16176 17092 16182
rect 17040 16118 17092 16124
rect 16816 15320 17080 15348
rect 16764 15302 16816 15308
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16946 15192 17002 15201
rect 16946 15127 16948 15136
rect 17000 15127 17002 15136
rect 16948 15098 17000 15104
rect 16396 14884 16448 14890
rect 16396 14826 16448 14832
rect 16396 14612 16448 14618
rect 16396 14554 16448 14560
rect 16302 14512 16358 14521
rect 16302 14447 16358 14456
rect 16210 14376 16266 14385
rect 16120 14340 16172 14346
rect 16210 14311 16266 14320
rect 16120 14282 16172 14288
rect 15948 13790 16068 13818
rect 15844 12912 15896 12918
rect 15844 12854 15896 12860
rect 15948 12434 15976 13790
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 16040 13326 16068 13670
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 16224 12986 16252 14311
rect 16212 12980 16264 12986
rect 16212 12922 16264 12928
rect 15764 12406 15884 12434
rect 15948 12406 16068 12434
rect 15660 12232 15712 12238
rect 15660 12174 15712 12180
rect 15672 11898 15700 12174
rect 15660 11892 15712 11898
rect 15660 11834 15712 11840
rect 15476 11552 15528 11558
rect 15476 11494 15528 11500
rect 15384 11280 15436 11286
rect 15384 11222 15436 11228
rect 15292 8968 15344 8974
rect 15396 8945 15424 11222
rect 15488 8974 15516 11494
rect 15658 10296 15714 10305
rect 15658 10231 15714 10240
rect 15672 10198 15700 10231
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15476 8968 15528 8974
rect 15292 8910 15344 8916
rect 15382 8936 15438 8945
rect 15476 8910 15528 8916
rect 15382 8871 15438 8880
rect 15384 8832 15436 8838
rect 15212 8758 15332 8786
rect 15384 8774 15436 8780
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15212 8498 15240 8570
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15304 8276 15332 8758
rect 15396 8498 15424 8774
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 15488 8362 15516 8570
rect 15660 8560 15712 8566
rect 15660 8502 15712 8508
rect 15476 8356 15528 8362
rect 15476 8298 15528 8304
rect 15212 8248 15332 8276
rect 15568 8288 15620 8294
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15016 7200 15068 7206
rect 14844 7160 15016 7188
rect 15016 7142 15068 7148
rect 14752 6854 14872 6882
rect 14844 6798 14872 6854
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14648 5364 14700 5370
rect 14648 5306 14700 5312
rect 14660 5234 14688 5306
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14660 3058 14688 4519
rect 14752 3534 14780 4762
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14844 3097 14872 6394
rect 14922 5128 14978 5137
rect 14922 5063 14978 5072
rect 14936 5030 14964 5063
rect 14924 5024 14976 5030
rect 14924 4966 14976 4972
rect 14922 4856 14978 4865
rect 14922 4791 14924 4800
rect 14976 4791 14978 4800
rect 14924 4762 14976 4768
rect 15028 3602 15056 7142
rect 15120 4826 15148 7822
rect 15212 7410 15240 8248
rect 15568 8230 15620 8236
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15304 6798 15332 7754
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15292 6792 15344 6798
rect 15292 6734 15344 6740
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15212 4214 15240 6666
rect 15382 6488 15438 6497
rect 15292 6452 15344 6458
rect 15488 6458 15516 7686
rect 15580 7342 15608 8230
rect 15672 7818 15700 8502
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15568 7336 15620 7342
rect 15568 7278 15620 7284
rect 15382 6423 15438 6432
rect 15476 6452 15528 6458
rect 15292 6394 15344 6400
rect 15304 6322 15332 6394
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15304 5914 15332 6258
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15290 5536 15346 5545
rect 15290 5471 15346 5480
rect 15200 4208 15252 4214
rect 15200 4150 15252 4156
rect 15304 4146 15332 5471
rect 15396 5234 15424 6423
rect 15476 6394 15528 6400
rect 15474 6352 15530 6361
rect 15474 6287 15530 6296
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15396 4214 15424 4626
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15292 4140 15344 4146
rect 15292 4082 15344 4088
rect 15382 4040 15438 4049
rect 15382 3975 15438 3984
rect 15016 3596 15068 3602
rect 15016 3538 15068 3544
rect 15396 3534 15424 3975
rect 15488 3534 15516 6287
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 15672 5914 15700 6190
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15580 4554 15608 5646
rect 15764 5234 15792 8774
rect 15856 8362 15884 12406
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15948 9586 15976 9998
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9178 15976 9522
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 15948 8634 15976 9114
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 15948 8090 15976 8570
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15948 7546 15976 8026
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15752 5228 15804 5234
rect 15752 5170 15804 5176
rect 15752 5024 15804 5030
rect 15752 4966 15804 4972
rect 15568 4548 15620 4554
rect 15568 4490 15620 4496
rect 15580 4146 15608 4490
rect 15764 4282 15792 4966
rect 15752 4276 15804 4282
rect 15752 4218 15804 4224
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15856 3992 15884 6190
rect 15948 5386 15976 7142
rect 16040 6662 16068 12406
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16132 8362 16160 9114
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16224 8242 16252 8774
rect 16132 8214 16252 8242
rect 16028 6656 16080 6662
rect 16028 6598 16080 6604
rect 16040 5817 16068 6598
rect 16026 5808 16082 5817
rect 16026 5743 16082 5752
rect 16132 5545 16160 8214
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16224 7410 16252 7686
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16224 6361 16252 7346
rect 16316 6458 16344 14447
rect 16408 13258 16436 14554
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 17052 13530 17080 15320
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16210 6352 16266 6361
rect 16210 6287 16266 6296
rect 16408 6186 16436 12786
rect 16960 12374 16988 13466
rect 17144 12753 17172 18022
rect 17328 16250 17356 19858
rect 17500 19712 17552 19718
rect 17500 19654 17552 19660
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17512 19417 17540 19654
rect 17604 19514 17632 19654
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17696 19446 17724 20198
rect 17788 19922 17816 20402
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 19536 20058 19564 20402
rect 20444 20256 20496 20262
rect 20444 20198 20496 20204
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 17776 19916 17828 19922
rect 17776 19858 17828 19864
rect 18880 19916 18932 19922
rect 18880 19858 18932 19864
rect 17958 19816 18014 19825
rect 17868 19780 17920 19786
rect 17958 19751 18014 19760
rect 17868 19722 17920 19728
rect 17880 19446 17908 19722
rect 17684 19440 17736 19446
rect 17498 19408 17554 19417
rect 17684 19382 17736 19388
rect 17868 19440 17920 19446
rect 17868 19382 17920 19388
rect 17498 19343 17554 19352
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17776 19236 17828 19242
rect 17776 19178 17828 19184
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17408 18352 17460 18358
rect 17408 18294 17460 18300
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17224 15700 17276 15706
rect 17224 15642 17276 15648
rect 17236 15026 17264 15642
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17130 12744 17186 12753
rect 17130 12679 17186 12688
rect 17236 12594 17264 14962
rect 17052 12566 17264 12594
rect 17052 12434 17080 12566
rect 17328 12434 17356 16050
rect 17420 14278 17448 18294
rect 17592 18216 17644 18222
rect 17592 18158 17644 18164
rect 17604 17542 17632 18158
rect 17592 17536 17644 17542
rect 17592 17478 17644 17484
rect 17500 16992 17552 16998
rect 17500 16934 17552 16940
rect 17512 16726 17540 16934
rect 17696 16726 17724 18362
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17684 16720 17736 16726
rect 17684 16662 17736 16668
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17052 12406 17172 12434
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16868 12186 16896 12242
rect 17038 12200 17094 12209
rect 16868 12170 16988 12186
rect 16856 12164 16988 12170
rect 16908 12158 16988 12164
rect 16856 12106 16908 12112
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16488 11620 16540 11626
rect 16488 11562 16540 11568
rect 16500 11268 16528 11562
rect 16580 11280 16632 11286
rect 16500 11240 16580 11268
rect 16580 11222 16632 11228
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16500 8838 16528 8910
rect 16488 8832 16540 8838
rect 16488 8774 16540 8780
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16960 8090 16988 12158
rect 17038 12135 17094 12144
rect 17052 12102 17080 12135
rect 17040 12096 17092 12102
rect 17040 12038 17092 12044
rect 17052 9382 17080 12038
rect 17144 10538 17172 12406
rect 17236 12406 17356 12434
rect 17132 10532 17184 10538
rect 17132 10474 17184 10480
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7579 16852 7588
rect 16960 7478 16988 7822
rect 16948 7472 17000 7478
rect 16948 7414 17000 7420
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16396 6180 16448 6186
rect 16396 6122 16448 6128
rect 16212 5840 16264 5846
rect 16212 5782 16264 5788
rect 16118 5536 16174 5545
rect 16118 5471 16174 5480
rect 15948 5358 16160 5386
rect 16028 5024 16080 5030
rect 15934 4992 15990 5001
rect 16028 4966 16080 4972
rect 15934 4927 15990 4936
rect 15948 4554 15976 4927
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15936 4004 15988 4010
rect 15856 3964 15936 3992
rect 15936 3946 15988 3952
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 14830 3088 14886 3097
rect 14648 3052 14700 3058
rect 14830 3023 14886 3032
rect 14648 2994 14700 3000
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14660 2106 14688 2382
rect 14648 2100 14700 2106
rect 14648 2042 14700 2048
rect 14556 1692 14608 1698
rect 14556 1634 14608 1640
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 14752 800 14780 2858
rect 14844 2774 14872 3023
rect 15108 2916 15160 2922
rect 15108 2858 15160 2864
rect 14844 2746 15056 2774
rect 15028 2514 15056 2746
rect 15016 2508 15068 2514
rect 15016 2450 15068 2456
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 14832 2304 14884 2310
rect 14832 2246 14884 2252
rect 14844 1970 14872 2246
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 14936 1902 14964 2382
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 15120 800 15148 2858
rect 16040 2650 16068 4966
rect 16132 3913 16160 5358
rect 16118 3904 16174 3913
rect 16118 3839 16174 3848
rect 16224 3641 16252 5782
rect 16868 5574 16896 6394
rect 16960 5760 16988 6598
rect 17052 5794 17080 8774
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 17144 6322 17172 7414
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17052 5766 17172 5794
rect 16951 5732 16988 5760
rect 16951 5624 16979 5732
rect 17144 5642 17172 5766
rect 17132 5636 17184 5642
rect 16951 5596 16988 5624
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16764 5364 16816 5370
rect 16764 5306 16816 5312
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16776 4978 16804 5306
rect 16960 5234 16988 5596
rect 17132 5578 17184 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16948 5228 17000 5234
rect 16948 5170 17000 5176
rect 16408 4622 16436 4966
rect 16776 4950 16988 4978
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16210 3632 16266 3641
rect 16210 3567 16266 3576
rect 16028 2644 16080 2650
rect 16028 2586 16080 2592
rect 15476 2576 15528 2582
rect 15476 2518 15528 2524
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15212 1766 15240 2382
rect 15200 1760 15252 1766
rect 15200 1702 15252 1708
rect 15488 800 15516 2518
rect 16316 2514 16344 3878
rect 16684 3738 16712 4082
rect 16960 4049 16988 4950
rect 16946 4040 17002 4049
rect 16946 3975 17002 3984
rect 16672 3732 16724 3738
rect 16672 3674 16724 3680
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16304 2508 16356 2514
rect 16304 2450 16356 2456
rect 16212 2372 16264 2378
rect 16212 2314 16264 2320
rect 15844 2304 15896 2310
rect 15844 2246 15896 2252
rect 15856 800 15884 2246
rect 16224 800 16252 2314
rect 16408 1630 16436 3538
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16948 3188 17000 3194
rect 17052 3176 17080 5510
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17144 3602 17172 5306
rect 17236 3738 17264 12406
rect 17316 12096 17368 12102
rect 17316 12038 17368 12044
rect 17328 11694 17356 12038
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 11558 17356 11630
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11150 17356 11494
rect 17420 11150 17448 14214
rect 17512 13530 17540 16662
rect 17696 16590 17724 16662
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17592 16244 17644 16250
rect 17592 16186 17644 16192
rect 17604 13954 17632 16186
rect 17684 15972 17736 15978
rect 17684 15914 17736 15920
rect 17696 15706 17724 15914
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17684 15496 17736 15502
rect 17684 15438 17736 15444
rect 17696 15094 17724 15438
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17604 13926 17724 13954
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17512 12968 17540 13466
rect 17604 13326 17632 13806
rect 17592 13320 17644 13326
rect 17592 13262 17644 13268
rect 17512 12940 17632 12968
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17328 10810 17356 11086
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17420 9722 17448 9862
rect 17408 9716 17460 9722
rect 17408 9658 17460 9664
rect 17512 9466 17540 12786
rect 17604 10470 17632 12940
rect 17696 10810 17724 13926
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17788 10742 17816 19178
rect 17880 19174 17908 19246
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17972 18970 18000 19751
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 19514 18276 19654
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18236 19304 18288 19310
rect 18236 19246 18288 19252
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17868 18420 17920 18426
rect 17868 18362 17920 18368
rect 17880 17882 17908 18362
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17868 17740 17920 17746
rect 17868 17682 17920 17688
rect 17880 17542 17908 17682
rect 17972 17678 18000 18566
rect 18156 18290 18184 18906
rect 18144 18284 18196 18290
rect 18144 18226 18196 18232
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 18086 18092 18158
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 17868 17536 17920 17542
rect 17868 17478 17920 17484
rect 17868 17332 17920 17338
rect 17868 17274 17920 17280
rect 17880 14006 17908 17274
rect 18064 16114 18092 17614
rect 18248 17610 18276 19246
rect 18708 18970 18736 19314
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18892 18902 18920 19858
rect 19708 19508 19760 19514
rect 19708 19450 19760 19456
rect 19720 19334 19748 19450
rect 20076 19372 20128 19378
rect 19720 19306 19840 19334
rect 20076 19314 20128 19320
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18696 18828 18748 18834
rect 18696 18770 18748 18776
rect 18604 18352 18656 18358
rect 18604 18294 18656 18300
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18248 17270 18276 17546
rect 18236 17264 18288 17270
rect 18236 17206 18288 17212
rect 18524 16250 18552 18022
rect 18616 17542 18644 18294
rect 18604 17536 18656 17542
rect 18602 17504 18604 17513
rect 18656 17504 18658 17513
rect 18602 17439 18658 17448
rect 18604 16992 18656 16998
rect 18604 16934 18656 16940
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 17868 14000 17920 14006
rect 17868 13942 17920 13948
rect 18064 12730 18092 16050
rect 18616 13841 18644 16934
rect 18708 16697 18736 18770
rect 19432 18692 19484 18698
rect 19484 18652 19564 18680
rect 19432 18634 19484 18640
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18972 18148 19024 18154
rect 18972 18090 19024 18096
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18694 16688 18750 16697
rect 18694 16623 18750 16632
rect 18800 16590 18828 18022
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18892 16454 18920 17138
rect 18696 16448 18748 16454
rect 18696 16390 18748 16396
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18708 15026 18736 16390
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18696 14816 18748 14822
rect 18696 14758 18748 14764
rect 18602 13832 18658 13841
rect 18602 13767 18658 13776
rect 18512 13728 18564 13734
rect 18512 13670 18564 13676
rect 18418 13288 18474 13297
rect 18524 13274 18552 13670
rect 18474 13246 18552 13274
rect 18418 13223 18420 13232
rect 18472 13223 18474 13232
rect 18420 13194 18472 13200
rect 18328 13184 18380 13190
rect 18380 13132 18460 13138
rect 18328 13126 18460 13132
rect 18340 13110 18460 13126
rect 18064 12702 18184 12730
rect 18156 12646 18184 12702
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18064 12186 18092 12582
rect 18156 12434 18184 12582
rect 18432 12434 18460 13110
rect 18156 12406 18276 12434
rect 18064 12158 18184 12186
rect 18156 12102 18184 12158
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18248 11762 18276 12406
rect 18340 12406 18460 12434
rect 18604 12436 18656 12442
rect 18052 11756 18104 11762
rect 18052 11698 18104 11704
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18064 11150 18092 11698
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17592 10464 17644 10470
rect 17592 10406 17644 10412
rect 17696 10266 17724 10610
rect 17684 10260 17736 10266
rect 17684 10202 17736 10208
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17328 9438 17540 9466
rect 17328 5370 17356 9438
rect 17500 9376 17552 9382
rect 17500 9318 17552 9324
rect 17408 8968 17460 8974
rect 17408 8910 17460 8916
rect 17420 8430 17448 8910
rect 17512 8838 17540 9318
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17408 8424 17460 8430
rect 17408 8366 17460 8372
rect 17420 8294 17448 8366
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17420 7886 17448 8230
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17420 5710 17448 7822
rect 17512 7410 17540 8434
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17500 6112 17552 6118
rect 17500 6054 17552 6060
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17316 5364 17368 5370
rect 17316 5306 17368 5312
rect 17408 5024 17460 5030
rect 17408 4966 17460 4972
rect 17316 4480 17368 4486
rect 17316 4422 17368 4428
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17132 3596 17184 3602
rect 17132 3538 17184 3544
rect 17000 3148 17080 3176
rect 16948 3130 17000 3136
rect 17328 2990 17356 4422
rect 17316 2984 17368 2990
rect 17316 2926 17368 2932
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 17040 2100 17092 2106
rect 17040 2042 17092 2048
rect 16580 1760 16632 1766
rect 16580 1702 16632 1708
rect 16396 1624 16448 1630
rect 16396 1566 16448 1572
rect 16592 800 16620 1702
rect 17052 898 17080 2042
rect 17236 1834 17264 2382
rect 17316 2032 17368 2038
rect 17316 1974 17368 1980
rect 17224 1828 17276 1834
rect 17224 1770 17276 1776
rect 16960 870 17080 898
rect 16960 800 16988 870
rect 17328 800 17356 1974
rect 17420 1970 17448 4966
rect 17512 4146 17540 6054
rect 17604 5234 17632 9862
rect 17788 9738 17816 10678
rect 17696 9710 17816 9738
rect 17696 5914 17724 9710
rect 17880 9586 17908 10746
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17776 9580 17828 9586
rect 17776 9522 17828 9528
rect 17868 9580 17920 9586
rect 17868 9522 17920 9528
rect 17788 9178 17816 9522
rect 17972 9518 18000 10066
rect 17960 9512 18012 9518
rect 17960 9454 18012 9460
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17880 9058 17908 9318
rect 17788 9042 17908 9058
rect 17776 9036 17908 9042
rect 17828 9030 17908 9036
rect 17776 8978 17828 8984
rect 17868 8900 17920 8906
rect 17868 8842 17920 8848
rect 17880 8498 17908 8842
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8634 18092 8774
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 18052 8492 18104 8498
rect 18104 8452 18184 8480
rect 18052 8434 18104 8440
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17788 5710 17816 8298
rect 17880 7857 17908 8434
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 8016 18012 8022
rect 17960 7958 18012 7964
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 17972 6730 18000 7958
rect 18064 7886 18092 8026
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18156 7546 18184 8452
rect 18144 7540 18196 7546
rect 18144 7482 18196 7488
rect 18142 7440 18198 7449
rect 18142 7375 18198 7384
rect 18050 6896 18106 6905
rect 18050 6831 18052 6840
rect 18104 6831 18106 6840
rect 18052 6802 18104 6808
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 18156 6458 18184 7375
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 6180 18012 6186
rect 17960 6122 18012 6128
rect 17776 5704 17828 5710
rect 17776 5646 17828 5652
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17696 5522 17724 5578
rect 17696 5494 17816 5522
rect 17592 5228 17644 5234
rect 17592 5170 17644 5176
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17512 3058 17540 4082
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17408 1964 17460 1970
rect 17408 1906 17460 1912
rect 17604 1902 17632 4966
rect 17696 4185 17724 5170
rect 17682 4176 17738 4185
rect 17682 4111 17738 4120
rect 17788 4078 17816 5494
rect 17972 5137 18000 6122
rect 17958 5128 18014 5137
rect 17958 5063 18014 5072
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17972 4185 18000 4966
rect 18064 4282 18092 6326
rect 18248 4570 18276 8570
rect 18340 7426 18368 12406
rect 18604 12378 18656 12384
rect 18616 12073 18644 12378
rect 18602 12064 18658 12073
rect 18602 11999 18658 12008
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18432 9489 18460 9998
rect 18418 9480 18474 9489
rect 18418 9415 18474 9424
rect 18418 8936 18474 8945
rect 18418 8871 18474 8880
rect 18432 7954 18460 8871
rect 18616 8004 18644 11222
rect 18708 8072 18736 14758
rect 18892 12850 18920 15982
rect 18984 14074 19012 18090
rect 19076 17882 19104 18158
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19536 17354 19564 18652
rect 19616 18624 19668 18630
rect 19616 18566 19668 18572
rect 19628 18193 19656 18566
rect 19614 18184 19670 18193
rect 19614 18119 19670 18128
rect 19708 17536 19760 17542
rect 19708 17478 19760 17484
rect 19536 17326 19656 17354
rect 19628 17270 19656 17326
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19536 16794 19564 17138
rect 19720 16810 19748 17478
rect 19524 16788 19576 16794
rect 19524 16730 19576 16736
rect 19628 16782 19748 16810
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19524 15496 19576 15502
rect 19524 15438 19576 15444
rect 19536 15366 19564 15438
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 18972 14068 19024 14074
rect 18972 14010 19024 14016
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18984 12434 19012 14010
rect 19444 13818 19472 14282
rect 19536 13977 19564 15302
rect 19522 13968 19578 13977
rect 19522 13903 19578 13912
rect 19444 13790 19564 13818
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19340 13184 19392 13190
rect 19340 13126 19392 13132
rect 19352 12918 19380 13126
rect 19340 12912 19392 12918
rect 19340 12854 19392 12860
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 18892 12406 19012 12434
rect 18786 11112 18842 11121
rect 18786 11047 18842 11056
rect 18800 10062 18828 11047
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18892 8566 18920 12406
rect 19536 12374 19564 13790
rect 19524 12368 19576 12374
rect 19524 12310 19576 12316
rect 19536 11558 19564 12310
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 18972 11348 19024 11354
rect 18972 11290 19024 11296
rect 18984 9602 19012 11290
rect 19536 11286 19564 11494
rect 19524 11280 19576 11286
rect 19524 11222 19576 11228
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19536 10130 19564 10406
rect 19628 10266 19656 16782
rect 19812 16776 19840 19306
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 19904 16969 19932 17682
rect 19996 17338 20024 18702
rect 20088 17882 20116 19314
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18834 20300 19110
rect 20260 18828 20312 18834
rect 20260 18770 20312 18776
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 18290 20300 18566
rect 20456 18290 20484 20198
rect 20548 19990 20576 20402
rect 20640 19990 20668 20839
rect 21742 20700 22050 20709
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 21180 20528 21232 20534
rect 21180 20470 21232 20476
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 20097 20760 20198
rect 20718 20088 20774 20097
rect 21100 20058 21128 20402
rect 20718 20023 20774 20032
rect 21088 20052 21140 20058
rect 21088 19994 21140 20000
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20628 19984 20680 19990
rect 20628 19926 20680 19932
rect 20536 19848 20588 19854
rect 20536 19790 20588 19796
rect 20548 19514 20576 19790
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20640 19281 20668 19450
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20626 19272 20682 19281
rect 20626 19207 20682 19216
rect 20812 18896 20864 18902
rect 20812 18838 20864 18844
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20444 18284 20496 18290
rect 20444 18226 20496 18232
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20260 17672 20312 17678
rect 20260 17614 20312 17620
rect 20640 17626 20668 18566
rect 20720 18080 20772 18086
rect 20718 18048 20720 18057
rect 20772 18048 20774 18057
rect 20718 17983 20774 17992
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19984 17332 20036 17338
rect 19984 17274 20036 17280
rect 19890 16960 19946 16969
rect 19890 16895 19946 16904
rect 19812 16748 20024 16776
rect 19798 16688 19854 16697
rect 19798 16623 19854 16632
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 19720 15162 19748 15642
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19812 14958 19840 16623
rect 19890 16552 19946 16561
rect 19890 16487 19946 16496
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19904 14906 19932 16487
rect 19996 16114 20024 16748
rect 20088 16538 20116 17546
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20180 16833 20208 16934
rect 20166 16824 20222 16833
rect 20166 16759 20222 16768
rect 20088 16510 20208 16538
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19708 14612 19760 14618
rect 19812 14600 19840 14894
rect 19904 14878 20024 14906
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19760 14572 19840 14600
rect 19708 14554 19760 14560
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12442 19748 13126
rect 19904 12850 19932 14758
rect 19996 14006 20024 14878
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13530 20024 13806
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19892 12844 19944 12850
rect 19892 12786 19944 12792
rect 19812 12753 19840 12786
rect 19798 12744 19854 12753
rect 20088 12714 20116 16390
rect 20180 13734 20208 16510
rect 20168 13728 20220 13734
rect 20168 13670 20220 13676
rect 20272 13512 20300 17614
rect 20640 17598 20760 17626
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20628 17536 20680 17542
rect 20628 17478 20680 17484
rect 20352 16992 20404 16998
rect 20352 16934 20404 16940
rect 20364 16590 20392 16934
rect 20456 16658 20484 17478
rect 20640 16697 20668 17478
rect 20626 16688 20682 16697
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20536 16652 20588 16658
rect 20626 16623 20682 16632
rect 20536 16594 20588 16600
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 15978 20392 16390
rect 20548 16266 20576 16594
rect 20732 16574 20760 17598
rect 20824 17338 20852 18838
rect 20916 17814 20944 19314
rect 21088 18624 21140 18630
rect 21088 18566 21140 18572
rect 20996 18148 21048 18154
rect 20996 18090 21048 18096
rect 20904 17808 20956 17814
rect 20904 17750 20956 17756
rect 20904 17672 20956 17678
rect 20904 17614 20956 17620
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20916 17218 20944 17614
rect 20456 16238 20576 16266
rect 20640 16546 20760 16574
rect 20824 17190 20944 17218
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20352 15428 20404 15434
rect 20352 15370 20404 15376
rect 20364 14074 20392 15370
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20352 13728 20404 13734
rect 20352 13670 20404 13676
rect 20180 13484 20300 13512
rect 20180 13308 20208 13484
rect 20180 13280 20300 13308
rect 19798 12679 19854 12688
rect 20076 12708 20128 12714
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19812 11898 19840 12679
rect 20076 12650 20128 12656
rect 19984 12164 20036 12170
rect 19984 12106 20036 12112
rect 19996 11898 20024 12106
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 19800 11620 19852 11626
rect 19800 11562 19852 11568
rect 19812 10742 19840 11562
rect 19800 10736 19852 10742
rect 20180 10713 20208 11698
rect 19800 10678 19852 10684
rect 20166 10704 20222 10713
rect 20166 10639 20222 10648
rect 20166 10296 20222 10305
rect 19616 10260 19668 10266
rect 20166 10231 20222 10240
rect 19616 10202 19668 10208
rect 19524 10124 19576 10130
rect 19524 10066 19576 10072
rect 18984 9586 19288 9602
rect 18984 9580 19300 9586
rect 18984 9574 19248 9580
rect 19248 9522 19300 9528
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18880 8560 18932 8566
rect 18880 8502 18932 8508
rect 18788 8084 18840 8090
rect 18708 8044 18788 8072
rect 18788 8026 18840 8032
rect 18616 7976 18736 8004
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18708 7886 18736 7976
rect 18786 7984 18842 7993
rect 18786 7919 18842 7928
rect 18512 7880 18564 7886
rect 18512 7822 18564 7828
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18340 7398 18460 7426
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 18340 6798 18368 7278
rect 18328 6792 18380 6798
rect 18432 6769 18460 7398
rect 18328 6734 18380 6740
rect 18418 6760 18474 6769
rect 18418 6695 18474 6704
rect 18420 6656 18472 6662
rect 18420 6598 18472 6604
rect 18432 6458 18460 6598
rect 18420 6452 18472 6458
rect 18420 6394 18472 6400
rect 18524 6118 18552 7822
rect 18800 7818 18828 7919
rect 18788 7812 18840 7818
rect 18788 7754 18840 7760
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18708 7410 18736 7686
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18696 7404 18748 7410
rect 18696 7346 18748 7352
rect 18604 6724 18656 6730
rect 18604 6666 18656 6672
rect 18420 6112 18472 6118
rect 18420 6054 18472 6060
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18432 5817 18460 6054
rect 18418 5808 18474 5817
rect 18418 5743 18474 5752
rect 18512 5568 18564 5574
rect 18616 5545 18644 6666
rect 18512 5510 18564 5516
rect 18602 5536 18658 5545
rect 18420 5296 18472 5302
rect 18340 5244 18420 5250
rect 18340 5238 18472 5244
rect 18340 5222 18460 5238
rect 18340 5137 18368 5222
rect 18326 5128 18382 5137
rect 18326 5063 18382 5072
rect 18156 4554 18276 4570
rect 18144 4548 18276 4554
rect 18196 4542 18276 4548
rect 18144 4490 18196 4496
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 17958 4176 18014 4185
rect 17958 4111 18014 4120
rect 17776 4072 17828 4078
rect 17776 4014 17828 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17776 3392 17828 3398
rect 17776 3334 17828 3340
rect 17788 3194 17816 3334
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17880 2938 17908 3946
rect 18064 3126 18092 4218
rect 18144 4140 18196 4146
rect 18144 4082 18196 4088
rect 18156 3738 18184 4082
rect 18144 3732 18196 3738
rect 18144 3674 18196 3680
rect 18052 3120 18104 3126
rect 18144 3120 18196 3126
rect 18052 3062 18104 3068
rect 18142 3088 18144 3097
rect 18196 3088 18198 3097
rect 18142 3023 18198 3032
rect 18248 2990 18276 4542
rect 18340 3466 18368 5063
rect 18524 4622 18552 5510
rect 18602 5471 18658 5480
rect 18604 5160 18656 5166
rect 18602 5128 18604 5137
rect 18656 5128 18658 5137
rect 18602 5063 18658 5072
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 18236 2984 18288 2990
rect 17880 2910 18184 2938
rect 18236 2926 18288 2932
rect 17960 2848 18012 2854
rect 17880 2796 17960 2802
rect 17880 2790 18012 2796
rect 17880 2774 18000 2790
rect 17880 2553 17908 2774
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17866 2544 17922 2553
rect 17866 2479 17922 2488
rect 17972 2428 18000 2586
rect 18156 2514 18184 2910
rect 18234 2544 18290 2553
rect 18144 2508 18196 2514
rect 18234 2479 18290 2488
rect 18144 2450 18196 2456
rect 17696 2400 18000 2428
rect 17592 1896 17644 1902
rect 17592 1838 17644 1844
rect 17696 800 17724 2400
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 17958 1728 18014 1737
rect 17958 1663 18014 1672
rect 17972 1562 18000 1663
rect 17960 1556 18012 1562
rect 17960 1498 18012 1504
rect 18064 800 18092 2314
rect 18248 1698 18276 2479
rect 18236 1692 18288 1698
rect 18236 1634 18288 1640
rect 18432 800 18460 4422
rect 18604 3936 18656 3942
rect 18604 3878 18656 3884
rect 18616 3602 18644 3878
rect 18604 3596 18656 3602
rect 18604 3538 18656 3544
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18524 1766 18552 2246
rect 18708 2009 18736 7346
rect 18892 7342 18920 7482
rect 18880 7336 18932 7342
rect 18880 7278 18932 7284
rect 18786 7168 18842 7177
rect 18786 7103 18842 7112
rect 18800 6798 18828 7103
rect 18788 6792 18840 6798
rect 18788 6734 18840 6740
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 5681 18828 6598
rect 18878 6216 18934 6225
rect 18878 6151 18934 6160
rect 18892 5710 18920 6151
rect 18880 5704 18932 5710
rect 18786 5672 18842 5681
rect 18880 5646 18932 5652
rect 18786 5607 18842 5616
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18694 2000 18750 2009
rect 18694 1935 18750 1944
rect 18512 1760 18564 1766
rect 18512 1702 18564 1708
rect 18800 800 18828 4966
rect 18892 4729 18920 5170
rect 18878 4720 18934 4729
rect 18878 4655 18934 4664
rect 18878 3904 18934 3913
rect 18878 3839 18934 3848
rect 18892 3602 18920 3839
rect 18880 3596 18932 3602
rect 18880 3538 18932 3544
rect 18984 3466 19012 8842
rect 19064 8288 19116 8294
rect 19064 8230 19116 8236
rect 19076 7546 19104 8230
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8123 19451 8132
rect 19248 7948 19300 7954
rect 19248 7890 19300 7896
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19156 7472 19208 7478
rect 19154 7440 19156 7449
rect 19208 7440 19210 7449
rect 19260 7410 19288 7890
rect 19154 7375 19210 7384
rect 19248 7404 19300 7410
rect 19248 7346 19300 7352
rect 19536 7154 19564 10066
rect 20180 9994 20208 10231
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19708 9512 19760 9518
rect 19706 9480 19708 9489
rect 19760 9480 19762 9489
rect 19706 9415 19762 9424
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19628 8294 19656 8978
rect 19616 8288 19668 8294
rect 19616 8230 19668 8236
rect 19628 7818 19656 8230
rect 19812 7954 19840 9862
rect 19996 9178 20024 9862
rect 20180 9586 20208 9930
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19984 8832 20036 8838
rect 19984 8774 20036 8780
rect 20168 8832 20220 8838
rect 20168 8774 20220 8780
rect 19800 7948 19852 7954
rect 19800 7890 19852 7896
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 19616 7812 19668 7818
rect 19616 7754 19668 7760
rect 19798 7576 19854 7585
rect 19798 7511 19854 7520
rect 19812 7478 19840 7511
rect 19800 7472 19852 7478
rect 19800 7414 19852 7420
rect 19536 7126 19656 7154
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19628 6984 19656 7126
rect 19536 6956 19656 6984
rect 19338 6896 19394 6905
rect 19338 6831 19394 6840
rect 19432 6860 19484 6866
rect 19246 6760 19302 6769
rect 19246 6695 19302 6704
rect 19260 6662 19288 6695
rect 19248 6656 19300 6662
rect 19248 6598 19300 6604
rect 19352 6390 19380 6831
rect 19536 6848 19564 6956
rect 19484 6820 19564 6848
rect 19614 6896 19670 6905
rect 19614 6831 19616 6840
rect 19432 6802 19484 6808
rect 19536 6497 19564 6820
rect 19668 6831 19670 6840
rect 19798 6896 19854 6905
rect 19798 6831 19854 6840
rect 19616 6802 19668 6808
rect 19616 6724 19668 6730
rect 19616 6666 19668 6672
rect 19522 6488 19578 6497
rect 19522 6423 19578 6432
rect 19340 6384 19392 6390
rect 19062 6352 19118 6361
rect 19340 6326 19392 6332
rect 19524 6384 19576 6390
rect 19524 6326 19576 6332
rect 19062 6287 19118 6296
rect 19076 3720 19104 6287
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19340 4140 19392 4146
rect 19536 4128 19564 6326
rect 19392 4100 19564 4128
rect 19340 4082 19392 4088
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19628 3738 19656 6666
rect 19708 5840 19760 5846
rect 19812 5828 19840 6831
rect 19760 5800 19840 5828
rect 19708 5782 19760 5788
rect 19720 5370 19748 5782
rect 19708 5364 19760 5370
rect 19708 5306 19760 5312
rect 19720 5166 19748 5306
rect 19708 5160 19760 5166
rect 19708 5102 19760 5108
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19720 4593 19748 4762
rect 19904 4706 19932 7822
rect 19996 6202 20024 8774
rect 20076 7812 20128 7818
rect 20076 7754 20128 7760
rect 20088 7478 20116 7754
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 20074 7304 20130 7313
rect 20074 7239 20130 7248
rect 20088 6338 20116 7239
rect 20180 6866 20208 8774
rect 20168 6860 20220 6866
rect 20168 6802 20220 6808
rect 20272 6662 20300 13280
rect 20364 7002 20392 13670
rect 20456 11626 20484 16238
rect 20536 16108 20588 16114
rect 20536 16050 20588 16056
rect 20548 15706 20576 16050
rect 20536 15700 20588 15706
rect 20536 15642 20588 15648
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20548 14346 20576 15098
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20534 13288 20590 13297
rect 20534 13223 20590 13232
rect 20548 12986 20576 13223
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20548 12345 20576 12718
rect 20640 12442 20668 16546
rect 20718 16416 20774 16425
rect 20718 16351 20774 16360
rect 20732 16250 20760 16351
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20718 16008 20774 16017
rect 20718 15943 20720 15952
rect 20772 15943 20774 15952
rect 20720 15914 20772 15920
rect 20824 15450 20852 17190
rect 20904 17060 20956 17066
rect 20904 17002 20956 17008
rect 20916 16114 20944 17002
rect 21008 16590 21036 18090
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20824 15422 20944 15450
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15088 20772 15094
rect 20824 15065 20852 15302
rect 20720 15030 20772 15036
rect 20810 15056 20866 15065
rect 20732 14414 20760 15030
rect 20810 14991 20866 15000
rect 20720 14408 20772 14414
rect 20720 14350 20772 14356
rect 20732 14006 20760 14350
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20732 13326 20760 13942
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20534 12336 20590 12345
rect 20534 12271 20590 12280
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20548 11801 20576 12106
rect 20534 11792 20590 11801
rect 20534 11727 20590 11736
rect 20444 11620 20496 11626
rect 20444 11562 20496 11568
rect 20732 10674 20760 13262
rect 20916 11898 20944 15422
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 13258 21036 14758
rect 21100 14414 21128 18566
rect 21192 17678 21220 20470
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21284 19825 21312 20198
rect 21270 19816 21326 19825
rect 21270 19751 21326 19760
rect 21364 19712 21416 19718
rect 21364 19654 21416 19660
rect 21272 19168 21324 19174
rect 21272 19110 21324 19116
rect 21284 18329 21312 19110
rect 21376 18873 21404 19654
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21362 18864 21418 18873
rect 21362 18799 21418 18808
rect 21364 18624 21416 18630
rect 21364 18566 21416 18572
rect 21270 18320 21326 18329
rect 21270 18255 21326 18264
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21284 17241 21312 18022
rect 21376 17649 21404 18566
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21362 17640 21418 17649
rect 21362 17575 21418 17584
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 21180 17128 21232 17134
rect 21180 17070 21232 17076
rect 21192 14822 21220 17070
rect 21456 16720 21508 16726
rect 21456 16662 21508 16668
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15609 21312 16390
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21270 15600 21326 15609
rect 21270 15535 21326 15544
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21180 14816 21232 14822
rect 21180 14758 21232 14764
rect 21088 14408 21140 14414
rect 21284 14385 21312 15302
rect 21376 14793 21404 15846
rect 21362 14784 21418 14793
rect 21362 14719 21418 14728
rect 21088 14350 21140 14356
rect 21270 14376 21326 14385
rect 21270 14311 21326 14320
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13977 21312 14214
rect 21270 13968 21326 13977
rect 21270 13903 21326 13912
rect 21270 13560 21326 13569
rect 21270 13495 21272 13504
rect 21324 13495 21326 13504
rect 21272 13466 21324 13472
rect 20996 13252 21048 13258
rect 20996 13194 21048 13200
rect 21468 12850 21496 16662
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 21742 14172 22050 14181
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21742 13084 22050 13093
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 20916 11778 20944 11834
rect 20824 11750 20944 11778
rect 20720 10668 20772 10674
rect 20720 10610 20772 10616
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20548 10033 20576 10066
rect 20628 10056 20680 10062
rect 20534 10024 20590 10033
rect 20628 9998 20680 10004
rect 20534 9959 20590 9968
rect 20442 9616 20498 9625
rect 20442 9551 20498 9560
rect 20456 7818 20484 9551
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 20548 9081 20576 9454
rect 20534 9072 20590 9081
rect 20534 9007 20590 9016
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20442 7576 20498 7585
rect 20442 7511 20498 7520
rect 20352 6996 20404 7002
rect 20352 6938 20404 6944
rect 20260 6656 20312 6662
rect 20260 6598 20312 6604
rect 20258 6488 20314 6497
rect 20258 6423 20314 6432
rect 20088 6310 20208 6338
rect 19996 6174 20116 6202
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19996 5370 20024 6054
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 19812 4678 19932 4706
rect 19706 4584 19762 4593
rect 19706 4519 19762 4528
rect 19616 3732 19668 3738
rect 19076 3692 19196 3720
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 19076 1442 19104 3470
rect 19168 2961 19196 3692
rect 19616 3674 19668 3680
rect 19720 3670 19748 4519
rect 19812 4214 19840 4678
rect 19892 4548 19944 4554
rect 19892 4490 19944 4496
rect 19800 4208 19852 4214
rect 19800 4150 19852 4156
rect 19904 4146 19932 4490
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19708 3664 19760 3670
rect 19708 3606 19760 3612
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19260 3126 19288 3538
rect 19800 3528 19852 3534
rect 19800 3470 19852 3476
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19248 3120 19300 3126
rect 19340 3120 19392 3126
rect 19248 3062 19300 3068
rect 19338 3088 19340 3097
rect 19392 3088 19394 3097
rect 19338 3023 19394 3032
rect 19248 2984 19300 2990
rect 19154 2952 19210 2961
rect 19352 2938 19380 3023
rect 19300 2932 19380 2938
rect 19248 2926 19380 2932
rect 19260 2910 19380 2926
rect 19154 2887 19210 2896
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19432 2304 19484 2310
rect 19432 2246 19484 2252
rect 19444 2106 19472 2246
rect 19432 2100 19484 2106
rect 19432 2042 19484 2048
rect 19076 1414 19196 1442
rect 19168 800 19196 1414
rect 19536 800 19564 3130
rect 19812 2774 19840 3470
rect 19904 2990 19932 4082
rect 19984 3392 20036 3398
rect 19984 3334 20036 3340
rect 19996 3058 20024 3334
rect 20088 3126 20116 6174
rect 20180 5710 20208 6310
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 20272 5216 20300 6423
rect 20456 5642 20484 7511
rect 20536 7404 20588 7410
rect 20536 7346 20588 7352
rect 20548 7041 20576 7346
rect 20534 7032 20590 7041
rect 20534 6967 20590 6976
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20444 5636 20496 5642
rect 20444 5578 20496 5584
rect 20350 5400 20406 5409
rect 20350 5335 20352 5344
rect 20404 5335 20406 5344
rect 20352 5306 20404 5312
rect 20180 5188 20300 5216
rect 20180 4826 20208 5188
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20076 3120 20128 3126
rect 20076 3062 20128 3068
rect 20166 3088 20222 3097
rect 19984 3052 20036 3058
rect 20166 3023 20168 3032
rect 19984 2994 20036 3000
rect 20220 3023 20222 3032
rect 20168 2994 20220 3000
rect 19892 2984 19944 2990
rect 19892 2926 19944 2932
rect 19812 2746 19932 2774
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 19812 1970 19840 2382
rect 19800 1964 19852 1970
rect 19800 1906 19852 1912
rect 19904 800 19932 2746
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19996 2038 20024 2246
rect 19984 2032 20036 2038
rect 19984 1974 20036 1980
rect 20272 800 20300 5034
rect 20456 3233 20484 5578
rect 20548 4078 20576 6258
rect 20640 5370 20668 9998
rect 20732 9450 20760 10610
rect 20720 9444 20772 9450
rect 20720 9386 20772 9392
rect 20824 9042 20852 11750
rect 20904 11620 20956 11626
rect 20904 11562 20956 11568
rect 20916 11082 20944 11562
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20996 11144 21048 11150
rect 20996 11086 21048 11092
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20916 10810 20944 11018
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 21008 10674 21036 11086
rect 20996 10668 21048 10674
rect 20996 10610 21048 10616
rect 20902 10160 20958 10169
rect 21100 10130 21128 11494
rect 21192 10810 21220 12174
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21284 11898 21312 12038
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21270 11520 21326 11529
rect 21270 11455 21326 11464
rect 21284 11354 21312 11455
rect 21272 11348 21324 11354
rect 21272 11290 21324 11296
rect 21180 10804 21232 10810
rect 21180 10746 21232 10752
rect 21364 10668 21416 10674
rect 21364 10610 21416 10616
rect 20902 10095 20958 10104
rect 21088 10124 21140 10130
rect 20812 9036 20864 9042
rect 20812 8978 20864 8984
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 6390 20760 7686
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20732 5710 20760 6190
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20628 5160 20680 5166
rect 20628 5102 20680 5108
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20548 3602 20576 4014
rect 20640 3738 20668 5102
rect 20732 4622 20760 5646
rect 20824 4729 20852 6394
rect 20916 6066 20944 10095
rect 21088 10066 21140 10072
rect 20996 9716 21048 9722
rect 20996 9658 21048 9664
rect 21008 9042 21036 9658
rect 21180 9444 21232 9450
rect 21180 9386 21232 9392
rect 20996 9036 21048 9042
rect 20996 8978 21048 8984
rect 21008 6338 21036 8978
rect 21192 8498 21220 9386
rect 21272 9104 21324 9110
rect 21272 9046 21324 9052
rect 21284 8537 21312 9046
rect 21270 8528 21326 8537
rect 21180 8492 21232 8498
rect 21270 8463 21326 8472
rect 21180 8434 21232 8440
rect 21284 7886 21312 8463
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21088 7812 21140 7818
rect 21088 7754 21140 7760
rect 21100 7721 21128 7754
rect 21086 7712 21142 7721
rect 21086 7647 21142 7656
rect 21376 7546 21404 10610
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21468 7410 21496 11698
rect 21456 7404 21508 7410
rect 21456 7346 21508 7352
rect 21008 6310 21128 6338
rect 21100 6254 21128 6310
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21088 6248 21140 6254
rect 21140 6196 21220 6202
rect 21088 6190 21220 6196
rect 21100 6174 21220 6190
rect 20916 6038 21036 6066
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 20810 4720 20866 4729
rect 20810 4655 20866 4664
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20720 4208 20772 4214
rect 20720 4150 20772 4156
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20732 3505 20760 4150
rect 20824 4146 20852 4655
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20718 3496 20774 3505
rect 20718 3431 20774 3440
rect 20442 3224 20498 3233
rect 20442 3159 20498 3168
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20364 1902 20392 2382
rect 20352 1896 20404 1902
rect 20352 1838 20404 1844
rect 20640 800 20668 2994
rect 20916 2446 20944 5850
rect 21008 5846 21036 6038
rect 20996 5840 21048 5846
rect 20996 5782 21048 5788
rect 21086 5264 21142 5273
rect 21086 5199 21142 5208
rect 21100 4758 21128 5199
rect 21192 5166 21220 6174
rect 21270 5808 21326 5817
rect 21270 5743 21326 5752
rect 21180 5160 21232 5166
rect 21180 5102 21232 5108
rect 21088 4752 21140 4758
rect 21088 4694 21140 4700
rect 21192 4554 21220 5102
rect 21284 4622 21312 5743
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 20904 2440 20956 2446
rect 21376 2417 21404 6258
rect 21468 5370 21496 7346
rect 21560 6458 21588 12106
rect 21742 11996 22050 12005
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21742 10908 22050 10917
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21548 6452 21600 6458
rect 21548 6394 21600 6400
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21456 5364 21508 5370
rect 21456 5306 21508 5312
rect 21468 3534 21496 5306
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21456 3528 21508 3534
rect 21456 3470 21508 3476
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 20904 2382 20956 2388
rect 21362 2408 21418 2417
rect 21362 2343 21418 2352
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21742 2139 22050 2148
rect 14108 734 14320 762
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15106 0 15162 800
rect 15474 0 15530 800
rect 15842 0 15898 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18050 0 18106 800
rect 18418 0 18474 800
rect 18786 0 18842 800
rect 19154 0 19210 800
rect 19522 0 19578 800
rect 19890 0 19946 800
rect 20258 0 20314 800
rect 20626 0 20682 800
<< via2 >>
rect 2962 21256 3018 21312
rect 1950 20848 2006 20904
rect 1306 20304 1362 20360
rect 1122 19760 1178 19816
rect 938 19488 994 19544
rect 938 17720 994 17776
rect 938 2932 940 2952
rect 940 2932 992 2952
rect 992 2932 994 2952
rect 938 2896 994 2932
rect 1490 20032 1546 20088
rect 2042 20440 2098 20496
rect 5262 20440 5318 20496
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 18694 21256 18750 21312
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 4526 20340 4528 20360
rect 4528 20340 4580 20360
rect 4580 20340 4582 20360
rect 2686 19488 2742 19544
rect 1490 18808 1546 18864
rect 1490 18400 1546 18456
rect 2042 19236 2098 19272
rect 2042 19216 2044 19236
rect 2044 19216 2096 19236
rect 2096 19216 2098 19236
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1398 15972 1454 16008
rect 1398 15952 1400 15972
rect 1400 15952 1452 15972
rect 1452 15952 1454 15972
rect 1490 15544 1546 15600
rect 1490 15136 1546 15192
rect 1490 14320 1546 14376
rect 1490 13504 1546 13560
rect 1490 11600 1546 11656
rect 2042 17584 2098 17640
rect 1674 14492 1676 14512
rect 1676 14492 1728 14512
rect 1728 14492 1730 14512
rect 1674 14456 1730 14492
rect 1766 13368 1822 13424
rect 1858 12144 1914 12200
rect 2134 14764 2136 14784
rect 2136 14764 2188 14784
rect 2188 14764 2190 14784
rect 2134 14728 2190 14764
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 4526 20304 4582 20340
rect 4526 19780 4582 19816
rect 4526 19760 4528 19780
rect 4528 19760 4580 19780
rect 4580 19760 4582 19780
rect 3698 19508 3754 19544
rect 3698 19488 3700 19508
rect 3700 19488 3752 19508
rect 3752 19488 3754 19508
rect 3882 19488 3938 19544
rect 4066 19488 4122 19544
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 2134 13912 2190 13968
rect 1950 11756 2006 11792
rect 1950 11736 1952 11756
rect 1952 11736 2004 11756
rect 2004 11736 2006 11756
rect 2226 12280 2282 12336
rect 2226 11872 2282 11928
rect 2226 11464 2282 11520
rect 1950 9560 2006 9616
rect 1490 7520 1546 7576
rect 2226 10512 2282 10568
rect 2226 9832 2282 9888
rect 2226 9580 2282 9616
rect 2226 9560 2228 9580
rect 2228 9560 2280 9580
rect 2280 9560 2282 9580
rect 2226 9424 2282 9480
rect 2134 8608 2190 8664
rect 2686 14864 2742 14920
rect 1490 7404 1546 7440
rect 1490 7384 1492 7404
rect 1492 7384 1544 7404
rect 1544 7384 1546 7404
rect 1490 6976 1546 7032
rect 1858 7692 1860 7712
rect 1860 7692 1912 7712
rect 1912 7692 1914 7712
rect 1858 7656 1914 7692
rect 1490 5480 1546 5536
rect 1398 4936 1454 4992
rect 2226 8200 2282 8256
rect 2318 5616 2374 5672
rect 2226 5092 2282 5128
rect 2226 5072 2228 5092
rect 2228 5072 2280 5092
rect 2280 5072 2282 5092
rect 2226 4564 2228 4584
rect 2228 4564 2280 4584
rect 2280 4564 2282 4584
rect 2226 4528 2282 4564
rect 2870 13132 2872 13152
rect 2872 13132 2924 13152
rect 2924 13132 2926 13152
rect 2870 13096 2926 13132
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3422 16496 3478 16552
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 2962 12416 3018 12472
rect 2778 10240 2834 10296
rect 2778 10104 2834 10160
rect 2962 10648 3018 10704
rect 3790 15136 3846 15192
rect 3146 12688 3202 12744
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 4894 19660 4896 19680
rect 4896 19660 4948 19680
rect 4948 19660 4950 19680
rect 4894 19624 4950 19660
rect 4250 17720 4306 17776
rect 4434 17040 4490 17096
rect 4250 16632 4306 16688
rect 3882 12280 3938 12336
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3790 11092 3792 11112
rect 3792 11092 3844 11112
rect 3844 11092 3846 11112
rect 3790 11056 3846 11092
rect 4158 12824 4214 12880
rect 16854 20460 16910 20496
rect 20626 20848 20682 20904
rect 16854 20440 16856 20460
rect 16856 20440 16908 20460
rect 16908 20440 16910 20460
rect 20166 20440 20222 20496
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5814 19488 5870 19544
rect 5722 18672 5778 18728
rect 4434 13232 4490 13288
rect 3238 10104 3294 10160
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3146 9016 3202 9072
rect 2778 7792 2834 7848
rect 3054 7928 3110 7984
rect 3606 9560 3662 9616
rect 3882 9424 3938 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 2962 6296 3018 6352
rect 3146 6976 3202 7032
rect 3054 6160 3110 6216
rect 3238 6704 3294 6760
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3422 5752 3478 5808
rect 3330 5616 3386 5672
rect 3146 5344 3202 5400
rect 3974 8200 4030 8256
rect 4434 11600 4490 11656
rect 5446 18128 5502 18184
rect 5446 17584 5502 17640
rect 4986 11092 4988 11112
rect 4988 11092 5040 11112
rect 5040 11092 5042 11112
rect 4986 11056 5042 11092
rect 3238 4820 3294 4856
rect 3238 4800 3240 4820
rect 3240 4800 3292 4820
rect 3292 4800 3294 4820
rect 3238 3440 3294 3496
rect 2870 3304 2926 3360
rect 2594 2896 2650 2952
rect 2778 2760 2834 2816
rect 2962 1672 3018 1728
rect 3882 5072 3938 5128
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3698 4528 3754 4584
rect 3514 4256 3570 4312
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3698 3440 3754 3496
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4342 6180 4398 6216
rect 4342 6160 4344 6180
rect 4344 6160 4396 6180
rect 4396 6160 4398 6180
rect 4618 6704 4674 6760
rect 4434 5752 4490 5808
rect 4342 4256 4398 4312
rect 4066 4120 4122 4176
rect 4802 8880 4858 8936
rect 4802 6296 4858 6352
rect 5354 15988 5356 16008
rect 5356 15988 5408 16008
rect 5408 15988 5410 16008
rect 5354 15952 5410 15988
rect 5630 18128 5686 18184
rect 7562 19352 7618 19408
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 5998 18264 6054 18320
rect 5906 17176 5962 17232
rect 5814 14728 5870 14784
rect 5722 13776 5778 13832
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6458 16516 6514 16552
rect 6458 16496 6460 16516
rect 6460 16496 6512 16516
rect 6512 16496 6514 16516
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6734 15816 6790 15872
rect 7102 17484 7104 17504
rect 7104 17484 7156 17504
rect 7156 17484 7158 17504
rect 7102 17448 7158 17484
rect 6918 16088 6974 16144
rect 6642 14864 6698 14920
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6550 14048 6606 14104
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5906 12724 5908 12744
rect 5908 12724 5960 12744
rect 5960 12724 5962 12744
rect 5906 12688 5962 12724
rect 5630 12416 5686 12472
rect 5538 12280 5594 12336
rect 5630 11328 5686 11384
rect 5814 10104 5870 10160
rect 6642 12416 6698 12472
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6550 11872 6606 11928
rect 6550 11464 6606 11520
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 4526 4664 4582 4720
rect 4158 3032 4214 3088
rect 3974 2352 4030 2408
rect 3974 2100 4030 2136
rect 3974 2080 3976 2100
rect 3976 2080 4028 2100
rect 4028 2080 4030 2100
rect 4986 4256 5042 4312
rect 5078 4004 5134 4040
rect 5078 3984 5080 4004
rect 5080 3984 5132 4004
rect 5132 3984 5134 4004
rect 5538 5752 5594 5808
rect 5170 2896 5226 2952
rect 5078 2624 5134 2680
rect 4802 1672 4858 1728
rect 4434 1536 4490 1592
rect 5722 5752 5778 5808
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 7470 17756 7472 17776
rect 7472 17756 7524 17776
rect 7524 17756 7526 17776
rect 7470 17720 7526 17756
rect 7562 16496 7618 16552
rect 7470 15816 7526 15872
rect 7102 13504 7158 13560
rect 6918 12008 6974 12064
rect 6918 9968 6974 10024
rect 6826 9424 6882 9480
rect 5998 7928 6054 7984
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6182 6704 6238 6760
rect 5998 6568 6054 6624
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6182 5888 6238 5944
rect 5998 5752 6054 5808
rect 5814 3848 5870 3904
rect 5814 3596 5870 3632
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6734 5344 6790 5400
rect 6642 4800 6698 4856
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6182 3848 6238 3904
rect 5814 3576 5816 3596
rect 5816 3576 5868 3596
rect 5868 3576 5870 3596
rect 5446 2508 5502 2544
rect 5446 2488 5448 2508
rect 5448 2488 5500 2508
rect 5500 2488 5502 2508
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6734 3168 6790 3224
rect 5630 2760 5686 2816
rect 5722 1672 5778 1728
rect 6366 2896 6422 2952
rect 7378 12300 7434 12336
rect 7378 12280 7380 12300
rect 7380 12280 7432 12300
rect 7432 12280 7434 12300
rect 7746 16360 7802 16416
rect 7930 16396 7932 16416
rect 7932 16396 7984 16416
rect 7984 16396 7986 16416
rect 7930 16360 7986 16396
rect 7930 16088 7986 16144
rect 7654 13776 7710 13832
rect 7470 8880 7526 8936
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 9034 17604 9090 17640
rect 9034 17584 9036 17604
rect 9036 17584 9088 17604
rect 9088 17584 9090 17604
rect 8298 17076 8300 17096
rect 8300 17076 8352 17096
rect 8352 17076 8354 17096
rect 8298 17040 8354 17076
rect 8942 17060 8998 17096
rect 8942 17040 8944 17060
rect 8944 17040 8996 17060
rect 8996 17040 8998 17060
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8574 16632 8630 16688
rect 8298 13368 8354 13424
rect 8298 12824 8354 12880
rect 8298 12588 8300 12608
rect 8300 12588 8352 12608
rect 8352 12588 8354 12608
rect 8298 12552 8354 12588
rect 8206 10804 8262 10840
rect 8206 10784 8208 10804
rect 8208 10784 8260 10804
rect 8260 10784 8262 10804
rect 8022 10648 8078 10704
rect 8206 10648 8262 10704
rect 8022 10512 8078 10568
rect 6918 5480 6974 5536
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7102 5344 7158 5400
rect 7378 5072 7434 5128
rect 6642 1808 6698 1864
rect 7746 7964 7748 7984
rect 7748 7964 7800 7984
rect 7800 7964 7802 7984
rect 7746 7928 7802 7964
rect 8114 8628 8170 8664
rect 8114 8608 8116 8628
rect 8116 8608 8168 8628
rect 8168 8608 8170 8628
rect 8114 6160 8170 6216
rect 8114 5480 8170 5536
rect 8114 3984 8170 4040
rect 7654 3032 7710 3088
rect 7654 2388 7656 2408
rect 7656 2388 7708 2408
rect 7708 2388 7710 2408
rect 7654 2352 7710 2388
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9770 15408 9826 15464
rect 9678 15156 9734 15192
rect 9678 15136 9680 15156
rect 9680 15136 9732 15156
rect 9732 15136 9734 15156
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8482 6432 8538 6488
rect 8666 10648 8722 10704
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8390 5344 8446 5400
rect 8206 3440 8262 3496
rect 8574 5480 8630 5536
rect 8574 3576 8630 3632
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 9034 7792 9090 7848
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9126 5888 9182 5944
rect 9494 10512 9550 10568
rect 9678 13912 9734 13968
rect 10414 17076 10416 17096
rect 10416 17076 10468 17096
rect 10468 17076 10470 17096
rect 10414 17040 10470 17076
rect 9954 13504 10010 13560
rect 9770 12552 9826 12608
rect 10322 15136 10378 15192
rect 9126 5616 9182 5672
rect 8758 5072 8814 5128
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8942 4156 8944 4176
rect 8944 4156 8996 4176
rect 8996 4156 8998 4176
rect 8942 4120 8998 4156
rect 9126 4120 9182 4176
rect 8942 4020 8944 4040
rect 8944 4020 8996 4040
rect 8996 4020 8998 4040
rect 8942 3984 8998 4020
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8942 3440 8998 3496
rect 8206 2896 8262 2952
rect 8298 2216 8354 2272
rect 8666 3188 8722 3224
rect 8666 3168 8668 3188
rect 8668 3168 8720 3188
rect 8720 3168 8722 3188
rect 9310 4004 9366 4040
rect 9310 3984 9312 4004
rect 9312 3984 9364 4004
rect 9364 3984 9366 4004
rect 9402 3440 9458 3496
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 8574 2624 8630 2680
rect 9586 4528 9642 4584
rect 9678 2896 9734 2952
rect 10046 4664 10102 4720
rect 11794 19760 11850 19816
rect 10690 17484 10692 17504
rect 10692 17484 10744 17504
rect 10744 17484 10746 17504
rect 10690 17448 10746 17484
rect 10414 11872 10470 11928
rect 10414 11600 10470 11656
rect 10598 12144 10654 12200
rect 10598 11600 10654 11656
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11518 17584 11574 17640
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11794 17076 11796 17096
rect 11796 17076 11848 17096
rect 11848 17076 11850 17096
rect 11794 17040 11850 17076
rect 10782 12144 10838 12200
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11150 12008 11206 12064
rect 11978 15580 11980 15600
rect 11980 15580 12032 15600
rect 12032 15580 12034 15600
rect 11978 15544 12034 15580
rect 11886 15308 11888 15328
rect 11888 15308 11940 15328
rect 11940 15308 11942 15328
rect 11886 15272 11942 15308
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11978 13776 12034 13832
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11518 12552 11574 12608
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 9770 2624 9826 2680
rect 10782 8880 10838 8936
rect 10506 5752 10562 5808
rect 10690 5072 10746 5128
rect 10966 5788 10968 5808
rect 10968 5788 11020 5808
rect 11020 5788 11022 5808
rect 10966 5752 11022 5788
rect 10782 4392 10838 4448
rect 11794 12824 11850 12880
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11702 9424 11758 9480
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11794 8336 11850 8392
rect 11794 6432 11850 6488
rect 11702 6160 11758 6216
rect 11794 6024 11850 6080
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11334 4972 11336 4992
rect 11336 4972 11388 4992
rect 11388 4972 11390 4992
rect 11334 4936 11390 4972
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 10598 2488 10654 2544
rect 11978 9560 12034 9616
rect 11978 9016 12034 9072
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12346 13096 12402 13152
rect 12714 13776 12770 13832
rect 12530 11736 12586 11792
rect 12346 8880 12402 8936
rect 12162 7248 12218 7304
rect 11978 1944 12034 2000
rect 12346 3576 12402 3632
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 14370 19508 14426 19544
rect 14370 19488 14372 19508
rect 14372 19488 14424 19508
rect 14424 19488 14426 19508
rect 14554 19352 14610 19408
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 12990 14456 13046 14512
rect 13082 13504 13138 13560
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 12990 12416 13046 12472
rect 12806 6024 12862 6080
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 12990 5616 13046 5672
rect 12806 4936 12862 4992
rect 12714 2624 12770 2680
rect 13266 5752 13322 5808
rect 13358 5616 13414 5672
rect 13358 3712 13414 3768
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14554 15272 14610 15328
rect 15106 17312 15162 17368
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 14278 9424 14334 9480
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13726 6160 13782 6216
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13542 4664 13598 4720
rect 14554 11600 14610 11656
rect 14370 7248 14426 7304
rect 14462 7112 14518 7168
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13910 4120 13966 4176
rect 13358 2896 13414 2952
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14370 3732 14426 3768
rect 14370 3712 14372 3732
rect 14372 3712 14424 3732
rect 14424 3712 14426 3732
rect 13174 2488 13230 2544
rect 12254 2080 12310 2136
rect 12254 1808 12310 1864
rect 13726 2896 13782 2952
rect 13910 3188 13966 3224
rect 13910 3168 13912 3188
rect 13912 3168 13964 3188
rect 13964 3168 13966 3188
rect 14094 3068 14096 3088
rect 14096 3068 14148 3088
rect 14148 3068 14150 3088
rect 14094 3032 14150 3068
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15658 17992 15714 18048
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 17038 19116 17040 19136
rect 17040 19116 17092 19136
rect 17092 19116 17094 19136
rect 17038 19080 17094 19116
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16210 18128 16266 18184
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 15842 14864 15898 14920
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16946 15156 17002 15192
rect 16946 15136 16948 15156
rect 16948 15136 17000 15156
rect 17000 15136 17002 15156
rect 16302 14456 16358 14512
rect 16210 14320 16266 14376
rect 15658 10240 15714 10296
rect 15382 8880 15438 8936
rect 14646 4528 14702 4584
rect 14922 5072 14978 5128
rect 14922 4820 14978 4856
rect 14922 4800 14924 4820
rect 14924 4800 14976 4820
rect 14976 4800 14978 4820
rect 15382 6432 15438 6488
rect 15290 5480 15346 5536
rect 15474 6296 15530 6352
rect 15382 3984 15438 4040
rect 16026 5752 16082 5808
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16210 6296 16266 6352
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 17958 19760 18014 19816
rect 17498 19352 17554 19408
rect 17130 12688 17186 12744
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 17038 12144 17094 12200
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16118 5480 16174 5536
rect 15934 4936 15990 4992
rect 14830 3032 14886 3088
rect 16118 3848 16174 3904
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16210 3576 16266 3632
rect 16946 3984 17002 4040
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 18602 17484 18604 17504
rect 18604 17484 18656 17504
rect 18656 17484 18658 17504
rect 18602 17448 18658 17484
rect 18694 16632 18750 16688
rect 18602 13776 18658 13832
rect 18418 13252 18474 13288
rect 18418 13232 18420 13252
rect 18420 13232 18472 13252
rect 18472 13232 18474 13252
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17866 7792 17922 7848
rect 18142 7384 18198 7440
rect 18050 6860 18106 6896
rect 18050 6840 18052 6860
rect 18052 6840 18104 6860
rect 18104 6840 18106 6860
rect 17682 4120 17738 4176
rect 17958 5072 18014 5128
rect 18602 12008 18658 12064
rect 18418 9424 18474 9480
rect 18418 8880 18474 8936
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19614 18128 19670 18184
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19522 13912 19578 13968
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18786 11056 18842 11112
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 20718 20032 20774 20088
rect 20626 19216 20682 19272
rect 20718 18028 20720 18048
rect 20720 18028 20772 18048
rect 20772 18028 20774 18048
rect 20718 17992 20774 18028
rect 19890 16904 19946 16960
rect 19798 16632 19854 16688
rect 19890 16496 19946 16552
rect 20166 16768 20222 16824
rect 19798 12688 19854 12744
rect 20626 16632 20682 16688
rect 20166 10648 20222 10704
rect 20166 10240 20222 10296
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 18786 7928 18842 7984
rect 18418 6704 18474 6760
rect 18418 5752 18474 5808
rect 18326 5072 18382 5128
rect 17958 4120 18014 4176
rect 18142 3068 18144 3088
rect 18144 3068 18196 3088
rect 18196 3068 18198 3088
rect 18142 3032 18198 3068
rect 18602 5480 18658 5536
rect 18602 5108 18604 5128
rect 18604 5108 18656 5128
rect 18656 5108 18658 5128
rect 18602 5072 18658 5108
rect 17866 2488 17922 2544
rect 18234 2488 18290 2544
rect 17958 1672 18014 1728
rect 18786 7112 18842 7168
rect 18878 6160 18934 6216
rect 18786 5616 18842 5672
rect 18694 1944 18750 2000
rect 18878 4664 18934 4720
rect 18878 3848 18934 3904
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19154 7420 19156 7440
rect 19156 7420 19208 7440
rect 19208 7420 19210 7440
rect 19154 7384 19210 7420
rect 19706 9460 19708 9480
rect 19708 9460 19760 9480
rect 19760 9460 19762 9480
rect 19706 9424 19762 9460
rect 19798 7520 19854 7576
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19338 6840 19394 6896
rect 19246 6704 19302 6760
rect 19614 6860 19670 6896
rect 19614 6840 19616 6860
rect 19616 6840 19668 6860
rect 19668 6840 19670 6860
rect 19798 6840 19854 6896
rect 19522 6432 19578 6488
rect 19062 6296 19118 6352
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 20074 7248 20130 7304
rect 20534 13232 20590 13288
rect 20718 16360 20774 16416
rect 20718 15972 20774 16008
rect 20718 15952 20720 15972
rect 20720 15952 20772 15972
rect 20772 15952 20774 15972
rect 20810 15000 20866 15056
rect 20534 12280 20590 12336
rect 20534 11736 20590 11792
rect 21270 19760 21326 19816
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21362 18808 21418 18864
rect 21270 18264 21326 18320
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21362 17584 21418 17640
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 21270 17176 21326 17232
rect 21270 15544 21326 15600
rect 21362 14728 21418 14784
rect 21270 14320 21326 14376
rect 21270 13912 21326 13968
rect 21270 13524 21326 13560
rect 21270 13504 21272 13524
rect 21272 13504 21324 13524
rect 21324 13504 21326 13524
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 20534 9968 20590 10024
rect 20442 9560 20498 9616
rect 20534 9016 20590 9072
rect 20442 7520 20498 7576
rect 20258 6432 20314 6488
rect 19706 4528 19762 4584
rect 19338 3068 19340 3088
rect 19340 3068 19392 3088
rect 19392 3068 19394 3088
rect 19338 3032 19394 3068
rect 19154 2896 19210 2952
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20534 6976 20590 7032
rect 20350 5364 20406 5400
rect 20350 5344 20352 5364
rect 20352 5344 20404 5364
rect 20404 5344 20406 5364
rect 20166 3052 20222 3088
rect 20166 3032 20168 3052
rect 20168 3032 20220 3052
rect 20220 3032 20222 3052
rect 20902 10104 20958 10160
rect 21270 11464 21326 11520
rect 21270 8472 21326 8528
rect 21086 7656 21142 7712
rect 20810 4664 20866 4720
rect 20718 3440 20774 3496
rect 20442 3168 20498 3224
rect 21086 5208 21142 5264
rect 21270 5752 21326 5808
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21362 2352 21418 2408
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
<< metal3 >>
rect 0 21314 800 21344
rect 2957 21314 3023 21317
rect 0 21312 3023 21314
rect 0 21256 2962 21312
rect 3018 21256 3023 21312
rect 0 21254 3023 21256
rect 0 21224 800 21254
rect 2957 21251 3023 21254
rect 18689 21314 18755 21317
rect 22200 21314 23000 21344
rect 18689 21312 23000 21314
rect 18689 21256 18694 21312
rect 18750 21256 23000 21312
rect 18689 21254 23000 21256
rect 18689 21251 18755 21254
rect 22200 21224 23000 21254
rect 0 20906 800 20936
rect 1945 20906 2011 20909
rect 0 20904 2011 20906
rect 0 20848 1950 20904
rect 2006 20848 2011 20904
rect 0 20846 2011 20848
rect 0 20816 800 20846
rect 1945 20843 2011 20846
rect 20621 20906 20687 20909
rect 22200 20906 23000 20936
rect 20621 20904 23000 20906
rect 20621 20848 20626 20904
rect 20682 20848 23000 20904
rect 20621 20846 23000 20848
rect 20621 20843 20687 20846
rect 22200 20816 23000 20846
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 21738 20639 22054 20640
rect 0 20498 800 20528
rect 2037 20498 2103 20501
rect 0 20496 2103 20498
rect 0 20440 2042 20496
rect 2098 20440 2103 20496
rect 0 20438 2103 20440
rect 0 20408 800 20438
rect 2037 20435 2103 20438
rect 5257 20498 5323 20501
rect 16849 20498 16915 20501
rect 17166 20498 17172 20500
rect 5257 20496 17172 20498
rect 5257 20440 5262 20496
rect 5318 20440 16854 20496
rect 16910 20440 17172 20496
rect 5257 20438 17172 20440
rect 5257 20435 5323 20438
rect 16849 20435 16915 20438
rect 17166 20436 17172 20438
rect 17236 20436 17242 20500
rect 20161 20498 20227 20501
rect 22200 20498 23000 20528
rect 20161 20496 23000 20498
rect 20161 20440 20166 20496
rect 20222 20440 23000 20496
rect 20161 20438 23000 20440
rect 20161 20435 20227 20438
rect 22200 20408 23000 20438
rect 1301 20362 1367 20365
rect 4521 20362 4587 20365
rect 1301 20360 4587 20362
rect 1301 20304 1306 20360
rect 1362 20304 4526 20360
rect 4582 20304 4587 20360
rect 1301 20302 4587 20304
rect 1301 20299 1367 20302
rect 4521 20299 4587 20302
rect 3545 20160 3861 20161
rect 0 20090 800 20120
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 19139 20095 19455 20096
rect 1485 20090 1551 20093
rect 0 20088 1551 20090
rect 0 20032 1490 20088
rect 1546 20032 1551 20088
rect 0 20030 1551 20032
rect 0 20000 800 20030
rect 1485 20027 1551 20030
rect 20713 20090 20779 20093
rect 22200 20090 23000 20120
rect 20713 20088 23000 20090
rect 20713 20032 20718 20088
rect 20774 20032 23000 20088
rect 20713 20030 23000 20032
rect 20713 20027 20779 20030
rect 22200 20000 23000 20030
rect 1117 19818 1183 19821
rect 4521 19818 4587 19821
rect 1117 19816 4587 19818
rect 1117 19760 1122 19816
rect 1178 19760 4526 19816
rect 4582 19760 4587 19816
rect 1117 19758 4587 19760
rect 1117 19755 1183 19758
rect 4521 19755 4587 19758
rect 11789 19818 11855 19821
rect 17953 19818 18019 19821
rect 11789 19816 18019 19818
rect 11789 19760 11794 19816
rect 11850 19760 17958 19816
rect 18014 19760 18019 19816
rect 11789 19758 18019 19760
rect 11789 19755 11855 19758
rect 17953 19755 18019 19758
rect 21265 19818 21331 19821
rect 21265 19816 22202 19818
rect 21265 19760 21270 19816
rect 21326 19760 22202 19816
rect 21265 19758 22202 19760
rect 21265 19755 21331 19758
rect 22142 19712 22202 19758
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 4889 19682 4955 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 1718 19680 4955 19682
rect 1718 19624 4894 19680
rect 4950 19624 4955 19680
rect 1718 19622 4955 19624
rect 22142 19622 23000 19712
rect 933 19546 999 19549
rect 1718 19546 1778 19622
rect 4889 19619 4955 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22200 19592 23000 19622
rect 21738 19551 22054 19552
rect 933 19544 1778 19546
rect 933 19488 938 19544
rect 994 19488 1778 19544
rect 933 19486 1778 19488
rect 2681 19546 2747 19549
rect 3693 19546 3759 19549
rect 3877 19548 3943 19549
rect 3877 19546 3924 19548
rect 2681 19544 3759 19546
rect 2681 19488 2686 19544
rect 2742 19488 3698 19544
rect 3754 19488 3759 19544
rect 2681 19486 3759 19488
rect 3832 19544 3924 19546
rect 3832 19488 3882 19544
rect 3832 19486 3924 19488
rect 933 19483 999 19486
rect 2681 19483 2747 19486
rect 3693 19483 3759 19486
rect 3877 19484 3924 19486
rect 3988 19484 3994 19548
rect 4061 19546 4127 19549
rect 5809 19546 5875 19549
rect 4061 19544 5875 19546
rect 4061 19488 4066 19544
rect 4122 19488 5814 19544
rect 5870 19488 5875 19544
rect 4061 19486 5875 19488
rect 3877 19483 3943 19484
rect 4061 19483 4127 19486
rect 5809 19483 5875 19486
rect 14365 19546 14431 19549
rect 14590 19546 14596 19548
rect 14365 19544 14596 19546
rect 14365 19488 14370 19544
rect 14426 19488 14596 19544
rect 14365 19486 14596 19488
rect 14365 19483 14431 19486
rect 14590 19484 14596 19486
rect 14660 19484 14666 19548
rect 1158 19348 1164 19412
rect 1228 19410 1234 19412
rect 7557 19410 7623 19413
rect 1228 19408 7623 19410
rect 1228 19352 7562 19408
rect 7618 19352 7623 19408
rect 1228 19350 7623 19352
rect 1228 19348 1234 19350
rect 7557 19347 7623 19350
rect 14406 19348 14412 19412
rect 14476 19410 14482 19412
rect 14549 19410 14615 19413
rect 14476 19408 14615 19410
rect 14476 19352 14554 19408
rect 14610 19352 14615 19408
rect 14476 19350 14615 19352
rect 14476 19348 14482 19350
rect 14549 19347 14615 19350
rect 17493 19412 17559 19413
rect 17493 19408 17540 19412
rect 17604 19410 17610 19412
rect 17493 19352 17498 19408
rect 17493 19348 17540 19352
rect 17604 19350 17650 19410
rect 17604 19348 17610 19350
rect 17493 19347 17559 19348
rect 0 19274 800 19304
rect 2037 19274 2103 19277
rect 0 19272 2103 19274
rect 0 19216 2042 19272
rect 2098 19216 2103 19272
rect 0 19214 2103 19216
rect 0 19184 800 19214
rect 2037 19211 2103 19214
rect 20621 19274 20687 19277
rect 22200 19274 23000 19304
rect 20621 19272 23000 19274
rect 20621 19216 20626 19272
rect 20682 19216 23000 19272
rect 20621 19214 23000 19216
rect 20621 19211 20687 19214
rect 22200 19184 23000 19214
rect 17033 19140 17099 19141
rect 16982 19076 16988 19140
rect 17052 19138 17099 19140
rect 17052 19136 17144 19138
rect 17094 19080 17144 19136
rect 17052 19078 17144 19080
rect 17052 19076 17099 19078
rect 17033 19075 17099 19076
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 19139 19007 19455 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 21357 18866 21423 18869
rect 22200 18866 23000 18896
rect 21357 18864 23000 18866
rect 21357 18808 21362 18864
rect 21418 18808 23000 18864
rect 21357 18806 23000 18808
rect 21357 18803 21423 18806
rect 22200 18776 23000 18806
rect 4654 18668 4660 18732
rect 4724 18730 4730 18732
rect 5717 18730 5783 18733
rect 4724 18728 5783 18730
rect 4724 18672 5722 18728
rect 5778 18672 5783 18728
rect 4724 18670 5783 18672
rect 4724 18668 4730 18670
rect 5717 18667 5783 18670
rect 6144 18528 6460 18529
rect 0 18458 800 18488
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 21738 18463 22054 18464
rect 1485 18458 1551 18461
rect 22200 18458 23000 18488
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 22142 18368 23000 18458
rect 5758 18260 5764 18324
rect 5828 18322 5834 18324
rect 5993 18322 6059 18325
rect 5828 18320 6059 18322
rect 5828 18264 5998 18320
rect 6054 18264 6059 18320
rect 5828 18262 6059 18264
rect 5828 18260 5834 18262
rect 5993 18259 6059 18262
rect 21265 18322 21331 18325
rect 22142 18322 22202 18368
rect 21265 18320 22202 18322
rect 21265 18264 21270 18320
rect 21326 18264 22202 18320
rect 21265 18262 22202 18264
rect 21265 18259 21331 18262
rect 2078 18124 2084 18188
rect 2148 18186 2154 18188
rect 5441 18186 5507 18189
rect 2148 18184 5507 18186
rect 2148 18128 5446 18184
rect 5502 18128 5507 18184
rect 2148 18126 5507 18128
rect 2148 18124 2154 18126
rect 5441 18123 5507 18126
rect 5625 18186 5691 18189
rect 9990 18186 9996 18188
rect 5625 18184 9996 18186
rect 5625 18128 5630 18184
rect 5686 18128 9996 18184
rect 5625 18126 9996 18128
rect 5625 18123 5691 18126
rect 9990 18124 9996 18126
rect 10060 18186 10066 18188
rect 16205 18186 16271 18189
rect 19609 18186 19675 18189
rect 10060 18184 16271 18186
rect 10060 18128 16210 18184
rect 16266 18128 16271 18184
rect 10060 18126 16271 18128
rect 10060 18124 10066 18126
rect 16205 18123 16271 18126
rect 18094 18184 19675 18186
rect 18094 18128 19614 18184
rect 19670 18128 19675 18184
rect 18094 18126 19675 18128
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 15510 17988 15516 18052
rect 15580 18050 15586 18052
rect 15653 18050 15719 18053
rect 15580 18048 15719 18050
rect 15580 17992 15658 18048
rect 15714 17992 15719 18048
rect 15580 17990 15719 17992
rect 15580 17988 15586 17990
rect 15653 17987 15719 17990
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 933 17778 999 17781
rect 4245 17778 4311 17781
rect 933 17776 4311 17778
rect 933 17720 938 17776
rect 994 17720 4250 17776
rect 4306 17720 4311 17776
rect 933 17718 4311 17720
rect 933 17715 999 17718
rect 4245 17715 4311 17718
rect 7465 17778 7531 17781
rect 18094 17778 18154 18126
rect 19609 18123 19675 18126
rect 20713 18050 20779 18053
rect 22200 18050 23000 18080
rect 20713 18048 23000 18050
rect 20713 17992 20718 18048
rect 20774 17992 23000 18048
rect 20713 17990 23000 17992
rect 20713 17987 20779 17990
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22200 17960 23000 17990
rect 19139 17919 19455 17920
rect 7465 17776 18154 17778
rect 7465 17720 7470 17776
rect 7526 17720 18154 17776
rect 7465 17718 18154 17720
rect 7465 17715 7531 17718
rect 0 17642 800 17672
rect 2037 17642 2103 17645
rect 0 17640 2103 17642
rect 0 17584 2042 17640
rect 2098 17584 2103 17640
rect 0 17582 2103 17584
rect 0 17552 800 17582
rect 2037 17579 2103 17582
rect 5441 17642 5507 17645
rect 9029 17642 9095 17645
rect 5441 17640 9095 17642
rect 5441 17584 5446 17640
rect 5502 17584 9034 17640
rect 9090 17584 9095 17640
rect 5441 17582 9095 17584
rect 5441 17579 5507 17582
rect 9029 17579 9095 17582
rect 11094 17580 11100 17644
rect 11164 17642 11170 17644
rect 11513 17642 11579 17645
rect 11164 17640 11579 17642
rect 11164 17584 11518 17640
rect 11574 17584 11579 17640
rect 11164 17582 11579 17584
rect 11164 17580 11170 17582
rect 11513 17579 11579 17582
rect 21357 17642 21423 17645
rect 22200 17642 23000 17672
rect 21357 17640 23000 17642
rect 21357 17584 21362 17640
rect 21418 17584 23000 17640
rect 21357 17582 23000 17584
rect 21357 17579 21423 17582
rect 22200 17552 23000 17582
rect 7097 17506 7163 17509
rect 10685 17508 10751 17509
rect 18597 17508 18663 17509
rect 7782 17506 7788 17508
rect 7097 17504 7788 17506
rect 7097 17448 7102 17504
rect 7158 17448 7788 17504
rect 7097 17446 7788 17448
rect 7097 17443 7163 17446
rect 7782 17444 7788 17446
rect 7852 17444 7858 17508
rect 10685 17506 10732 17508
rect 10640 17504 10732 17506
rect 10640 17448 10690 17504
rect 10640 17446 10732 17448
rect 10685 17444 10732 17446
rect 10796 17444 10802 17508
rect 18597 17506 18644 17508
rect 18552 17504 18644 17506
rect 18552 17448 18602 17504
rect 18552 17446 18644 17448
rect 18597 17444 18644 17446
rect 18708 17444 18714 17508
rect 10685 17443 10751 17444
rect 18597 17443 18663 17444
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 21738 17375 22054 17376
rect 14958 17308 14964 17372
rect 15028 17370 15034 17372
rect 15101 17370 15167 17373
rect 15028 17368 15167 17370
rect 15028 17312 15106 17368
rect 15162 17312 15167 17368
rect 15028 17310 15167 17312
rect 15028 17308 15034 17310
rect 15101 17307 15167 17310
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 5901 17234 5967 17237
rect 9806 17234 9812 17236
rect 5901 17232 9812 17234
rect 5901 17176 5906 17232
rect 5962 17176 9812 17232
rect 5901 17174 9812 17176
rect 5901 17171 5967 17174
rect 9806 17172 9812 17174
rect 9876 17172 9882 17236
rect 21265 17234 21331 17237
rect 22200 17234 23000 17264
rect 21265 17232 23000 17234
rect 21265 17176 21270 17232
rect 21326 17176 23000 17232
rect 21265 17174 23000 17176
rect 21265 17171 21331 17174
rect 22200 17144 23000 17174
rect 3182 17036 3188 17100
rect 3252 17098 3258 17100
rect 4429 17098 4495 17101
rect 3252 17096 4495 17098
rect 3252 17040 4434 17096
rect 4490 17040 4495 17096
rect 3252 17038 4495 17040
rect 3252 17036 3258 17038
rect 4429 17035 4495 17038
rect 8293 17098 8359 17101
rect 8937 17098 9003 17101
rect 8293 17096 9003 17098
rect 8293 17040 8298 17096
rect 8354 17040 8942 17096
rect 8998 17040 9003 17096
rect 8293 17038 9003 17040
rect 8293 17035 8359 17038
rect 8937 17035 9003 17038
rect 10409 17098 10475 17101
rect 11789 17098 11855 17101
rect 10409 17096 11855 17098
rect 10409 17040 10414 17096
rect 10470 17040 11794 17096
rect 11850 17040 11855 17096
rect 10409 17038 11855 17040
rect 10409 17035 10475 17038
rect 11789 17035 11855 17038
rect 19885 16962 19951 16965
rect 19885 16960 19994 16962
rect 19885 16904 19890 16960
rect 19946 16904 19994 16960
rect 19885 16899 19994 16904
rect 3545 16896 3861 16897
rect 0 16826 800 16856
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 19139 16831 19455 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 2998 16628 3004 16692
rect 3068 16690 3074 16692
rect 4245 16690 4311 16693
rect 8569 16692 8635 16693
rect 8518 16690 8524 16692
rect 3068 16688 4311 16690
rect 3068 16632 4250 16688
rect 4306 16632 4311 16688
rect 3068 16630 4311 16632
rect 8478 16630 8524 16690
rect 8588 16688 8635 16692
rect 8630 16632 8635 16688
rect 3068 16628 3074 16630
rect 4245 16627 4311 16630
rect 8518 16628 8524 16630
rect 8588 16628 8635 16632
rect 8569 16627 8635 16628
rect 18689 16690 18755 16693
rect 19793 16690 19859 16693
rect 18689 16688 19859 16690
rect 18689 16632 18694 16688
rect 18750 16632 19798 16688
rect 19854 16632 19859 16688
rect 18689 16630 19859 16632
rect 18689 16627 18755 16630
rect 19793 16627 19859 16630
rect 19934 16557 19994 16899
rect 20161 16826 20227 16829
rect 22200 16826 23000 16856
rect 20161 16824 23000 16826
rect 20161 16768 20166 16824
rect 20222 16768 23000 16824
rect 20161 16766 23000 16768
rect 20161 16763 20227 16766
rect 22200 16736 23000 16766
rect 20478 16628 20484 16692
rect 20548 16690 20554 16692
rect 20621 16690 20687 16693
rect 20548 16688 20687 16690
rect 20548 16632 20626 16688
rect 20682 16632 20687 16688
rect 20548 16630 20687 16632
rect 20548 16628 20554 16630
rect 20621 16627 20687 16630
rect 2630 16492 2636 16556
rect 2700 16554 2706 16556
rect 3417 16554 3483 16557
rect 2700 16552 3483 16554
rect 2700 16496 3422 16552
rect 3478 16496 3483 16552
rect 2700 16494 3483 16496
rect 2700 16492 2706 16494
rect 3417 16491 3483 16494
rect 6453 16554 6519 16557
rect 7557 16554 7623 16557
rect 6453 16552 7623 16554
rect 6453 16496 6458 16552
rect 6514 16496 7562 16552
rect 7618 16496 7623 16552
rect 6453 16494 7623 16496
rect 6453 16491 6519 16494
rect 7557 16491 7623 16494
rect 19885 16552 19994 16557
rect 19885 16496 19890 16552
rect 19946 16496 19994 16552
rect 19885 16494 19994 16496
rect 20854 16494 22202 16554
rect 19885 16491 19951 16494
rect 0 16418 800 16448
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 7598 16356 7604 16420
rect 7668 16418 7674 16420
rect 7741 16418 7807 16421
rect 7925 16418 7991 16421
rect 7668 16416 7991 16418
rect 7668 16360 7746 16416
rect 7802 16360 7930 16416
rect 7986 16360 7991 16416
rect 7668 16358 7991 16360
rect 7668 16356 7674 16358
rect 7741 16355 7807 16358
rect 7925 16355 7991 16358
rect 20713 16418 20779 16421
rect 20854 16418 20914 16494
rect 20713 16416 20914 16418
rect 20713 16360 20718 16416
rect 20774 16360 20914 16416
rect 20713 16358 20914 16360
rect 22142 16448 22202 16494
rect 22142 16358 23000 16448
rect 20713 16355 20779 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22200 16328 23000 16358
rect 21738 16287 22054 16288
rect 5206 16084 5212 16148
rect 5276 16146 5282 16148
rect 6913 16146 6979 16149
rect 7925 16146 7991 16149
rect 5276 16144 7991 16146
rect 5276 16088 6918 16144
rect 6974 16088 7930 16144
rect 7986 16088 7991 16144
rect 5276 16086 7991 16088
rect 5276 16084 5282 16086
rect 6913 16083 6979 16086
rect 7925 16083 7991 16086
rect 0 16010 800 16040
rect 1393 16010 1459 16013
rect 0 16008 1459 16010
rect 0 15952 1398 16008
rect 1454 15952 1459 16008
rect 0 15950 1459 15952
rect 0 15920 800 15950
rect 1393 15947 1459 15950
rect 5349 16010 5415 16013
rect 7782 16010 7788 16012
rect 5349 16008 7788 16010
rect 5349 15952 5354 16008
rect 5410 15952 7788 16008
rect 5349 15950 7788 15952
rect 5349 15947 5415 15950
rect 7782 15948 7788 15950
rect 7852 15948 7858 16012
rect 20713 16010 20779 16013
rect 22200 16010 23000 16040
rect 20713 16008 23000 16010
rect 20713 15952 20718 16008
rect 20774 15952 23000 16008
rect 20713 15950 23000 15952
rect 20713 15947 20779 15950
rect 22200 15920 23000 15950
rect 6729 15874 6795 15877
rect 7465 15874 7531 15877
rect 6729 15872 7531 15874
rect 6729 15816 6734 15872
rect 6790 15816 7470 15872
rect 7526 15816 7531 15872
rect 6729 15814 7531 15816
rect 6729 15811 6795 15814
rect 7465 15811 7531 15814
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 19139 15743 19455 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 11973 15602 12039 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 1718 15600 12039 15602
rect 1718 15544 11978 15600
rect 12034 15544 12039 15600
rect 1718 15542 12039 15544
rect 974 15404 980 15468
rect 1044 15466 1050 15468
rect 1718 15466 1778 15542
rect 11973 15539 12039 15542
rect 21265 15602 21331 15605
rect 22200 15602 23000 15632
rect 21265 15600 23000 15602
rect 21265 15544 21270 15600
rect 21326 15544 23000 15600
rect 21265 15542 23000 15544
rect 21265 15539 21331 15542
rect 22200 15512 23000 15542
rect 9765 15466 9831 15469
rect 1044 15406 1778 15466
rect 4294 15464 9831 15466
rect 4294 15408 9770 15464
rect 9826 15408 9831 15464
rect 4294 15406 9831 15408
rect 1044 15404 1050 15406
rect 0 15194 800 15224
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 3785 15194 3851 15197
rect 4294 15196 4354 15406
rect 9765 15403 9831 15406
rect 11881 15330 11947 15333
rect 12198 15330 12204 15332
rect 11881 15328 12204 15330
rect 11881 15272 11886 15328
rect 11942 15272 12204 15328
rect 11881 15270 12204 15272
rect 11881 15267 11947 15270
rect 12198 15268 12204 15270
rect 12268 15268 12274 15332
rect 14549 15330 14615 15333
rect 15326 15330 15332 15332
rect 14549 15328 15332 15330
rect 14549 15272 14554 15328
rect 14610 15272 15332 15328
rect 14549 15270 15332 15272
rect 14549 15267 14615 15270
rect 15326 15268 15332 15270
rect 15396 15268 15402 15332
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 21738 15199 22054 15200
rect 4286 15194 4292 15196
rect 3785 15192 4292 15194
rect 3785 15136 3790 15192
rect 3846 15136 4292 15192
rect 3785 15134 4292 15136
rect 3785 15131 3851 15134
rect 4286 15132 4292 15134
rect 4356 15132 4362 15196
rect 9673 15194 9739 15197
rect 10317 15194 10383 15197
rect 9673 15192 10383 15194
rect 9673 15136 9678 15192
rect 9734 15136 10322 15192
rect 10378 15136 10383 15192
rect 9673 15134 10383 15136
rect 9673 15131 9739 15134
rect 10317 15131 10383 15134
rect 10726 15132 10732 15196
rect 10796 15194 10802 15196
rect 16941 15194 17007 15197
rect 17166 15194 17172 15196
rect 10796 15134 11162 15194
rect 10796 15132 10802 15134
rect 11102 15058 11162 15134
rect 16941 15192 17172 15194
rect 16941 15136 16946 15192
rect 17002 15136 17172 15192
rect 16941 15134 17172 15136
rect 16941 15131 17007 15134
rect 17166 15132 17172 15134
rect 17236 15132 17242 15196
rect 22200 15194 23000 15224
rect 22142 15104 23000 15194
rect 19006 15058 19012 15060
rect 11102 14998 19012 15058
rect 19006 14996 19012 14998
rect 19076 14996 19082 15060
rect 20805 15058 20871 15061
rect 22142 15058 22202 15104
rect 20805 15056 22202 15058
rect 20805 15000 20810 15056
rect 20866 15000 22202 15056
rect 20805 14998 22202 15000
rect 20805 14995 20871 14998
rect 2446 14860 2452 14924
rect 2516 14922 2522 14924
rect 2681 14922 2747 14925
rect 6637 14922 6703 14925
rect 15837 14922 15903 14925
rect 2516 14920 5090 14922
rect 2516 14864 2686 14920
rect 2742 14864 5090 14920
rect 2516 14862 5090 14864
rect 2516 14860 2522 14862
rect 2681 14859 2747 14862
rect 0 14786 800 14816
rect 2129 14786 2195 14789
rect 0 14784 2195 14786
rect 0 14728 2134 14784
rect 2190 14728 2195 14784
rect 0 14726 2195 14728
rect 5030 14786 5090 14862
rect 6637 14920 15903 14922
rect 6637 14864 6642 14920
rect 6698 14864 15842 14920
rect 15898 14864 15903 14920
rect 6637 14862 15903 14864
rect 6637 14859 6703 14862
rect 15837 14859 15903 14862
rect 5809 14786 5875 14789
rect 6678 14786 6684 14788
rect 5030 14784 6684 14786
rect 5030 14728 5814 14784
rect 5870 14728 6684 14784
rect 5030 14726 6684 14728
rect 0 14696 800 14726
rect 2129 14723 2195 14726
rect 5809 14723 5875 14726
rect 6678 14724 6684 14726
rect 6748 14724 6754 14788
rect 21357 14786 21423 14789
rect 22200 14786 23000 14816
rect 21357 14784 23000 14786
rect 21357 14728 21362 14784
rect 21418 14728 23000 14784
rect 21357 14726 23000 14728
rect 21357 14723 21423 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22200 14696 23000 14726
rect 19139 14655 19455 14656
rect 1669 14514 1735 14517
rect 12985 14514 13051 14517
rect 1669 14512 13051 14514
rect 1669 14456 1674 14512
rect 1730 14456 12990 14512
rect 13046 14456 13051 14512
rect 1669 14454 13051 14456
rect 1669 14451 1735 14454
rect 12985 14451 13051 14454
rect 16297 14514 16363 14517
rect 17534 14514 17540 14516
rect 16297 14512 17540 14514
rect 16297 14456 16302 14512
rect 16358 14456 17540 14512
rect 16297 14454 17540 14456
rect 16297 14451 16363 14454
rect 17534 14452 17540 14454
rect 17604 14452 17610 14516
rect 0 14378 800 14408
rect 1485 14378 1551 14381
rect 0 14376 1551 14378
rect 0 14320 1490 14376
rect 1546 14320 1551 14376
rect 0 14318 1551 14320
rect 0 14288 800 14318
rect 1485 14315 1551 14318
rect 7598 14316 7604 14380
rect 7668 14378 7674 14380
rect 16205 14378 16271 14381
rect 7668 14376 16271 14378
rect 7668 14320 16210 14376
rect 16266 14320 16271 14376
rect 7668 14318 16271 14320
rect 7668 14316 7674 14318
rect 16205 14315 16271 14318
rect 21265 14378 21331 14381
rect 22200 14378 23000 14408
rect 21265 14376 23000 14378
rect 21265 14320 21270 14376
rect 21326 14320 23000 14376
rect 21265 14318 23000 14320
rect 21265 14315 21331 14318
rect 22200 14288 23000 14318
rect 8334 14180 8340 14244
rect 8404 14242 8410 14244
rect 11094 14242 11100 14244
rect 8404 14182 11100 14242
rect 8404 14180 8410 14182
rect 11094 14180 11100 14182
rect 11164 14180 11170 14244
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 21738 14111 22054 14112
rect 6545 14106 6611 14109
rect 7046 14106 7052 14108
rect 6545 14104 7052 14106
rect 6545 14048 6550 14104
rect 6606 14048 7052 14104
rect 6545 14046 7052 14048
rect 6545 14043 6611 14046
rect 7046 14044 7052 14046
rect 7116 14106 7122 14108
rect 7116 14046 9874 14106
rect 7116 14044 7122 14046
rect 0 13970 800 14000
rect 2129 13970 2195 13973
rect 0 13968 2195 13970
rect 0 13912 2134 13968
rect 2190 13912 2195 13968
rect 0 13910 2195 13912
rect 0 13880 800 13910
rect 2129 13907 2195 13910
rect 5574 13908 5580 13972
rect 5644 13970 5650 13972
rect 9673 13970 9739 13973
rect 5644 13968 9739 13970
rect 5644 13912 9678 13968
rect 9734 13912 9739 13968
rect 5644 13910 9739 13912
rect 9814 13970 9874 14046
rect 19517 13970 19583 13973
rect 9814 13968 19583 13970
rect 9814 13912 19522 13968
rect 19578 13912 19583 13968
rect 9814 13910 19583 13912
rect 5644 13908 5650 13910
rect 9673 13907 9739 13910
rect 19517 13907 19583 13910
rect 21265 13970 21331 13973
rect 22200 13970 23000 14000
rect 21265 13968 23000 13970
rect 21265 13912 21270 13968
rect 21326 13912 23000 13968
rect 21265 13910 23000 13912
rect 21265 13907 21331 13910
rect 22200 13880 23000 13910
rect 3918 13772 3924 13836
rect 3988 13772 3994 13836
rect 4102 13772 4108 13836
rect 4172 13834 4178 13836
rect 5717 13834 5783 13837
rect 4172 13832 5783 13834
rect 4172 13776 5722 13832
rect 5778 13776 5783 13832
rect 4172 13774 5783 13776
rect 4172 13772 4178 13774
rect 3926 13698 3986 13772
rect 5717 13771 5783 13774
rect 7649 13834 7715 13837
rect 11973 13836 12039 13837
rect 12709 13836 12775 13837
rect 7966 13834 7972 13836
rect 7649 13832 7972 13834
rect 7649 13776 7654 13832
rect 7710 13776 7972 13832
rect 7649 13774 7972 13776
rect 7649 13771 7715 13774
rect 7966 13772 7972 13774
rect 8036 13772 8042 13836
rect 11973 13832 12020 13836
rect 12084 13834 12090 13836
rect 11973 13776 11978 13832
rect 11973 13772 12020 13776
rect 12084 13774 12130 13834
rect 12709 13832 12756 13836
rect 12820 13834 12826 13836
rect 18597 13834 18663 13837
rect 20110 13834 20116 13836
rect 12709 13776 12714 13832
rect 12084 13772 12090 13774
rect 12709 13772 12756 13776
rect 12820 13774 12866 13834
rect 18597 13832 20116 13834
rect 18597 13776 18602 13832
rect 18658 13776 20116 13832
rect 18597 13774 20116 13776
rect 12820 13772 12826 13774
rect 11973 13771 12039 13772
rect 12709 13771 12775 13772
rect 18597 13771 18663 13774
rect 20110 13772 20116 13774
rect 20180 13772 20186 13836
rect 3926 13638 8586 13698
rect 3545 13632 3861 13633
rect 0 13562 800 13592
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 1485 13562 1551 13565
rect 7097 13562 7163 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 4294 13560 7163 13562
rect 4294 13504 7102 13560
rect 7158 13504 7163 13560
rect 4294 13502 7163 13504
rect 1761 13426 1827 13429
rect 4294 13426 4354 13502
rect 7097 13499 7163 13502
rect 1761 13424 4354 13426
rect 1761 13368 1766 13424
rect 1822 13368 4354 13424
rect 1761 13366 4354 13368
rect 1761 13363 1827 13366
rect 4470 13364 4476 13428
rect 4540 13426 4546 13428
rect 8293 13426 8359 13429
rect 4540 13424 8359 13426
rect 4540 13368 8298 13424
rect 8354 13368 8359 13424
rect 4540 13366 8359 13368
rect 8526 13426 8586 13638
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 19139 13567 19455 13568
rect 9949 13562 10015 13565
rect 13077 13562 13143 13565
rect 9949 13560 13143 13562
rect 9949 13504 9954 13560
rect 10010 13504 13082 13560
rect 13138 13504 13143 13560
rect 9949 13502 13143 13504
rect 9949 13499 10015 13502
rect 13077 13499 13143 13502
rect 21265 13562 21331 13565
rect 22200 13562 23000 13592
rect 21265 13560 23000 13562
rect 21265 13504 21270 13560
rect 21326 13504 23000 13560
rect 21265 13502 23000 13504
rect 21265 13499 21331 13502
rect 22200 13472 23000 13502
rect 8526 13366 12450 13426
rect 4540 13364 4546 13366
rect 8293 13363 8359 13366
rect 4429 13290 4495 13293
rect 12390 13290 12450 13366
rect 18413 13290 18479 13293
rect 4429 13288 11898 13290
rect 4429 13232 4434 13288
rect 4490 13232 11898 13288
rect 4429 13230 11898 13232
rect 12390 13288 18479 13290
rect 12390 13232 18418 13288
rect 18474 13232 18479 13288
rect 12390 13230 18479 13232
rect 4429 13227 4495 13230
rect 0 13154 800 13184
rect 2865 13154 2931 13157
rect 0 13152 2931 13154
rect 0 13096 2870 13152
rect 2926 13096 2931 13152
rect 0 13094 2931 13096
rect 11838 13154 11898 13230
rect 18413 13227 18479 13230
rect 20529 13290 20595 13293
rect 20529 13288 22202 13290
rect 20529 13232 20534 13288
rect 20590 13232 22202 13288
rect 20529 13230 22202 13232
rect 20529 13227 20595 13230
rect 22142 13184 22202 13230
rect 12341 13154 12407 13157
rect 11838 13152 12407 13154
rect 11838 13096 12346 13152
rect 12402 13096 12407 13152
rect 11838 13094 12407 13096
rect 22142 13094 23000 13184
rect 0 13064 800 13094
rect 2865 13091 2931 13094
rect 12341 13091 12407 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22200 13064 23000 13094
rect 21738 13023 22054 13024
rect 3366 12820 3372 12884
rect 3436 12882 3442 12884
rect 4153 12882 4219 12885
rect 3436 12880 4219 12882
rect 3436 12824 4158 12880
rect 4214 12824 4219 12880
rect 3436 12822 4219 12824
rect 3436 12820 3442 12822
rect 4153 12819 4219 12822
rect 8293 12882 8359 12885
rect 11789 12884 11855 12885
rect 8293 12880 10426 12882
rect 8293 12824 8298 12880
rect 8354 12824 10426 12880
rect 8293 12822 10426 12824
rect 8293 12819 8359 12822
rect 0 12746 800 12776
rect 3141 12746 3207 12749
rect 0 12744 3207 12746
rect 0 12688 3146 12744
rect 3202 12688 3207 12744
rect 0 12686 3207 12688
rect 0 12656 800 12686
rect 3141 12683 3207 12686
rect 5901 12746 5967 12749
rect 10174 12746 10180 12748
rect 5901 12744 10180 12746
rect 5901 12688 5906 12744
rect 5962 12688 10180 12744
rect 5901 12686 10180 12688
rect 5901 12683 5967 12686
rect 10174 12684 10180 12686
rect 10244 12684 10250 12748
rect 10366 12746 10426 12822
rect 11789 12880 11836 12884
rect 11900 12882 11906 12884
rect 11789 12824 11794 12880
rect 11789 12820 11836 12824
rect 11900 12822 11946 12882
rect 11900 12820 11906 12822
rect 11789 12819 11855 12820
rect 17125 12746 17191 12749
rect 10366 12744 17191 12746
rect 10366 12688 17130 12744
rect 17186 12688 17191 12744
rect 10366 12686 17191 12688
rect 17125 12683 17191 12686
rect 19793 12746 19859 12749
rect 22200 12746 23000 12776
rect 19793 12744 23000 12746
rect 19793 12688 19798 12744
rect 19854 12688 23000 12744
rect 19793 12686 23000 12688
rect 19793 12683 19859 12686
rect 22200 12656 23000 12686
rect 5942 12548 5948 12612
rect 6012 12610 6018 12612
rect 8293 12610 8359 12613
rect 6012 12608 8359 12610
rect 6012 12552 8298 12608
rect 8354 12552 8359 12608
rect 6012 12550 8359 12552
rect 6012 12548 6018 12550
rect 8293 12547 8359 12550
rect 9765 12610 9831 12613
rect 11513 12610 11579 12613
rect 9765 12608 11579 12610
rect 9765 12552 9770 12608
rect 9826 12552 11518 12608
rect 11574 12552 11579 12608
rect 9765 12550 11579 12552
rect 9765 12547 9831 12550
rect 11513 12547 11579 12550
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 19139 12479 19455 12480
rect 2957 12472 3023 12477
rect 2957 12416 2962 12472
rect 3018 12416 3023 12472
rect 2957 12411 3023 12416
rect 5390 12412 5396 12476
rect 5460 12474 5466 12476
rect 5625 12474 5691 12477
rect 5460 12472 5691 12474
rect 5460 12416 5630 12472
rect 5686 12416 5691 12472
rect 5460 12414 5691 12416
rect 5460 12412 5466 12414
rect 5625 12411 5691 12414
rect 6637 12474 6703 12477
rect 12985 12476 13051 12477
rect 8150 12474 8156 12476
rect 6637 12472 8156 12474
rect 6637 12416 6642 12472
rect 6698 12416 8156 12472
rect 6637 12414 8156 12416
rect 6637 12411 6703 12414
rect 8150 12412 8156 12414
rect 8220 12412 8226 12476
rect 12934 12474 12940 12476
rect 12894 12414 12940 12474
rect 13004 12472 13051 12476
rect 13046 12416 13051 12472
rect 12934 12412 12940 12414
rect 13004 12412 13051 12416
rect 12985 12411 13051 12412
rect 0 12338 800 12368
rect 2221 12338 2287 12341
rect 0 12336 2287 12338
rect 0 12280 2226 12336
rect 2282 12280 2287 12336
rect 0 12278 2287 12280
rect 2960 12338 3020 12411
rect 3877 12338 3943 12341
rect 2960 12336 3943 12338
rect 2960 12280 3882 12336
rect 3938 12280 3943 12336
rect 2960 12278 3943 12280
rect 0 12248 800 12278
rect 2221 12275 2287 12278
rect 3877 12275 3943 12278
rect 5390 12276 5396 12340
rect 5460 12338 5466 12340
rect 5533 12338 5599 12341
rect 5460 12336 5599 12338
rect 5460 12280 5538 12336
rect 5594 12280 5599 12336
rect 5460 12278 5599 12280
rect 5460 12276 5466 12278
rect 5533 12275 5599 12278
rect 6678 12276 6684 12340
rect 6748 12338 6754 12340
rect 7373 12338 7439 12341
rect 6748 12336 7439 12338
rect 6748 12280 7378 12336
rect 7434 12280 7439 12336
rect 6748 12278 7439 12280
rect 6748 12276 6754 12278
rect 7373 12275 7439 12278
rect 8150 12276 8156 12340
rect 8220 12338 8226 12340
rect 9254 12338 9260 12340
rect 8220 12278 9260 12338
rect 8220 12276 8226 12278
rect 9254 12276 9260 12278
rect 9324 12276 9330 12340
rect 20529 12338 20595 12341
rect 22200 12338 23000 12368
rect 20529 12336 23000 12338
rect 20529 12280 20534 12336
rect 20590 12280 23000 12336
rect 20529 12278 23000 12280
rect 20529 12275 20595 12278
rect 22200 12248 23000 12278
rect 1853 12202 1919 12205
rect 10593 12202 10659 12205
rect 1853 12200 10659 12202
rect 1853 12144 1858 12200
rect 1914 12144 10598 12200
rect 10654 12144 10659 12200
rect 1853 12142 10659 12144
rect 1853 12139 1919 12142
rect 10593 12139 10659 12142
rect 10777 12202 10843 12205
rect 17033 12202 17099 12205
rect 10777 12200 17099 12202
rect 10777 12144 10782 12200
rect 10838 12144 17038 12200
rect 17094 12144 17099 12200
rect 10777 12142 17099 12144
rect 10777 12139 10843 12142
rect 17033 12139 17099 12142
rect 6913 12066 6979 12069
rect 11145 12066 11211 12069
rect 6913 12064 11211 12066
rect 6913 12008 6918 12064
rect 6974 12008 11150 12064
rect 11206 12008 11211 12064
rect 6913 12006 11211 12008
rect 6913 12003 6979 12006
rect 11145 12003 11211 12006
rect 18597 12068 18663 12069
rect 18597 12064 18644 12068
rect 18708 12066 18714 12068
rect 18597 12008 18602 12064
rect 18597 12004 18644 12008
rect 18708 12006 18754 12066
rect 18708 12004 18714 12006
rect 18597 12003 18663 12004
rect 6144 12000 6460 12001
rect 0 11930 800 11960
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 21738 11935 22054 11936
rect 2221 11930 2287 11933
rect 0 11928 2287 11930
rect 0 11872 2226 11928
rect 2282 11872 2287 11928
rect 0 11870 2287 11872
rect 0 11840 800 11870
rect 2221 11867 2287 11870
rect 6545 11930 6611 11933
rect 10409 11930 10475 11933
rect 22200 11930 23000 11960
rect 6545 11928 10475 11930
rect 6545 11872 6550 11928
rect 6606 11872 10414 11928
rect 10470 11872 10475 11928
rect 6545 11870 10475 11872
rect 6545 11867 6611 11870
rect 10409 11867 10475 11870
rect 22142 11840 23000 11930
rect 1945 11794 2011 11797
rect 12525 11794 12591 11797
rect 1945 11792 12591 11794
rect 1945 11736 1950 11792
rect 2006 11736 12530 11792
rect 12586 11736 12591 11792
rect 1945 11734 12591 11736
rect 1945 11731 2011 11734
rect 12525 11731 12591 11734
rect 20529 11794 20595 11797
rect 22142 11794 22202 11840
rect 20529 11792 22202 11794
rect 20529 11736 20534 11792
rect 20590 11736 22202 11792
rect 20529 11734 22202 11736
rect 20529 11731 20595 11734
rect 1485 11658 1551 11661
rect 4429 11658 4495 11661
rect 10409 11658 10475 11661
rect 1485 11656 4354 11658
rect 1485 11600 1490 11656
rect 1546 11600 4354 11656
rect 1485 11598 4354 11600
rect 1485 11595 1551 11598
rect 0 11522 800 11552
rect 2221 11522 2287 11525
rect 0 11520 2287 11522
rect 0 11464 2226 11520
rect 2282 11464 2287 11520
rect 0 11462 2287 11464
rect 4294 11522 4354 11598
rect 4429 11656 10475 11658
rect 4429 11600 4434 11656
rect 4490 11600 10414 11656
rect 10470 11600 10475 11656
rect 4429 11598 10475 11600
rect 4429 11595 4495 11598
rect 10409 11595 10475 11598
rect 10593 11658 10659 11661
rect 14549 11658 14615 11661
rect 10593 11656 14615 11658
rect 10593 11600 10598 11656
rect 10654 11600 14554 11656
rect 14610 11600 14615 11656
rect 10593 11598 14615 11600
rect 10593 11595 10659 11598
rect 14549 11595 14615 11598
rect 6545 11522 6611 11525
rect 4294 11520 6611 11522
rect 4294 11464 6550 11520
rect 6606 11464 6611 11520
rect 4294 11462 6611 11464
rect 0 11432 800 11462
rect 2221 11459 2287 11462
rect 6545 11459 6611 11462
rect 21265 11522 21331 11525
rect 22200 11522 23000 11552
rect 21265 11520 23000 11522
rect 21265 11464 21270 11520
rect 21326 11464 23000 11520
rect 21265 11462 23000 11464
rect 21265 11459 21331 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22200 11432 23000 11462
rect 19139 11391 19455 11392
rect 5625 11386 5691 11389
rect 6678 11386 6684 11388
rect 5625 11384 6684 11386
rect 5625 11328 5630 11384
rect 5686 11328 6684 11384
rect 5625 11326 6684 11328
rect 5625 11323 5691 11326
rect 6678 11324 6684 11326
rect 6748 11324 6754 11388
rect 0 11114 800 11144
rect 3785 11114 3851 11117
rect 0 11112 3851 11114
rect 0 11056 3790 11112
rect 3846 11056 3851 11112
rect 0 11054 3851 11056
rect 0 11024 800 11054
rect 3785 11051 3851 11054
rect 4286 11052 4292 11116
rect 4356 11114 4362 11116
rect 4838 11114 4844 11116
rect 4356 11054 4844 11114
rect 4356 11052 4362 11054
rect 4838 11052 4844 11054
rect 4908 11114 4914 11116
rect 4981 11114 5047 11117
rect 4908 11112 5047 11114
rect 4908 11056 4986 11112
rect 5042 11056 5047 11112
rect 4908 11054 5047 11056
rect 4908 11052 4914 11054
rect 4981 11051 5047 11054
rect 18781 11114 18847 11117
rect 22200 11114 23000 11144
rect 18781 11112 23000 11114
rect 18781 11056 18786 11112
rect 18842 11056 23000 11112
rect 18781 11054 23000 11056
rect 18781 11051 18847 11054
rect 22200 11024 23000 11054
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 21738 10847 22054 10848
rect 8201 10842 8267 10845
rect 9438 10842 9444 10844
rect 8201 10840 9444 10842
rect 8201 10784 8206 10840
rect 8262 10784 9444 10840
rect 8201 10782 9444 10784
rect 8201 10779 8267 10782
rect 9438 10780 9444 10782
rect 9508 10780 9514 10844
rect 0 10706 800 10736
rect 2957 10706 3023 10709
rect 0 10704 3023 10706
rect 0 10648 2962 10704
rect 3018 10648 3023 10704
rect 0 10646 3023 10648
rect 0 10616 800 10646
rect 2957 10643 3023 10646
rect 8017 10706 8083 10709
rect 8201 10706 8267 10709
rect 8017 10704 8267 10706
rect 8017 10648 8022 10704
rect 8078 10648 8206 10704
rect 8262 10648 8267 10704
rect 8017 10646 8267 10648
rect 8017 10643 8083 10646
rect 8201 10643 8267 10646
rect 8661 10706 8727 10709
rect 16982 10706 16988 10708
rect 8661 10704 16988 10706
rect 8661 10648 8666 10704
rect 8722 10648 16988 10704
rect 8661 10646 16988 10648
rect 8661 10643 8727 10646
rect 16982 10644 16988 10646
rect 17052 10644 17058 10708
rect 20161 10706 20227 10709
rect 22200 10706 23000 10736
rect 20161 10704 23000 10706
rect 20161 10648 20166 10704
rect 20222 10648 23000 10704
rect 20161 10646 23000 10648
rect 20161 10643 20227 10646
rect 22200 10616 23000 10646
rect 2221 10570 2287 10573
rect 8017 10570 8083 10573
rect 2221 10568 8083 10570
rect 2221 10512 2226 10568
rect 2282 10512 8022 10568
rect 8078 10512 8083 10568
rect 2221 10510 8083 10512
rect 2221 10507 2287 10510
rect 8017 10507 8083 10510
rect 8150 10508 8156 10572
rect 8220 10570 8226 10572
rect 9489 10570 9555 10573
rect 8220 10568 9555 10570
rect 8220 10512 9494 10568
rect 9550 10512 9555 10568
rect 8220 10510 9555 10512
rect 8220 10508 8226 10510
rect 9489 10507 9555 10510
rect 3545 10368 3861 10369
rect 0 10298 800 10328
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 19139 10303 19455 10304
rect 2773 10298 2839 10301
rect 0 10296 2839 10298
rect 0 10240 2778 10296
rect 2834 10240 2839 10296
rect 0 10238 2839 10240
rect 0 10208 800 10238
rect 2773 10235 2839 10238
rect 15326 10236 15332 10300
rect 15396 10298 15402 10300
rect 15653 10298 15719 10301
rect 15396 10296 15719 10298
rect 15396 10240 15658 10296
rect 15714 10240 15719 10296
rect 15396 10238 15719 10240
rect 15396 10236 15402 10238
rect 15653 10235 15719 10238
rect 20161 10298 20227 10301
rect 22200 10298 23000 10328
rect 20161 10296 23000 10298
rect 20161 10240 20166 10296
rect 20222 10240 23000 10296
rect 20161 10238 23000 10240
rect 20161 10235 20227 10238
rect 22200 10208 23000 10238
rect 2773 10162 2839 10165
rect 3233 10162 3299 10165
rect 2773 10160 3299 10162
rect 2773 10104 2778 10160
rect 2834 10104 3238 10160
rect 3294 10104 3299 10160
rect 2773 10102 3299 10104
rect 2773 10099 2839 10102
rect 3233 10099 3299 10102
rect 5809 10162 5875 10165
rect 20897 10162 20963 10165
rect 5809 10160 20963 10162
rect 5809 10104 5814 10160
rect 5870 10104 20902 10160
rect 20958 10104 20963 10160
rect 5809 10102 20963 10104
rect 5809 10099 5875 10102
rect 20897 10099 20963 10102
rect 6913 10026 6979 10029
rect 7046 10026 7052 10028
rect 6913 10024 7052 10026
rect 6913 9968 6918 10024
rect 6974 9968 7052 10024
rect 6913 9966 7052 9968
rect 6913 9963 6979 9966
rect 7046 9964 7052 9966
rect 7116 9964 7122 10028
rect 20529 10026 20595 10029
rect 20529 10024 22202 10026
rect 20529 9968 20534 10024
rect 20590 9968 22202 10024
rect 20529 9966 22202 9968
rect 20529 9963 20595 9966
rect 22142 9920 22202 9966
rect 0 9890 800 9920
rect 2221 9890 2287 9893
rect 0 9888 2287 9890
rect 0 9832 2226 9888
rect 2282 9832 2287 9888
rect 0 9830 2287 9832
rect 22142 9830 23000 9920
rect 0 9800 800 9830
rect 2221 9827 2287 9830
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22200 9800 23000 9830
rect 21738 9759 22054 9760
rect 1945 9618 2011 9621
rect 2078 9618 2084 9620
rect 1945 9616 2084 9618
rect 1945 9560 1950 9616
rect 2006 9560 2084 9616
rect 1945 9558 2084 9560
rect 1945 9555 2011 9558
rect 2078 9556 2084 9558
rect 2148 9556 2154 9620
rect 2221 9618 2287 9621
rect 2630 9618 2636 9620
rect 2221 9616 2636 9618
rect 2221 9560 2226 9616
rect 2282 9560 2636 9616
rect 2221 9558 2636 9560
rect 2221 9555 2287 9558
rect 2630 9556 2636 9558
rect 2700 9556 2706 9620
rect 3601 9618 3667 9621
rect 5758 9618 5764 9620
rect 3601 9616 5764 9618
rect 3601 9560 3606 9616
rect 3662 9560 5764 9616
rect 3601 9558 5764 9560
rect 3601 9555 3667 9558
rect 5758 9556 5764 9558
rect 5828 9556 5834 9620
rect 11973 9618 12039 9621
rect 20437 9618 20503 9621
rect 11973 9616 20503 9618
rect 11973 9560 11978 9616
rect 12034 9560 20442 9616
rect 20498 9560 20503 9616
rect 11973 9558 20503 9560
rect 11973 9555 12039 9558
rect 20437 9555 20503 9558
rect 0 9482 800 9512
rect 2221 9482 2287 9485
rect 0 9480 2287 9482
rect 0 9424 2226 9480
rect 2282 9424 2287 9480
rect 0 9422 2287 9424
rect 0 9392 800 9422
rect 2221 9419 2287 9422
rect 3877 9482 3943 9485
rect 6821 9482 6887 9485
rect 3877 9480 6887 9482
rect 3877 9424 3882 9480
rect 3938 9424 6826 9480
rect 6882 9424 6887 9480
rect 3877 9422 6887 9424
rect 3877 9419 3943 9422
rect 6821 9419 6887 9422
rect 11697 9482 11763 9485
rect 14273 9482 14339 9485
rect 11697 9480 14339 9482
rect 11697 9424 11702 9480
rect 11758 9424 14278 9480
rect 14334 9424 14339 9480
rect 11697 9422 14339 9424
rect 11697 9419 11763 9422
rect 14273 9419 14339 9422
rect 18413 9482 18479 9485
rect 19701 9482 19767 9485
rect 22200 9482 23000 9512
rect 18413 9480 23000 9482
rect 18413 9424 18418 9480
rect 18474 9424 19706 9480
rect 19762 9424 23000 9480
rect 18413 9422 23000 9424
rect 18413 9419 18479 9422
rect 19701 9419 19767 9422
rect 22200 9392 23000 9422
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 19139 9215 19455 9216
rect 0 9074 800 9104
rect 3141 9074 3207 9077
rect 0 9072 3207 9074
rect 0 9016 3146 9072
rect 3202 9016 3207 9072
rect 0 9014 3207 9016
rect 0 8984 800 9014
rect 3141 9011 3207 9014
rect 4838 9012 4844 9076
rect 4908 9074 4914 9076
rect 11973 9074 12039 9077
rect 4908 9072 12039 9074
rect 4908 9016 11978 9072
rect 12034 9016 12039 9072
rect 4908 9014 12039 9016
rect 4908 9012 4914 9014
rect 11973 9011 12039 9014
rect 20529 9074 20595 9077
rect 22200 9074 23000 9104
rect 20529 9072 23000 9074
rect 20529 9016 20534 9072
rect 20590 9016 23000 9072
rect 20529 9014 23000 9016
rect 20529 9011 20595 9014
rect 22200 8984 23000 9014
rect 4797 8938 4863 8941
rect 7465 8938 7531 8941
rect 4797 8936 7531 8938
rect 4797 8880 4802 8936
rect 4858 8880 7470 8936
rect 7526 8880 7531 8936
rect 4797 8878 7531 8880
rect 4797 8875 4863 8878
rect 7465 8875 7531 8878
rect 10174 8876 10180 8940
rect 10244 8938 10250 8940
rect 10777 8938 10843 8941
rect 12341 8938 12407 8941
rect 10244 8936 12407 8938
rect 10244 8880 10782 8936
rect 10838 8880 12346 8936
rect 12402 8880 12407 8936
rect 10244 8878 12407 8880
rect 10244 8876 10250 8878
rect 10777 8875 10843 8878
rect 12341 8875 12407 8878
rect 15377 8938 15443 8941
rect 18413 8938 18479 8941
rect 15377 8936 18479 8938
rect 15377 8880 15382 8936
rect 15438 8880 18418 8936
rect 18474 8880 18479 8936
rect 15377 8878 18479 8880
rect 15377 8875 15443 8878
rect 18413 8875 18479 8878
rect 6144 8736 6460 8737
rect 0 8666 800 8696
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 21738 8671 22054 8672
rect 2129 8666 2195 8669
rect 0 8664 2195 8666
rect 0 8608 2134 8664
rect 2190 8608 2195 8664
rect 0 8606 2195 8608
rect 0 8576 800 8606
rect 2129 8603 2195 8606
rect 8109 8666 8175 8669
rect 8334 8666 8340 8668
rect 8109 8664 8340 8666
rect 8109 8608 8114 8664
rect 8170 8608 8340 8664
rect 8109 8606 8340 8608
rect 8109 8603 8175 8606
rect 8334 8604 8340 8606
rect 8404 8604 8410 8668
rect 22200 8666 23000 8696
rect 22142 8576 23000 8666
rect 21265 8530 21331 8533
rect 22142 8530 22202 8576
rect 21265 8528 22202 8530
rect 21265 8472 21270 8528
rect 21326 8472 22202 8528
rect 21265 8470 22202 8472
rect 21265 8467 21331 8470
rect 6862 8332 6868 8396
rect 6932 8394 6938 8396
rect 11789 8394 11855 8397
rect 6932 8392 11855 8394
rect 6932 8336 11794 8392
rect 11850 8336 11855 8392
rect 6932 8334 11855 8336
rect 6932 8332 6938 8334
rect 11789 8331 11855 8334
rect 0 8258 800 8288
rect 2221 8258 2287 8261
rect 0 8256 2287 8258
rect 0 8200 2226 8256
rect 2282 8200 2287 8256
rect 0 8198 2287 8200
rect 0 8168 800 8198
rect 2221 8195 2287 8198
rect 3969 8258 4035 8261
rect 8150 8258 8156 8260
rect 3969 8256 8156 8258
rect 3969 8200 3974 8256
rect 4030 8200 8156 8256
rect 3969 8198 8156 8200
rect 3969 8195 4035 8198
rect 8150 8196 8156 8198
rect 8220 8196 8226 8260
rect 22200 8258 23000 8288
rect 19566 8198 23000 8258
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 3049 7986 3115 7989
rect 4102 7986 4108 7988
rect 3049 7984 4108 7986
rect 3049 7928 3054 7984
rect 3110 7928 4108 7984
rect 3049 7926 4108 7928
rect 3049 7923 3115 7926
rect 4102 7924 4108 7926
rect 4172 7924 4178 7988
rect 5758 7924 5764 7988
rect 5828 7986 5834 7988
rect 5993 7986 6059 7989
rect 5828 7984 6059 7986
rect 5828 7928 5998 7984
rect 6054 7928 6059 7984
rect 5828 7926 6059 7928
rect 5828 7924 5834 7926
rect 5993 7923 6059 7926
rect 7741 7986 7807 7989
rect 9806 7986 9812 7988
rect 7741 7984 9812 7986
rect 7741 7928 7746 7984
rect 7802 7928 9812 7984
rect 7741 7926 9812 7928
rect 7741 7923 7807 7926
rect 9806 7924 9812 7926
rect 9876 7924 9882 7988
rect 18781 7986 18847 7989
rect 19566 7986 19626 8198
rect 22200 8168 23000 8198
rect 18781 7984 19626 7986
rect 18781 7928 18786 7984
rect 18842 7928 19626 7984
rect 18781 7926 19626 7928
rect 18781 7923 18847 7926
rect 0 7850 800 7880
rect 2773 7850 2839 7853
rect 9029 7850 9095 7853
rect 0 7848 9095 7850
rect 0 7792 2778 7848
rect 2834 7792 9034 7848
rect 9090 7792 9095 7848
rect 0 7790 9095 7792
rect 0 7760 800 7790
rect 2773 7787 2839 7790
rect 9029 7787 9095 7790
rect 17861 7850 17927 7853
rect 22200 7850 23000 7880
rect 17861 7848 23000 7850
rect 17861 7792 17866 7848
rect 17922 7792 23000 7848
rect 17861 7790 23000 7792
rect 17861 7787 17927 7790
rect 22200 7760 23000 7790
rect 1853 7714 1919 7717
rect 1853 7712 5458 7714
rect 1853 7656 1858 7712
rect 1914 7656 5458 7712
rect 1853 7654 5458 7656
rect 1853 7651 1919 7654
rect 1485 7578 1551 7581
rect 2630 7578 2636 7580
rect 1485 7576 2636 7578
rect 1485 7520 1490 7576
rect 1546 7520 2636 7576
rect 1485 7518 2636 7520
rect 1485 7515 1551 7518
rect 2630 7516 2636 7518
rect 2700 7516 2706 7580
rect 0 7442 800 7472
rect 1485 7442 1551 7445
rect 0 7440 1551 7442
rect 0 7384 1490 7440
rect 1546 7384 1551 7440
rect 0 7382 1551 7384
rect 5398 7442 5458 7654
rect 19006 7652 19012 7716
rect 19076 7714 19082 7716
rect 21081 7714 21147 7717
rect 19076 7712 21147 7714
rect 19076 7656 21086 7712
rect 21142 7656 21147 7712
rect 19076 7654 21147 7656
rect 19076 7652 19082 7654
rect 21081 7651 21147 7654
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 18638 7516 18644 7580
rect 18708 7578 18714 7580
rect 19793 7578 19859 7581
rect 20437 7578 20503 7581
rect 18708 7576 20503 7578
rect 18708 7520 19798 7576
rect 19854 7520 20442 7576
rect 20498 7520 20503 7576
rect 18708 7518 20503 7520
rect 18708 7516 18714 7518
rect 19793 7515 19859 7518
rect 20437 7515 20503 7518
rect 6678 7442 6684 7444
rect 5398 7382 6684 7442
rect 0 7352 800 7382
rect 1485 7379 1551 7382
rect 6678 7380 6684 7382
rect 6748 7380 6754 7444
rect 18137 7442 18203 7445
rect 19149 7442 19215 7445
rect 22200 7442 23000 7472
rect 18137 7440 19215 7442
rect 18137 7384 18142 7440
rect 18198 7384 19154 7440
rect 19210 7384 19215 7440
rect 18137 7382 19215 7384
rect 18137 7379 18203 7382
rect 19149 7379 19215 7382
rect 20118 7382 23000 7442
rect 20118 7309 20178 7382
rect 22200 7352 23000 7382
rect 12157 7306 12223 7309
rect 2730 7304 12223 7306
rect 2730 7248 12162 7304
rect 12218 7248 12223 7304
rect 2730 7246 12223 7248
rect 0 7034 800 7064
rect 1485 7034 1551 7037
rect 2730 7034 2790 7246
rect 12157 7243 12223 7246
rect 14365 7306 14431 7309
rect 20069 7306 20178 7309
rect 14365 7304 20178 7306
rect 14365 7248 14370 7304
rect 14426 7248 20074 7304
rect 20130 7248 20178 7304
rect 14365 7246 20178 7248
rect 14365 7243 14431 7246
rect 20069 7243 20135 7246
rect 14457 7170 14523 7173
rect 18781 7170 18847 7173
rect 14457 7168 18847 7170
rect 14457 7112 14462 7168
rect 14518 7112 18786 7168
rect 18842 7112 18847 7168
rect 14457 7110 18847 7112
rect 14457 7107 14523 7110
rect 18781 7107 18847 7110
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 3141 7036 3207 7037
rect 3141 7034 3188 7036
rect 0 7032 2790 7034
rect 0 6976 1490 7032
rect 1546 6976 2790 7032
rect 0 6974 2790 6976
rect 3096 7032 3188 7034
rect 3096 6976 3146 7032
rect 3096 6974 3188 6976
rect 0 6944 800 6974
rect 1485 6971 1551 6974
rect 3141 6972 3188 6974
rect 3252 6972 3258 7036
rect 20529 7034 20595 7037
rect 22200 7034 23000 7064
rect 20529 7032 23000 7034
rect 20529 6976 20534 7032
rect 20590 6976 23000 7032
rect 20529 6974 23000 6976
rect 3141 6971 3207 6972
rect 20529 6971 20595 6974
rect 22200 6944 23000 6974
rect 12198 6898 12204 6900
rect 2730 6838 12204 6898
rect 0 6626 800 6656
rect 1526 6626 1532 6628
rect 0 6566 1532 6626
rect 0 6536 800 6566
rect 1526 6564 1532 6566
rect 1596 6626 1602 6628
rect 2730 6626 2790 6838
rect 12198 6836 12204 6838
rect 12268 6836 12274 6900
rect 18045 6898 18111 6901
rect 19333 6898 19399 6901
rect 18045 6896 19399 6898
rect 18045 6840 18050 6896
rect 18106 6840 19338 6896
rect 19394 6840 19399 6896
rect 18045 6838 19399 6840
rect 18045 6835 18111 6838
rect 19333 6835 19399 6838
rect 19609 6898 19675 6901
rect 19793 6898 19859 6901
rect 19609 6896 19859 6898
rect 19609 6840 19614 6896
rect 19670 6840 19798 6896
rect 19854 6840 19859 6896
rect 19609 6838 19859 6840
rect 19609 6835 19675 6838
rect 19793 6835 19859 6838
rect 3233 6762 3299 6765
rect 1596 6566 2790 6626
rect 3006 6760 3299 6762
rect 3006 6704 3238 6760
rect 3294 6704 3299 6760
rect 3006 6702 3299 6704
rect 1596 6564 1602 6566
rect 3006 6357 3066 6702
rect 3233 6699 3299 6702
rect 4613 6762 4679 6765
rect 4838 6762 4844 6764
rect 4613 6760 4844 6762
rect 4613 6704 4618 6760
rect 4674 6704 4844 6760
rect 4613 6702 4844 6704
rect 4613 6699 4679 6702
rect 4838 6700 4844 6702
rect 4908 6700 4914 6764
rect 5942 6700 5948 6764
rect 6012 6762 6018 6764
rect 6177 6762 6243 6765
rect 6012 6760 6243 6762
rect 6012 6704 6182 6760
rect 6238 6704 6243 6760
rect 6012 6702 6243 6704
rect 6012 6700 6018 6702
rect 6177 6699 6243 6702
rect 18413 6762 18479 6765
rect 19241 6762 19307 6765
rect 18413 6760 22202 6762
rect 18413 6704 18418 6760
rect 18474 6704 19246 6760
rect 19302 6704 22202 6760
rect 18413 6702 22202 6704
rect 18413 6699 18479 6702
rect 19241 6699 19307 6702
rect 22142 6656 22202 6702
rect 5758 6564 5764 6628
rect 5828 6626 5834 6628
rect 5993 6626 6059 6629
rect 5828 6624 6059 6626
rect 5828 6568 5998 6624
rect 6054 6568 6059 6624
rect 5828 6566 6059 6568
rect 22142 6566 23000 6656
rect 5828 6564 5834 6566
rect 5993 6563 6059 6566
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22200 6536 23000 6566
rect 21738 6495 22054 6496
rect 7414 6428 7420 6492
rect 7484 6490 7490 6492
rect 8477 6490 8543 6493
rect 9438 6490 9444 6492
rect 7484 6488 9444 6490
rect 7484 6432 8482 6488
rect 8538 6432 9444 6488
rect 7484 6430 9444 6432
rect 7484 6428 7490 6430
rect 8477 6427 8543 6430
rect 9438 6428 9444 6430
rect 9508 6428 9514 6492
rect 11789 6490 11855 6493
rect 15377 6490 15443 6493
rect 11789 6488 15443 6490
rect 11789 6432 11794 6488
rect 11850 6432 15382 6488
rect 15438 6432 15443 6488
rect 11789 6430 15443 6432
rect 11789 6427 11855 6430
rect 15377 6427 15443 6430
rect 19517 6490 19583 6493
rect 20253 6490 20319 6493
rect 19517 6488 20319 6490
rect 19517 6432 19522 6488
rect 19578 6432 20258 6488
rect 20314 6432 20319 6488
rect 19517 6430 20319 6432
rect 19517 6427 19583 6430
rect 20253 6427 20319 6430
rect 2957 6352 3066 6357
rect 2957 6296 2962 6352
rect 3018 6296 3066 6352
rect 2957 6294 3066 6296
rect 4797 6354 4863 6357
rect 15469 6354 15535 6357
rect 4797 6352 15535 6354
rect 4797 6296 4802 6352
rect 4858 6296 15474 6352
rect 15530 6296 15535 6352
rect 4797 6294 15535 6296
rect 2957 6291 3023 6294
rect 4797 6291 4863 6294
rect 15469 6291 15535 6294
rect 16205 6354 16271 6357
rect 19057 6354 19123 6357
rect 16205 6352 19123 6354
rect 16205 6296 16210 6352
rect 16266 6296 19062 6352
rect 19118 6296 19123 6352
rect 16205 6294 19123 6296
rect 16205 6291 16271 6294
rect 19057 6291 19123 6294
rect 0 6218 800 6248
rect 3049 6218 3115 6221
rect 0 6216 3115 6218
rect 0 6160 3054 6216
rect 3110 6160 3115 6216
rect 0 6158 3115 6160
rect 0 6128 800 6158
rect 3049 6155 3115 6158
rect 3918 6156 3924 6220
rect 3988 6218 3994 6220
rect 4337 6218 4403 6221
rect 3988 6216 4403 6218
rect 3988 6160 4342 6216
rect 4398 6160 4403 6216
rect 3988 6158 4403 6160
rect 3988 6156 3994 6158
rect 4337 6155 4403 6158
rect 8109 6218 8175 6221
rect 11697 6218 11763 6221
rect 8109 6216 11763 6218
rect 8109 6160 8114 6216
rect 8170 6160 11702 6216
rect 11758 6160 11763 6216
rect 8109 6158 11763 6160
rect 8109 6155 8175 6158
rect 11697 6155 11763 6158
rect 13721 6218 13787 6221
rect 18873 6218 18939 6221
rect 22200 6218 23000 6248
rect 13721 6216 23000 6218
rect 13721 6160 13726 6216
rect 13782 6160 18878 6216
rect 18934 6160 23000 6216
rect 13721 6158 23000 6160
rect 13721 6155 13787 6158
rect 18873 6155 18939 6158
rect 22200 6128 23000 6158
rect 11789 6082 11855 6085
rect 12801 6082 12867 6085
rect 11789 6080 12867 6082
rect 11789 6024 11794 6080
rect 11850 6024 12806 6080
rect 12862 6024 12867 6080
rect 11789 6022 12867 6024
rect 11789 6019 11855 6022
rect 12801 6019 12867 6022
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 19139 5951 19455 5952
rect 5942 5884 5948 5948
rect 6012 5946 6018 5948
rect 6177 5946 6243 5949
rect 6012 5944 6243 5946
rect 6012 5888 6182 5944
rect 6238 5888 6243 5944
rect 6012 5886 6243 5888
rect 6012 5884 6018 5886
rect 6177 5883 6243 5886
rect 9121 5946 9187 5949
rect 9438 5946 9444 5948
rect 9121 5944 9444 5946
rect 9121 5888 9126 5944
rect 9182 5888 9444 5944
rect 9121 5886 9444 5888
rect 9121 5883 9187 5886
rect 9438 5884 9444 5886
rect 9508 5884 9514 5948
rect 0 5810 800 5840
rect 2998 5810 3004 5812
rect 0 5750 3004 5810
rect 0 5720 800 5750
rect 2998 5748 3004 5750
rect 3068 5810 3074 5812
rect 3417 5810 3483 5813
rect 4429 5812 4495 5813
rect 4429 5810 4476 5812
rect 3068 5808 3483 5810
rect 3068 5752 3422 5808
rect 3478 5752 3483 5808
rect 3068 5750 3483 5752
rect 4384 5808 4476 5810
rect 4384 5752 4434 5808
rect 4384 5750 4476 5752
rect 3068 5748 3074 5750
rect 3417 5747 3483 5750
rect 4429 5748 4476 5750
rect 4540 5748 4546 5812
rect 5533 5810 5599 5813
rect 5717 5810 5783 5813
rect 5533 5808 5783 5810
rect 5533 5752 5538 5808
rect 5594 5752 5722 5808
rect 5778 5752 5783 5808
rect 5533 5750 5783 5752
rect 4429 5747 4495 5748
rect 5533 5747 5599 5750
rect 5717 5747 5783 5750
rect 5993 5810 6059 5813
rect 10501 5810 10567 5813
rect 10961 5810 11027 5813
rect 5993 5808 11027 5810
rect 5993 5752 5998 5808
rect 6054 5752 10506 5808
rect 10562 5752 10966 5808
rect 11022 5752 11027 5808
rect 5993 5750 11027 5752
rect 5993 5747 6059 5750
rect 10501 5747 10567 5750
rect 10961 5747 11027 5750
rect 13261 5810 13327 5813
rect 16021 5810 16087 5813
rect 13261 5808 16087 5810
rect 13261 5752 13266 5808
rect 13322 5752 16026 5808
rect 16082 5752 16087 5808
rect 13261 5750 16087 5752
rect 13261 5747 13327 5750
rect 16021 5747 16087 5750
rect 18413 5810 18479 5813
rect 21265 5810 21331 5813
rect 22200 5810 23000 5840
rect 18413 5808 23000 5810
rect 18413 5752 18418 5808
rect 18474 5752 21270 5808
rect 21326 5752 23000 5808
rect 18413 5750 23000 5752
rect 18413 5747 18479 5750
rect 21265 5747 21331 5750
rect 22200 5720 23000 5750
rect 2313 5674 2379 5677
rect 3325 5674 3391 5677
rect 9121 5674 9187 5677
rect 12985 5674 13051 5677
rect 13353 5674 13419 5677
rect 18781 5674 18847 5677
rect 2313 5672 13232 5674
rect 2313 5616 2318 5672
rect 2374 5616 3330 5672
rect 3386 5616 9126 5672
rect 9182 5616 12990 5672
rect 13046 5616 13232 5672
rect 2313 5614 13232 5616
rect 2313 5611 2379 5614
rect 3325 5611 3391 5614
rect 9121 5611 9187 5614
rect 12985 5611 13051 5614
rect 1485 5540 1551 5541
rect 1485 5538 1532 5540
rect 1440 5536 1532 5538
rect 1440 5480 1490 5536
rect 1440 5478 1532 5480
rect 1485 5476 1532 5478
rect 1596 5476 1602 5540
rect 6678 5476 6684 5540
rect 6748 5538 6754 5540
rect 6913 5538 6979 5541
rect 6748 5536 6979 5538
rect 6748 5480 6918 5536
rect 6974 5480 6979 5536
rect 6748 5478 6979 5480
rect 6748 5476 6754 5478
rect 1485 5475 1551 5476
rect 6913 5475 6979 5478
rect 7966 5476 7972 5540
rect 8036 5538 8042 5540
rect 8109 5538 8175 5541
rect 8569 5540 8635 5541
rect 8518 5538 8524 5540
rect 8036 5536 8175 5538
rect 8036 5480 8114 5536
rect 8170 5480 8175 5536
rect 8036 5478 8175 5480
rect 8478 5478 8524 5538
rect 8588 5536 8635 5540
rect 8630 5480 8635 5536
rect 8036 5476 8042 5478
rect 8109 5475 8175 5478
rect 8518 5476 8524 5478
rect 8588 5476 8635 5480
rect 13172 5538 13232 5614
rect 13353 5672 18847 5674
rect 13353 5616 13358 5672
rect 13414 5616 18786 5672
rect 18842 5616 18847 5672
rect 13353 5614 18847 5616
rect 13353 5611 13419 5614
rect 18781 5611 18847 5614
rect 15285 5538 15351 5541
rect 16113 5538 16179 5541
rect 13172 5536 16179 5538
rect 13172 5480 15290 5536
rect 15346 5480 16118 5536
rect 16174 5480 16179 5536
rect 13172 5478 16179 5480
rect 8569 5475 8635 5476
rect 15285 5475 15351 5478
rect 16113 5475 16179 5478
rect 18597 5538 18663 5541
rect 18597 5536 21282 5538
rect 18597 5480 18602 5536
rect 18658 5480 21282 5536
rect 18597 5478 21282 5480
rect 18597 5475 18663 5478
rect 6144 5472 6460 5473
rect 0 5402 800 5432
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 3141 5402 3207 5405
rect 0 5400 3207 5402
rect 0 5344 3146 5400
rect 3202 5344 3207 5400
rect 0 5342 3207 5344
rect 0 5312 800 5342
rect 3141 5339 3207 5342
rect 6729 5402 6795 5405
rect 6862 5402 6868 5404
rect 6729 5400 6868 5402
rect 6729 5344 6734 5400
rect 6790 5344 6868 5400
rect 6729 5342 6868 5344
rect 6729 5339 6795 5342
rect 6862 5340 6868 5342
rect 6932 5340 6938 5404
rect 7097 5402 7163 5405
rect 8385 5402 8451 5405
rect 7097 5400 8451 5402
rect 7097 5344 7102 5400
rect 7158 5344 8390 5400
rect 8446 5344 8451 5400
rect 7097 5342 8451 5344
rect 7097 5339 7163 5342
rect 8385 5339 8451 5342
rect 20345 5402 20411 5405
rect 20478 5402 20484 5404
rect 20345 5400 20484 5402
rect 20345 5344 20350 5400
rect 20406 5344 20484 5400
rect 20345 5342 20484 5344
rect 20345 5339 20411 5342
rect 20478 5340 20484 5342
rect 20548 5340 20554 5404
rect 21081 5266 21147 5269
rect 2730 5264 21147 5266
rect 2730 5208 21086 5264
rect 21142 5208 21147 5264
rect 2730 5206 21147 5208
rect 21222 5266 21282 5478
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 22200 5402 23000 5432
rect 22142 5312 23000 5402
rect 22142 5266 22202 5312
rect 21222 5206 22202 5266
rect 2221 5130 2287 5133
rect 2446 5130 2452 5132
rect 2221 5128 2452 5130
rect 2221 5072 2226 5128
rect 2282 5072 2452 5128
rect 2221 5070 2452 5072
rect 2221 5067 2287 5070
rect 2446 5068 2452 5070
rect 2516 5130 2522 5132
rect 2730 5130 2790 5206
rect 21081 5203 21147 5206
rect 2516 5070 2790 5130
rect 3877 5130 3943 5133
rect 4654 5130 4660 5132
rect 3877 5128 4660 5130
rect 3877 5072 3882 5128
rect 3938 5072 4660 5128
rect 3877 5070 4660 5072
rect 2516 5068 2522 5070
rect 3877 5067 3943 5070
rect 4654 5068 4660 5070
rect 4724 5068 4730 5132
rect 7373 5130 7439 5133
rect 8753 5130 8819 5133
rect 7373 5128 8819 5130
rect 7373 5072 7378 5128
rect 7434 5072 8758 5128
rect 8814 5072 8819 5128
rect 7373 5070 8819 5072
rect 7373 5067 7439 5070
rect 8753 5067 8819 5070
rect 10685 5130 10751 5133
rect 14917 5130 14983 5133
rect 17953 5130 18019 5133
rect 18321 5130 18387 5133
rect 10685 5128 14842 5130
rect 10685 5072 10690 5128
rect 10746 5072 14842 5128
rect 10685 5070 14842 5072
rect 10685 5067 10751 5070
rect 0 4994 800 5024
rect 974 4994 980 4996
rect 0 4934 980 4994
rect 0 4904 800 4934
rect 974 4932 980 4934
rect 1044 4994 1050 4996
rect 1393 4994 1459 4997
rect 1044 4992 1459 4994
rect 1044 4936 1398 4992
rect 1454 4936 1459 4992
rect 1044 4934 1459 4936
rect 1044 4932 1050 4934
rect 1393 4931 1459 4934
rect 11329 4994 11395 4997
rect 12801 4994 12867 4997
rect 11329 4992 12867 4994
rect 11329 4936 11334 4992
rect 11390 4936 12806 4992
rect 12862 4936 12867 4992
rect 11329 4934 12867 4936
rect 14782 4994 14842 5070
rect 14917 5128 18387 5130
rect 14917 5072 14922 5128
rect 14978 5072 17958 5128
rect 18014 5072 18326 5128
rect 18382 5072 18387 5128
rect 14917 5070 18387 5072
rect 14917 5067 14983 5070
rect 17953 5067 18019 5070
rect 18321 5067 18387 5070
rect 18597 5130 18663 5133
rect 18597 5128 19626 5130
rect 18597 5072 18602 5128
rect 18658 5072 19626 5128
rect 18597 5070 19626 5072
rect 18597 5067 18663 5070
rect 15929 4994 15995 4997
rect 14782 4992 15995 4994
rect 14782 4936 15934 4992
rect 15990 4936 15995 4992
rect 14782 4934 15995 4936
rect 19566 4994 19626 5070
rect 22200 4994 23000 5024
rect 19566 4934 23000 4994
rect 11329 4931 11395 4934
rect 12801 4931 12867 4934
rect 15929 4931 15995 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22200 4904 23000 4934
rect 19139 4863 19455 4864
rect 3233 4858 3299 4861
rect 6637 4860 6703 4861
rect 3366 4858 3372 4860
rect 3233 4856 3372 4858
rect 3233 4800 3238 4856
rect 3294 4800 3372 4856
rect 3233 4798 3372 4800
rect 3233 4795 3299 4798
rect 3366 4796 3372 4798
rect 3436 4796 3442 4860
rect 6637 4856 6684 4860
rect 6748 4858 6754 4860
rect 14917 4858 14983 4861
rect 6637 4800 6642 4856
rect 6637 4796 6684 4800
rect 6748 4798 6794 4858
rect 14917 4856 19074 4858
rect 14917 4800 14922 4856
rect 14978 4800 19074 4856
rect 14917 4798 19074 4800
rect 6748 4796 6754 4798
rect 6637 4795 6703 4796
rect 14917 4795 14983 4798
rect 4521 4722 4587 4725
rect 10041 4722 10107 4725
rect 4521 4720 10107 4722
rect 4521 4664 4526 4720
rect 4582 4664 10046 4720
rect 10102 4664 10107 4720
rect 4521 4662 10107 4664
rect 4521 4659 4587 4662
rect 10041 4659 10107 4662
rect 13537 4722 13603 4725
rect 18873 4722 18939 4725
rect 13537 4720 18939 4722
rect 13537 4664 13542 4720
rect 13598 4664 18878 4720
rect 18934 4664 18939 4720
rect 13537 4662 18939 4664
rect 19014 4722 19074 4798
rect 20805 4722 20871 4725
rect 19014 4720 20871 4722
rect 19014 4664 20810 4720
rect 20866 4664 20871 4720
rect 19014 4662 20871 4664
rect 13537 4659 13603 4662
rect 18873 4659 18939 4662
rect 20805 4659 20871 4662
rect 0 4586 800 4616
rect 2221 4586 2287 4589
rect 0 4584 2287 4586
rect 0 4528 2226 4584
rect 2282 4528 2287 4584
rect 0 4526 2287 4528
rect 0 4496 800 4526
rect 2221 4523 2287 4526
rect 3693 4586 3759 4589
rect 9581 4586 9647 4589
rect 14641 4586 14707 4589
rect 3693 4584 9506 4586
rect 3693 4528 3698 4584
rect 3754 4528 9506 4584
rect 3693 4526 9506 4528
rect 3693 4523 3759 4526
rect 9446 4450 9506 4526
rect 9581 4584 14707 4586
rect 9581 4528 9586 4584
rect 9642 4528 14646 4584
rect 14702 4528 14707 4584
rect 9581 4526 14707 4528
rect 9581 4523 9647 4526
rect 14641 4523 14707 4526
rect 19701 4586 19767 4589
rect 22200 4586 23000 4616
rect 19701 4584 23000 4586
rect 19701 4528 19706 4584
rect 19762 4528 23000 4584
rect 19701 4526 23000 4528
rect 19701 4523 19767 4526
rect 22200 4496 23000 4526
rect 10777 4450 10843 4453
rect 9446 4448 10843 4450
rect 9446 4392 10782 4448
rect 10838 4392 10843 4448
rect 9446 4390 10843 4392
rect 10777 4387 10843 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 21738 4319 22054 4320
rect 3509 4314 3575 4317
rect 4337 4314 4403 4317
rect 4981 4314 5047 4317
rect 5574 4314 5580 4316
rect 3509 4312 4484 4314
rect 3509 4256 3514 4312
rect 3570 4256 4342 4312
rect 4398 4256 4484 4312
rect 3509 4254 4484 4256
rect 4981 4312 5580 4314
rect 4981 4256 4986 4312
rect 5042 4256 5580 4312
rect 4981 4254 5580 4256
rect 3509 4251 3575 4254
rect 4294 4251 4403 4254
rect 4981 4251 5047 4254
rect 5574 4252 5580 4254
rect 5644 4252 5650 4316
rect 0 4178 800 4208
rect 4061 4178 4127 4181
rect 0 4176 4127 4178
rect 0 4120 4066 4176
rect 4122 4120 4127 4176
rect 0 4118 4127 4120
rect 4294 4178 4354 4251
rect 8937 4178 9003 4181
rect 4294 4176 9003 4178
rect 4294 4120 8942 4176
rect 8998 4120 9003 4176
rect 4294 4118 9003 4120
rect 0 4088 800 4118
rect 4061 4115 4127 4118
rect 8937 4115 9003 4118
rect 9121 4178 9187 4181
rect 9622 4178 9628 4180
rect 9121 4176 9628 4178
rect 9121 4120 9126 4176
rect 9182 4120 9628 4176
rect 9121 4118 9628 4120
rect 9121 4115 9187 4118
rect 9622 4116 9628 4118
rect 9692 4116 9698 4180
rect 13905 4178 13971 4181
rect 17677 4178 17743 4181
rect 13905 4176 17743 4178
rect 13905 4120 13910 4176
rect 13966 4120 17682 4176
rect 17738 4120 17743 4176
rect 13905 4118 17743 4120
rect 13905 4115 13971 4118
rect 17677 4115 17743 4118
rect 17953 4178 18019 4181
rect 22200 4178 23000 4208
rect 17953 4176 23000 4178
rect 17953 4120 17958 4176
rect 18014 4120 23000 4176
rect 17953 4118 23000 4120
rect 17953 4115 18019 4118
rect 22200 4088 23000 4118
rect 1158 3980 1164 4044
rect 1228 4042 1234 4044
rect 5073 4042 5139 4045
rect 5206 4042 5212 4044
rect 1228 3982 4354 4042
rect 1228 3980 1234 3982
rect 4294 3906 4354 3982
rect 5073 4040 5212 4042
rect 5073 3984 5078 4040
rect 5134 3984 5212 4040
rect 5073 3982 5212 3984
rect 5073 3979 5139 3982
rect 5206 3980 5212 3982
rect 5276 3980 5282 4044
rect 7782 3980 7788 4044
rect 7852 4042 7858 4044
rect 8109 4042 8175 4045
rect 8937 4042 9003 4045
rect 7852 4040 8175 4042
rect 7852 3984 8114 4040
rect 8170 3984 8175 4040
rect 7852 3982 8175 3984
rect 7852 3980 7858 3982
rect 8109 3979 8175 3982
rect 8342 4040 9003 4042
rect 8342 3984 8942 4040
rect 8998 3984 9003 4040
rect 8342 3982 9003 3984
rect 5809 3906 5875 3909
rect 4294 3904 5875 3906
rect 4294 3848 5814 3904
rect 5870 3848 5875 3904
rect 4294 3846 5875 3848
rect 5809 3843 5875 3846
rect 6177 3906 6243 3909
rect 8342 3906 8402 3982
rect 8937 3979 9003 3982
rect 9305 4042 9371 4045
rect 14958 4042 14964 4044
rect 9305 4040 14964 4042
rect 9305 3984 9310 4040
rect 9366 3984 14964 4040
rect 9305 3982 14964 3984
rect 9305 3979 9371 3982
rect 14958 3980 14964 3982
rect 15028 3980 15034 4044
rect 15377 4042 15443 4045
rect 15510 4042 15516 4044
rect 15377 4040 15516 4042
rect 15377 3984 15382 4040
rect 15438 3984 15516 4040
rect 15377 3982 15516 3984
rect 15377 3979 15443 3982
rect 15510 3980 15516 3982
rect 15580 3980 15586 4044
rect 16941 4042 17007 4045
rect 16941 4040 19626 4042
rect 16941 3984 16946 4040
rect 17002 3984 19626 4040
rect 16941 3982 19626 3984
rect 16941 3979 17007 3982
rect 6177 3904 8402 3906
rect 6177 3848 6182 3904
rect 6238 3848 8402 3904
rect 6177 3846 8402 3848
rect 6177 3843 6243 3846
rect 11094 3844 11100 3908
rect 11164 3906 11170 3908
rect 11830 3906 11836 3908
rect 11164 3846 11836 3906
rect 11164 3844 11170 3846
rect 11830 3844 11836 3846
rect 11900 3844 11906 3908
rect 16113 3906 16179 3909
rect 18873 3906 18939 3909
rect 16113 3904 18939 3906
rect 16113 3848 16118 3904
rect 16174 3848 18878 3904
rect 18934 3848 18939 3904
rect 16113 3846 18939 3848
rect 16113 3843 16179 3846
rect 18873 3843 18939 3846
rect 3545 3840 3861 3841
rect 0 3770 800 3800
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 6862 3770 6868 3772
rect 0 3710 2790 3770
rect 0 3680 800 3710
rect 2730 3634 2790 3710
rect 3926 3710 6868 3770
rect 3926 3634 3986 3710
rect 6862 3708 6868 3710
rect 6932 3708 6938 3772
rect 9438 3708 9444 3772
rect 9508 3770 9514 3772
rect 13353 3770 13419 3773
rect 9508 3768 13419 3770
rect 9508 3712 13358 3768
rect 13414 3712 13419 3768
rect 9508 3710 13419 3712
rect 9508 3708 9514 3710
rect 13353 3707 13419 3710
rect 14365 3770 14431 3773
rect 14590 3770 14596 3772
rect 14365 3768 14596 3770
rect 14365 3712 14370 3768
rect 14426 3712 14596 3768
rect 14365 3710 14596 3712
rect 14365 3707 14431 3710
rect 14590 3708 14596 3710
rect 14660 3708 14666 3772
rect 19566 3770 19626 3982
rect 22200 3770 23000 3800
rect 19566 3710 23000 3770
rect 22200 3680 23000 3710
rect 2730 3574 3986 3634
rect 5809 3634 5875 3637
rect 8569 3634 8635 3637
rect 12341 3634 12407 3637
rect 5809 3632 8635 3634
rect 5809 3576 5814 3632
rect 5870 3576 8574 3632
rect 8630 3576 8635 3632
rect 5809 3574 8635 3576
rect 5809 3571 5875 3574
rect 8569 3571 8635 3574
rect 8710 3632 12407 3634
rect 8710 3576 12346 3632
rect 12402 3576 12407 3632
rect 8710 3574 12407 3576
rect 3233 3498 3299 3501
rect 3693 3498 3759 3501
rect 8201 3498 8267 3501
rect 8710 3498 8770 3574
rect 12341 3571 12407 3574
rect 16205 3634 16271 3637
rect 16205 3632 20914 3634
rect 16205 3576 16210 3632
rect 16266 3576 20914 3632
rect 16205 3574 20914 3576
rect 16205 3571 16271 3574
rect 3233 3496 6700 3498
rect 3233 3440 3238 3496
rect 3294 3440 3698 3496
rect 3754 3440 6700 3496
rect 3233 3438 6700 3440
rect 3233 3435 3299 3438
rect 3693 3435 3759 3438
rect 0 3362 800 3392
rect 2865 3362 2931 3365
rect 0 3360 2931 3362
rect 0 3304 2870 3360
rect 2926 3304 2931 3360
rect 0 3302 2931 3304
rect 6640 3362 6700 3438
rect 8201 3496 8770 3498
rect 8201 3440 8206 3496
rect 8262 3440 8770 3496
rect 8201 3438 8770 3440
rect 8937 3498 9003 3501
rect 9254 3498 9260 3500
rect 8937 3496 9260 3498
rect 8937 3440 8942 3496
rect 8998 3440 9260 3496
rect 8937 3438 9260 3440
rect 8201 3435 8267 3438
rect 8937 3435 9003 3438
rect 9254 3436 9260 3438
rect 9324 3436 9330 3500
rect 9397 3498 9463 3501
rect 20713 3498 20779 3501
rect 9397 3496 20779 3498
rect 9397 3440 9402 3496
rect 9458 3440 20718 3496
rect 20774 3440 20779 3496
rect 9397 3438 20779 3440
rect 20854 3498 20914 3574
rect 20854 3438 22202 3498
rect 9397 3435 9463 3438
rect 20713 3435 20779 3438
rect 22142 3392 22202 3438
rect 11094 3362 11100 3364
rect 6640 3302 11100 3362
rect 0 3272 800 3302
rect 2865 3299 2931 3302
rect 11094 3300 11100 3302
rect 11164 3300 11170 3364
rect 22142 3302 23000 3392
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22200 3272 23000 3302
rect 21738 3231 22054 3232
rect 6729 3226 6795 3229
rect 8661 3226 8727 3229
rect 6729 3224 8727 3226
rect 6729 3168 6734 3224
rect 6790 3168 8666 3224
rect 8722 3168 8727 3224
rect 6729 3166 8727 3168
rect 6729 3163 6795 3166
rect 8661 3163 8727 3166
rect 13905 3226 13971 3229
rect 14406 3226 14412 3228
rect 13905 3224 14412 3226
rect 13905 3168 13910 3224
rect 13966 3168 14412 3224
rect 13905 3166 14412 3168
rect 13905 3163 13971 3166
rect 14406 3164 14412 3166
rect 14476 3164 14482 3228
rect 19006 3164 19012 3228
rect 19076 3226 19082 3228
rect 20437 3226 20503 3229
rect 19076 3224 20503 3226
rect 19076 3168 20442 3224
rect 20498 3168 20503 3224
rect 19076 3166 20503 3168
rect 19076 3164 19082 3166
rect 20437 3163 20503 3166
rect 4153 3090 4219 3093
rect 7414 3090 7420 3092
rect 4153 3088 7420 3090
rect 4153 3032 4158 3088
rect 4214 3032 7420 3088
rect 4153 3030 7420 3032
rect 4153 3027 4219 3030
rect 7414 3028 7420 3030
rect 7484 3028 7490 3092
rect 7649 3090 7715 3093
rect 14089 3090 14155 3093
rect 7649 3088 14155 3090
rect 7649 3032 7654 3088
rect 7710 3032 14094 3088
rect 14150 3032 14155 3088
rect 7649 3030 14155 3032
rect 7649 3027 7715 3030
rect 14089 3027 14155 3030
rect 14825 3090 14891 3093
rect 18137 3090 18203 3093
rect 19333 3090 19399 3093
rect 20161 3092 20227 3093
rect 14825 3088 18203 3090
rect 14825 3032 14830 3088
rect 14886 3032 18142 3088
rect 18198 3032 18203 3088
rect 14825 3030 18203 3032
rect 14825 3027 14891 3030
rect 18137 3027 18203 3030
rect 18278 3088 19399 3090
rect 18278 3032 19338 3088
rect 19394 3032 19399 3088
rect 18278 3030 19399 3032
rect 0 2954 800 2984
rect 933 2954 999 2957
rect 0 2952 999 2954
rect 0 2896 938 2952
rect 994 2896 999 2952
rect 0 2894 999 2896
rect 0 2864 800 2894
rect 933 2891 999 2894
rect 2589 2954 2655 2957
rect 5165 2954 5231 2957
rect 2589 2952 5231 2954
rect 2589 2896 2594 2952
rect 2650 2896 5170 2952
rect 5226 2896 5231 2952
rect 2589 2894 5231 2896
rect 2589 2891 2655 2894
rect 5165 2891 5231 2894
rect 6361 2954 6427 2957
rect 6678 2954 6684 2956
rect 6361 2952 6684 2954
rect 6361 2896 6366 2952
rect 6422 2896 6684 2952
rect 6361 2894 6684 2896
rect 6361 2891 6427 2894
rect 6678 2892 6684 2894
rect 6748 2892 6754 2956
rect 8201 2954 8267 2957
rect 9673 2954 9739 2957
rect 8201 2952 9739 2954
rect 8201 2896 8206 2952
rect 8262 2896 9678 2952
rect 9734 2896 9739 2952
rect 8201 2894 9739 2896
rect 8201 2891 8267 2894
rect 9673 2891 9739 2894
rect 13353 2954 13419 2957
rect 13721 2954 13787 2957
rect 18278 2954 18338 3030
rect 19333 3027 19399 3030
rect 20110 3028 20116 3092
rect 20180 3090 20227 3092
rect 20180 3088 20272 3090
rect 20222 3032 20272 3088
rect 20180 3030 20272 3032
rect 20180 3028 20227 3030
rect 20161 3027 20227 3028
rect 13353 2952 18338 2954
rect 13353 2896 13358 2952
rect 13414 2896 13726 2952
rect 13782 2896 18338 2952
rect 13353 2894 18338 2896
rect 19149 2954 19215 2957
rect 22200 2954 23000 2984
rect 19149 2952 23000 2954
rect 19149 2896 19154 2952
rect 19210 2896 23000 2952
rect 19149 2894 23000 2896
rect 13353 2891 13419 2894
rect 13721 2891 13787 2894
rect 19149 2891 19215 2894
rect 22200 2864 23000 2894
rect 2630 2756 2636 2820
rect 2700 2818 2706 2820
rect 2773 2818 2839 2821
rect 5625 2818 5691 2821
rect 2700 2816 2839 2818
rect 2700 2760 2778 2816
rect 2834 2760 2839 2816
rect 2700 2758 2839 2760
rect 2700 2756 2706 2758
rect 2773 2755 2839 2758
rect 4110 2816 5691 2818
rect 4110 2760 5630 2816
rect 5686 2760 5691 2816
rect 4110 2758 5691 2760
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 0 2546 800 2576
rect 4110 2546 4170 2758
rect 5625 2755 5691 2758
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 19139 2687 19455 2688
rect 5073 2682 5139 2685
rect 8569 2682 8635 2685
rect 5073 2680 8635 2682
rect 5073 2624 5078 2680
rect 5134 2624 8574 2680
rect 8630 2624 8635 2680
rect 5073 2622 8635 2624
rect 5073 2619 5139 2622
rect 8569 2619 8635 2622
rect 9765 2682 9831 2685
rect 9990 2682 9996 2684
rect 9765 2680 9996 2682
rect 9765 2624 9770 2680
rect 9826 2624 9996 2680
rect 9765 2622 9996 2624
rect 9765 2619 9831 2622
rect 9990 2620 9996 2622
rect 10060 2620 10066 2684
rect 12709 2682 12775 2685
rect 12390 2680 12775 2682
rect 12390 2624 12714 2680
rect 12770 2624 12775 2680
rect 12390 2622 12775 2624
rect 0 2486 4170 2546
rect 5441 2546 5507 2549
rect 5758 2546 5764 2548
rect 5441 2544 5764 2546
rect 5441 2488 5446 2544
rect 5502 2488 5764 2544
rect 5441 2486 5764 2488
rect 0 2456 800 2486
rect 5441 2483 5507 2486
rect 5758 2484 5764 2486
rect 5828 2484 5834 2548
rect 10593 2546 10659 2549
rect 12390 2546 12450 2622
rect 12709 2619 12775 2622
rect 5904 2544 12450 2546
rect 5904 2488 10598 2544
rect 10654 2488 12450 2544
rect 5904 2486 12450 2488
rect 13169 2546 13235 2549
rect 17861 2546 17927 2549
rect 13169 2544 17927 2546
rect 13169 2488 13174 2544
rect 13230 2488 17866 2544
rect 17922 2488 17927 2544
rect 13169 2486 17927 2488
rect 3969 2410 4035 2413
rect 5904 2410 5964 2486
rect 10593 2483 10659 2486
rect 13169 2483 13235 2486
rect 17861 2483 17927 2486
rect 18229 2546 18295 2549
rect 22200 2546 23000 2576
rect 18229 2544 23000 2546
rect 18229 2488 18234 2544
rect 18290 2488 23000 2544
rect 18229 2486 23000 2488
rect 18229 2483 18295 2486
rect 22200 2456 23000 2486
rect 3969 2408 5964 2410
rect 3969 2352 3974 2408
rect 4030 2352 5964 2408
rect 3969 2350 5964 2352
rect 7649 2410 7715 2413
rect 7782 2410 7788 2412
rect 7649 2408 7788 2410
rect 7649 2352 7654 2408
rect 7710 2352 7788 2408
rect 7649 2350 7788 2352
rect 3969 2347 4035 2350
rect 7649 2347 7715 2350
rect 7782 2348 7788 2350
rect 7852 2410 7858 2412
rect 21357 2410 21423 2413
rect 7852 2408 21423 2410
rect 7852 2352 21362 2408
rect 21418 2352 21423 2408
rect 7852 2350 21423 2352
rect 7852 2348 7858 2350
rect 21357 2347 21423 2350
rect 8293 2274 8359 2277
rect 9438 2274 9444 2276
rect 8293 2272 9444 2274
rect 8293 2216 8298 2272
rect 8354 2216 9444 2272
rect 8293 2214 9444 2216
rect 8293 2211 8359 2214
rect 9438 2212 9444 2214
rect 9508 2212 9514 2276
rect 6144 2208 6460 2209
rect 0 2138 800 2168
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 21738 2143 22054 2144
rect 3969 2138 4035 2141
rect 0 2136 4035 2138
rect 0 2080 3974 2136
rect 4030 2080 4035 2136
rect 0 2078 4035 2080
rect 0 2048 800 2078
rect 3969 2075 4035 2078
rect 12249 2138 12315 2141
rect 12750 2138 12756 2140
rect 12249 2136 12756 2138
rect 12249 2080 12254 2136
rect 12310 2080 12756 2136
rect 12249 2078 12756 2080
rect 12249 2075 12315 2078
rect 12750 2076 12756 2078
rect 12820 2076 12826 2140
rect 19006 2138 19012 2140
rect 16990 2078 19012 2138
rect 9622 1940 9628 2004
rect 9692 2002 9698 2004
rect 11973 2002 12039 2005
rect 16990 2002 17050 2078
rect 19006 2076 19012 2078
rect 19076 2076 19082 2140
rect 22200 2138 23000 2168
rect 22142 2048 23000 2138
rect 9692 2000 17050 2002
rect 9692 1944 11978 2000
rect 12034 1944 17050 2000
rect 9692 1942 17050 1944
rect 18689 2002 18755 2005
rect 22142 2002 22202 2048
rect 18689 2000 22202 2002
rect 18689 1944 18694 2000
rect 18750 1944 22202 2000
rect 18689 1942 22202 1944
rect 9692 1940 9698 1942
rect 11973 1939 12039 1942
rect 18689 1939 18755 1942
rect 6637 1866 6703 1869
rect 12249 1866 12315 1869
rect 12934 1866 12940 1868
rect 6637 1864 12315 1866
rect 6637 1808 6642 1864
rect 6698 1808 12254 1864
rect 12310 1808 12315 1864
rect 6637 1806 12315 1808
rect 6637 1803 6703 1806
rect 12249 1803 12315 1806
rect 12390 1806 12940 1866
rect 0 1730 800 1760
rect 2957 1730 3023 1733
rect 0 1728 3023 1730
rect 0 1672 2962 1728
rect 3018 1672 3023 1728
rect 0 1670 3023 1672
rect 0 1640 800 1670
rect 2957 1667 3023 1670
rect 4797 1730 4863 1733
rect 5717 1730 5783 1733
rect 12014 1730 12020 1732
rect 4797 1728 12020 1730
rect 4797 1672 4802 1728
rect 4858 1672 5722 1728
rect 5778 1672 12020 1728
rect 4797 1670 12020 1672
rect 4797 1667 4863 1670
rect 5717 1667 5783 1670
rect 12014 1668 12020 1670
rect 12084 1668 12090 1732
rect 4429 1594 4495 1597
rect 12390 1594 12450 1806
rect 12934 1804 12940 1806
rect 13004 1804 13010 1868
rect 17953 1730 18019 1733
rect 22200 1730 23000 1760
rect 17953 1728 23000 1730
rect 17953 1672 17958 1728
rect 18014 1672 23000 1728
rect 17953 1670 23000 1672
rect 17953 1667 18019 1670
rect 22200 1640 23000 1670
rect 4429 1592 12450 1594
rect 4429 1536 4434 1592
rect 4490 1536 12450 1592
rect 4429 1534 12450 1536
rect 4429 1531 4495 1534
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 17172 20436 17236 20500
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3924 19544 3988 19548
rect 3924 19488 3938 19544
rect 3938 19488 3988 19544
rect 3924 19484 3988 19488
rect 14596 19484 14660 19548
rect 1164 19348 1228 19412
rect 14412 19348 14476 19412
rect 17540 19408 17604 19412
rect 17540 19352 17554 19408
rect 17554 19352 17604 19408
rect 17540 19348 17604 19352
rect 16988 19136 17052 19140
rect 16988 19080 17038 19136
rect 17038 19080 17052 19136
rect 16988 19076 17052 19080
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 4660 18668 4724 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 5764 18260 5828 18324
rect 2084 18124 2148 18188
rect 9996 18124 10060 18188
rect 15516 17988 15580 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 11100 17580 11164 17644
rect 7788 17444 7852 17508
rect 10732 17504 10796 17508
rect 10732 17448 10746 17504
rect 10746 17448 10796 17504
rect 10732 17444 10796 17448
rect 18644 17504 18708 17508
rect 18644 17448 18658 17504
rect 18658 17448 18708 17504
rect 18644 17444 18708 17448
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 14964 17308 15028 17372
rect 9812 17172 9876 17236
rect 3188 17036 3252 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 3004 16628 3068 16692
rect 8524 16688 8588 16692
rect 8524 16632 8574 16688
rect 8574 16632 8588 16688
rect 8524 16628 8588 16632
rect 20484 16628 20548 16692
rect 2636 16492 2700 16556
rect 7604 16356 7668 16420
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 5212 16084 5276 16148
rect 7788 15948 7852 16012
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 980 15404 1044 15468
rect 12204 15268 12268 15332
rect 15332 15268 15396 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 4292 15132 4356 15196
rect 10732 15132 10796 15196
rect 17172 15132 17236 15196
rect 19012 14996 19076 15060
rect 2452 14860 2516 14924
rect 6684 14724 6748 14788
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 17540 14452 17604 14516
rect 7604 14316 7668 14380
rect 8340 14180 8404 14244
rect 11100 14180 11164 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 7052 14044 7116 14108
rect 5580 13908 5644 13972
rect 3924 13772 3988 13836
rect 4108 13772 4172 13836
rect 7972 13772 8036 13836
rect 12020 13832 12084 13836
rect 12020 13776 12034 13832
rect 12034 13776 12084 13832
rect 12020 13772 12084 13776
rect 12756 13832 12820 13836
rect 12756 13776 12770 13832
rect 12770 13776 12820 13832
rect 12756 13772 12820 13776
rect 20116 13772 20180 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 4476 13364 4540 13428
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 3372 12820 3436 12884
rect 10180 12684 10244 12748
rect 11836 12880 11900 12884
rect 11836 12824 11850 12880
rect 11850 12824 11900 12880
rect 11836 12820 11900 12824
rect 5948 12548 6012 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 5396 12412 5460 12476
rect 8156 12412 8220 12476
rect 12940 12472 13004 12476
rect 12940 12416 12990 12472
rect 12990 12416 13004 12472
rect 12940 12412 13004 12416
rect 5396 12276 5460 12340
rect 6684 12276 6748 12340
rect 8156 12276 8220 12340
rect 9260 12276 9324 12340
rect 18644 12064 18708 12068
rect 18644 12008 18658 12064
rect 18658 12008 18708 12064
rect 18644 12004 18708 12008
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6684 11324 6748 11388
rect 4292 11052 4356 11116
rect 4844 11052 4908 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 9444 10780 9508 10844
rect 16988 10644 17052 10708
rect 8156 10508 8220 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 15332 10236 15396 10300
rect 7052 9964 7116 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 2084 9556 2148 9620
rect 2636 9556 2700 9620
rect 5764 9556 5828 9620
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 4844 9012 4908 9076
rect 10180 8876 10244 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 8340 8604 8404 8668
rect 6868 8332 6932 8396
rect 8156 8196 8220 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 4108 7924 4172 7988
rect 5764 7924 5828 7988
rect 9812 7924 9876 7988
rect 2636 7516 2700 7580
rect 19012 7652 19076 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 18644 7516 18708 7580
rect 6684 7380 6748 7444
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 3188 7032 3252 7036
rect 3188 6976 3202 7032
rect 3202 6976 3252 7032
rect 3188 6972 3252 6976
rect 1532 6564 1596 6628
rect 12204 6836 12268 6900
rect 4844 6700 4908 6764
rect 5948 6700 6012 6764
rect 5764 6564 5828 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 7420 6428 7484 6492
rect 9444 6428 9508 6492
rect 3924 6156 3988 6220
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 5948 5884 6012 5948
rect 9444 5884 9508 5948
rect 3004 5748 3068 5812
rect 4476 5808 4540 5812
rect 4476 5752 4490 5808
rect 4490 5752 4540 5808
rect 4476 5748 4540 5752
rect 1532 5536 1596 5540
rect 1532 5480 1546 5536
rect 1546 5480 1596 5536
rect 1532 5476 1596 5480
rect 6684 5476 6748 5540
rect 7972 5476 8036 5540
rect 8524 5536 8588 5540
rect 8524 5480 8574 5536
rect 8574 5480 8588 5536
rect 8524 5476 8588 5480
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 6868 5340 6932 5404
rect 20484 5340 20548 5404
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 2452 5068 2516 5132
rect 4660 5068 4724 5132
rect 980 4932 1044 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 3372 4796 3436 4860
rect 6684 4856 6748 4860
rect 6684 4800 6698 4856
rect 6698 4800 6748 4856
rect 6684 4796 6748 4800
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 5580 4252 5644 4316
rect 9628 4116 9692 4180
rect 1164 3980 1228 4044
rect 5212 3980 5276 4044
rect 7788 3980 7852 4044
rect 14964 3980 15028 4044
rect 15516 3980 15580 4044
rect 11100 3844 11164 3908
rect 11836 3844 11900 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6868 3708 6932 3772
rect 9444 3708 9508 3772
rect 14596 3708 14660 3772
rect 9260 3436 9324 3500
rect 11100 3300 11164 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 14412 3164 14476 3228
rect 19012 3164 19076 3228
rect 7420 3028 7484 3092
rect 6684 2892 6748 2956
rect 20116 3088 20180 3092
rect 20116 3032 20166 3088
rect 20166 3032 20180 3088
rect 20116 3028 20180 3032
rect 2636 2756 2700 2820
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 9996 2620 10060 2684
rect 5764 2484 5828 2548
rect 7788 2348 7852 2412
rect 9444 2212 9508 2276
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 12756 2076 12820 2140
rect 9628 1940 9692 2004
rect 19012 2076 19076 2140
rect 12020 1668 12084 1732
rect 12940 1804 13004 1868
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 1163 19412 1229 19413
rect 1163 19348 1164 19412
rect 1228 19348 1229 19412
rect 1163 19347 1229 19348
rect 979 15468 1045 15469
rect 979 15404 980 15468
rect 1044 15404 1045 15468
rect 979 15403 1045 15404
rect 982 4997 1042 15403
rect 979 4996 1045 4997
rect 979 4932 980 4996
rect 1044 4932 1045 4996
rect 979 4931 1045 4932
rect 1166 4045 1226 19347
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 3923 19548 3989 19549
rect 3923 19484 3924 19548
rect 3988 19484 3989 19548
rect 3923 19483 3989 19484
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 2083 18188 2149 18189
rect 2083 18124 2084 18188
rect 2148 18124 2149 18188
rect 2083 18123 2149 18124
rect 2086 9621 2146 18123
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3187 17100 3253 17101
rect 3187 17036 3188 17100
rect 3252 17036 3253 17100
rect 3187 17035 3253 17036
rect 3003 16692 3069 16693
rect 3003 16628 3004 16692
rect 3068 16628 3069 16692
rect 3003 16627 3069 16628
rect 2635 16556 2701 16557
rect 2635 16492 2636 16556
rect 2700 16492 2701 16556
rect 2635 16491 2701 16492
rect 2451 14924 2517 14925
rect 2451 14860 2452 14924
rect 2516 14860 2517 14924
rect 2451 14859 2517 14860
rect 2083 9620 2149 9621
rect 2083 9556 2084 9620
rect 2148 9556 2149 9620
rect 2083 9555 2149 9556
rect 1531 6628 1597 6629
rect 1531 6564 1532 6628
rect 1596 6564 1597 6628
rect 1531 6563 1597 6564
rect 1534 5541 1594 6563
rect 1531 5540 1597 5541
rect 1531 5476 1532 5540
rect 1596 5476 1597 5540
rect 1531 5475 1597 5476
rect 2454 5133 2514 14859
rect 2638 9621 2698 16491
rect 2635 9620 2701 9621
rect 2635 9556 2636 9620
rect 2700 9556 2701 9620
rect 2635 9555 2701 9556
rect 2635 7580 2701 7581
rect 2635 7516 2636 7580
rect 2700 7516 2701 7580
rect 2635 7515 2701 7516
rect 2451 5132 2517 5133
rect 2451 5068 2452 5132
rect 2516 5068 2517 5132
rect 2451 5067 2517 5068
rect 1163 4044 1229 4045
rect 1163 3980 1164 4044
rect 1228 3980 1229 4044
rect 1163 3979 1229 3980
rect 2638 2821 2698 7515
rect 3006 5813 3066 16627
rect 3190 7037 3250 17035
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3926 13837 3986 19483
rect 4659 18732 4725 18733
rect 4659 18668 4660 18732
rect 4724 18668 4725 18732
rect 4659 18667 4725 18668
rect 4291 15196 4357 15197
rect 4291 15132 4292 15196
rect 4356 15132 4357 15196
rect 4291 15131 4357 15132
rect 3923 13836 3989 13837
rect 3923 13772 3924 13836
rect 3988 13772 3989 13836
rect 3923 13771 3989 13772
rect 4107 13836 4173 13837
rect 4107 13772 4108 13836
rect 4172 13772 4173 13836
rect 4107 13771 4173 13772
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3371 12884 3437 12885
rect 3371 12820 3372 12884
rect 3436 12820 3437 12884
rect 3371 12819 3437 12820
rect 3187 7036 3253 7037
rect 3187 6972 3188 7036
rect 3252 6972 3253 7036
rect 3187 6971 3253 6972
rect 3003 5812 3069 5813
rect 3003 5748 3004 5812
rect 3068 5748 3069 5812
rect 3003 5747 3069 5748
rect 3374 4861 3434 12819
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3926 6221 3986 13771
rect 4110 7989 4170 13771
rect 4294 11117 4354 15131
rect 4475 13428 4541 13429
rect 4475 13364 4476 13428
rect 4540 13364 4541 13428
rect 4475 13363 4541 13364
rect 4291 11116 4357 11117
rect 4291 11052 4292 11116
rect 4356 11052 4357 11116
rect 4291 11051 4357 11052
rect 4107 7988 4173 7989
rect 4107 7924 4108 7988
rect 4172 7924 4173 7988
rect 4107 7923 4173 7924
rect 3923 6220 3989 6221
rect 3923 6156 3924 6220
rect 3988 6156 3989 6220
rect 3923 6155 3989 6156
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 4478 5813 4538 13363
rect 4475 5812 4541 5813
rect 4475 5748 4476 5812
rect 4540 5748 4541 5812
rect 4475 5747 4541 5748
rect 4662 5133 4722 18667
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5763 18324 5829 18325
rect 5763 18260 5764 18324
rect 5828 18260 5829 18324
rect 5763 18259 5829 18260
rect 5211 16148 5277 16149
rect 5211 16084 5212 16148
rect 5276 16084 5277 16148
rect 5211 16083 5277 16084
rect 4843 11116 4909 11117
rect 4843 11052 4844 11116
rect 4908 11052 4909 11116
rect 4843 11051 4909 11052
rect 4846 9077 4906 11051
rect 4843 9076 4909 9077
rect 4843 9012 4844 9076
rect 4908 9012 4909 9076
rect 4843 9011 4909 9012
rect 4846 6765 4906 9011
rect 4843 6764 4909 6765
rect 4843 6700 4844 6764
rect 4908 6700 4909 6764
rect 4843 6699 4909 6700
rect 4659 5132 4725 5133
rect 4659 5068 4660 5132
rect 4724 5068 4725 5132
rect 4659 5067 4725 5068
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3371 4860 3437 4861
rect 3371 4796 3372 4860
rect 3436 4796 3437 4860
rect 3371 4795 3437 4796
rect 3543 3840 3863 4864
rect 5214 4045 5274 16083
rect 5579 13972 5645 13973
rect 5579 13908 5580 13972
rect 5644 13908 5645 13972
rect 5579 13907 5645 13908
rect 5395 12476 5461 12477
rect 5395 12412 5396 12476
rect 5460 12412 5461 12476
rect 5395 12411 5461 12412
rect 5398 12341 5458 12411
rect 5395 12340 5461 12341
rect 5395 12276 5396 12340
rect 5460 12276 5461 12340
rect 5395 12275 5461 12276
rect 5582 4317 5642 13907
rect 5766 9621 5826 18259
rect 6142 17440 6462 18464
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 9995 18188 10061 18189
rect 9995 18124 9996 18188
rect 10060 18124 10061 18188
rect 9995 18123 10061 18124
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 7787 17508 7853 17509
rect 7787 17444 7788 17508
rect 7852 17444 7853 17508
rect 7787 17443 7853 17444
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 7603 16420 7669 16421
rect 7603 16356 7604 16420
rect 7668 16356 7669 16420
rect 7603 16355 7669 16356
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6683 14788 6749 14789
rect 6683 14724 6684 14788
rect 6748 14724 6749 14788
rect 6683 14723 6749 14724
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 5947 12612 6013 12613
rect 5947 12548 5948 12612
rect 6012 12548 6013 12612
rect 5947 12547 6013 12548
rect 5763 9620 5829 9621
rect 5763 9556 5764 9620
rect 5828 9556 5829 9620
rect 5763 9555 5829 9556
rect 5763 7988 5829 7989
rect 5763 7924 5764 7988
rect 5828 7924 5829 7988
rect 5763 7923 5829 7924
rect 5766 6629 5826 7923
rect 5950 6765 6010 12547
rect 6142 12000 6462 13024
rect 6686 12341 6746 14723
rect 7606 14381 7666 16355
rect 7790 16013 7850 17443
rect 8741 16896 9061 17920
rect 9811 17236 9877 17237
rect 9811 17172 9812 17236
rect 9876 17172 9877 17236
rect 9811 17171 9877 17172
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 7787 16012 7853 16013
rect 7787 15948 7788 16012
rect 7852 15948 7853 16012
rect 7787 15947 7853 15948
rect 7603 14380 7669 14381
rect 7603 14316 7604 14380
rect 7668 14316 7669 14380
rect 7603 14315 7669 14316
rect 7051 14108 7117 14109
rect 7051 14044 7052 14108
rect 7116 14044 7117 14108
rect 7051 14043 7117 14044
rect 6683 12340 6749 12341
rect 6683 12276 6684 12340
rect 6748 12276 6749 12340
rect 6683 12275 6749 12276
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6683 11388 6749 11389
rect 6683 11324 6684 11388
rect 6748 11324 6749 11388
rect 6683 11323 6749 11324
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5947 6764 6013 6765
rect 5947 6700 5948 6764
rect 6012 6700 6013 6764
rect 5947 6699 6013 6700
rect 5763 6628 5829 6629
rect 5763 6564 5764 6628
rect 5828 6564 5829 6628
rect 5763 6563 5829 6564
rect 5579 4316 5645 4317
rect 5579 4252 5580 4316
rect 5644 4252 5645 4316
rect 5579 4251 5645 4252
rect 5211 4044 5277 4045
rect 5211 3980 5212 4044
rect 5276 3980 5277 4044
rect 5211 3979 5277 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 2635 2820 2701 2821
rect 2635 2756 2636 2820
rect 2700 2756 2701 2820
rect 2635 2755 2701 2756
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 5766 2549 5826 6563
rect 5950 5949 6010 6699
rect 6142 6560 6462 7584
rect 6686 7445 6746 11323
rect 7054 10029 7114 14043
rect 7051 10028 7117 10029
rect 7051 9964 7052 10028
rect 7116 9964 7117 10028
rect 7051 9963 7117 9964
rect 6867 8396 6933 8397
rect 6867 8332 6868 8396
rect 6932 8332 6933 8396
rect 6867 8331 6933 8332
rect 6683 7444 6749 7445
rect 6683 7380 6684 7444
rect 6748 7380 6749 7444
rect 6683 7379 6749 7380
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 5947 5948 6013 5949
rect 5947 5884 5948 5948
rect 6012 5884 6013 5948
rect 5947 5883 6013 5884
rect 6142 5472 6462 6496
rect 6686 5541 6746 7379
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6870 5405 6930 8331
rect 7419 6492 7485 6493
rect 7419 6428 7420 6492
rect 7484 6428 7485 6492
rect 7419 6427 7485 6428
rect 6867 5404 6933 5405
rect 6867 5340 6868 5404
rect 6932 5340 6933 5404
rect 6867 5339 6933 5340
rect 6683 4860 6749 4861
rect 6683 4796 6684 4860
rect 6748 4796 6749 4860
rect 6683 4795 6749 4796
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5763 2548 5829 2549
rect 5763 2484 5764 2548
rect 5828 2484 5829 2548
rect 5763 2483 5829 2484
rect 6142 2208 6462 3232
rect 6686 2957 6746 4795
rect 6870 3773 6930 5339
rect 6867 3772 6933 3773
rect 6867 3708 6868 3772
rect 6932 3708 6933 3772
rect 6867 3707 6933 3708
rect 7422 3093 7482 6427
rect 7419 3092 7485 3093
rect 7419 3028 7420 3092
rect 7484 3028 7485 3092
rect 7419 3027 7485 3028
rect 6683 2956 6749 2957
rect 6683 2892 6684 2956
rect 6748 2892 6749 2956
rect 6683 2891 6749 2892
rect 7606 2790 7666 14315
rect 7790 4045 7850 15947
rect 8339 14244 8405 14245
rect 8339 14180 8340 14244
rect 8404 14180 8405 14244
rect 8339 14179 8405 14180
rect 7971 13836 8037 13837
rect 7971 13772 7972 13836
rect 8036 13772 8037 13836
rect 7971 13771 8037 13772
rect 7974 5541 8034 13771
rect 8155 12476 8221 12477
rect 8155 12412 8156 12476
rect 8220 12412 8221 12476
rect 8155 12411 8221 12412
rect 8158 12341 8218 12411
rect 8155 12340 8221 12341
rect 8155 12276 8156 12340
rect 8220 12276 8221 12340
rect 8155 12275 8221 12276
rect 8155 10572 8221 10573
rect 8155 10508 8156 10572
rect 8220 10508 8221 10572
rect 8155 10507 8221 10508
rect 8158 8261 8218 10507
rect 8342 8669 8402 14179
rect 8339 8668 8405 8669
rect 8339 8604 8340 8668
rect 8404 8604 8405 8668
rect 8339 8603 8405 8604
rect 8155 8260 8221 8261
rect 8155 8196 8156 8260
rect 8220 8196 8221 8260
rect 8155 8195 8221 8196
rect 8526 5541 8586 16627
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 9259 12340 9325 12341
rect 9259 12276 9260 12340
rect 9324 12276 9325 12340
rect 9259 12275 9325 12276
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 7971 5540 8037 5541
rect 7971 5476 7972 5540
rect 8036 5476 8037 5540
rect 7971 5475 8037 5476
rect 8523 5540 8589 5541
rect 8523 5476 8524 5540
rect 8588 5476 8589 5540
rect 8523 5475 8589 5476
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 7787 4044 7853 4045
rect 7787 3980 7788 4044
rect 7852 3980 7853 4044
rect 7787 3979 7853 3980
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7606 2730 7850 2790
rect 7790 2413 7850 2730
rect 8741 2752 9061 3776
rect 9262 3501 9322 12275
rect 9443 10844 9509 10845
rect 9443 10780 9444 10844
rect 9508 10780 9509 10844
rect 9443 10779 9509 10780
rect 9446 6493 9506 10779
rect 9814 7989 9874 17171
rect 9811 7988 9877 7989
rect 9811 7924 9812 7988
rect 9876 7924 9877 7988
rect 9811 7923 9877 7924
rect 9443 6492 9509 6493
rect 9443 6428 9444 6492
rect 9508 6428 9509 6492
rect 9443 6427 9509 6428
rect 9443 5948 9509 5949
rect 9443 5884 9444 5948
rect 9508 5884 9509 5948
rect 9443 5883 9509 5884
rect 9446 3773 9506 5883
rect 9627 4180 9693 4181
rect 9627 4116 9628 4180
rect 9692 4116 9693 4180
rect 9627 4115 9693 4116
rect 9443 3772 9509 3773
rect 9443 3708 9444 3772
rect 9508 3708 9509 3772
rect 9443 3707 9509 3708
rect 9259 3500 9325 3501
rect 9259 3436 9260 3500
rect 9324 3436 9325 3500
rect 9259 3435 9325 3436
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 7787 2412 7853 2413
rect 7787 2348 7788 2412
rect 7852 2348 7853 2412
rect 7787 2347 7853 2348
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9446 2277 9506 3707
rect 9443 2276 9509 2277
rect 9443 2212 9444 2276
rect 9508 2212 9509 2276
rect 9443 2211 9509 2212
rect 9630 2005 9690 4115
rect 9998 2685 10058 18123
rect 11099 17644 11165 17645
rect 11099 17580 11100 17644
rect 11164 17580 11165 17644
rect 11099 17579 11165 17580
rect 10731 17508 10797 17509
rect 10731 17444 10732 17508
rect 10796 17444 10797 17508
rect 10731 17443 10797 17444
rect 10734 15197 10794 17443
rect 10731 15196 10797 15197
rect 10731 15132 10732 15196
rect 10796 15132 10797 15196
rect 10731 15131 10797 15132
rect 11102 14245 11162 17579
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 17171 20500 17237 20501
rect 17171 20436 17172 20500
rect 17236 20436 17237 20500
rect 17171 20435 17237 20436
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 14595 19548 14661 19549
rect 14595 19484 14596 19548
rect 14660 19484 14661 19548
rect 14595 19483 14661 19484
rect 14411 19412 14477 19413
rect 14411 19348 14412 19412
rect 14476 19348 14477 19412
rect 14411 19347 14477 19348
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 12203 15332 12269 15333
rect 12203 15268 12204 15332
rect 12268 15268 12269 15332
rect 12203 15267 12269 15268
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11099 14244 11165 14245
rect 11099 14180 11100 14244
rect 11164 14180 11165 14244
rect 11099 14179 11165 14180
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 12019 13836 12085 13837
rect 12019 13772 12020 13836
rect 12084 13772 12085 13836
rect 12019 13771 12085 13772
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 10179 12748 10245 12749
rect 10179 12684 10180 12748
rect 10244 12684 10245 12748
rect 10179 12683 10245 12684
rect 10182 8941 10242 12683
rect 11340 12000 11660 13024
rect 11835 12884 11901 12885
rect 11835 12820 11836 12884
rect 11900 12820 11901 12884
rect 11835 12819 11901 12820
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 10179 8940 10245 8941
rect 10179 8876 10180 8940
rect 10244 8876 10245 8940
rect 10179 8875 10245 8876
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11099 3908 11165 3909
rect 11099 3844 11100 3908
rect 11164 3844 11165 3908
rect 11099 3843 11165 3844
rect 11102 3365 11162 3843
rect 11099 3364 11165 3365
rect 11099 3300 11100 3364
rect 11164 3300 11165 3364
rect 11099 3299 11165 3300
rect 11340 3296 11660 4320
rect 11838 3909 11898 12819
rect 11835 3908 11901 3909
rect 11835 3844 11836 3908
rect 11900 3844 11901 3908
rect 11835 3843 11901 3844
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9995 2684 10061 2685
rect 9995 2620 9996 2684
rect 10060 2620 10061 2684
rect 9995 2619 10061 2620
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 9627 2004 9693 2005
rect 9627 1940 9628 2004
rect 9692 1940 9693 2004
rect 9627 1939 9693 1940
rect 12022 1733 12082 13771
rect 12206 6901 12266 15267
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 12755 13836 12821 13837
rect 12755 13772 12756 13836
rect 12820 13772 12821 13836
rect 12755 13771 12821 13772
rect 12203 6900 12269 6901
rect 12203 6836 12204 6900
rect 12268 6836 12269 6900
rect 12203 6835 12269 6836
rect 12758 2141 12818 13771
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 12939 12476 13005 12477
rect 12939 12412 12940 12476
rect 13004 12412 13005 12476
rect 12939 12411 13005 12412
rect 12755 2140 12821 2141
rect 12755 2076 12756 2140
rect 12820 2076 12821 2140
rect 12755 2075 12821 2076
rect 12942 1869 13002 12411
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 14414 3229 14474 19347
rect 14598 3773 14658 19483
rect 16538 18528 16858 19552
rect 16987 19140 17053 19141
rect 16987 19076 16988 19140
rect 17052 19076 17053 19140
rect 16987 19075 17053 19076
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 15515 18052 15581 18053
rect 15515 17988 15516 18052
rect 15580 17988 15581 18052
rect 15515 17987 15581 17988
rect 14963 17372 15029 17373
rect 14963 17308 14964 17372
rect 15028 17308 15029 17372
rect 14963 17307 15029 17308
rect 14966 4045 15026 17307
rect 15331 15332 15397 15333
rect 15331 15268 15332 15332
rect 15396 15268 15397 15332
rect 15331 15267 15397 15268
rect 15334 10301 15394 15267
rect 15331 10300 15397 10301
rect 15331 10236 15332 10300
rect 15396 10236 15397 10300
rect 15331 10235 15397 10236
rect 15518 4045 15578 17987
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16990 10709 17050 19075
rect 17174 15197 17234 20435
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 17539 19412 17605 19413
rect 17539 19348 17540 19412
rect 17604 19348 17605 19412
rect 17539 19347 17605 19348
rect 17171 15196 17237 15197
rect 17171 15132 17172 15196
rect 17236 15132 17237 15196
rect 17171 15131 17237 15132
rect 17542 14517 17602 19347
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 18643 17508 18709 17509
rect 18643 17444 18644 17508
rect 18708 17444 18709 17508
rect 18643 17443 18709 17444
rect 17539 14516 17605 14517
rect 17539 14452 17540 14516
rect 17604 14452 17605 14516
rect 17539 14451 17605 14452
rect 18646 12069 18706 17443
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 21736 20704 22056 20720
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 20483 16692 20549 16693
rect 20483 16628 20484 16692
rect 20548 16628 20549 16692
rect 20483 16627 20549 16628
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19011 15060 19077 15061
rect 19011 14996 19012 15060
rect 19076 14996 19077 15060
rect 19011 14995 19077 14996
rect 18643 12068 18709 12069
rect 18643 12004 18644 12068
rect 18708 12004 18709 12068
rect 18643 12003 18709 12004
rect 16987 10708 17053 10709
rect 16987 10644 16988 10708
rect 17052 10644 17053 10708
rect 16987 10643 17053 10644
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 18646 7581 18706 12003
rect 19014 7717 19074 14995
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 20115 13836 20181 13837
rect 20115 13772 20116 13836
rect 20180 13772 20181 13836
rect 20115 13771 20181 13772
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19011 7716 19077 7717
rect 19011 7652 19012 7716
rect 19076 7652 19077 7716
rect 19011 7651 19077 7652
rect 18643 7580 18709 7581
rect 18643 7516 18644 7580
rect 18708 7516 18709 7580
rect 18643 7515 18709 7516
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 15515 4044 15581 4045
rect 15515 3980 15516 4044
rect 15580 3980 15581 4044
rect 15515 3979 15581 3980
rect 14595 3772 14661 3773
rect 14595 3708 14596 3772
rect 14660 3708 14661 3772
rect 14595 3707 14661 3708
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 14411 3228 14477 3229
rect 14411 3164 14412 3228
rect 14476 3164 14477 3228
rect 14411 3163 14477 3164
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 2208 16858 3232
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19011 3228 19077 3229
rect 19011 3164 19012 3228
rect 19076 3164 19077 3228
rect 19011 3163 19077 3164
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19014 2141 19074 3163
rect 19137 2752 19457 3776
rect 20118 3093 20178 13771
rect 20486 5405 20546 16627
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 20483 5404 20549 5405
rect 20483 5340 20484 5404
rect 20548 5340 20549 5404
rect 20483 5339 20549 5340
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 20115 3092 20181 3093
rect 20115 3028 20116 3092
rect 20180 3028 20181 3092
rect 20115 3027 20181 3028
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19011 2140 19077 2141
rect 19011 2076 19012 2140
rect 19076 2076 19077 2140
rect 19137 2128 19457 2688
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 2128 22056 2144
rect 19011 2075 19077 2076
rect 12939 1868 13005 1869
rect 12939 1804 12940 1868
rect 13004 1804 13005 1868
rect 12939 1803 13005 1804
rect 12019 1732 12085 1733
rect 12019 1668 12020 1732
rect 12084 1668 12085 1732
rect 12019 1667 12085 1668
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform 1 0 3404 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform 1 0 3772 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 4140 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform -1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 20424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform -1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform -1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform 1 0 18768 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform -1 0 12512 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 5060 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 12512 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 4968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 3220 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 5152 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 6624 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 6164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 4416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 9200 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 15824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 12604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 4692 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 10948 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 10120 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 9844 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 9476 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 9016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 6900 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 13156 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 8464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 5888 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 4324 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11224 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 17204 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17572 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 15272 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3__D
timestamp 1649977179
transform 1 0 17204 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 16284 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11868 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 10948 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18308 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 16836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform 1 0 15640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18768 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16744 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 15456 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3__CLK
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 17112 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 15272 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0__CLK
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1__CLK
timestamp 1649977179
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2__CLK
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5520 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4140 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8280 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7544 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9568 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 4876 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_0__S
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l3_in_1__S
timestamp 1649977179
transform -1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l4_in_0__S
timestamp 1649977179
transform -1 0 5152 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8004 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 6072 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_3__S
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__S
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 6440 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 6532 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 16744 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l3_in_1__A1
timestamp 1649977179
transform -1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8280 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 12972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__S
timestamp 1649977179
transform -1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 17572 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__S
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 7544 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__S
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 6532 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 16192 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 15732 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 15272 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__S
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__S
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 17204 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__S
timestamp 1649977179
transform -1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_115
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_219
timestamp 1649977179
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_24
timestamp 1649977179
transform 1 0 3312 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_47
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_66
timestamp 1649977179
transform 1 0 7176 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_71
timestamp 1649977179
transform 1 0 7636 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_86
timestamp 1649977179
transform 1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_91
timestamp 1649977179
transform 1 0 9476 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_129
timestamp 1649977179
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_140
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_200
timestamp 1649977179
transform 1 0 19504 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_204
timestamp 1649977179
transform 1 0 19872 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_50
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_62
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_67
timestamp 1649977179
transform 1 0 7268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_72
timestamp 1649977179
transform 1 0 7728 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_125
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_130
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_134
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_158
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_166
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_172
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_183
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_210
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_10
timestamp 1649977179
transform 1 0 2024 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_24
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1649977179
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_67
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_79
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_117
timestamp 1649977179
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_126
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 1649977179
transform 1 0 13064 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_135
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_140
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_163
timestamp 1649977179
transform 1 0 16100 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_172
timestamp 1649977179
transform 1 0 16928 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_183
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_187
timestamp 1649977179
transform 1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_218
timestamp 1649977179
transform 1 0 21160 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_222
timestamp 1649977179
transform 1 0 21528 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_36
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_46
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_58
timestamp 1649977179
transform 1 0 6440 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_63
timestamp 1649977179
transform 1 0 6900 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_68
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_73
timestamp 1649977179
transform 1 0 7820 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_80
timestamp 1649977179
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_98
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_117
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1649977179
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_145
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_168
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_187
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1649977179
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_215
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_11
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_26
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_30
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_60
timestamp 1649977179
transform 1 0 6624 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_64
timestamp 1649977179
transform 1 0 6992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_68
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_73
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_79
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_84
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_88
timestamp 1649977179
transform 1 0 9200 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_106
timestamp 1649977179
transform 1 0 10856 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_115
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_119
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_139
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_143
timestamp 1649977179
transform 1 0 14260 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_147
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 1649977179
transform 1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_162
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_172
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_177
timestamp 1649977179
transform 1 0 17388 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_182
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_186
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_191
timestamp 1649977179
transform 1 0 18676 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_197
timestamp 1649977179
transform 1 0 19228 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_32
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_60
timestamp 1649977179
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_75
timestamp 1649977179
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 1649977179
transform 1 0 9384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_108
timestamp 1649977179
transform 1 0 11040 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_112
timestamp 1649977179
transform 1 0 11408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_122
timestamp 1649977179
transform 1 0 12328 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_127
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_158
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_162
timestamp 1649977179
transform 1 0 16008 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_179
timestamp 1649977179
transform 1 0 17572 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_184
timestamp 1649977179
transform 1 0 18032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_14
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_25
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_41
timestamp 1649977179
transform 1 0 4876 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_64
timestamp 1649977179
transform 1 0 6992 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 1649977179
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_90
timestamp 1649977179
transform 1 0 9384 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_96
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_108
timestamp 1649977179
transform 1 0 11040 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_135
timestamp 1649977179
transform 1 0 13524 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_139
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_150
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1649977179
transform 1 0 17848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_210
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_7
timestamp 1649977179
transform 1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_12
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_104
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_108
timestamp 1649977179
transform 1 0 11040 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_112
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_117
timestamp 1649977179
transform 1 0 11868 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_143
timestamp 1649977179
transform 1 0 14260 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_170
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_181
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_18
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_44
timestamp 1649977179
transform 1 0 5152 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_59
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_77
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1649977179
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_133
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_152
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_160
timestamp 1649977179
transform 1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp 1649977179
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_36
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_44
timestamp 1649977179
transform 1 0 5152 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_69
timestamp 1649977179
transform 1 0 7452 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_119
timestamp 1649977179
transform 1 0 12052 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_123
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_127
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_130
timestamp 1649977179
transform 1 0 13064 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_134
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_145
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_149
timestamp 1649977179
transform 1 0 14812 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_161
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_188
timestamp 1649977179
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_203
timestamp 1649977179
transform 1 0 19780 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_214
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 1649977179
transform 1 0 3312 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_29
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_35
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_50
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_63
timestamp 1649977179
transform 1 0 6900 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_67
timestamp 1649977179
transform 1 0 7268 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_85
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_94
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_98
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_115
timestamp 1649977179
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_119
timestamp 1649977179
transform 1 0 12052 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_127
timestamp 1649977179
transform 1 0 12788 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_131
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_135
timestamp 1649977179
transform 1 0 13524 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_139
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_173
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_201
timestamp 1649977179
transform 1 0 19596 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_19
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_69
timestamp 1649977179
transform 1 0 7452 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_79
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_143
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_152
timestamp 1649977179
transform 1 0 15088 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1649977179
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_208
timestamp 1649977179
transform 1 0 20240 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_28
timestamp 1649977179
transform 1 0 3680 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_53
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_60
timestamp 1649977179
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_115
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_144
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_173
timestamp 1649977179
transform 1 0 17020 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_177
timestamp 1649977179
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_199
timestamp 1649977179
transform 1 0 19412 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_209
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_13
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_32
timestamp 1649977179
transform 1 0 4048 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_50
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_60
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_76
timestamp 1649977179
transform 1 0 8096 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_87
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_107
timestamp 1649977179
transform 1 0 10948 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_111
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_119
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_148
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_152
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_156
timestamp 1649977179
transform 1 0 15456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_160
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_182
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_35
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_43
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_67
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_78
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_15_129
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_148
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_152
timestamp 1649977179
transform 1 0 15088 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_162
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_172
timestamp 1649977179
transform 1 0 16928 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_176
timestamp 1649977179
transform 1 0 17296 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_180
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_198
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_21
timestamp 1649977179
transform 1 0 3036 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_47
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_69
timestamp 1649977179
transform 1 0 7452 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_125
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_131
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_155
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_215
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_42
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_61
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_72
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_76
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_80
timestamp 1649977179
transform 1 0 8464 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_132
timestamp 1649977179
transform 1 0 13248 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_136
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_140
timestamp 1649977179
transform 1 0 13984 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_173
timestamp 1649977179
transform 1 0 17020 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_177
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_199
timestamp 1649977179
transform 1 0 19412 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_209
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 1649977179
transform 1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_13
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_24
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_39
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_43
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_47
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_51
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_56
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_60
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_72
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_78
timestamp 1649977179
transform 1 0 8280 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_104
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_122
timestamp 1649977179
transform 1 0 12328 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_152
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_156
timestamp 1649977179
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_178
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_182
timestamp 1649977179
transform 1 0 17848 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_203
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_18
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_33
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_38
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_42
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_76
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_138
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_157
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_172
timestamp 1649977179
transform 1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_176
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_180
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 1649977179
transform 1 0 19320 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 1649977179
transform 1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_209
timestamp 1649977179
transform 1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_21
timestamp 1649977179
transform 1 0 3036 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_42
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_45
timestamp 1649977179
transform 1 0 5244 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_67
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_78
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_106
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_110
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_114
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_118
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_122
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_126
timestamp 1649977179
transform 1 0 12696 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_130
timestamp 1649977179
transform 1 0 13064 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_146
timestamp 1649977179
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_152
timestamp 1649977179
transform 1 0 15088 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_156
timestamp 1649977179
transform 1 0 15456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_160
timestamp 1649977179
transform 1 0 15824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1649977179
transform 1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_214
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_20
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_40
timestamp 1649977179
transform 1 0 4784 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_44
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_49
timestamp 1649977179
transform 1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_67
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_73
timestamp 1649977179
transform 1 0 7820 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_77
timestamp 1649977179
transform 1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_85
timestamp 1649977179
transform 1 0 8924 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_104
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_117
timestamp 1649977179
transform 1 0 11868 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_144
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_173
timestamp 1649977179
transform 1 0 17020 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_195
timestamp 1649977179
transform 1 0 19044 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_202
timestamp 1649977179
transform 1 0 19688 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_19
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1649977179
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_56
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_76
timestamp 1649977179
transform 1 0 8096 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_80
timestamp 1649977179
transform 1 0 8464 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_91
timestamp 1649977179
transform 1 0 9476 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_95
timestamp 1649977179
transform 1 0 9844 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_13
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_18
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_23
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_31
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_47
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_61
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_80
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_84
timestamp 1649977179
transform 1 0 8832 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_115
timestamp 1649977179
transform 1 0 11684 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_119
timestamp 1649977179
transform 1 0 12052 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_123
timestamp 1649977179
transform 1 0 12420 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_131
timestamp 1649977179
transform 1 0 13156 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_154
timestamp 1649977179
transform 1 0 15272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_159
timestamp 1649977179
transform 1 0 15732 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_189
timestamp 1649977179
transform 1 0 18492 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_195
timestamp 1649977179
transform 1 0 19044 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_202
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_220
timestamp 1649977179
transform 1 0 21344 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_21
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_33
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_50
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_54
timestamp 1649977179
transform 1 0 6072 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_64
timestamp 1649977179
transform 1 0 6992 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_68
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_78
timestamp 1649977179
transform 1 0 8280 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_104
timestamp 1649977179
transform 1 0 10672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_112
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_116
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_124 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12512 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_169
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_173
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_199
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_204
timestamp 1649977179
transform 1 0 19872 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_22
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_26
timestamp 1649977179
transform 1 0 3496 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_41
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_52
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_79
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_83
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_103
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_107
timestamp 1649977179
transform 1 0 10948 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_115
timestamp 1649977179
transform 1 0 11684 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_127 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_133
timestamp 1649977179
transform 1 0 13340 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_136
timestamp 1649977179
transform 1 0 13616 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_147
timestamp 1649977179
transform 1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_172
timestamp 1649977179
transform 1 0 16928 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_201
timestamp 1649977179
transform 1 0 19596 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_209
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_12
timestamp 1649977179
transform 1 0 2208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_16
timestamp 1649977179
transform 1 0 2576 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_20
timestamp 1649977179
transform 1 0 2944 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_55
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_59
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_63
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_67
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_70
timestamp 1649977179
transform 1 0 7544 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_89
timestamp 1649977179
transform 1 0 9292 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_93
timestamp 1649977179
transform 1 0 9660 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_104
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_119
timestamp 1649977179
transform 1 0 12052 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_26_134
timestamp 1649977179
transform 1 0 13432 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_159
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1649977179
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_214
timestamp 1649977179
transform 1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_17
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_37
timestamp 1649977179
transform 1 0 4508 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_48
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_68
timestamp 1649977179
transform 1 0 7360 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_95
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_99
timestamp 1649977179
transform 1 0 10212 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_128 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_154
timestamp 1649977179
transform 1 0 15272 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_172
timestamp 1649977179
transform 1 0 16928 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 1649977179
transform 1 0 17296 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_180
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1649977179
transform 1 0 18400 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_191
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_196
timestamp 1649977179
transform 1 0 19136 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_201
timestamp 1649977179
transform 1 0 19596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_218
timestamp 1649977179
transform 1 0 21160 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_222
timestamp 1649977179
transform 1 0 21528 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_13
timestamp 1649977179
transform 1 0 2300 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_32
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_36
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_47
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_58
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_70
timestamp 1649977179
transform 1 0 7544 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1649977179
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_88
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_105
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_111
timestamp 1649977179
transform 1 0 11316 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_131
timestamp 1649977179
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_149
timestamp 1649977179
transform 1 0 14812 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_164
timestamp 1649977179
transform 1 0 16192 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_169
timestamp 1649977179
transform 1 0 16652 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_173
timestamp 1649977179
transform 1 0 17020 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_188
timestamp 1649977179
transform 1 0 18400 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1649977179
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_60
timestamp 1649977179
transform 1 0 6624 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_67
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1649977179
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_99
timestamp 1649977179
transform 1 0 10212 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_107
timestamp 1649977179
transform 1 0 10948 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1649977179
transform 1 0 12420 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_128
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_143
timestamp 1649977179
transform 1 0 14260 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_163
timestamp 1649977179
transform 1 0 16100 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_171
timestamp 1649977179
transform 1 0 16836 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_175
timestamp 1649977179
transform 1 0 17204 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_179
timestamp 1649977179
transform 1 0 17572 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_190
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_54
timestamp 1649977179
transform 1 0 6072 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_59
timestamp 1649977179
transform 1 0 6532 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_63
timestamp 1649977179
transform 1 0 6900 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_67
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_79
timestamp 1649977179
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_92
timestamp 1649977179
transform 1 0 9568 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_104
timestamp 1649977179
transform 1 0 10672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_110
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_132
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_155
timestamp 1649977179
transform 1 0 15364 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_166
timestamp 1649977179
transform 1 0 16376 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_186
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_190
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1649977179
transform 1 0 20056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_31
timestamp 1649977179
transform 1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 1649977179
transform 1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1649977179
transform 1 0 5520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_59
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_67
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_79
timestamp 1649977179
transform 1 0 8372 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_102
timestamp 1649977179
transform 1 0 10488 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1649977179
transform 1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_129
timestamp 1649977179
transform 1 0 12972 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_150
timestamp 1649977179
transform 1 0 14904 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_154
timestamp 1649977179
transform 1 0 15272 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_157
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1649977179
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_171
timestamp 1649977179
transform 1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1649977179
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_190
timestamp 1649977179
transform 1 0 18584 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_199
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_204
timestamp 1649977179
transform 1 0 19872 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_18
timestamp 1649977179
transform 1 0 2760 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_35
timestamp 1649977179
transform 1 0 4324 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_39
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_93
timestamp 1649977179
transform 1 0 9660 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_120
timestamp 1649977179
transform 1 0 12144 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_132
timestamp 1649977179
transform 1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_150
timestamp 1649977179
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_172
timestamp 1649977179
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_200
timestamp 1649977179
transform 1 0 19504 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_204
timestamp 1649977179
transform 1 0 19872 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_32_208
timestamp 1649977179
transform 1 0 20240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_18
timestamp 1649977179
transform 1 0 2760 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_23
timestamp 1649977179
transform 1 0 3220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_31
timestamp 1649977179
transform 1 0 3956 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_35
timestamp 1649977179
transform 1 0 4324 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_71
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_76
timestamp 1649977179
transform 1 0 8096 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_124
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_136
timestamp 1649977179
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_158
timestamp 1649977179
transform 1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp 1649977179
transform 1 0 16008 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_186
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_190
timestamp 1649977179
transform 1 0 18584 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _056_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13984 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform -1 0 2760 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 3128 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 2852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 19780 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 19688 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 19872 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 16928 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 20332 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 19780 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 16652 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 20240 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 12788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 7268 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 7268 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 8188 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 16100 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 17388 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 17848 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 18032 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 18492 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 13524 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 13064 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 4876 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 14168 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 5796 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 3036 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 2300 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 4416 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform -1 0 2300 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 20516 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 20332 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 20332 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 18952 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 20332 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform 1 0 20516 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 16468 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 20516 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 21436 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 17940 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 18952 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 8372 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 8280 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform 1 0 12052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 8004 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 7912 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform 1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform 1 0 6808 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input74
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input78
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform -1 0 3220 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input81
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1649977179
transform -1 0 14628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 15088 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1649977179
transform -1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19412 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13892 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13524 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11040 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12052 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13340 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10580 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10212 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14536 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16652 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19964 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20424 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18032 0 1 7616
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12144 0 1 3264
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13708 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11868 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10672 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12788 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10672 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9384 0 1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13248 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16008 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20884 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21344 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17572 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21252 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18308 0 1 4352
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16560 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17940 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19504 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20884 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 19872 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20792 0 1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17572 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4324 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2668 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l1_in_3__172 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4324 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3864 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l1_in_3__182
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4968 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5336 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6440 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7360 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l1_in_3__155
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3312 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_7.mux_l1_in_3__156
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5980 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6624 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9016 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_1__157
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8280 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_11.mux_l2_in_1__173
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8556 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8832 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_13.mux_l1_in_1__174
timestamp 1649977179
transform -1 0 6716 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_15.mux_l1_in_1__175
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l1_in_1__176
timestamp 1649977179
transform 1 0 6992 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7360 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_19.mux_l1_in_1__177
timestamp 1649977179
transform 1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9936 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_21.mux_l1_in_1__178
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12420 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13432 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10672 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_23.mux_l1_in_1__179
timestamp 1649977179
transform 1 0 12328 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11684 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__180
timestamp 1649977179
transform 1 0 14996 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15732 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_27.mux_l2_in_0__181
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4876 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__158
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4416 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2576 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7452 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2392 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__161
timestamp 1649977179
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2944 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2760 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 3496 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform -1 0 2392 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform -1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_3__163
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 1656 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2484 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3680 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__164
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4692 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_3__159
timestamp 1649977179
transform 1 0 3220 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5244 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_3__160
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform -1 0 3588 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3864 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 3680 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_1__162
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20424 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 9384 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__165
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 16192 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 18768 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18584 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__167
timestamp 1649977179
transform 1 0 12512 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8556 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20240 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 20608 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 18768 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 12696 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform -1 0 18584 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20332 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 20424 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 17940 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_3__170
timestamp 1649977179
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 18308 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19136 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21344 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20516 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7544 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6992 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__171
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 12420 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13708 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16560 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_3__166
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14628 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_3__168
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14536 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15364 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17112 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_1__169
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 16836 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 2300 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 2300 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 20516 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 14720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  repeater151
timestamp 1649977179
transform -1 0 19780 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater152
timestamp 1649977179
transform -1 0 20240 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater153
timestamp 1649977179
transform -1 0 2852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater154
timestamp 1649977179
transform -1 0 11868 0 -1 4352
box -38 -48 406 592
<< labels >>
flabel metal2 s 19890 0 19946 800 0 FreeSans 224 90 0 0 SC_IN_BOT
port 0 nsew signal input
flabel metal2 s 20258 0 20314 800 0 FreeSans 224 90 0 0 SC_OUT_BOT
port 1 nsew signal tristate
flabel metal4 s 6142 2128 6462 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 11340 2128 11660 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 16538 2128 16858 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 21736 2128 22056 20720 0 FreeSans 1920 90 0 0 VGND
port 2 nsew ground bidirectional
flabel metal4 s 3543 2128 3863 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 8741 2128 9061 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 13939 2128 14259 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal4 s 19137 2128 19457 20720 0 FreeSans 1920 90 0 0 VPWR
port 3 nsew power bidirectional
flabel metal2 s 2226 0 2282 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_42_
port 4 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_43_
port 5 nsew signal input
flabel metal2 s 2962 0 3018 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_44_
port 6 nsew signal input
flabel metal2 s 3330 0 3386 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_45_
port 7 nsew signal input
flabel metal2 s 3698 0 3754 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_46_
port 8 nsew signal input
flabel metal2 s 4066 0 4122 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_47_
port 9 nsew signal input
flabel metal2 s 4434 0 4490 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_48_
port 10 nsew signal input
flabel metal2 s 4802 0 4858 800 0 FreeSans 224 90 0 0 bottom_left_grid_pin_49_
port 11 nsew signal input
flabel metal2 s 5722 22200 5778 23000 0 FreeSans 224 90 0 0 ccff_head
port 12 nsew signal input
flabel metal2 s 17222 22200 17278 23000 0 FreeSans 224 90 0 0 ccff_tail
port 13 nsew signal tristate
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 chanx_left_in[0]
port 14 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 chanx_left_in[10]
port 15 nsew signal input
flabel metal3 s 0 9392 800 9512 0 FreeSans 480 0 0 0 chanx_left_in[11]
port 16 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 chanx_left_in[12]
port 17 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 chanx_left_in[13]
port 18 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 chanx_left_in[14]
port 19 nsew signal input
flabel metal3 s 0 11024 800 11144 0 FreeSans 480 0 0 0 chanx_left_in[15]
port 20 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 chanx_left_in[16]
port 21 nsew signal input
flabel metal3 s 0 11840 800 11960 0 FreeSans 480 0 0 0 chanx_left_in[17]
port 22 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 chanx_left_in[18]
port 23 nsew signal input
flabel metal3 s 0 12656 800 12776 0 FreeSans 480 0 0 0 chanx_left_in[19]
port 24 nsew signal input
flabel metal3 s 0 5312 800 5432 0 FreeSans 480 0 0 0 chanx_left_in[1]
port 25 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 chanx_left_in[2]
port 26 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 chanx_left_in[3]
port 27 nsew signal input
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 chanx_left_in[4]
port 28 nsew signal input
flabel metal3 s 0 6944 800 7064 0 FreeSans 480 0 0 0 chanx_left_in[5]
port 29 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 chanx_left_in[6]
port 30 nsew signal input
flabel metal3 s 0 7760 800 7880 0 FreeSans 480 0 0 0 chanx_left_in[7]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 chanx_left_in[8]
port 32 nsew signal input
flabel metal3 s 0 8576 800 8696 0 FreeSans 480 0 0 0 chanx_left_in[9]
port 33 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 chanx_left_out[0]
port 34 nsew signal tristate
flabel metal3 s 0 17144 800 17264 0 FreeSans 480 0 0 0 chanx_left_out[10]
port 35 nsew signal tristate
flabel metal3 s 0 17552 800 17672 0 FreeSans 480 0 0 0 chanx_left_out[11]
port 36 nsew signal tristate
flabel metal3 s 0 17960 800 18080 0 FreeSans 480 0 0 0 chanx_left_out[12]
port 37 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 chanx_left_out[13]
port 38 nsew signal tristate
flabel metal3 s 0 18776 800 18896 0 FreeSans 480 0 0 0 chanx_left_out[14]
port 39 nsew signal tristate
flabel metal3 s 0 19184 800 19304 0 FreeSans 480 0 0 0 chanx_left_out[15]
port 40 nsew signal tristate
flabel metal3 s 0 19592 800 19712 0 FreeSans 480 0 0 0 chanx_left_out[16]
port 41 nsew signal tristate
flabel metal3 s 0 20000 800 20120 0 FreeSans 480 0 0 0 chanx_left_out[17]
port 42 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 chanx_left_out[18]
port 43 nsew signal tristate
flabel metal3 s 0 20816 800 20936 0 FreeSans 480 0 0 0 chanx_left_out[19]
port 44 nsew signal tristate
flabel metal3 s 0 13472 800 13592 0 FreeSans 480 0 0 0 chanx_left_out[1]
port 45 nsew signal tristate
flabel metal3 s 0 13880 800 14000 0 FreeSans 480 0 0 0 chanx_left_out[2]
port 46 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 chanx_left_out[3]
port 47 nsew signal tristate
flabel metal3 s 0 14696 800 14816 0 FreeSans 480 0 0 0 chanx_left_out[4]
port 48 nsew signal tristate
flabel metal3 s 0 15104 800 15224 0 FreeSans 480 0 0 0 chanx_left_out[5]
port 49 nsew signal tristate
flabel metal3 s 0 15512 800 15632 0 FreeSans 480 0 0 0 chanx_left_out[6]
port 50 nsew signal tristate
flabel metal3 s 0 15920 800 16040 0 FreeSans 480 0 0 0 chanx_left_out[7]
port 51 nsew signal tristate
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 chanx_left_out[8]
port 52 nsew signal tristate
flabel metal3 s 0 16736 800 16856 0 FreeSans 480 0 0 0 chanx_left_out[9]
port 53 nsew signal tristate
flabel metal3 s 22200 4904 23000 5024 0 FreeSans 480 0 0 0 chanx_right_in[0]
port 54 nsew signal input
flabel metal3 s 22200 8984 23000 9104 0 FreeSans 480 0 0 0 chanx_right_in[10]
port 55 nsew signal input
flabel metal3 s 22200 9392 23000 9512 0 FreeSans 480 0 0 0 chanx_right_in[11]
port 56 nsew signal input
flabel metal3 s 22200 9800 23000 9920 0 FreeSans 480 0 0 0 chanx_right_in[12]
port 57 nsew signal input
flabel metal3 s 22200 10208 23000 10328 0 FreeSans 480 0 0 0 chanx_right_in[13]
port 58 nsew signal input
flabel metal3 s 22200 10616 23000 10736 0 FreeSans 480 0 0 0 chanx_right_in[14]
port 59 nsew signal input
flabel metal3 s 22200 11024 23000 11144 0 FreeSans 480 0 0 0 chanx_right_in[15]
port 60 nsew signal input
flabel metal3 s 22200 11432 23000 11552 0 FreeSans 480 0 0 0 chanx_right_in[16]
port 61 nsew signal input
flabel metal3 s 22200 11840 23000 11960 0 FreeSans 480 0 0 0 chanx_right_in[17]
port 62 nsew signal input
flabel metal3 s 22200 12248 23000 12368 0 FreeSans 480 0 0 0 chanx_right_in[18]
port 63 nsew signal input
flabel metal3 s 22200 12656 23000 12776 0 FreeSans 480 0 0 0 chanx_right_in[19]
port 64 nsew signal input
flabel metal3 s 22200 5312 23000 5432 0 FreeSans 480 0 0 0 chanx_right_in[1]
port 65 nsew signal input
flabel metal3 s 22200 5720 23000 5840 0 FreeSans 480 0 0 0 chanx_right_in[2]
port 66 nsew signal input
flabel metal3 s 22200 6128 23000 6248 0 FreeSans 480 0 0 0 chanx_right_in[3]
port 67 nsew signal input
flabel metal3 s 22200 6536 23000 6656 0 FreeSans 480 0 0 0 chanx_right_in[4]
port 68 nsew signal input
flabel metal3 s 22200 6944 23000 7064 0 FreeSans 480 0 0 0 chanx_right_in[5]
port 69 nsew signal input
flabel metal3 s 22200 7352 23000 7472 0 FreeSans 480 0 0 0 chanx_right_in[6]
port 70 nsew signal input
flabel metal3 s 22200 7760 23000 7880 0 FreeSans 480 0 0 0 chanx_right_in[7]
port 71 nsew signal input
flabel metal3 s 22200 8168 23000 8288 0 FreeSans 480 0 0 0 chanx_right_in[8]
port 72 nsew signal input
flabel metal3 s 22200 8576 23000 8696 0 FreeSans 480 0 0 0 chanx_right_in[9]
port 73 nsew signal input
flabel metal3 s 22200 13064 23000 13184 0 FreeSans 480 0 0 0 chanx_right_out[0]
port 74 nsew signal tristate
flabel metal3 s 22200 17144 23000 17264 0 FreeSans 480 0 0 0 chanx_right_out[10]
port 75 nsew signal tristate
flabel metal3 s 22200 17552 23000 17672 0 FreeSans 480 0 0 0 chanx_right_out[11]
port 76 nsew signal tristate
flabel metal3 s 22200 17960 23000 18080 0 FreeSans 480 0 0 0 chanx_right_out[12]
port 77 nsew signal tristate
flabel metal3 s 22200 18368 23000 18488 0 FreeSans 480 0 0 0 chanx_right_out[13]
port 78 nsew signal tristate
flabel metal3 s 22200 18776 23000 18896 0 FreeSans 480 0 0 0 chanx_right_out[14]
port 79 nsew signal tristate
flabel metal3 s 22200 19184 23000 19304 0 FreeSans 480 0 0 0 chanx_right_out[15]
port 80 nsew signal tristate
flabel metal3 s 22200 19592 23000 19712 0 FreeSans 480 0 0 0 chanx_right_out[16]
port 81 nsew signal tristate
flabel metal3 s 22200 20000 23000 20120 0 FreeSans 480 0 0 0 chanx_right_out[17]
port 82 nsew signal tristate
flabel metal3 s 22200 20408 23000 20528 0 FreeSans 480 0 0 0 chanx_right_out[18]
port 83 nsew signal tristate
flabel metal3 s 22200 20816 23000 20936 0 FreeSans 480 0 0 0 chanx_right_out[19]
port 84 nsew signal tristate
flabel metal3 s 22200 13472 23000 13592 0 FreeSans 480 0 0 0 chanx_right_out[1]
port 85 nsew signal tristate
flabel metal3 s 22200 13880 23000 14000 0 FreeSans 480 0 0 0 chanx_right_out[2]
port 86 nsew signal tristate
flabel metal3 s 22200 14288 23000 14408 0 FreeSans 480 0 0 0 chanx_right_out[3]
port 87 nsew signal tristate
flabel metal3 s 22200 14696 23000 14816 0 FreeSans 480 0 0 0 chanx_right_out[4]
port 88 nsew signal tristate
flabel metal3 s 22200 15104 23000 15224 0 FreeSans 480 0 0 0 chanx_right_out[5]
port 89 nsew signal tristate
flabel metal3 s 22200 15512 23000 15632 0 FreeSans 480 0 0 0 chanx_right_out[6]
port 90 nsew signal tristate
flabel metal3 s 22200 15920 23000 16040 0 FreeSans 480 0 0 0 chanx_right_out[7]
port 91 nsew signal tristate
flabel metal3 s 22200 16328 23000 16448 0 FreeSans 480 0 0 0 chanx_right_out[8]
port 92 nsew signal tristate
flabel metal3 s 22200 16736 23000 16856 0 FreeSans 480 0 0 0 chanx_right_out[9]
port 93 nsew signal tristate
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 chany_bottom_in[0]
port 94 nsew signal input
flabel metal2 s 8850 0 8906 800 0 FreeSans 224 90 0 0 chany_bottom_in[10]
port 95 nsew signal input
flabel metal2 s 9218 0 9274 800 0 FreeSans 224 90 0 0 chany_bottom_in[11]
port 96 nsew signal input
flabel metal2 s 9586 0 9642 800 0 FreeSans 224 90 0 0 chany_bottom_in[12]
port 97 nsew signal input
flabel metal2 s 9954 0 10010 800 0 FreeSans 224 90 0 0 chany_bottom_in[13]
port 98 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 chany_bottom_in[14]
port 99 nsew signal input
flabel metal2 s 10690 0 10746 800 0 FreeSans 224 90 0 0 chany_bottom_in[15]
port 100 nsew signal input
flabel metal2 s 11058 0 11114 800 0 FreeSans 224 90 0 0 chany_bottom_in[16]
port 101 nsew signal input
flabel metal2 s 11426 0 11482 800 0 FreeSans 224 90 0 0 chany_bottom_in[17]
port 102 nsew signal input
flabel metal2 s 11794 0 11850 800 0 FreeSans 224 90 0 0 chany_bottom_in[18]
port 103 nsew signal input
flabel metal2 s 12162 0 12218 800 0 FreeSans 224 90 0 0 chany_bottom_in[19]
port 104 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 chany_bottom_in[1]
port 105 nsew signal input
flabel metal2 s 5906 0 5962 800 0 FreeSans 224 90 0 0 chany_bottom_in[2]
port 106 nsew signal input
flabel metal2 s 6274 0 6330 800 0 FreeSans 224 90 0 0 chany_bottom_in[3]
port 107 nsew signal input
flabel metal2 s 6642 0 6698 800 0 FreeSans 224 90 0 0 chany_bottom_in[4]
port 108 nsew signal input
flabel metal2 s 7010 0 7066 800 0 FreeSans 224 90 0 0 chany_bottom_in[5]
port 109 nsew signal input
flabel metal2 s 7378 0 7434 800 0 FreeSans 224 90 0 0 chany_bottom_in[6]
port 110 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 chany_bottom_in[7]
port 111 nsew signal input
flabel metal2 s 8114 0 8170 800 0 FreeSans 224 90 0 0 chany_bottom_in[8]
port 112 nsew signal input
flabel metal2 s 8482 0 8538 800 0 FreeSans 224 90 0 0 chany_bottom_in[9]
port 113 nsew signal input
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 chany_bottom_out[0]
port 114 nsew signal tristate
flabel metal2 s 16210 0 16266 800 0 FreeSans 224 90 0 0 chany_bottom_out[10]
port 115 nsew signal tristate
flabel metal2 s 16578 0 16634 800 0 FreeSans 224 90 0 0 chany_bottom_out[11]
port 116 nsew signal tristate
flabel metal2 s 16946 0 17002 800 0 FreeSans 224 90 0 0 chany_bottom_out[12]
port 117 nsew signal tristate
flabel metal2 s 17314 0 17370 800 0 FreeSans 224 90 0 0 chany_bottom_out[13]
port 118 nsew signal tristate
flabel metal2 s 17682 0 17738 800 0 FreeSans 224 90 0 0 chany_bottom_out[14]
port 119 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 chany_bottom_out[15]
port 120 nsew signal tristate
flabel metal2 s 18418 0 18474 800 0 FreeSans 224 90 0 0 chany_bottom_out[16]
port 121 nsew signal tristate
flabel metal2 s 18786 0 18842 800 0 FreeSans 224 90 0 0 chany_bottom_out[17]
port 122 nsew signal tristate
flabel metal2 s 19154 0 19210 800 0 FreeSans 224 90 0 0 chany_bottom_out[18]
port 123 nsew signal tristate
flabel metal2 s 19522 0 19578 800 0 FreeSans 224 90 0 0 chany_bottom_out[19]
port 124 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 chany_bottom_out[1]
port 125 nsew signal tristate
flabel metal2 s 13266 0 13322 800 0 FreeSans 224 90 0 0 chany_bottom_out[2]
port 126 nsew signal tristate
flabel metal2 s 13634 0 13690 800 0 FreeSans 224 90 0 0 chany_bottom_out[3]
port 127 nsew signal tristate
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 chany_bottom_out[4]
port 128 nsew signal tristate
flabel metal2 s 14370 0 14426 800 0 FreeSans 224 90 0 0 chany_bottom_out[5]
port 129 nsew signal tristate
flabel metal2 s 14738 0 14794 800 0 FreeSans 224 90 0 0 chany_bottom_out[6]
port 130 nsew signal tristate
flabel metal2 s 15106 0 15162 800 0 FreeSans 224 90 0 0 chany_bottom_out[7]
port 131 nsew signal tristate
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 chany_bottom_out[8]
port 132 nsew signal tristate
flabel metal2 s 15842 0 15898 800 0 FreeSans 224 90 0 0 chany_bottom_out[9]
port 133 nsew signal tristate
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 left_bottom_grid_pin_34_
port 134 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 left_bottom_grid_pin_35_
port 135 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 left_bottom_grid_pin_36_
port 136 nsew signal input
flabel metal3 s 0 2864 800 2984 0 FreeSans 480 0 0 0 left_bottom_grid_pin_37_
port 137 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 left_bottom_grid_pin_38_
port 138 nsew signal input
flabel metal3 s 0 3680 800 3800 0 FreeSans 480 0 0 0 left_bottom_grid_pin_39_
port 139 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 left_bottom_grid_pin_40_
port 140 nsew signal input
flabel metal3 s 0 4496 800 4616 0 FreeSans 480 0 0 0 left_bottom_grid_pin_41_
port 141 nsew signal input
flabel metal3 s 0 21224 800 21344 0 FreeSans 480 0 0 0 left_top_grid_pin_1_
port 142 nsew signal input
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 prog_clk_0_S_in
port 143 nsew signal input
flabel metal3 s 22200 1640 23000 1760 0 FreeSans 480 0 0 0 right_bottom_grid_pin_34_
port 144 nsew signal input
flabel metal3 s 22200 2048 23000 2168 0 FreeSans 480 0 0 0 right_bottom_grid_pin_35_
port 145 nsew signal input
flabel metal3 s 22200 2456 23000 2576 0 FreeSans 480 0 0 0 right_bottom_grid_pin_36_
port 146 nsew signal input
flabel metal3 s 22200 2864 23000 2984 0 FreeSans 480 0 0 0 right_bottom_grid_pin_37_
port 147 nsew signal input
flabel metal3 s 22200 3272 23000 3392 0 FreeSans 480 0 0 0 right_bottom_grid_pin_38_
port 148 nsew signal input
flabel metal3 s 22200 3680 23000 3800 0 FreeSans 480 0 0 0 right_bottom_grid_pin_39_
port 149 nsew signal input
flabel metal3 s 22200 4088 23000 4208 0 FreeSans 480 0 0 0 right_bottom_grid_pin_40_
port 150 nsew signal input
flabel metal3 s 22200 4496 23000 4616 0 FreeSans 480 0 0 0 right_bottom_grid_pin_41_
port 151 nsew signal input
flabel metal3 s 22200 21224 23000 21344 0 FreeSans 480 0 0 0 right_top_grid_pin_1_
port 152 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
