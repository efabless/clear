* NGSPICE file created from cbx_1__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_4 abstract view
.subckt sky130_fd_sc_hd__ebufn_4 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

.subckt cbx_1__2_ IO_ISOL_N SC_IN_BOT SC_IN_TOP SC_OUT_BOT SC_OUT_TOP VGND VPWR bottom_grid_pin_0_
+ bottom_grid_pin_10_ bottom_grid_pin_11_ bottom_grid_pin_12_ bottom_grid_pin_13_
+ bottom_grid_pin_14_ bottom_grid_pin_15_ bottom_grid_pin_1_ bottom_grid_pin_2_ bottom_grid_pin_3_
+ bottom_grid_pin_4_ bottom_grid_pin_5_ bottom_grid_pin_6_ bottom_grid_pin_7_ bottom_grid_pin_8_
+ bottom_grid_pin_9_ bottom_width_0_height_0__pin_0_ bottom_width_0_height_0__pin_1_lower
+ bottom_width_0_height_0__pin_1_upper ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chanx_right_in[0] chanx_right_in[10]
+ chanx_right_in[11] chanx_right_in[12] chanx_right_in[13] chanx_right_in[14] chanx_right_in[15]
+ chanx_right_in[16] chanx_right_in[17] chanx_right_in[18] chanx_right_in[19] chanx_right_in[1]
+ chanx_right_in[2] chanx_right_in[3] chanx_right_in[4] chanx_right_in[5] chanx_right_in[6]
+ chanx_right_in[7] chanx_right_in[8] chanx_right_in[9] chanx_right_out[0] chanx_right_out[10]
+ chanx_right_out[11] chanx_right_out[12] chanx_right_out[13] chanx_right_out[14]
+ chanx_right_out[15] chanx_right_out[16] chanx_right_out[17] chanx_right_out[18]
+ chanx_right_out[19] chanx_right_out[1] chanx_right_out[2] chanx_right_out[3] chanx_right_out[4]
+ chanx_right_out[5] chanx_right_out[6] chanx_right_out[7] chanx_right_out[8] chanx_right_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ prog_clk_0_S_in prog_clk_0_W_out top_grid_pin_0_
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_13.mux_l3_in_0_ mux_top_ipin_13.mux_l2_in_1_/X mux_top_ipin_13.mux_l2_in_0_/X
+ mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_66_ chanx_left_in[9] VGND VGND VPWR VPWR chanx_right_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_6.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_6.mux_l1_in_0_/X mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_49_ chanx_right_in[12] VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_3.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D ccff_head VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_1.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_65_ chanx_left_in[8] VGND VGND VPWR VPWR chanx_right_out[8] sky130_fd_sc_hd__buf_2
XFILLER_5_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_prog_clk_0_W_FTB01_A prog_clk_0_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_48_ chanx_right_in[11] VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_13.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_13.mux_l1_in_0_/X mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_6.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_0.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_bottom_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_64_ chanx_left_in[7] VGND VGND VPWR VPWR chanx_right_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_4_ sky130_fd_sc_hd__buf_4
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_47_ chanx_right_in[10] VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_top_ipin_14.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_12.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_bottom_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_63_ chanx_left_in[6] VGND VGND VPWR VPWR chanx_right_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xprog_clk_0_FTB00 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
X_46_ chanx_right_in[9] VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_29_ VGND VGND VPWR VPWR _29_/HI _29_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_11.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_11_ sky130_fd_sc_hd__buf_4
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_bottom_ipin_0.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR top_grid_pin_0_ sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_bottom_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_11.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l2_in_3_ _32_/HI chanx_right_in[15] mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_62_ chanx_left_in[5] VGND VGND VPWR VPWR chanx_right_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_4.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
+ gfpga_pad_EMBEDDED_IO_HD_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_45_ chanx_right_in[8] VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_2.mux_l4_in_0_ mux_top_ipin_2.mux_l3_in_1_/X mux_top_ipin_2.mux_l3_in_0_/X
+ mux_top_ipin_2.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_28_ VGND VGND VPWR VPWR _28_/HI _28_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_3_ _20_/HI chanx_right_in[18] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_2.mux_l3_in_1_ mux_top_ipin_2.mux_l2_in_3_/X mux_top_ipin_2.mux_l2_in_2_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_2.mux_l2_in_2__A1 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X ccff_head VGND VGND
+ VPWR VPWR mux_bottom_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_7.mux_l4_in_0_ mux_top_ipin_7.mux_l3_in_1_/X mux_top_ipin_7.mux_l3_in_0_/X
+ mux_top_ipin_7.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_61_ chanx_left_in[4] VGND VGND VPWR VPWR chanx_right_out[4] sky130_fd_sc_hd__buf_2
XFILLER_5_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_0.mux_l4_in_0__S mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l3_in_1_ mux_top_ipin_7.mux_l2_in_3_/X mux_top_ipin_7.mux_l2_in_2_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_44_ chanx_right_in[7] VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_27_ VGND VGND VPWR VPWR _27_/HI _27_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_7.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[12] mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__34__A SC_IN_TOP VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_9.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l3_in_0_ mux_top_ipin_2.mux_l2_in_1_/X mux_top_ipin_2.mux_l2_in_0_/X
+ mux_top_ipin_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_14.mux_l2_in_3_ _30_/HI chanx_right_in[19] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_13.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l4_in_0_ mux_top_ipin_14.mux_l3_in_1_/X mux_top_ipin_14.mux_l3_in_0_/X
+ mux_top_ipin_14.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_60_ chanx_left_in[3] VGND VGND VPWR VPWR chanx_right_out[3] sky130_fd_sc_hd__buf_2
XANTENNA__42__A chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A0 chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l3_in_0_ mux_top_ipin_7.mux_l2_in_1_/X mux_top_ipin_7.mux_l2_in_0_/X
+ mux_top_ipin_7.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__37__A chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_7.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_7_ sky130_fd_sc_hd__buf_4
X_43_ chanx_right_in[6] VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_14.mux_l3_in_1_ mux_top_ipin_14.mux_l2_in_3_/X mux_top_ipin_14.mux_l2_in_2_/X
+ mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_7.mux_l1_in_2_/X mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_26_ VGND VGND VPWR VPWR _26_/HI _26_/LO sky130_fd_sc_hd__conb_1
XFILLER_1_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__50__A chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2__D mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__45__A chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_7.mux_l1_in_2_ chanx_right_in[8] chanx_left_in[8] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_2.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_2.mux_l1_in_0_/X mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_11.mux_l2_in_2__A1 chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XANTENNA_mux_top_ipin_6.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_1__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__53__A chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_42_ chanx_right_in[5] VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__48__A chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l3_in_0_ mux_top_ipin_14.mux_l2_in_1_/X mux_top_ipin_14.mux_l2_in_0_/X
+ mux_top_ipin_14.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_11.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_7.mux_l2_in_0_ mux_top_ipin_7.mux_l1_in_1_/X mux_top_ipin_7.mux_l1_in_0_/X
+ mux_top_ipin_7.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_25_ VGND VGND VPWR VPWR _25_/HI _25_/LO sky130_fd_sc_hd__conb_1
XFILLER_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_14.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_14.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_14_ sky130_fd_sc_hd__buf_4
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__61__A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__56__A chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_14.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_2.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_41_ chanx_right_in[4] VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
XANTENNA__64__A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_24_ VGND VGND VPWR VPWR _24_/HI _24_/LO sky130_fd_sc_hd__conb_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_15.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__59__A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_14.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_14.mux_l1_in_0_/X mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_0_ sky130_fd_sc_hd__buf_4
XFILLER_21_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_7.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__72__A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__67__A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_14.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_40_ chanx_right_in[3] VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_23_ VGND VGND VPWR VPWR _23_/HI _23_/LO sky130_fd_sc_hd__conb_1
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__75__A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_13.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_73 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_14.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_14.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_22_ VGND VGND VPWR VPWR _22_/HI _22_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_10.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_7.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE gfpga_pad_EMBEDDED_IO_HD_SOC_IN
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR bottom_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_4
XFILLER_21_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_13.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_14.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_3.mux_l2_in_3_ _33_/HI chanx_right_in[14] mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_10.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_21_ VGND VGND VPWR VPWR _21_/HI _21_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_3.mux_l2_in_2__A1 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_7.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_3.mux_l4_in_0_ mux_top_ipin_3.mux_l3_in_1_/X mux_top_ipin_3.mux_l3_in_0_/X
+ mux_top_ipin_3.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_21_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l2_in_3_ _21_/HI chanx_right_in[19] mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l3_in_1_ mux_top_ipin_3.mux_l2_in_3_/X mux_top_ipin_3.mux_l2_in_2_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[8] mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l4_in_0_ mux_top_ipin_8.mux_l3_in_1_/X mux_top_ipin_8.mux_l3_in_0_/X
+ mux_top_ipin_8.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_3_ _26_/HI chanx_right_in[15] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_20_ VGND VGND VPWR VPWR _20_/HI _20_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_8.mux_l3_in_1_ mux_top_ipin_8.mux_l2_in_3_/X mux_top_ipin_8.mux_l2_in_2_/X
+ mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_14.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A0 chanx_right_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_8.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[13] mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l4_in_0_ mux_top_ipin_10.mux_l3_in_1_/X mux_top_ipin_10.mux_l3_in_0_/X
+ mux_top_ipin_10.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_3.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_3_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_3.mux_l3_in_0_ mux_top_ipin_3.mux_l2_in_1_/X mux_top_ipin_3.mux_l2_in_0_/X
+ mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_7.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l2_in_3_ _31_/HI chanx_right_in[16] mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l3_in_1_ mux_top_ipin_10.mux_l2_in_3_/X mux_top_ipin_10.mux_l2_in_2_/X
+ mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_3.mux_l2_in_1_ chanx_left_in[8] mux_top_ipin_3.mux_l1_in_2_/X mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[7] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l4_in_0_ mux_top_ipin_15.mux_l3_in_1_/X mux_top_ipin_15.mux_l3_in_0_/X
+ mux_top_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l3_in_0_ mux_top_ipin_8.mux_l2_in_1_/X mux_top_ipin_8.mux_l2_in_0_/X
+ mux_top_ipin_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_9.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_7.mux_l1_in_2__A1 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l3_in_1_ mux_top_ipin_15.mux_l2_in_3_/X mux_top_ipin_15.mux_l2_in_2_/X
+ mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_8.mux_l1_in_2_/X mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_12.mux_l2_in_2__A1 chanx_right_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l1_in_2_ chanx_right_in[9] chanx_left_in[9] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l3_in_0_ mux_top_ipin_10.mux_l2_in_1_/X mux_top_ipin_10.mux_l2_in_0_/X
+ mux_top_ipin_10.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_3.mux_l2_in_0_ mux_top_ipin_3.mux_l1_in_1_/X mux_top_ipin_3.mux_l1_in_0_/X
+ mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_10.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_10_ sky130_fd_sc_hd__buf_4
XANTENNA_mux_top_ipin_5.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_10.mux_l2_in_1_ chanx_left_in[7] chanx_right_in[3] mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_3.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A0 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l3_in_0_ mux_top_ipin_15.mux_l2_in_1_/X mux_top_ipin_15.mux_l2_in_0_/X
+ mux_top_ipin_15.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l2_in_0_ mux_top_ipin_8.mux_l1_in_1_/X mux_top_ipin_8.mux_l1_in_0_/X
+ mux_top_ipin_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_15.mux_l2_in_1_ chanx_left_in[10] mux_top_ipin_15.mux_l1_in_2_/X mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_4.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_15.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_top_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_10.mux_l2_in_0_ chanx_left_in[3] mux_top_ipin_10.mux_l1_in_0_/X mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_ipin_3.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_1__A1 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0__CLK
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l2_in_3__A1 chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_15.mux_l2_in_0_ mux_top_ipin_15.mux_l1_in_1_/X mux_top_ipin_15.mux_l1_in_0_/X
+ mux_top_ipin_15.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_8.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_76_ chanx_left_in[19] VGND VGND VPWR VPWR chanx_right_out[19] sky130_fd_sc_hd__buf_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_ipin_10.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_9.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_59_ chanx_left_in[2] VGND VGND VPWR VPWR chanx_right_out[2] sky130_fd_sc_hd__buf_2
XFILLER_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A0 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_6.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_6_ sky130_fd_sc_hd__buf_4
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_11.mux_l2_in_1__A0 chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_6.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_15.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_75_ chanx_left_in[18] VGND VGND VPWR VPWR chanx_right_out[18] sky130_fd_sc_hd__buf_2
XFILLER_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_13.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__40__A chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_58_ chanx_left_in[1] VGND VGND VPWR VPWR chanx_right_out[1] sky130_fd_sc_hd__buf_2
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__35__A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_ipin_11.mux_l1_in_2__A1 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_13.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_13_ sky130_fd_sc_hd__buf_4
XANTENNA__43__A chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_4.mux_l2_in_2__A1 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__38__A chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_3_ _17_/HI chanx_right_in[15] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_74_ chanx_left_in[17] VGND VGND VPWR VPWR chanx_right_out[17] sky130_fd_sc_hd__buf_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_ipin_0.mux_l2_in_3_ _23_/HI chanx_right_in[16] mux_bottom_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_57_ chanx_left_in[0] VGND VGND VPWR VPWR chanx_right_out[0] sky130_fd_sc_hd__buf_2
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__D mux_top_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__51__A chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE bottom_width_0_height_0__pin_0_
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ sky130_fd_sc_hd__ebufn_4
Xmux_top_ipin_4.mux_l4_in_0_ mux_top_ipin_4.mux_l3_in_1_/X mux_top_ipin_4.mux_l3_in_0_/X
+ mux_top_ipin_4.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__46__A chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_0__A0 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
+ bottom_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_0.mux_l4_in_0_ mux_bottom_ipin_0.mux_l3_in_1_/X mux_bottom_ipin_0.mux_l3_in_0_/X
+ mux_bottom_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_9.mux_l2_in_3_ _22_/HI chanx_right_in[14] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_4.mux_l3_in_1_ mux_top_ipin_4.mux_l2_in_3_/X mux_top_ipin_4.mux_l2_in_2_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_10.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_2__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_ipin_0.mux_l3_in_1_ mux_bottom_ipin_0.mux_l2_in_3_/X mux_bottom_ipin_0.mux_l2_in_2_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__54__A chanx_right_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_2_ chanx_left_in[15] chanx_right_in[9] mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_73_ chanx_left_in[16] VGND VGND VPWR VPWR chanx_right_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A0 chanx_right_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l4_in_0_ mux_top_ipin_9.mux_l3_in_1_/X mux_top_ipin_9.mux_l3_in_0_/X
+ mux_top_ipin_9.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__49__A chanx_right_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xprog_clk_0_W_FTB01 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_W_out sky130_fd_sc_hd__buf_4
Xmux_bottom_ipin_0.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[10] mux_bottom_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l2_in_3_ _27_/HI chanx_right_in[16] mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
X_56_ chanx_right_in[19] VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_8.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_9.mux_l3_in_1_ mux_top_ipin_9.mux_l2_in_3_/X mux_top_ipin_9.mux_l2_in_2_/X
+ mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_39_ chanx_right_in[2] VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_13.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__62__A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_9.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l4_in_0_ mux_top_ipin_11.mux_l3_in_1_/X mux_top_ipin_11.mux_l3_in_0_/X
+ mux_top_ipin_11.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__57__A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l3_in_0_ mux_top_ipin_4.mux_l2_in_1_/X mux_top_ipin_4.mux_l2_in_0_/X
+ mux_top_ipin_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_10.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_ipin_0.mux_l3_in_0_ mux_bottom_ipin_0.mux_l2_in_1_/X mux_bottom_ipin_0.mux_l2_in_0_/X
+ mux_bottom_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l3_in_1_ mux_top_ipin_11.mux_l2_in_3_/X mux_top_ipin_11.mux_l2_in_2_/X
+ mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__70__A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_72_ chanx_left_in[15] VGND VGND VPWR VPWR chanx_right_out[15] sky130_fd_sc_hd__buf_2
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l1_in_2__A1 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l2_in_1_ chanx_left_in[9] mux_top_ipin_4.mux_l1_in_2_/X mux_top_ipin_4.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__65__A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_11.mux_l2_in_2_ chanx_left_in[16] chanx_right_in[12] mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_0.mux_l2_in_1_ chanx_left_in[10] mux_bottom_ipin_0.mux_l1_in_2_/X
+ mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_55_ chanx_right_in[18] VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_13.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_4.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_9.mux_l3_in_0_ mux_top_ipin_9.mux_l2_in_1_/X mux_top_ipin_9.mux_l2_in_0_/X
+ mux_top_ipin_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_20_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_38_ chanx_right_in[1] VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmux_bottom_ipin_0.mux_l1_in_2_ chanx_right_in[4] chanx_left_in[4] mux_bottom_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_6.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_9.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_9.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_9_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_9.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__73__A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_10.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_10.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__68__A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_11.mux_l3_in_0_ mux_top_ipin_11.mux_l2_in_1_/X mux_top_ipin_11.mux_l2_in_0_/X
+ mux_top_ipin_11.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_71_ chanx_left_in[14] VGND VGND VPWR VPWR chanx_right_out[14] sky130_fd_sc_hd__buf_2
XFILLER_19_18 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_4.mux_l2_in_0_ mux_top_ipin_4.mux_l1_in_1_/X mux_top_ipin_4.mux_l1_in_0_/X
+ mux_top_ipin_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_3.mux_l2_in_1__A0 chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_54_ chanx_right_in[17] VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l2_in_1_ chanx_left_in[12] mux_top_ipin_11.mux_l1_in_2_/X mux_top_ipin_11.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_0.mux_l2_in_0_ mux_bottom_ipin_0.mux_l1_in_1_/X mux_bottom_ipin_0.mux_l1_in_0_/X
+ mux_bottom_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_3.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l3_in_0__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_4.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__76__A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_166 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_13.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_37_ chanx_right_in[0] VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_11.mux_l1_in_2_ chanx_right_in[6] chanx_left_in[6] mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_ipin_0.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_bottom_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_bottom_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_5.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_9.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_10.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_9.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_9.mux_l1_in_0_/X mux_top_ipin_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_6.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
X_70_ chanx_left_in[13] VGND VGND VPWR VPWR chanx_right_out[13] sky130_fd_sc_hd__buf_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_ipin_11.mux_l2_in_0_ mux_top_ipin_11.mux_l1_in_1_/X mux_top_ipin_11.mux_l1_in_0_/X
+ mux_top_ipin_11.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_11.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_3.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
X_53_ chanx_right_in[16] VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_4.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_4.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_1.mux_l2_in_3__A1 chanx_right_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_178 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_36_ bottom_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR bottom_width_0_height_0__pin_1_upper
+ sky130_fd_sc_hd__buf_2
Xmem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_12.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_ipin_0.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_bottom_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_11.mux_l1_in_1_ chanx_right_in[2] chanx_left_in[2] mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_19_ VGND VGND VPWR VPWR _19_/HI _19_/LO sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_2_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_9.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_9.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A0 chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_52_ chanx_right_in[15] VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_35_ SC_IN_BOT VGND VGND VPWR VPWR SC_OUT_TOP sky130_fd_sc_hd__buf_2
XFILLER_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_top_ipin_12.mux_l2_in_1__A0 chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_0.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_11.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_11.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ prog_clk_0_FTB00/X mux_top_ipin_15.mux_l4_in_0_/S VGND VGND VPWR VPWR ccff_tail
+ sky130_fd_sc_hd__dfxtp_1
X_18_ VGND VGND VPWR VPWR _18_/HI _18_/LO sky130_fd_sc_hd__conb_1
Xmem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_9.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
+ IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A0 chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_12.mux_l1_in_2__A1 chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_51_ chanx_right_in[14] VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_ipin_7.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_34_ SC_IN_TOP VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
XFILLER_22_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17_ VGND VGND VPWR VPWR _17_/HI _17_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_10.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_3_ _24_/HI chanx_right_in[17] mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_0.mux_l4_in_0_ mux_top_ipin_0.mux_l3_in_1_/X mux_top_ipin_0.mux_l3_in_0_/X
+ mux_top_ipin_0.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_50_ chanx_right_in[13] VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_2.mux_l2_in_0__A0 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_33_ VGND VGND VPWR VPWR _33_/HI _33_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l2_in_3_ _18_/HI chanx_right_in[18] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A0 chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l3_in_1_ mux_top_ipin_0.mux_l2_in_3_/X mux_top_ipin_0.mux_l2_in_2_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[11] mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l4_in_0_ mux_top_ipin_5.mux_l3_in_1_/X mux_top_ipin_5.mux_l3_in_0_/X
+ mux_top_ipin_5.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l3_in_1_ mux_top_ipin_5.mux_l2_in_3_/X mux_top_ipin_5.mux_l2_in_2_/X
+ mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A0 chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_5.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_32_ VGND VGND VPWR VPWR _32_/HI _32_/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_ipin_0.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l3_in_0_ mux_top_ipin_0.mux_l2_in_1_/X mux_top_ipin_0.mux_l2_in_0_/X
+ mux_top_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.mux_l2_in_3_ _28_/HI chanx_right_in[17] mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l2_in_1_ chanx_left_in[11] mux_top_ipin_0.mux_l1_in_2_/X mux_top_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l4_in_0_ mux_top_ipin_12.mux_l3_in_1_/X mux_top_ipin_12.mux_l3_in_0_/X
+ mux_top_ipin_12.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0__D mux_top_ipin_0.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_14.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_2_ chanx_right_in[5] chanx_left_in[5] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_5.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_5_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_5.mux_l3_in_0_ mux_top_ipin_5.mux_l2_in_1_/X mux_top_ipin_5.mux_l2_in_0_/X
+ mux_top_ipin_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_9.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l3_in_1_ mux_top_ipin_12.mux_l2_in_3_/X mux_top_ipin_12.mux_l2_in_2_/X
+ mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_7.mux_l2_in_3__A1 chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_5.mux_l2_in_1_ chanx_left_in[10] chanx_right_in[2] mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
X_31_ VGND VGND VPWR VPWR _31_/HI _31_/LO sky130_fd_sc_hd__conb_1
XFILLER_22_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l2_in_2_ chanx_left_in[17] chanx_right_in[13] mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A0 chanx_right_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l2_in_0_ mux_top_ipin_0.mux_l1_in_1_/X mux_top_ipin_0.mux_l1_in_0_/X
+ mux_top_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_4.mux_l2_in_1__A0 chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_0.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l3_in_0_ mux_top_ipin_12.mux_l2_in_1_/X mux_top_ipin_12.mux_l2_in_0_/X
+ mux_top_ipin_12.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_11.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_30_ VGND VGND VPWR VPWR _30_/HI _30_/LO sky130_fd_sc_hd__conb_1
Xmux_top_ipin_5.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_5.mux_l1_in_0_/X mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_6.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_12.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_12_ sky130_fd_sc_hd__buf_4
Xmux_top_ipin_12.mux_l2_in_1_ chanx_left_in[13] mux_top_ipin_12.mux_l1_in_2_/X mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_4.mux_l1_in_2__A1 chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_12.mux_l1_in_2_ chanx_right_in[7] chanx_left_in[7] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_0.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_0.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_2.mux_l2_in_3__A1 chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__41__A chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__36__A bottom_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l2_in_0_ mux_top_ipin_12.mux_l1_in_1_/X mux_top_ipin_12.mux_l1_in_0_/X
+ mux_top_ipin_12.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_ipin_5.mux_l1_in_0_ chanx_right_in[0] chanx_left_in[0] mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_ipin_12.mux_l1_in_1_ chanx_right_in[3] chanx_left_in[3] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__44__A chanx_right_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__39__A chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_3.mux_l2_in_0__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__52__A chanx_right_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A0 chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__47__A chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0 chanx_right_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_15.mux_l1_in_0__A1 chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_12.mux_l1_in_0_ chanx_right_in[1] chanx_left_in[1] mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__60__A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_3.mux_l2_in_3__S mux_top_ipin_3.mux_l2_in_3_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_8.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_12.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_8_ sky130_fd_sc_hd__buf_4
XANTENNA__55__A chanx_right_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_13.mux_l2_in_1__A1 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE ccff_tail
+ IO_ISOL_N VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR sky130_fd_sc_hd__or2b_4
XANTENNA_mux_top_ipin_11.mux_l2_in_3__A1 chanx_right_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A0 chanx_right_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_6.mux_l2_in_2__A1 chanx_right_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA__63__A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1 chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__58__A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_15.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A0 chanx_right_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_1.mux_l2_in_3_ _25_/HI chanx_right_in[14] mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_12.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_16_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__71__A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__66__A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A0 chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l3_in_1_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l4_in_0_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_10.mux_l1_in_0__A1 chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l4_in_0_ mux_top_ipin_1.mux_l3_in_1_/X mux_top_ipin_1.mux_l3_in_0_/X
+ mux_top_ipin_1.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_15.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_15_ sky130_fd_sc_hd__buf_4
XANTENNA_mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
X_69_ chanx_left_in[12] VGND VGND VPWR VPWR chanx_right_out[12] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l2_in_3_ _19_/HI chanx_right_in[19] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_1.mux_l3_in_1_ mux_top_ipin_1.mux_l2_in_3_/X mux_top_ipin_1.mux_l2_in_2_/X
+ mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_15.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_3.mux_l1_in_1__A1 chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__74__A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_2.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A0 chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__69__A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l2_in_2_ chanx_left_in[14] chanx_right_in[6] mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_ipin_6.mux_l4_in_0_ mux_top_ipin_6.mux_l3_in_1_/X mux_top_ipin_6.mux_l3_in_0_/X
+ mux_top_ipin_6.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_12.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_ipin_1.mux_l2_in_2__A1 chanx_right_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l3_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_1_ mux_top_ipin_6.mux_l2_in_3_/X mux_top_ipin_6.mux_l2_in_2_/X
+ mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_3.mux_l3_in_1__S mux_top_ipin_3.mux_l3_in_1_/S VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_ mux_top_ipin_1.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR bottom_grid_pin_1_ sky130_fd_sc_hd__buf_4
X_68_ chanx_left_in[11] VGND VGND VPWR VPWR chanx_right_out[11] sky130_fd_sc_hd__buf_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_5.mux_l1_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_3_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_6.mux_l2_in_2_ chanx_left_in[19] chanx_right_in[11] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_1.mux_l3_in_0_ mux_top_ipin_1.mux_l2_in_1_/X mux_top_ipin_1.mux_l2_in_0_/X
+ mux_top_ipin_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_15.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_13.mux_l2_in_3_ _29_/HI chanx_right_in[18] mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_1.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_2.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_ipin_15.mux_l2_in_2__A1 chanx_right_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_1.mux_l2_in_1_ chanx_left_in[6] chanx_right_in[2] mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_11.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_12.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A0 chanx_right_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_top_ipin_8.mux_l2_in_3__A1 chanx_right_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l4_in_0_ mux_top_ipin_13.mux_l3_in_1_/X mux_top_ipin_13.mux_l3_in_0_/X
+ mux_top_ipin_13.mux_l4_in_0_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l4_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_ipin_7.mux_l1_in_0__A0 chanx_right_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_ prog_clk_0_FTB00/X mux_top_ipin_8.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_ipin_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_ipin_6.mux_l3_in_0_ mux_top_ipin_6.mux_l2_in_1_/X mux_top_ipin_6.mux_l2_in_0_/X
+ mux_top_ipin_6.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_6.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_ipin_13.mux_l3_in_1_ mux_top_ipin_13.mux_l2_in_3_/X mux_top_ipin_13.mux_l2_in_2_/X
+ mux_top_ipin_13.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_ipin_13.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_10.mux_l2_in_2__A0 chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_4.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_5.mux_l1_in_0_/S sky130_fd_sc_hd__dfxtp_1
X_67_ chanx_left_in[10] VGND VGND VPWR VPWR chanx_right_out[10] sky130_fd_sc_hd__buf_2
Xmux_top_ipin_6.mux_l2_in_1_ chanx_left_in[11] chanx_right_in[3] mux_top_ipin_6.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_ipin_5.mux_l2_in_1__A0 chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_ prog_clk_0_FTB00/X mux_top_ipin_14.mux_l4_in_0_/S
+ VGND VGND VPWR VPWR mux_top_ipin_15.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND
+ VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_ipin_13.mux_l2_in_2_ chanx_left_in[18] chanx_right_in[10] mux_top_ipin_13.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_13.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_ipin_1.mux_l2_in_0_ chanx_left_in[2] mux_top_ipin_1.mux_l1_in_0_/X mux_top_ipin_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_ipin_1.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_ipin_12.mux_l1_in_1__A1 chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1__CLK prog_clk_0_FTB00/X VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

